module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 ;
  assign n256 = ( x106 & ~x124 ) | ( x106 & x182 ) | ( ~x124 & x182 ) ;
  assign n257 = ( x102 & ~x137 ) | ( x102 & x251 ) | ( ~x137 & x251 ) ;
  assign n258 = x213 ^ x195 ^ x104 ;
  assign n259 = x130 ^ x82 ^ x77 ;
  assign n260 = x144 & x233 ;
  assign n261 = n260 ^ x130 ^ 1'b0 ;
  assign n262 = x226 ^ x162 ^ x9 ;
  assign n263 = x68 ^ x1 ^ 1'b0 ;
  assign n264 = x116 & n263 ;
  assign n265 = x82 ^ x69 ^ 1'b0 ;
  assign n266 = x147 & n265 ;
  assign n267 = x44 & x128 ;
  assign n268 = ~x149 & n267 ;
  assign n269 = ( x10 & ~x228 ) | ( x10 & n264 ) | ( ~x228 & n264 ) ;
  assign n270 = x86 & x90 ;
  assign n271 = ~x189 & n270 ;
  assign n272 = x252 ^ x183 ^ x151 ;
  assign n273 = x105 & x231 ;
  assign n274 = n273 ^ x5 ^ 1'b0 ;
  assign n275 = x122 & ~n274 ;
  assign n276 = n275 ^ x59 ^ 1'b0 ;
  assign n277 = ( x0 & x36 ) | ( x0 & ~x180 ) | ( x36 & ~x180 ) ;
  assign n278 = x8 & x53 ;
  assign n279 = ~n277 & n278 ;
  assign n280 = x224 ^ x6 ^ 1'b0 ;
  assign n281 = ( x51 & ~x199 ) | ( x51 & x247 ) | ( ~x199 & x247 ) ;
  assign n282 = ( x82 & ~x161 ) | ( x82 & n281 ) | ( ~x161 & n281 ) ;
  assign n283 = x77 & x174 ;
  assign n284 = ~x81 & n283 ;
  assign n285 = ( x60 & x152 ) | ( x60 & n284 ) | ( x152 & n284 ) ;
  assign n286 = x2 & x246 ;
  assign n287 = n286 ^ x124 ^ 1'b0 ;
  assign n288 = x30 & x182 ;
  assign n289 = ~x87 & n288 ;
  assign n290 = x244 ^ x87 ^ 1'b0 ;
  assign n291 = x231 ^ x80 ^ 1'b0 ;
  assign n292 = x186 ^ x96 ^ 1'b0 ;
  assign n293 = x126 & n292 ;
  assign n294 = x39 & ~x211 ;
  assign n295 = ( x0 & ~x51 ) | ( x0 & x182 ) | ( ~x51 & x182 ) ;
  assign n296 = x156 & n295 ;
  assign n297 = n296 ^ x77 ^ 1'b0 ;
  assign n298 = x2 & ~n297 ;
  assign n299 = n298 ^ x146 ^ 1'b0 ;
  assign n300 = x243 & ~n299 ;
  assign n301 = n300 ^ x200 ^ 1'b0 ;
  assign n302 = x85 ^ x64 ^ 1'b0 ;
  assign n303 = n257 & n302 ;
  assign n304 = x132 & n303 ;
  assign n305 = ~x4 & n304 ;
  assign n306 = ( x5 & x61 ) | ( x5 & ~x130 ) | ( x61 & ~x130 ) ;
  assign n307 = x228 ^ x182 ^ 1'b0 ;
  assign n308 = x60 ^ x23 ^ 1'b0 ;
  assign n309 = x64 & n308 ;
  assign n310 = ( ~x0 & x141 ) | ( ~x0 & n309 ) | ( x141 & n309 ) ;
  assign n311 = x189 ^ x121 ^ x33 ;
  assign n312 = n311 ^ x64 ^ 1'b0 ;
  assign n313 = x222 & ~n312 ;
  assign n314 = x201 ^ x37 ^ x2 ;
  assign n315 = ( ~x150 & x250 ) | ( ~x150 & x253 ) | ( x250 & x253 ) ;
  assign n316 = n315 ^ x220 ^ x36 ;
  assign n317 = n316 ^ x174 ^ x78 ;
  assign n318 = ( ~x122 & n314 ) | ( ~x122 & n317 ) | ( n314 & n317 ) ;
  assign n319 = x226 ^ x195 ^ 1'b0 ;
  assign n320 = x201 & n319 ;
  assign n321 = ( x30 & n282 ) | ( x30 & ~n320 ) | ( n282 & ~n320 ) ;
  assign n322 = n307 ^ x200 ^ x131 ;
  assign n323 = x149 & ~n271 ;
  assign n324 = n323 ^ x170 ^ 1'b0 ;
  assign n325 = ( ~x17 & x87 ) | ( ~x17 & n324 ) | ( x87 & n324 ) ;
  assign n326 = n258 ^ x226 ^ x0 ;
  assign n327 = ~x247 & n326 ;
  assign n328 = x129 ^ x1 ^ 1'b0 ;
  assign n329 = x57 & n328 ;
  assign n330 = n309 ^ x149 ^ x134 ;
  assign n331 = ( x21 & n329 ) | ( x21 & n330 ) | ( n329 & n330 ) ;
  assign n332 = x116 & n331 ;
  assign n333 = ( ~x86 & x157 ) | ( ~x86 & x170 ) | ( x157 & x170 ) ;
  assign n334 = ~x114 & x226 ;
  assign n335 = n334 ^ n326 ^ x85 ;
  assign n336 = n316 ^ x197 ^ x132 ;
  assign n337 = ( x7 & ~x208 ) | ( x7 & x210 ) | ( ~x208 & x210 ) ;
  assign n338 = n336 ^ n333 ^ 1'b0 ;
  assign n339 = x16 & n338 ;
  assign n340 = ~x65 & n339 ;
  assign n341 = x235 & x242 ;
  assign n342 = x136 ^ x40 ^ 1'b0 ;
  assign n343 = x84 & n342 ;
  assign n344 = n343 ^ x99 ^ 1'b0 ;
  assign n345 = x129 & n344 ;
  assign n346 = n309 ^ x228 ^ x40 ;
  assign n347 = n274 ^ x253 ^ 1'b0 ;
  assign n348 = x88 & ~n347 ;
  assign n352 = ~x83 & x252 ;
  assign n349 = x9 & x76 ;
  assign n350 = ~x178 & n349 ;
  assign n351 = x165 & ~n350 ;
  assign n353 = n352 ^ n351 ^ 1'b0 ;
  assign n354 = x105 & n322 ;
  assign n355 = ( ~x108 & x191 ) | ( ~x108 & x247 ) | ( x191 & x247 ) ;
  assign n356 = x131 & ~n284 ;
  assign n357 = ~x9 & n356 ;
  assign n358 = ( ~x38 & x200 ) | ( ~x38 & x241 ) | ( x200 & x241 ) ;
  assign n359 = n290 & n358 ;
  assign n360 = n357 & n359 ;
  assign n361 = x224 & n360 ;
  assign n362 = x127 ^ x29 ^ x11 ;
  assign n363 = n362 ^ x186 ^ x47 ;
  assign n364 = n363 ^ x234 ^ 1'b0 ;
  assign n365 = x85 & n364 ;
  assign n366 = ( x95 & ~x128 ) | ( x95 & x135 ) | ( ~x128 & x135 ) ;
  assign n367 = ( ~x61 & x222 ) | ( ~x61 & x225 ) | ( x222 & x225 ) ;
  assign n368 = ( ~x113 & x171 ) | ( ~x113 & x209 ) | ( x171 & x209 ) ;
  assign n369 = n367 & n368 ;
  assign n370 = ~n366 & n369 ;
  assign n371 = x70 & x212 ;
  assign n372 = ~x45 & n371 ;
  assign n373 = ( x26 & x118 ) | ( x26 & ~x120 ) | ( x118 & ~x120 ) ;
  assign n376 = ( ~x239 & n279 ) | ( ~x239 & n329 ) | ( n279 & n329 ) ;
  assign n377 = n376 ^ x217 ^ 1'b0 ;
  assign n378 = x74 & ~n377 ;
  assign n374 = ( ~x15 & x234 ) | ( ~x15 & n293 ) | ( x234 & n293 ) ;
  assign n375 = x1 & n374 ;
  assign n379 = n378 ^ n375 ^ 1'b0 ;
  assign n380 = n262 ^ n259 ^ x208 ;
  assign n381 = n380 ^ n256 ^ x216 ;
  assign n382 = ( x133 & x254 ) | ( x133 & ~n381 ) | ( x254 & ~n381 ) ;
  assign n383 = x68 & x131 ;
  assign n384 = ~x254 & n383 ;
  assign n385 = x20 & ~n297 ;
  assign n386 = n385 ^ x189 ^ 1'b0 ;
  assign n387 = x149 & x197 ;
  assign n388 = ~x47 & n387 ;
  assign n389 = ( ~n284 & n333 ) | ( ~n284 & n388 ) | ( n333 & n388 ) ;
  assign n390 = n321 ^ x209 ^ 1'b0 ;
  assign n391 = x157 & n390 ;
  assign n392 = n280 ^ x228 ^ x81 ;
  assign n393 = x72 & ~n376 ;
  assign n394 = ( x126 & ~x197 ) | ( x126 & n368 ) | ( ~x197 & n368 ) ;
  assign n395 = n367 & n394 ;
  assign n396 = ~n307 & n395 ;
  assign n397 = ( x2 & x49 ) | ( x2 & ~x200 ) | ( x49 & ~x200 ) ;
  assign n398 = n397 ^ n368 ^ x109 ;
  assign n399 = n334 ^ n313 ^ 1'b0 ;
  assign n400 = x25 & n399 ;
  assign n401 = n378 & n400 ;
  assign n402 = ~x201 & n401 ;
  assign n403 = x158 & ~x214 ;
  assign n404 = n403 ^ n374 ^ n346 ;
  assign n405 = n388 ^ n366 ^ x79 ;
  assign n406 = ( x14 & x26 ) | ( x14 & ~x64 ) | ( x26 & ~x64 ) ;
  assign n407 = n406 ^ x21 ^ 1'b0 ;
  assign n408 = x252 & n407 ;
  assign n409 = ~x159 & n408 ;
  assign n412 = x164 & n264 ;
  assign n413 = ~x216 & n412 ;
  assign n411 = x11 & ~n314 ;
  assign n414 = n413 ^ n411 ^ 1'b0 ;
  assign n415 = x166 & x193 ;
  assign n416 = ~n414 & n415 ;
  assign n417 = ( x51 & ~x183 ) | ( x51 & x231 ) | ( ~x183 & x231 ) ;
  assign n418 = n282 & n417 ;
  assign n419 = n416 & n418 ;
  assign n410 = x144 ^ x12 ^ x10 ;
  assign n420 = n419 ^ n410 ^ x102 ;
  assign n421 = n320 & n420 ;
  assign n422 = x130 & n389 ;
  assign n423 = ~x68 & n422 ;
  assign n424 = ~n360 & n419 ;
  assign n425 = n424 ^ x8 ^ 1'b0 ;
  assign n426 = x11 & ~n425 ;
  assign n428 = ( x72 & x90 ) | ( x72 & ~x236 ) | ( x90 & ~x236 ) ;
  assign n427 = x186 & ~n361 ;
  assign n429 = n428 ^ n427 ^ 1'b0 ;
  assign n430 = n326 ^ x43 ^ 1'b0 ;
  assign n431 = n430 ^ x170 ^ x13 ;
  assign n432 = n431 ^ x217 ^ x67 ;
  assign n433 = x246 ^ x170 ^ 1'b0 ;
  assign n434 = ~n432 & n433 ;
  assign n435 = ( x9 & ~x93 ) | ( x9 & x172 ) | ( ~x93 & x172 ) ;
  assign n436 = ( ~x184 & x236 ) | ( ~x184 & n317 ) | ( x236 & n317 ) ;
  assign n437 = x232 ^ x47 ^ 1'b0 ;
  assign n438 = x161 & n437 ;
  assign n443 = ( x60 & n314 ) | ( x60 & n416 ) | ( n314 & n416 ) ;
  assign n440 = x1 & x251 ;
  assign n441 = n440 ^ x112 ^ 1'b0 ;
  assign n442 = x242 & ~n441 ;
  assign n444 = n443 ^ n442 ^ 1'b0 ;
  assign n439 = n294 & ~n370 ;
  assign n445 = n444 ^ n439 ^ 1'b0 ;
  assign n446 = ( x10 & ~x152 ) | ( x10 & x207 ) | ( ~x152 & x207 ) ;
  assign n447 = n446 ^ x252 ^ 1'b0 ;
  assign n449 = ( x46 & x67 ) | ( x46 & ~x211 ) | ( x67 & ~x211 ) ;
  assign n448 = n345 ^ n310 ^ x221 ;
  assign n450 = n449 ^ n448 ^ n317 ;
  assign n451 = x184 & ~n305 ;
  assign n452 = n451 ^ x141 ^ 1'b0 ;
  assign n453 = n309 & ~n452 ;
  assign n454 = n453 ^ n409 ^ 1'b0 ;
  assign n455 = x132 & x195 ;
  assign n456 = n454 & n455 ;
  assign n457 = n456 ^ x122 ^ 1'b0 ;
  assign n458 = x147 & n389 ;
  assign n459 = n458 ^ n346 ^ 1'b0 ;
  assign n460 = x36 & ~n413 ;
  assign n461 = n287 & n460 ;
  assign n462 = ( x54 & n416 ) | ( x54 & n461 ) | ( n416 & n461 ) ;
  assign n463 = x149 & n367 ;
  assign n464 = ~n317 & n463 ;
  assign n465 = n413 | n464 ;
  assign n466 = n465 ^ x158 ^ 1'b0 ;
  assign n467 = ~n462 & n466 ;
  assign n468 = n467 ^ n334 ^ 1'b0 ;
  assign n469 = n468 ^ n332 ^ x242 ;
  assign n470 = x235 & ~n303 ;
  assign n471 = x28 & ~x95 ;
  assign n472 = x242 & ~n471 ;
  assign n473 = n472 ^ x143 ^ 1'b0 ;
  assign n474 = ~x76 & x196 ;
  assign n475 = n269 ^ x223 ^ x16 ;
  assign n476 = n314 | n475 ;
  assign n477 = x225 & n476 ;
  assign n478 = n477 ^ x47 ^ 1'b0 ;
  assign n479 = ~n474 & n478 ;
  assign n480 = n462 ^ x132 ^ x85 ;
  assign n481 = ( ~x138 & x186 ) | ( ~x138 & x243 ) | ( x186 & x243 ) ;
  assign n482 = ( ~x171 & x250 ) | ( ~x171 & n481 ) | ( x250 & n481 ) ;
  assign n483 = n482 ^ x117 ^ 1'b0 ;
  assign n486 = ( x125 & ~x135 ) | ( x125 & x240 ) | ( ~x135 & x240 ) ;
  assign n484 = x38 & x201 ;
  assign n485 = n484 ^ x125 ^ 1'b0 ;
  assign n487 = n486 ^ n485 ^ 1'b0 ;
  assign n488 = ( x22 & x149 ) | ( x22 & ~x209 ) | ( x149 & ~x209 ) ;
  assign n489 = x167 ^ x54 ^ 1'b0 ;
  assign n490 = x112 & n489 ;
  assign n497 = x131 ^ x52 ^ x41 ;
  assign n491 = ( ~x132 & x177 ) | ( ~x132 & x189 ) | ( x177 & x189 ) ;
  assign n492 = ( x16 & ~x25 ) | ( x16 & x203 ) | ( ~x25 & x203 ) ;
  assign n493 = n492 ^ x141 ^ x33 ;
  assign n494 = n491 & ~n493 ;
  assign n495 = n494 ^ x246 ^ 1'b0 ;
  assign n496 = n495 ^ x254 ^ x131 ;
  assign n498 = n497 ^ n496 ^ 1'b0 ;
  assign n499 = n490 & ~n498 ;
  assign n500 = ( x35 & ~x118 ) | ( x35 & n499 ) | ( ~x118 & n499 ) ;
  assign n508 = n268 ^ x150 ^ x125 ;
  assign n509 = x98 & n508 ;
  assign n510 = ~x241 & n509 ;
  assign n501 = x171 & x208 ;
  assign n502 = ~x253 & n501 ;
  assign n503 = n502 ^ x101 ^ x64 ;
  assign n504 = ( ~x57 & n346 ) | ( ~x57 & n503 ) | ( n346 & n503 ) ;
  assign n505 = n504 ^ n271 ^ 1'b0 ;
  assign n506 = x65 & n505 ;
  assign n507 = x201 & n506 ;
  assign n511 = n510 ^ n507 ^ 1'b0 ;
  assign n512 = n500 ^ x178 ^ x155 ;
  assign n513 = x50 & x204 ;
  assign n514 = n513 ^ x112 ^ 1'b0 ;
  assign n515 = n514 ^ n502 ^ n340 ;
  assign n516 = ( x9 & x13 ) | ( x9 & ~x41 ) | ( x13 & ~x41 ) ;
  assign n517 = ~n430 & n516 ;
  assign n518 = n517 ^ x33 ^ 1'b0 ;
  assign n519 = n373 & n400 ;
  assign n520 = n519 ^ n261 ^ 1'b0 ;
  assign n521 = x175 & ~x186 ;
  assign n522 = n521 ^ x98 ^ 1'b0 ;
  assign n523 = x108 & n522 ;
  assign n524 = ( x106 & x157 ) | ( x106 & ~n523 ) | ( x157 & ~n523 ) ;
  assign n525 = x10 & n256 ;
  assign n526 = ~x153 & n525 ;
  assign n527 = n526 ^ n345 ^ 1'b0 ;
  assign n528 = x150 & ~n527 ;
  assign n529 = x170 & n528 ;
  assign n530 = n495 & n529 ;
  assign n531 = x93 & n434 ;
  assign n532 = n531 ^ x176 ^ 1'b0 ;
  assign n533 = n532 ^ n282 ^ x218 ;
  assign n534 = ( ~x41 & x154 ) | ( ~x41 & n533 ) | ( x154 & n533 ) ;
  assign n535 = x220 & x248 ;
  assign n536 = ~x2 & n535 ;
  assign n539 = x23 & x176 ;
  assign n540 = n539 ^ x236 ^ 1'b0 ;
  assign n541 = ~x39 & n331 ;
  assign n542 = ( ~x135 & n540 ) | ( ~x135 & n541 ) | ( n540 & n541 ) ;
  assign n537 = x85 ^ x9 ^ x8 ;
  assign n538 = n357 | n537 ;
  assign n543 = n542 ^ n538 ^ 1'b0 ;
  assign n544 = ( x32 & ~x243 ) | ( x32 & n382 ) | ( ~x243 & n382 ) ;
  assign n549 = x99 & x226 ;
  assign n550 = ~x246 & n549 ;
  assign n548 = x253 ^ x222 ^ x189 ;
  assign n547 = x188 ^ x29 ^ x23 ;
  assign n551 = n550 ^ n548 ^ n547 ;
  assign n552 = n551 ^ n446 ^ n388 ;
  assign n545 = ( x198 & x207 ) | ( x198 & ~n516 ) | ( x207 & ~n516 ) ;
  assign n546 = x196 & n545 ;
  assign n553 = n552 ^ n546 ^ 1'b0 ;
  assign n554 = n365 ^ x161 ^ x113 ;
  assign n555 = ( ~x23 & x36 ) | ( ~x23 & n495 ) | ( x36 & n495 ) ;
  assign n556 = x66 ^ x49 ^ 1'b0 ;
  assign n557 = n556 ^ x51 ^ 1'b0 ;
  assign n558 = x27 & n557 ;
  assign n559 = x132 & x173 ;
  assign n560 = n559 ^ x60 ^ 1'b0 ;
  assign n561 = n560 ^ x204 ^ x163 ;
  assign n562 = ~x153 & x222 ;
  assign n563 = x1 & x19 ;
  assign n564 = ~n562 & n563 ;
  assign n565 = x228 & x251 ;
  assign n566 = n565 ^ x62 ^ 1'b0 ;
  assign n567 = x191 ^ x130 ^ 1'b0 ;
  assign n568 = ~n566 & n567 ;
  assign n570 = ~x33 & x207 ;
  assign n571 = x217 ^ x37 ^ 1'b0 ;
  assign n572 = ~n570 & n571 ;
  assign n569 = ~n325 & n524 ;
  assign n573 = n572 ^ n569 ^ 1'b0 ;
  assign n574 = ( x84 & ~n537 ) | ( x84 & n573 ) | ( ~n537 & n573 ) ;
  assign n575 = ~x219 & n368 ;
  assign n576 = ( x91 & x210 ) | ( x91 & n526 ) | ( x210 & n526 ) ;
  assign n577 = ( ~x200 & n575 ) | ( ~x200 & n576 ) | ( n575 & n576 ) ;
  assign n578 = ( x90 & ~x136 ) | ( x90 & x232 ) | ( ~x136 & x232 ) ;
  assign n579 = ( x96 & n274 ) | ( x96 & n306 ) | ( n274 & n306 ) ;
  assign n580 = ( n417 & ~n578 ) | ( n417 & n579 ) | ( ~n578 & n579 ) ;
  assign n581 = x248 & ~n580 ;
  assign n582 = x42 & x164 ;
  assign n583 = ~x76 & n582 ;
  assign n584 = ~x67 & x110 ;
  assign n585 = n584 ^ n566 ^ x213 ;
  assign n586 = ( x9 & ~x31 ) | ( x9 & n585 ) | ( ~x31 & n585 ) ;
  assign n589 = x74 & x102 ;
  assign n590 = ~x185 & n589 ;
  assign n587 = n491 ^ x135 ^ x111 ;
  assign n588 = x220 & ~n587 ;
  assign n591 = n590 ^ n588 ^ 1'b0 ;
  assign n598 = x199 & ~n259 ;
  assign n592 = n428 ^ x244 ^ 1'b0 ;
  assign n593 = x39 & n592 ;
  assign n594 = ( n363 & n432 ) | ( n363 & ~n593 ) | ( n432 & ~n593 ) ;
  assign n595 = ( x195 & ~n410 ) | ( x195 & n594 ) | ( ~n410 & n594 ) ;
  assign n596 = n595 ^ x238 ^ 1'b0 ;
  assign n597 = n320 & n596 ;
  assign n599 = n598 ^ n597 ^ 1'b0 ;
  assign n600 = n348 & n599 ;
  assign n601 = n591 & n600 ;
  assign n602 = ~x207 & n601 ;
  assign n603 = x151 ^ x10 ^ 1'b0 ;
  assign n604 = x213 & n603 ;
  assign n605 = ( ~n261 & n410 ) | ( ~n261 & n604 ) | ( n410 & n604 ) ;
  assign n606 = ~n429 & n605 ;
  assign n607 = ~x246 & n606 ;
  assign n608 = ~x20 & x96 ;
  assign n609 = n335 ^ x234 ^ x133 ;
  assign n610 = x58 & ~n609 ;
  assign n611 = n610 ^ x32 ^ 1'b0 ;
  assign n612 = n447 | n611 ;
  assign n613 = n612 ^ n355 ^ 1'b0 ;
  assign n614 = ( x191 & n608 ) | ( x191 & n613 ) | ( n608 & n613 ) ;
  assign n615 = ( x42 & x98 ) | ( x42 & ~n486 ) | ( x98 & ~n486 ) ;
  assign n616 = n536 | n615 ;
  assign n617 = n545 ^ n365 ^ x120 ;
  assign n618 = n617 ^ x227 ^ x133 ;
  assign n619 = ( x20 & ~x143 ) | ( x20 & n374 ) | ( ~x143 & n374 ) ;
  assign n624 = x30 & x215 ;
  assign n625 = n624 ^ x173 ^ 1'b0 ;
  assign n626 = ( x226 & ~n322 ) | ( x226 & n625 ) | ( ~n322 & n625 ) ;
  assign n627 = n626 ^ x6 ^ 1'b0 ;
  assign n620 = x124 & ~n419 ;
  assign n621 = ~x182 & n620 ;
  assign n622 = x247 & ~n621 ;
  assign n623 = n622 ^ x117 ^ 1'b0 ;
  assign n628 = n627 ^ n623 ^ 1'b0 ;
  assign n629 = n619 & ~n628 ;
  assign n630 = n508 ^ x114 ^ 1'b0 ;
  assign n631 = n629 & n630 ;
  assign n632 = ( ~n341 & n495 ) | ( ~n341 & n631 ) | ( n495 & n631 ) ;
  assign n633 = ( x218 & ~x229 ) | ( x218 & x232 ) | ( ~x229 & x232 ) ;
  assign n634 = ( x144 & ~x253 ) | ( x144 & n261 ) | ( ~x253 & n261 ) ;
  assign n635 = x112 & ~n634 ;
  assign n636 = ~n633 & n635 ;
  assign n637 = n636 ^ n572 ^ n350 ;
  assign n638 = x21 & x36 ;
  assign n639 = n638 ^ x124 ^ 1'b0 ;
  assign n640 = n639 ^ n587 ^ n487 ;
  assign n641 = x36 & n640 ;
  assign n642 = n637 & n641 ;
  assign n643 = n585 ^ n393 ^ x171 ;
  assign n644 = ( ~x12 & x237 ) | ( ~x12 & x245 ) | ( x237 & x245 ) ;
  assign n645 = ~n643 & n644 ;
  assign n646 = x32 & x57 ;
  assign n647 = ~x205 & n646 ;
  assign n648 = n647 ^ x101 ^ x64 ;
  assign n649 = ( ~x115 & x138 ) | ( ~x115 & n541 ) | ( x138 & n541 ) ;
  assign n650 = ( ~n368 & n578 ) | ( ~n368 & n649 ) | ( n578 & n649 ) ;
  assign n651 = n650 ^ x51 ^ 1'b0 ;
  assign n652 = ~n396 & n651 ;
  assign n653 = x149 & n652 ;
  assign n654 = n653 ^ n587 ^ 1'b0 ;
  assign n655 = n654 ^ x235 ^ 1'b0 ;
  assign n656 = n648 & n655 ;
  assign n657 = n355 ^ n330 ^ 1'b0 ;
  assign n659 = x75 & ~n360 ;
  assign n658 = x21 & n392 ;
  assign n660 = n659 ^ n658 ^ 1'b0 ;
  assign n662 = n548 ^ n441 ^ x176 ;
  assign n661 = x177 & n648 ;
  assign n663 = n662 ^ n661 ^ 1'b0 ;
  assign n664 = n663 ^ n441 ^ 1'b0 ;
  assign n665 = n619 & ~n664 ;
  assign n666 = ( n282 & n406 ) | ( n282 & ~n665 ) | ( n406 & ~n665 ) ;
  assign n667 = n521 ^ x227 ^ 1'b0 ;
  assign n668 = x204 & n667 ;
  assign n669 = n547 ^ x99 ^ 1'b0 ;
  assign n670 = ~n487 & n490 ;
  assign n671 = n670 ^ x236 ^ 1'b0 ;
  assign n672 = x54 & ~n671 ;
  assign n673 = n672 ^ n591 ^ 1'b0 ;
  assign n674 = n634 ^ x7 ^ 1'b0 ;
  assign n675 = n578 & ~n674 ;
  assign n676 = ( ~x109 & x141 ) | ( ~x109 & n675 ) | ( x141 & n675 ) ;
  assign n677 = ~n310 & n676 ;
  assign n678 = n677 ^ n432 ^ x111 ;
  assign n679 = x253 ^ x234 ^ x137 ;
  assign n680 = n360 ^ n258 ^ x106 ;
  assign n681 = ( x147 & n679 ) | ( x147 & n680 ) | ( n679 & n680 ) ;
  assign n682 = n310 & n503 ;
  assign n683 = x234 ^ x171 ^ x96 ;
  assign n684 = n683 ^ x95 ^ 1'b0 ;
  assign n685 = n552 & ~n684 ;
  assign n686 = ~n682 & n685 ;
  assign n687 = n544 ^ x246 ^ x203 ;
  assign n688 = n343 | n462 ;
  assign n689 = n617 ^ n616 ^ x121 ;
  assign n690 = ( ~x56 & n379 ) | ( ~x56 & n481 ) | ( n379 & n481 ) ;
  assign n691 = x28 & ~n271 ;
  assign n692 = n691 ^ x96 ^ 1'b0 ;
  assign n693 = ( x228 & n690 ) | ( x228 & n692 ) | ( n690 & n692 ) ;
  assign n697 = x13 & x27 ;
  assign n698 = ~n294 & n697 ;
  assign n699 = n482 ^ n380 ^ x250 ;
  assign n700 = ( x20 & ~x25 ) | ( x20 & n399 ) | ( ~x25 & n399 ) ;
  assign n701 = n699 & ~n700 ;
  assign n702 = n698 & n701 ;
  assign n694 = n663 ^ x143 ^ 1'b0 ;
  assign n695 = x184 & n694 ;
  assign n696 = n503 & n695 ;
  assign n703 = n702 ^ n696 ^ 1'b0 ;
  assign n704 = n627 ^ x117 ^ 1'b0 ;
  assign n705 = n429 ^ x34 ^ 1'b0 ;
  assign n706 = n380 | n705 ;
  assign n707 = ( n264 & n704 ) | ( n264 & n706 ) | ( n704 & n706 ) ;
  assign n708 = n703 & n707 ;
  assign n709 = n708 ^ n586 ^ 1'b0 ;
  assign n710 = x204 ^ x27 ^ 1'b0 ;
  assign n711 = x140 & n710 ;
  assign n712 = x104 & n711 ;
  assign n713 = n536 & n712 ;
  assign n714 = x78 & n406 ;
  assign n715 = n714 ^ x21 ^ 1'b0 ;
  assign n716 = ( x220 & ~x251 ) | ( x220 & n479 ) | ( ~x251 & n479 ) ;
  assign n717 = ~n715 & n716 ;
  assign n718 = n717 ^ n337 ^ 1'b0 ;
  assign n719 = x115 & ~n718 ;
  assign n720 = n719 ^ x89 ^ 1'b0 ;
  assign n721 = x3 & n266 ;
  assign n722 = n721 ^ x33 ^ 1'b0 ;
  assign n723 = n297 | n722 ;
  assign n724 = n723 ^ x122 ^ x107 ;
  assign n725 = ( n353 & n378 ) | ( n353 & ~n724 ) | ( n378 & ~n724 ) ;
  assign n726 = n276 ^ x127 ^ 1'b0 ;
  assign n727 = n722 | n726 ;
  assign n728 = x94 | n727 ;
  assign n729 = x100 & n294 ;
  assign n730 = n729 ^ n315 ^ 1'b0 ;
  assign n731 = n730 ^ n623 ^ n548 ;
  assign n732 = n731 ^ n631 ^ x59 ;
  assign n733 = x236 & n374 ;
  assign n734 = ( ~x54 & x175 ) | ( ~x54 & n542 ) | ( x175 & n542 ) ;
  assign n735 = x157 & ~n305 ;
  assign n736 = n735 ^ x124 ^ 1'b0 ;
  assign n737 = ( ~n604 & n734 ) | ( ~n604 & n736 ) | ( n734 & n736 ) ;
  assign n738 = ( ~n325 & n426 ) | ( ~n325 & n737 ) | ( n426 & n737 ) ;
  assign n739 = x132 & ~n495 ;
  assign n740 = x228 ^ x213 ^ 1'b0 ;
  assign n741 = x252 & n740 ;
  assign n742 = n276 ^ x12 ^ 1'b0 ;
  assign n743 = n741 & ~n742 ;
  assign n744 = n743 ^ n279 ^ 1'b0 ;
  assign n745 = ( ~x19 & x96 ) | ( ~x19 & x228 ) | ( x96 & x228 ) ;
  assign n746 = x29 & ~n325 ;
  assign n747 = ~n600 & n746 ;
  assign n748 = n745 & ~n747 ;
  assign n749 = ( n739 & n744 ) | ( n739 & ~n748 ) | ( n744 & ~n748 ) ;
  assign n750 = ( ~x103 & x149 ) | ( ~x103 & n590 ) | ( x149 & n590 ) ;
  assign n751 = ( ~x222 & n257 ) | ( ~x222 & n750 ) | ( n257 & n750 ) ;
  assign n752 = x24 & x139 ;
  assign n753 = ~x112 & n752 ;
  assign n754 = n753 ^ n625 ^ 1'b0 ;
  assign n755 = x43 & n754 ;
  assign n756 = ( ~n259 & n455 ) | ( ~n259 & n542 ) | ( n455 & n542 ) ;
  assign n757 = x247 & n524 ;
  assign n758 = n745 ^ x48 ^ 1'b0 ;
  assign n759 = ( x73 & x90 ) | ( x73 & ~x102 ) | ( x90 & ~x102 ) ;
  assign n760 = x80 ^ x28 ^ 1'b0 ;
  assign n761 = n759 & n760 ;
  assign n762 = n496 & n761 ;
  assign n763 = ~n758 & n762 ;
  assign n767 = x153 ^ x137 ^ x70 ;
  assign n768 = n316 | n767 ;
  assign n764 = n315 ^ x226 ^ x93 ;
  assign n765 = n764 ^ n722 ^ 1'b0 ;
  assign n766 = ( ~x151 & n556 ) | ( ~x151 & n765 ) | ( n556 & n765 ) ;
  assign n769 = n768 ^ n766 ^ n459 ;
  assign n770 = n488 ^ n464 ^ x85 ;
  assign n771 = ( n289 & n406 ) | ( n289 & ~n770 ) | ( n406 & ~n770 ) ;
  assign n772 = x51 & x132 ;
  assign n773 = n772 ^ x212 ^ 1'b0 ;
  assign n774 = ~x171 & n366 ;
  assign n775 = x30 & n408 ;
  assign n776 = n775 ^ n388 ^ 1'b0 ;
  assign n777 = n378 ^ x228 ^ x217 ;
  assign n778 = x241 & ~n777 ;
  assign n779 = ~n776 & n778 ;
  assign n780 = ( x95 & ~x232 ) | ( x95 & n715 ) | ( ~x232 & n715 ) ;
  assign n781 = x102 & ~n532 ;
  assign n782 = n781 ^ n325 ^ 1'b0 ;
  assign n783 = ( ~n496 & n780 ) | ( ~n496 & n782 ) | ( n780 & n782 ) ;
  assign n784 = n779 | n783 ;
  assign n785 = n774 & ~n784 ;
  assign n786 = n419 ^ x83 ^ 1'b0 ;
  assign n787 = n325 | n786 ;
  assign n788 = x4 & n348 ;
  assign n789 = ~x96 & n788 ;
  assign n790 = ( x86 & ~n305 ) | ( x86 & n789 ) | ( ~n305 & n789 ) ;
  assign n791 = n787 & n790 ;
  assign n792 = x31 & ~n791 ;
  assign n793 = n792 ^ x56 ^ 1'b0 ;
  assign n794 = ~n287 & n394 ;
  assign n795 = n794 ^ n578 ^ 1'b0 ;
  assign n796 = n795 ^ n333 ^ x120 ;
  assign n797 = n758 & n796 ;
  assign n798 = ~n665 & n797 ;
  assign n799 = n798 ^ n594 ^ x44 ;
  assign n800 = n389 ^ n354 ^ x121 ;
  assign n801 = x115 & ~n623 ;
  assign n802 = n801 ^ x8 ^ 1'b0 ;
  assign n803 = n551 & ~n621 ;
  assign n804 = n803 ^ n279 ^ 1'b0 ;
  assign n805 = n576 & n804 ;
  assign n806 = n673 & n805 ;
  assign n807 = ( n290 & n334 ) | ( n290 & ~n417 ) | ( n334 & ~n417 ) ;
  assign n808 = n503 ^ x224 ^ 1'b0 ;
  assign n809 = ( x10 & x110 ) | ( x10 & ~n808 ) | ( x110 & ~n808 ) ;
  assign n811 = ~n376 & n490 ;
  assign n812 = n268 & n811 ;
  assign n813 = ( x56 & x141 ) | ( x56 & n812 ) | ( x141 & n812 ) ;
  assign n814 = n813 ^ n537 ^ n376 ;
  assign n810 = n566 ^ n386 ^ x78 ;
  assign n815 = n814 ^ n810 ^ 1'b0 ;
  assign n816 = x64 & n815 ;
  assign n818 = ( x84 & n396 ) | ( x84 & n469 ) | ( n396 & n469 ) ;
  assign n819 = x157 & ~n570 ;
  assign n820 = n818 & n819 ;
  assign n817 = ~n609 & n615 ;
  assign n821 = n820 ^ n817 ^ 1'b0 ;
  assign n824 = x118 & x220 ;
  assign n825 = ~n428 & n824 ;
  assign n826 = n508 | n825 ;
  assign n822 = x115 & n676 ;
  assign n823 = n449 & n822 ;
  assign n827 = n826 ^ n823 ^ 1'b0 ;
  assign n828 = x113 & ~n702 ;
  assign n829 = n828 ^ n550 ^ 1'b0 ;
  assign n831 = ( x147 & ~x187 ) | ( x147 & x243 ) | ( ~x187 & x243 ) ;
  assign n830 = x128 & ~n350 ;
  assign n832 = n831 ^ n830 ^ n767 ;
  assign n833 = x103 & n832 ;
  assign n834 = ~x209 & n833 ;
  assign n835 = x70 & ~x206 ;
  assign n836 = n835 ^ n370 ^ x225 ;
  assign n837 = n396 | n836 ;
  assign n838 = n837 ^ x137 ^ 1'b0 ;
  assign n839 = x149 & n838 ;
  assign n840 = n839 ^ x71 ^ 1'b0 ;
  assign n841 = x62 & ~x111 ;
  assign n842 = n358 & ~n730 ;
  assign n843 = ( n777 & n841 ) | ( n777 & n842 ) | ( n841 & n842 ) ;
  assign n844 = n470 ^ x243 ^ 1'b0 ;
  assign n845 = n419 | n844 ;
  assign n846 = x24 & x93 ;
  assign n847 = ~x209 & n846 ;
  assign n848 = n847 ^ n481 ^ 1'b0 ;
  assign n849 = n657 | n848 ;
  assign n850 = n272 | n849 ;
  assign n851 = n850 ^ n336 ^ 1'b0 ;
  assign n852 = n481 ^ n449 ^ 1'b0 ;
  assign n853 = ~n537 & n852 ;
  assign n854 = x89 & ~n570 ;
  assign n855 = ~x38 & n854 ;
  assign n856 = x116 & n436 ;
  assign n857 = ~n329 & n856 ;
  assign n858 = x175 & x248 ;
  assign n859 = n858 ^ x136 ^ 1'b0 ;
  assign n860 = x216 & ~n310 ;
  assign n861 = ( ~n570 & n859 ) | ( ~n570 & n860 ) | ( n859 & n860 ) ;
  assign n862 = x179 & ~n861 ;
  assign n863 = n857 & n862 ;
  assign n864 = n256 & ~n700 ;
  assign n865 = x44 & x191 ;
  assign n866 = ( x20 & ~x84 ) | ( x20 & x175 ) | ( ~x84 & x175 ) ;
  assign n867 = ~x51 & x224 ;
  assign n868 = ( n470 & ~n689 ) | ( n470 & n867 ) | ( ~n689 & n867 ) ;
  assign n869 = ( n575 & n866 ) | ( n575 & n868 ) | ( n866 & n868 ) ;
  assign n870 = n835 ^ n332 ^ x247 ;
  assign n871 = x46 & n870 ;
  assign n872 = ( n340 & n345 ) | ( n340 & n488 ) | ( n345 & n488 ) ;
  assign n873 = ( x47 & ~x164 ) | ( x47 & n706 ) | ( ~x164 & n706 ) ;
  assign n874 = n294 & ~n446 ;
  assign n875 = n874 ^ n594 ^ n410 ;
  assign n876 = x187 & ~n575 ;
  assign n877 = n876 ^ x247 ^ 1'b0 ;
  assign n878 = n750 | n877 ;
  assign n879 = x160 | n878 ;
  assign n880 = ( ~x71 & n409 ) | ( ~x71 & n879 ) | ( n409 & n879 ) ;
  assign n881 = n880 ^ x43 ^ 1'b0 ;
  assign n882 = x230 & n881 ;
  assign n883 = ~x116 & n882 ;
  assign n885 = ( x164 & x166 ) | ( x164 & n376 ) | ( x166 & n376 ) ;
  assign n884 = ( ~n309 & n830 ) | ( ~n309 & n835 ) | ( n830 & n835 ) ;
  assign n886 = n885 ^ n884 ^ 1'b0 ;
  assign n887 = n886 ^ n682 ^ n329 ;
  assign n888 = n887 ^ x124 ^ 1'b0 ;
  assign n889 = x106 & ~n888 ;
  assign n890 = n313 | n660 ;
  assign n891 = n890 ^ n480 ^ x8 ;
  assign n892 = n587 ^ x190 ^ x115 ;
  assign n893 = ( ~n343 & n516 ) | ( ~n343 & n892 ) | ( n516 & n892 ) ;
  assign n894 = ( x22 & ~x91 ) | ( x22 & n636 ) | ( ~x91 & n636 ) ;
  assign n900 = n812 ^ n461 ^ n293 ;
  assign n897 = n550 | n836 ;
  assign n898 = x232 | n897 ;
  assign n895 = n368 ^ n272 ^ x123 ;
  assign n896 = ~n271 & n895 ;
  assign n899 = n898 ^ n896 ^ 1'b0 ;
  assign n901 = n900 ^ n899 ^ x158 ;
  assign n902 = n884 | n901 ;
  assign n903 = x137 | n902 ;
  assign n904 = ( x72 & ~x210 ) | ( x72 & n767 ) | ( ~x210 & n767 ) ;
  assign n905 = n904 ^ n880 ^ 1'b0 ;
  assign n909 = x205 ^ x140 ^ 1'b0 ;
  assign n910 = n408 & n909 ;
  assign n906 = x6 & ~n380 ;
  assign n907 = n764 & n906 ;
  assign n908 = n613 | n907 ;
  assign n911 = n910 ^ n908 ^ 1'b0 ;
  assign n912 = ~n834 & n911 ;
  assign n913 = x116 & x161 ;
  assign n914 = ~x223 & n913 ;
  assign n915 = n914 ^ x206 ^ x3 ;
  assign n916 = x137 ^ x125 ^ x39 ;
  assign n917 = n916 ^ n388 ^ 1'b0 ;
  assign n918 = ~n647 & n917 ;
  assign n919 = ( x4 & x144 ) | ( x4 & ~n918 ) | ( x144 & ~n918 ) ;
  assign n920 = n915 & n919 ;
  assign n921 = n920 ^ n426 ^ 1'b0 ;
  assign n922 = n590 ^ n475 ^ 1'b0 ;
  assign n923 = x184 & n922 ;
  assign n924 = ~n720 & n923 ;
  assign n925 = ~n665 & n924 ;
  assign n928 = x35 & n604 ;
  assign n929 = ~x59 & n928 ;
  assign n926 = n636 ^ n566 ^ x173 ;
  assign n927 = n311 | n926 ;
  assign n930 = n929 ^ n927 ^ 1'b0 ;
  assign n931 = x112 & x206 ;
  assign n932 = ~x42 & n931 ;
  assign n933 = n408 ^ x152 ^ x16 ;
  assign n934 = ( ~x92 & x149 ) | ( ~x92 & n933 ) | ( x149 & n933 ) ;
  assign n935 = n932 | n934 ;
  assign n936 = n935 ^ n644 ^ 1'b0 ;
  assign n937 = n870 ^ n428 ^ n403 ;
  assign n938 = ( n447 & n545 ) | ( n447 & ~n937 ) | ( n545 & ~n937 ) ;
  assign n939 = ( x127 & ~n400 ) | ( x127 & n938 ) | ( ~n400 & n938 ) ;
  assign n940 = ( x162 & n424 ) | ( x162 & n755 ) | ( n424 & n755 ) ;
  assign n941 = x204 & ~n307 ;
  assign n942 = x165 & x217 ;
  assign n943 = n942 ^ x26 ^ 1'b0 ;
  assign n944 = n631 ^ n500 ^ n424 ;
  assign n945 = x75 & n944 ;
  assign n946 = ~n336 & n945 ;
  assign n947 = ( ~x55 & x189 ) | ( ~x55 & n946 ) | ( x189 & n946 ) ;
  assign n948 = ~n607 & n618 ;
  assign n949 = n947 & n948 ;
  assign n950 = n949 ^ x162 ^ 1'b0 ;
  assign n951 = n921 ^ n777 ^ x164 ;
  assign n953 = ~n380 & n499 ;
  assign n954 = ~x149 & n953 ;
  assign n952 = n291 & ~n330 ;
  assign n955 = n954 ^ n952 ^ n735 ;
  assign n963 = n345 ^ x171 ^ x169 ;
  assign n961 = n835 ^ n715 ^ n352 ;
  assign n958 = x238 & n291 ;
  assign n959 = x197 & n958 ;
  assign n960 = ~x126 & n959 ;
  assign n957 = n537 ^ n338 ^ n280 ;
  assign n962 = n961 ^ n960 ^ n957 ;
  assign n956 = n768 ^ n656 ^ n431 ;
  assign n964 = n963 ^ n962 ^ n956 ;
  assign n965 = n956 ^ x62 ^ 1'b0 ;
  assign n966 = ~n907 & n965 ;
  assign n967 = ( ~x85 & x94 ) | ( ~x85 & n289 ) | ( x94 & n289 ) ;
  assign n968 = x191 ^ x110 ^ 1'b0 ;
  assign n969 = x217 ^ x134 ^ x35 ;
  assign n970 = n969 ^ x243 ^ 1'b0 ;
  assign n971 = n877 | n970 ;
  assign n972 = n968 | n971 ;
  assign n973 = n326 | n972 ;
  assign n974 = n973 ^ x234 ^ x119 ;
  assign n975 = x2 & ~n421 ;
  assign n976 = n975 ^ x105 ^ 1'b0 ;
  assign n977 = ( n827 & n974 ) | ( n827 & ~n976 ) | ( n974 & ~n976 ) ;
  assign n978 = n438 ^ x125 ^ 1'b0 ;
  assign n979 = ~n977 & n978 ;
  assign n980 = ( x15 & ~x128 ) | ( x15 & n295 ) | ( ~x128 & n295 ) ;
  assign n981 = x95 & x218 ;
  assign n982 = n981 ^ x19 ^ 1'b0 ;
  assign n983 = n980 & ~n982 ;
  assign n984 = ( ~n550 & n556 ) | ( ~n550 & n841 ) | ( n556 & n841 ) ;
  assign n987 = ( x4 & n528 ) | ( x4 & n730 ) | ( n528 & n730 ) ;
  assign n986 = x221 & n508 ;
  assign n988 = n987 ^ n986 ^ 1'b0 ;
  assign n985 = ~n379 & n435 ;
  assign n989 = n988 ^ n985 ^ 1'b0 ;
  assign n990 = x48 & ~x117 ;
  assign n991 = n990 ^ n537 ^ 1'b0 ;
  assign n992 = x194 & n991 ;
  assign n993 = n992 ^ n893 ^ n879 ;
  assign n994 = n581 ^ x173 ^ 1'b0 ;
  assign n995 = n392 & ~n994 ;
  assign n996 = n605 ^ x205 ^ x87 ;
  assign n997 = n873 | n996 ;
  assign n998 = ( x151 & x186 ) | ( x151 & n997 ) | ( x186 & n997 ) ;
  assign n999 = x242 & ~n698 ;
  assign n1000 = n999 ^ n555 ^ 1'b0 ;
  assign n1001 = n354 | n1000 ;
  assign n1006 = ( ~x6 & x149 ) | ( ~x6 & n835 ) | ( x149 & n835 ) ;
  assign n1002 = n626 ^ x33 ^ 1'b0 ;
  assign n1003 = x237 & n1002 ;
  assign n1004 = n1003 ^ x156 ^ 1'b0 ;
  assign n1005 = x5 & ~n1004 ;
  assign n1007 = n1006 ^ n1005 ^ 1'b0 ;
  assign n1008 = n444 & n1007 ;
  assign n1009 = n1008 ^ x13 ^ 1'b0 ;
  assign n1010 = ( n413 & n479 ) | ( n413 & ~n548 ) | ( n479 & ~n548 ) ;
  assign n1011 = x106 & ~x130 ;
  assign n1012 = n1011 ^ n937 ^ n747 ;
  assign n1013 = n1010 & ~n1012 ;
  assign n1014 = n1013 ^ n707 ^ 1'b0 ;
  assign n1015 = x91 & x150 ;
  assign n1016 = n1015 ^ n503 ^ 1'b0 ;
  assign n1017 = ( ~n487 & n665 ) | ( ~n487 & n1016 ) | ( n665 & n1016 ) ;
  assign n1018 = x15 & n1017 ;
  assign n1021 = x80 & x145 ;
  assign n1022 = n1021 ^ x147 ^ 1'b0 ;
  assign n1023 = x232 & n295 ;
  assign n1024 = n1023 ^ x209 ^ 1'b0 ;
  assign n1025 = n1022 | n1024 ;
  assign n1026 = n1025 ^ x7 ^ 1'b0 ;
  assign n1019 = x155 & n733 ;
  assign n1020 = n1019 ^ n842 ^ 1'b0 ;
  assign n1027 = n1026 ^ n1020 ^ n504 ;
  assign n1028 = x233 | n1027 ;
  assign n1029 = n1028 ^ n720 ^ x182 ;
  assign n1030 = x211 & ~n403 ;
  assign n1031 = n806 ^ n745 ^ n429 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = n1032 ^ n268 ^ 1'b0 ;
  assign n1034 = n397 & n1033 ;
  assign n1035 = ( ~n264 & n540 ) | ( ~n264 & n579 ) | ( n540 & n579 ) ;
  assign n1036 = n448 | n1035 ;
  assign n1037 = x193 | n350 ;
  assign n1038 = n650 & n1037 ;
  assign n1039 = n693 & n1038 ;
  assign n1040 = ( x39 & n787 ) | ( x39 & n1039 ) | ( n787 & n1039 ) ;
  assign n1041 = n426 ^ x212 ^ 1'b0 ;
  assign n1042 = n809 | n1041 ;
  assign n1043 = ( ~x41 & n481 ) | ( ~x41 & n595 ) | ( n481 & n595 ) ;
  assign n1044 = n1043 ^ n1030 ^ n556 ;
  assign n1045 = n1044 ^ n336 ^ x143 ;
  assign n1046 = n1045 ^ n793 ^ 1'b0 ;
  assign n1047 = n820 ^ n259 ^ x143 ;
  assign n1048 = n346 & n643 ;
  assign n1049 = n864 | n1048 ;
  assign n1050 = n502 | n964 ;
  assign n1051 = n587 ^ n378 ^ x48 ;
  assign n1052 = ( x48 & ~x89 ) | ( x48 & n1051 ) | ( ~x89 & n1051 ) ;
  assign n1053 = ~n1014 & n1050 ;
  assign n1054 = n1010 ^ x166 ^ 1'b0 ;
  assign n1055 = x210 & x222 ;
  assign n1056 = n750 & n1055 ;
  assign n1057 = n1056 ^ n374 ^ x109 ;
  assign n1058 = ~n409 & n1057 ;
  assign n1059 = n1058 ^ x239 ^ 1'b0 ;
  assign n1060 = n1059 ^ x241 ^ 1'b0 ;
  assign n1061 = x26 & ~n1060 ;
  assign n1062 = ~x52 & n1061 ;
  assign n1063 = ( n765 & ~n1054 ) | ( n765 & n1062 ) | ( ~n1054 & n1062 ) ;
  assign n1064 = ( x71 & n495 ) | ( x71 & n825 ) | ( n495 & n825 ) ;
  assign n1066 = ( n271 & n446 ) | ( n271 & n968 ) | ( n446 & n968 ) ;
  assign n1065 = x130 & ~n932 ;
  assign n1067 = n1066 ^ n1065 ^ 1'b0 ;
  assign n1068 = n1064 & n1067 ;
  assign n1069 = x61 & x140 ;
  assign n1070 = n1069 ^ n1057 ^ 1'b0 ;
  assign n1071 = n318 ^ x171 ^ 1'b0 ;
  assign n1072 = x42 & ~n1071 ;
  assign n1073 = ~n877 & n1072 ;
  assign n1074 = n274 & n1073 ;
  assign n1075 = ( x103 & ~n1070 ) | ( x103 & n1074 ) | ( ~n1070 & n1074 ) ;
  assign n1076 = n1020 | n1075 ;
  assign n1077 = x237 | n1076 ;
  assign n1078 = ( x45 & x190 ) | ( x45 & ~x217 ) | ( x190 & ~x217 ) ;
  assign n1079 = n264 & n1078 ;
  assign n1080 = n1079 ^ x19 ^ 1'b0 ;
  assign n1081 = n633 ^ x62 ^ 1'b0 ;
  assign n1082 = n313 ^ x128 ^ 1'b0 ;
  assign n1083 = ~n476 & n1082 ;
  assign n1084 = ( ~x116 & n477 ) | ( ~x116 & n1083 ) | ( n477 & n1083 ) ;
  assign n1085 = n1081 & n1084 ;
  assign n1086 = n1080 & n1085 ;
  assign n1087 = n1086 ^ n938 ^ 1'b0 ;
  assign n1090 = ( ~x5 & x37 ) | ( ~x5 & n734 ) | ( x37 & n734 ) ;
  assign n1089 = x4 & x207 ;
  assign n1091 = n1090 ^ n1089 ^ 1'b0 ;
  assign n1088 = n331 ^ x149 ^ 1'b0 ;
  assign n1092 = n1091 ^ n1088 ^ n838 ;
  assign n1103 = n338 & ~n543 ;
  assign n1104 = ~n337 & n1103 ;
  assign n1105 = x144 & n1104 ;
  assign n1102 = n454 & ~n678 ;
  assign n1098 = n825 ^ n473 ^ x141 ;
  assign n1093 = ( ~x94 & x253 ) | ( ~x94 & n745 ) | ( x253 & n745 ) ;
  assign n1094 = ~n259 & n654 ;
  assign n1095 = n951 & n1094 ;
  assign n1096 = n1084 & ~n1095 ;
  assign n1097 = ~n1093 & n1096 ;
  assign n1099 = n1098 ^ n1097 ^ n262 ;
  assign n1100 = ~n673 & n1099 ;
  assign n1101 = n1100 ^ n413 ^ 1'b0 ;
  assign n1106 = n1105 ^ n1102 ^ n1101 ;
  assign n1107 = n715 ^ n335 ^ x20 ;
  assign n1108 = n594 | n1107 ;
  assign n1109 = n692 ^ n502 ^ n445 ;
  assign n1110 = n366 & n1109 ;
  assign n1111 = n1110 ^ n908 ^ 1'b0 ;
  assign n1112 = ( x158 & n548 ) | ( x158 & n1091 ) | ( n548 & n1091 ) ;
  assign n1113 = x188 ^ x157 ^ 1'b0 ;
  assign n1114 = n995 & ~n1113 ;
  assign n1115 = ~n723 & n1083 ;
  assign n1116 = n448 & n1115 ;
  assign n1117 = ( x73 & x112 ) | ( x73 & n1116 ) | ( x112 & n1116 ) ;
  assign n1118 = n1117 ^ x89 ^ 1'b0 ;
  assign n1119 = n962 ^ x138 ^ 1'b0 ;
  assign n1120 = n783 | n1119 ;
  assign n1121 = ( x224 & ~n294 ) | ( x224 & n554 ) | ( ~n294 & n554 ) ;
  assign n1122 = ~x11 & x38 ;
  assign n1123 = ( n357 & ~n1121 ) | ( n357 & n1122 ) | ( ~n1121 & n1122 ) ;
  assign n1124 = ~n671 & n1123 ;
  assign n1125 = x115 & n1124 ;
  assign n1126 = n1045 ^ x167 ^ 1'b0 ;
  assign n1127 = n718 | n1126 ;
  assign n1128 = n1127 ^ x98 ^ 1'b0 ;
  assign n1129 = n1128 ^ x67 ^ 1'b0 ;
  assign n1130 = n1030 | n1129 ;
  assign n1132 = x181 & n497 ;
  assign n1131 = x12 & ~x121 ;
  assign n1133 = n1132 ^ n1131 ^ 1'b0 ;
  assign n1134 = ( x65 & x85 ) | ( x65 & ~x141 ) | ( x85 & ~x141 ) ;
  assign n1135 = n1134 ^ n741 ^ n636 ;
  assign n1136 = n1135 ^ n268 ^ x253 ;
  assign n1137 = x54 & n423 ;
  assign n1139 = x85 & x205 ;
  assign n1140 = n1139 ^ n281 ^ 1'b0 ;
  assign n1141 = x37 ^ x36 ^ 1'b0 ;
  assign n1142 = ~n1140 & n1141 ;
  assign n1143 = n487 ^ x16 ^ 1'b0 ;
  assign n1144 = n1142 & ~n1143 ;
  assign n1138 = n340 | n976 ;
  assign n1145 = n1144 ^ n1138 ^ 1'b0 ;
  assign n1146 = n1145 ^ x123 ^ 1'b0 ;
  assign n1147 = x115 & n1146 ;
  assign n1148 = n1137 & n1147 ;
  assign n1149 = n682 | n698 ;
  assign n1150 = n1112 ^ n864 ^ x57 ;
  assign n1151 = n317 & n480 ;
  assign n1152 = n1056 & n1151 ;
  assign n1153 = n1152 ^ n552 ^ x27 ;
  assign n1156 = n566 ^ x220 ^ x211 ;
  assign n1154 = n293 ^ x222 ^ x32 ;
  assign n1155 = n796 & ~n1154 ;
  assign n1157 = n1156 ^ n1155 ^ 1'b0 ;
  assign n1158 = n831 & n1157 ;
  assign n1159 = n1064 ^ n618 ^ n584 ;
  assign n1160 = x24 & ~n461 ;
  assign n1161 = n1160 ^ x120 ^ 1'b0 ;
  assign n1162 = n1161 ^ n969 ^ x85 ;
  assign n1163 = ( n461 & ~n497 ) | ( n461 & n734 ) | ( ~n497 & n734 ) ;
  assign n1164 = ( x199 & ~n393 ) | ( x199 & n1163 ) | ( ~n393 & n1163 ) ;
  assign n1165 = n466 & n711 ;
  assign n1166 = x112 & n1062 ;
  assign n1167 = n1165 & n1166 ;
  assign n1168 = ~x91 & n1167 ;
  assign n1169 = ( x104 & ~n1164 ) | ( x104 & n1168 ) | ( ~n1164 & n1168 ) ;
  assign n1177 = x71 & ~n575 ;
  assign n1178 = n1177 ^ x164 ^ 1'b0 ;
  assign n1173 = n1134 ^ n735 ^ n271 ;
  assign n1174 = n1173 ^ x208 ^ x91 ;
  assign n1175 = ( ~x89 & n776 ) | ( ~x89 & n919 ) | ( n776 & n919 ) ;
  assign n1176 = n1174 & n1175 ;
  assign n1179 = n1178 ^ n1176 ^ n671 ;
  assign n1170 = n952 ^ n898 ^ 1'b0 ;
  assign n1171 = x69 & n1170 ;
  assign n1172 = n1026 & n1171 ;
  assign n1180 = n1179 ^ n1172 ^ 1'b0 ;
  assign n1181 = ( x208 & x221 ) | ( x208 & ~n711 ) | ( x221 & ~n711 ) ;
  assign n1182 = n1181 ^ n504 ^ 1'b0 ;
  assign n1183 = n722 | n1182 ;
  assign n1184 = ( x81 & ~n378 ) | ( x81 & n435 ) | ( ~n378 & n435 ) ;
  assign n1185 = n305 | n932 ;
  assign n1186 = n673 & ~n1185 ;
  assign n1187 = n332 & ~n941 ;
  assign n1188 = n367 | n877 ;
  assign n1189 = n526 ^ x232 ^ x41 ;
  assign n1190 = n1189 ^ n444 ^ 1'b0 ;
  assign n1191 = n1188 & n1190 ;
  assign n1192 = x161 & ~n933 ;
  assign n1193 = ~n388 & n1192 ;
  assign n1194 = n1193 ^ n963 ^ 1'b0 ;
  assign n1195 = n1194 ^ x142 ^ 1'b0 ;
  assign n1196 = ~n750 & n1195 ;
  assign n1197 = x137 & ~n1196 ;
  assign n1198 = ( x75 & n1191 ) | ( x75 & ~n1197 ) | ( n1191 & ~n1197 ) ;
  assign n1199 = n583 ^ x184 ^ 1'b0 ;
  assign n1200 = n814 | n835 ;
  assign n1201 = n1200 ^ x189 ^ 1'b0 ;
  assign n1202 = n1070 ^ n1003 ^ n971 ;
  assign n1203 = n1202 ^ n403 ^ 1'b0 ;
  assign n1204 = n1201 & ~n1203 ;
  assign n1205 = n700 ^ x147 ^ 1'b0 ;
  assign n1206 = n867 ^ n520 ^ n370 ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = x68 | n1207 ;
  assign n1209 = ( x112 & n423 ) | ( x112 & n1006 ) | ( n423 & n1006 ) ;
  assign n1210 = n869 ^ n682 ^ 1'b0 ;
  assign n1211 = n723 | n1210 ;
  assign n1212 = ( n892 & ~n1209 ) | ( n892 & n1211 ) | ( ~n1209 & n1211 ) ;
  assign n1213 = n836 ^ n305 ^ 1'b0 ;
  assign n1214 = x174 & n1213 ;
  assign n1215 = n739 ^ n731 ^ 1'b0 ;
  assign n1216 = ~n299 & n1215 ;
  assign n1217 = n1216 ^ n840 ^ n660 ;
  assign n1218 = ( ~n324 & n1214 ) | ( ~n324 & n1217 ) | ( n1214 & n1217 ) ;
  assign n1221 = x169 & n334 ;
  assign n1219 = ( x121 & n317 ) | ( x121 & n495 ) | ( n317 & n495 ) ;
  assign n1220 = ~n715 & n1219 ;
  assign n1222 = n1221 ^ n1220 ^ n470 ;
  assign n1223 = n1187 & ~n1222 ;
  assign n1224 = n795 ^ x5 ^ 1'b0 ;
  assign n1225 = n679 | n1224 ;
  assign n1226 = n1225 ^ n923 ^ n416 ;
  assign n1227 = n1226 ^ n330 ^ 1'b0 ;
  assign n1228 = x221 & n1227 ;
  assign n1231 = x41 & ~x213 ;
  assign n1232 = n1231 ^ n1173 ^ x177 ;
  assign n1229 = n916 ^ n758 ^ x210 ;
  assign n1230 = x235 & n1229 ;
  assign n1233 = n1232 ^ n1230 ^ 1'b0 ;
  assign n1234 = n639 | n1233 ;
  assign n1235 = n1016 & ~n1234 ;
  assign n1236 = x216 ^ x201 ^ x141 ;
  assign n1238 = ~n445 & n644 ;
  assign n1239 = n1238 ^ x200 ^ 1'b0 ;
  assign n1237 = n325 | n1173 ;
  assign n1240 = n1239 ^ n1237 ^ 1'b0 ;
  assign n1241 = x167 ^ x146 ^ x58 ;
  assign n1242 = n966 ^ n333 ^ 1'b0 ;
  assign n1243 = n404 & n1242 ;
  assign n1244 = x106 & x123 ;
  assign n1245 = ( ~x163 & n449 ) | ( ~x163 & n1244 ) | ( n449 & n1244 ) ;
  assign n1246 = n814 | n901 ;
  assign n1247 = ( ~n1007 & n1245 ) | ( ~n1007 & n1246 ) | ( n1245 & n1246 ) ;
  assign n1248 = n921 ^ n365 ^ 1'b0 ;
  assign n1249 = n564 | n1248 ;
  assign n1250 = n625 | n1219 ;
  assign n1251 = n855 | n1250 ;
  assign n1252 = n971 ^ n579 ^ 1'b0 ;
  assign n1253 = x232 & n1252 ;
  assign n1254 = n1253 ^ n732 ^ 1'b0 ;
  assign n1255 = n1254 ^ n849 ^ x117 ;
  assign n1256 = x54 & ~n345 ;
  assign n1257 = n1163 ^ x226 ^ 1'b0 ;
  assign n1258 = n583 | n1257 ;
  assign n1259 = n490 & ~n904 ;
  assign n1260 = n1259 ^ x41 ^ 1'b0 ;
  assign n1261 = ( ~x237 & n1081 ) | ( ~x237 & n1140 ) | ( n1081 & n1140 ) ;
  assign n1262 = n324 | n1261 ;
  assign n1263 = n782 | n1262 ;
  assign n1264 = ( n376 & ~n1260 ) | ( n376 & n1263 ) | ( ~n1260 & n1263 ) ;
  assign n1265 = n587 ^ x8 ^ 1'b0 ;
  assign n1266 = x228 & ~n1265 ;
  assign n1267 = ( n324 & ~n482 ) | ( n324 & n1165 ) | ( ~n482 & n1165 ) ;
  assign n1268 = ( x68 & ~x246 ) | ( x68 & n722 ) | ( ~x246 & n722 ) ;
  assign n1269 = ( ~n318 & n320 ) | ( ~n318 & n1268 ) | ( n320 & n1268 ) ;
  assign n1270 = ( n1059 & ~n1267 ) | ( n1059 & n1269 ) | ( ~n1267 & n1269 ) ;
  assign n1271 = x124 & ~n581 ;
  assign n1272 = n814 & n1271 ;
  assign n1273 = n1272 ^ n482 ^ x117 ;
  assign n1274 = n1273 ^ n613 ^ 1'b0 ;
  assign n1276 = x224 ^ x176 ^ x18 ;
  assign n1275 = x153 & n808 ;
  assign n1277 = n1276 ^ n1275 ^ 1'b0 ;
  assign n1278 = ( n444 & n530 ) | ( n444 & ~n1277 ) | ( n530 & ~n1277 ) ;
  assign n1279 = ( x146 & ~n1075 ) | ( x146 & n1278 ) | ( ~n1075 & n1278 ) ;
  assign n1284 = n361 ^ n331 ^ x19 ;
  assign n1280 = n528 ^ x16 ^ 1'b0 ;
  assign n1281 = n831 & n1202 ;
  assign n1282 = x140 & ~n1281 ;
  assign n1283 = n1280 & n1282 ;
  assign n1285 = n1284 ^ n1283 ^ n830 ;
  assign n1286 = n1285 ^ n1194 ^ 1'b0 ;
  assign n1287 = ~n642 & n1286 ;
  assign n1288 = n540 ^ n441 ^ 1'b0 ;
  assign n1289 = n665 & n1288 ;
  assign n1290 = n1289 ^ n761 ^ n404 ;
  assign n1291 = n634 | n1290 ;
  assign n1292 = x152 | n1291 ;
  assign n1293 = n903 ^ n495 ^ 1'b0 ;
  assign n1294 = n750 | n1293 ;
  assign n1295 = n528 & ~n1294 ;
  assign n1296 = ~n293 & n1295 ;
  assign n1297 = n461 | n702 ;
  assign n1298 = x26 & n764 ;
  assign n1299 = n1298 ^ n1244 ^ 1'b0 ;
  assign n1300 = x72 & n1299 ;
  assign n1301 = ( x207 & n614 ) | ( x207 & ~n903 ) | ( n614 & ~n903 ) ;
  assign n1302 = ~n632 & n1301 ;
  assign n1303 = ~n1300 & n1302 ;
  assign n1305 = x214 & ~n434 ;
  assign n1306 = n1305 ^ n1027 ^ 1'b0 ;
  assign n1307 = ~n584 & n1306 ;
  assign n1304 = ( ~x123 & x130 ) | ( ~x123 & n416 ) | ( x130 & n416 ) ;
  assign n1308 = n1307 ^ n1304 ^ 1'b0 ;
  assign n1309 = x139 & n679 ;
  assign n1310 = n914 | n1309 ;
  assign n1311 = n1310 ^ n554 ^ 1'b0 ;
  assign n1312 = ( x168 & ~n595 ) | ( x168 & n662 ) | ( ~n595 & n662 ) ;
  assign n1313 = n1312 ^ n796 ^ 1'b0 ;
  assign n1314 = n835 | n1313 ;
  assign n1315 = ( x10 & x54 ) | ( x10 & n770 ) | ( x54 & n770 ) ;
  assign n1316 = x196 & n1315 ;
  assign n1317 = n1316 ^ n1266 ^ 1'b0 ;
  assign n1321 = n692 ^ x197 ^ x26 ;
  assign n1318 = n515 ^ n504 ^ x27 ;
  assign n1319 = n1318 ^ n585 ^ 1'b0 ;
  assign n1320 = n898 & ~n1319 ;
  assign n1322 = n1321 ^ n1320 ^ 1'b0 ;
  assign n1323 = x17 & n1322 ;
  assign n1324 = n446 ^ x204 ^ 1'b0 ;
  assign n1325 = n1072 & n1121 ;
  assign n1326 = ~n570 & n1220 ;
  assign n1327 = ~n394 & n1326 ;
  assign n1328 = n1327 ^ n618 ^ n556 ;
  assign n1329 = x163 ^ x2 ^ 1'b0 ;
  assign n1330 = x192 & n1329 ;
  assign n1331 = n1330 ^ n1268 ^ n1267 ;
  assign n1332 = x84 & n414 ;
  assign n1333 = n1332 ^ n963 ^ 1'b0 ;
  assign n1334 = n680 ^ x90 ^ 1'b0 ;
  assign n1335 = n552 & ~n1334 ;
  assign n1336 = n1335 ^ n688 ^ 1'b0 ;
  assign n1337 = ~n1333 & n1336 ;
  assign n1338 = n373 & n389 ;
  assign n1339 = x84 & x156 ;
  assign n1340 = ~n1338 & n1339 ;
  assign n1341 = n365 & ~n1340 ;
  assign n1342 = n1337 & n1341 ;
  assign n1343 = x212 & n711 ;
  assign n1344 = n1343 ^ x88 ^ 1'b0 ;
  assign n1345 = n1304 & ~n1344 ;
  assign n1346 = n614 & n1345 ;
  assign n1347 = n995 ^ n757 ^ 1'b0 ;
  assign n1348 = n1347 ^ n908 ^ x129 ;
  assign n1349 = ( x152 & ~x180 ) | ( x152 & n731 ) | ( ~x180 & n731 ) ;
  assign n1350 = n879 ^ x254 ^ x34 ;
  assign n1351 = n1350 ^ n733 ^ 1'b0 ;
  assign n1352 = x56 ^ x5 ^ 1'b0 ;
  assign n1353 = ( n315 & ~n1003 ) | ( n315 & n1352 ) | ( ~n1003 & n1352 ) ;
  assign n1354 = n1353 ^ n890 ^ 1'b0 ;
  assign n1355 = n963 ^ n393 ^ 1'b0 ;
  assign n1356 = n1330 ^ n508 ^ x12 ;
  assign n1359 = ( x94 & n1057 ) | ( x94 & n1260 ) | ( n1057 & n1260 ) ;
  assign n1357 = n566 ^ n461 ^ x248 ;
  assign n1358 = n1357 ^ x251 ^ x206 ;
  assign n1360 = n1359 ^ n1358 ^ 1'b0 ;
  assign n1361 = n1360 ^ n1030 ^ x121 ;
  assign n1362 = ~n1356 & n1361 ;
  assign n1363 = n1359 ^ n613 ^ 1'b0 ;
  assign n1364 = n551 ^ x2 ^ 1'b0 ;
  assign n1365 = ~n1363 & n1364 ;
  assign n1366 = ( ~x154 & x162 ) | ( ~x154 & x186 ) | ( x162 & x186 ) ;
  assign n1367 = ( x114 & n320 ) | ( x114 & ~n1366 ) | ( n320 & ~n1366 ) ;
  assign n1368 = n1040 ^ n335 ^ 1'b0 ;
  assign n1369 = n1226 | n1368 ;
  assign n1370 = ( n686 & n1367 ) | ( n686 & ~n1369 ) | ( n1367 & ~n1369 ) ;
  assign n1371 = n758 ^ n281 ^ 1'b0 ;
  assign n1372 = x219 & n1371 ;
  assign n1373 = x69 & x131 ;
  assign n1374 = n1373 ^ n765 ^ 1'b0 ;
  assign n1375 = x79 & n1116 ;
  assign n1376 = n1375 ^ n464 ^ 1'b0 ;
  assign n1377 = ~n1374 & n1376 ;
  assign n1378 = n579 & n1377 ;
  assign n1379 = x49 & ~n1378 ;
  assign n1380 = n826 | n868 ;
  assign n1381 = n1380 ^ x247 ^ 1'b0 ;
  assign n1382 = n1105 & n1381 ;
  assign n1383 = n1382 ^ x60 ^ 1'b0 ;
  assign n1384 = ( n382 & n397 ) | ( n382 & n1278 ) | ( n397 & n1278 ) ;
  assign n1385 = x20 | n771 ;
  assign n1386 = n1324 ^ n480 ^ 1'b0 ;
  assign n1387 = n1385 & n1386 ;
  assign n1388 = n1281 ^ n903 ^ 1'b0 ;
  assign n1389 = ~n284 & n400 ;
  assign n1390 = ~x17 & n1389 ;
  assign n1391 = n591 | n1390 ;
  assign n1392 = x114 & n1391 ;
  assign n1393 = x218 ^ x127 ^ x71 ;
  assign n1394 = n279 | n812 ;
  assign n1395 = x18 | n1394 ;
  assign n1396 = n1393 | n1395 ;
  assign n1397 = n642 ^ n548 ^ 1'b0 ;
  assign n1398 = n944 & ~n1397 ;
  assign n1399 = n996 ^ n294 ^ 1'b0 ;
  assign n1400 = n1398 & ~n1399 ;
  assign n1401 = n1400 ^ n326 ^ x115 ;
  assign n1402 = n459 & n790 ;
  assign n1403 = n419 & n1402 ;
  assign n1404 = x231 & ~n929 ;
  assign n1405 = n1403 & n1404 ;
  assign n1406 = ( x221 & ~x226 ) | ( x221 & n880 ) | ( ~x226 & n880 ) ;
  assign n1407 = x186 & ~n1406 ;
  assign n1408 = n1405 & n1407 ;
  assign n1409 = n329 & ~n1146 ;
  assign n1410 = n1409 ^ n1297 ^ 1'b0 ;
  assign n1411 = ( ~n305 & n410 ) | ( ~n305 & n1104 ) | ( n410 & n1104 ) ;
  assign n1412 = n1411 ^ n504 ^ x39 ;
  assign n1413 = n493 | n849 ;
  assign n1414 = n1413 ^ n1239 ^ 1'b0 ;
  assign n1415 = ~n751 & n1414 ;
  assign n1416 = n939 & n1415 ;
  assign n1417 = ~n1201 & n1416 ;
  assign n1418 = n1035 ^ n631 ^ n362 ;
  assign n1419 = n1189 ^ n943 ^ 1'b0 ;
  assign n1420 = n1418 | n1419 ;
  assign n1421 = ( ~n330 & n373 ) | ( ~n330 & n577 ) | ( n373 & n577 ) ;
  assign n1422 = ( ~n999 & n1374 ) | ( ~n999 & n1421 ) | ( n1374 & n1421 ) ;
  assign n1423 = ( ~n873 & n1420 ) | ( ~n873 & n1422 ) | ( n1420 & n1422 ) ;
  assign n1427 = n757 ^ n388 ^ 1'b0 ;
  assign n1424 = ~n259 & n1084 ;
  assign n1425 = n1424 ^ n367 ^ 1'b0 ;
  assign n1426 = n1387 & ~n1425 ;
  assign n1428 = n1427 ^ n1426 ^ 1'b0 ;
  assign n1429 = n1074 & ~n1428 ;
  assign n1438 = ( x95 & n340 ) | ( x95 & n825 ) | ( n340 & n825 ) ;
  assign n1439 = n829 & ~n969 ;
  assign n1440 = n553 & n1439 ;
  assign n1441 = n1438 | n1440 ;
  assign n1442 = n301 & ~n1441 ;
  assign n1430 = ( ~x69 & x110 ) | ( ~x69 & x116 ) | ( x110 & x116 ) ;
  assign n1431 = ~x60 & x136 ;
  assign n1432 = x69 & ~n1431 ;
  assign n1433 = ~n466 & n1432 ;
  assign n1434 = n1433 ^ n493 ^ 1'b0 ;
  assign n1435 = ( x62 & n449 ) | ( x62 & ~n1434 ) | ( n449 & ~n1434 ) ;
  assign n1436 = ( ~n614 & n1430 ) | ( ~n614 & n1435 ) | ( n1430 & n1435 ) ;
  assign n1437 = n1436 ^ x179 ^ x132 ;
  assign n1443 = n1442 ^ n1437 ^ 1'b0 ;
  assign n1444 = n1318 ^ n1155 ^ n331 ;
  assign n1445 = x131 ^ x81 ^ 1'b0 ;
  assign n1449 = ( x90 & ~n633 ) | ( x90 & n711 ) | ( ~n633 & n711 ) ;
  assign n1446 = n774 ^ n550 ^ n317 ;
  assign n1447 = x79 & ~n1446 ;
  assign n1448 = ~n410 & n1447 ;
  assign n1450 = n1449 ^ n1448 ^ 1'b0 ;
  assign n1451 = ( ~n1078 & n1445 ) | ( ~n1078 & n1450 ) | ( n1445 & n1450 ) ;
  assign n1453 = n429 | n639 ;
  assign n1454 = x110 | n1453 ;
  assign n1455 = n820 ^ x20 ^ 1'b0 ;
  assign n1456 = n1454 & ~n1455 ;
  assign n1457 = n1456 ^ x136 ^ 1'b0 ;
  assign n1452 = n1244 ^ n352 ^ n290 ;
  assign n1458 = n1457 ^ n1452 ^ 1'b0 ;
  assign n1459 = n428 ^ n360 ^ 1'b0 ;
  assign n1460 = n1357 | n1459 ;
  assign n1461 = ( n542 & n1117 ) | ( n542 & n1134 ) | ( n1117 & n1134 ) ;
  assign n1462 = n1461 ^ n776 ^ n379 ;
  assign n1463 = n500 & n1462 ;
  assign n1464 = n1460 & n1463 ;
  assign n1465 = n590 ^ x91 ^ x5 ;
  assign n1466 = n1011 & n1465 ;
  assign n1467 = n1464 & n1466 ;
  assign n1468 = n1420 ^ n1357 ^ n633 ;
  assign n1469 = x175 ^ x156 ^ x124 ;
  assign n1470 = ~n1406 & n1469 ;
  assign n1474 = n562 ^ x17 ^ 1'b0 ;
  assign n1471 = n633 & ~n996 ;
  assign n1472 = n1471 ^ n367 ^ 1'b0 ;
  assign n1473 = n1472 ^ n1241 ^ n317 ;
  assign n1475 = n1474 ^ n1473 ^ n381 ;
  assign n1476 = ~x64 & x156 ;
  assign n1477 = n1476 ^ n832 ^ n773 ;
  assign n1478 = ( x4 & x244 ) | ( x4 & ~n294 ) | ( x244 & ~n294 ) ;
  assign n1479 = n403 & ~n687 ;
  assign n1480 = n1479 ^ x18 ^ 1'b0 ;
  assign n1481 = n1480 ^ n340 ^ 1'b0 ;
  assign n1482 = n1298 & n1481 ;
  assign n1483 = ( n1011 & ~n1478 ) | ( n1011 & n1482 ) | ( ~n1478 & n1482 ) ;
  assign n1484 = ( x194 & x212 ) | ( x194 & ~n987 ) | ( x212 & ~n987 ) ;
  assign n1485 = n734 ^ x239 ^ 1'b0 ;
  assign n1486 = n1485 ^ n468 ^ 1'b0 ;
  assign n1487 = x238 & ~n1486 ;
  assign n1488 = ( ~n870 & n1485 ) | ( ~n870 & n1487 ) | ( n1485 & n1487 ) ;
  assign n1489 = ( x230 & n631 ) | ( x230 & ~n1488 ) | ( n631 & ~n1488 ) ;
  assign n1490 = x247 & n408 ;
  assign n1491 = n1490 ^ x212 ^ 1'b0 ;
  assign n1492 = x213 ^ x167 ^ 1'b0 ;
  assign n1493 = n704 & n1492 ;
  assign n1494 = ( x42 & n1491 ) | ( x42 & ~n1493 ) | ( n1491 & ~n1493 ) ;
  assign n1495 = x89 & n285 ;
  assign n1496 = n1494 & n1495 ;
  assign n1497 = n812 ^ n713 ^ n372 ;
  assign n1498 = n790 & n1497 ;
  assign n1499 = n1173 & n1498 ;
  assign n1500 = ~n299 & n417 ;
  assign n1501 = ~x122 & n1500 ;
  assign n1502 = ( ~x23 & x125 ) | ( ~x23 & n1377 ) | ( x125 & n1377 ) ;
  assign n1503 = ( ~n362 & n1501 ) | ( ~n362 & n1502 ) | ( n1501 & n1502 ) ;
  assign n1504 = n553 ^ x214 ^ x22 ;
  assign n1505 = ~n1503 & n1504 ;
  assign n1506 = n771 ^ x247 ^ x87 ;
  assign n1511 = n939 ^ n426 ^ x57 ;
  assign n1507 = x241 & ~n1491 ;
  assign n1508 = n1507 ^ n841 ^ 1'b0 ;
  assign n1509 = n871 ^ n271 ^ 1'b0 ;
  assign n1510 = n1508 | n1509 ;
  assign n1512 = n1511 ^ n1510 ^ 1'b0 ;
  assign n1513 = ( n1469 & ~n1506 ) | ( n1469 & n1512 ) | ( ~n1506 & n1512 ) ;
  assign n1515 = x117 & x154 ;
  assign n1516 = n1515 ^ x99 ^ 1'b0 ;
  assign n1517 = ( ~n625 & n869 ) | ( ~n625 & n1516 ) | ( n869 & n1516 ) ;
  assign n1514 = x197 & ~n1022 ;
  assign n1518 = n1517 ^ n1514 ^ 1'b0 ;
  assign n1519 = x98 & x159 ;
  assign n1520 = n1519 ^ x4 ^ 1'b0 ;
  assign n1521 = ( x158 & ~n357 ) | ( x158 & n1520 ) | ( ~n357 & n1520 ) ;
  assign n1522 = n1521 ^ n1278 ^ 1'b0 ;
  assign n1523 = n1522 ^ n321 ^ 1'b0 ;
  assign n1524 = n506 & n1523 ;
  assign n1526 = ( x167 & ~n733 ) | ( x167 & n1113 ) | ( ~n733 & n1113 ) ;
  assign n1525 = n573 ^ n268 ^ x156 ;
  assign n1527 = n1526 ^ n1525 ^ 1'b0 ;
  assign n1528 = n1527 ^ n1268 ^ 1'b0 ;
  assign n1529 = n1003 & n1528 ;
  assign n1530 = n268 ^ x66 ^ 1'b0 ;
  assign n1531 = n590 | n1530 ;
  assign n1532 = n1531 ^ n1048 ^ n311 ;
  assign n1533 = ( n497 & n1443 ) | ( n497 & n1532 ) | ( n1443 & n1532 ) ;
  assign n1534 = n490 & n1264 ;
  assign n1535 = ~n397 & n1534 ;
  assign n1536 = x73 & x239 ;
  assign n1537 = n1536 ^ x1 ^ 1'b0 ;
  assign n1538 = ( ~x120 & n842 ) | ( ~x120 & n1537 ) | ( n842 & n1537 ) ;
  assign n1539 = n1538 ^ n490 ^ n320 ;
  assign n1540 = ~n271 & n1539 ;
  assign n1541 = n1535 & n1540 ;
  assign n1542 = ( ~x248 & n547 ) | ( ~x248 & n1044 ) | ( n547 & n1044 ) ;
  assign n1543 = n1542 ^ x130 ^ x51 ;
  assign n1544 = x96 & x250 ;
  assign n1545 = n1544 ^ n537 ^ 1'b0 ;
  assign n1546 = x76 & n1545 ;
  assign n1547 = n324 & n1546 ;
  assign n1548 = n1547 ^ x150 ^ x79 ;
  assign n1549 = n277 & n1548 ;
  assign n1550 = ~n1543 & n1549 ;
  assign n1551 = n1550 ^ n1184 ^ n1010 ;
  assign n1552 = n1418 ^ n859 ^ 1'b0 ;
  assign n1553 = n512 ^ x171 ^ 1'b0 ;
  assign n1554 = n1093 & ~n1553 ;
  assign n1555 = ( ~x204 & n1477 ) | ( ~x204 & n1554 ) | ( n1477 & n1554 ) ;
  assign n1556 = n1485 ^ n1247 ^ x73 ;
  assign n1557 = ( ~n647 & n802 ) | ( ~n647 & n1556 ) | ( n802 & n1556 ) ;
  assign n1558 = n1474 ^ n1417 ^ 1'b0 ;
  assign n1559 = n1543 ^ n1010 ^ n771 ;
  assign n1564 = n399 | n627 ;
  assign n1560 = ( x196 & n934 ) | ( x196 & n1004 ) | ( n934 & n1004 ) ;
  assign n1561 = n294 & ~n841 ;
  assign n1562 = n1560 & n1561 ;
  assign n1563 = n360 | n1562 ;
  assign n1565 = n1564 ^ n1563 ^ 1'b0 ;
  assign n1566 = x78 & ~n1565 ;
  assign n1567 = ~n1559 & n1566 ;
  assign n1568 = n793 & n1398 ;
  assign n1570 = n879 ^ n430 ^ 1'b0 ;
  assign n1569 = x202 & ~n335 ;
  assign n1571 = n1570 ^ n1569 ^ 1'b0 ;
  assign n1572 = n1571 ^ x126 ^ 1'b0 ;
  assign n1573 = n595 & n1572 ;
  assign n1574 = n301 & ~n780 ;
  assign n1575 = n791 ^ x223 ^ 1'b0 ;
  assign n1576 = n1454 & ~n1575 ;
  assign n1577 = n1452 & n1576 ;
  assign n1578 = ~n1574 & n1577 ;
  assign n1579 = n757 & ~n782 ;
  assign n1580 = ( x8 & n941 ) | ( x8 & n1579 ) | ( n941 & n1579 ) ;
  assign n1581 = n1194 ^ n1020 ^ 1'b0 ;
  assign n1582 = ~x33 & n1034 ;
  assign n1583 = n1582 ^ x46 ^ 1'b0 ;
  assign n1584 = x163 ^ x121 ^ 1'b0 ;
  assign n1585 = n1347 & ~n1584 ;
  assign n1590 = n731 ^ n486 ^ x1 ;
  assign n1586 = ( n963 & ~n1098 ) | ( n963 & n1178 ) | ( ~n1098 & n1178 ) ;
  assign n1587 = n1586 ^ n1245 ^ 1'b0 ;
  assign n1588 = n455 & ~n1587 ;
  assign n1589 = x188 & ~n1588 ;
  assign n1591 = n1590 ^ n1589 ^ n331 ;
  assign n1592 = n1374 ^ n1074 ^ x49 ;
  assign n1593 = n1592 ^ n1305 ^ n709 ;
  assign n1594 = ( ~n279 & n362 ) | ( ~n279 & n1040 ) | ( n362 & n1040 ) ;
  assign n1595 = ( x243 & n1593 ) | ( x243 & n1594 ) | ( n1593 & n1594 ) ;
  assign n1596 = x35 & ~n1595 ;
  assign n1597 = ~n1591 & n1596 ;
  assign n1598 = ( n621 & n1585 ) | ( n621 & ~n1597 ) | ( n1585 & ~n1597 ) ;
  assign n1600 = ( x92 & n1054 ) | ( x92 & n1118 ) | ( n1054 & n1118 ) ;
  assign n1599 = n1409 ^ x241 ^ x211 ;
  assign n1601 = n1600 ^ n1599 ^ 1'b0 ;
  assign n1603 = ( ~x207 & n381 ) | ( ~x207 & n397 ) | ( n381 & n397 ) ;
  assign n1604 = n1603 ^ n1064 ^ 1'b0 ;
  assign n1602 = n695 & ~n962 ;
  assign n1605 = n1604 ^ n1602 ^ 1'b0 ;
  assign n1606 = x175 & n1605 ;
  assign n1607 = n1606 ^ n343 ^ 1'b0 ;
  assign n1608 = n1607 ^ n926 ^ n293 ;
  assign n1609 = n534 & n1445 ;
  assign n1610 = n1609 ^ n406 ^ 1'b0 ;
  assign n1611 = ( ~x225 & n305 ) | ( ~x225 & n414 ) | ( n305 & n414 ) ;
  assign n1614 = x252 | n464 ;
  assign n1615 = ~n447 & n618 ;
  assign n1616 = n1614 & n1615 ;
  assign n1612 = x236 ^ x226 ^ x76 ;
  assign n1613 = n261 | n1612 ;
  assign n1617 = n1616 ^ n1613 ^ 1'b0 ;
  assign n1618 = n1611 | n1617 ;
  assign n1619 = n1610 & ~n1618 ;
  assign n1620 = x155 & ~n424 ;
  assign n1621 = n1620 ^ n1374 ^ 1'b0 ;
  assign n1622 = x31 & ~n1621 ;
  assign n1623 = ~n515 & n1443 ;
  assign n1624 = ( x188 & ~n598 ) | ( x188 & n1582 ) | ( ~n598 & n1582 ) ;
  assign n1625 = n307 ^ x116 ^ 1'b0 ;
  assign n1626 = n290 & n1625 ;
  assign n1627 = n1626 ^ n455 ^ 1'b0 ;
  assign n1628 = n1064 | n1357 ;
  assign n1629 = n1083 | n1628 ;
  assign n1630 = ( x199 & n457 ) | ( x199 & ~n1629 ) | ( n457 & ~n1629 ) ;
  assign n1631 = ( x143 & ~n1627 ) | ( x143 & n1630 ) | ( ~n1627 & n1630 ) ;
  assign n1632 = ( n751 & n1465 ) | ( n751 & n1631 ) | ( n1465 & n1631 ) ;
  assign n1633 = ~n1624 & n1632 ;
  assign n1634 = ~x183 & n1633 ;
  assign n1635 = n1594 ^ n1538 ^ n1350 ;
  assign n1636 = n881 & n1635 ;
  assign n1637 = n657 & n1636 ;
  assign n1638 = n616 & n1081 ;
  assign n1639 = n1638 ^ n629 ^ 1'b0 ;
  assign n1640 = ( x241 & ~n404 ) | ( x241 & n898 ) | ( ~n404 & n898 ) ;
  assign n1641 = n1051 & ~n1640 ;
  assign n1642 = n1011 & ~n1163 ;
  assign n1643 = n1642 ^ x3 ^ 1'b0 ;
  assign n1644 = n966 ^ n331 ^ 1'b0 ;
  assign n1645 = ( ~n720 & n767 ) | ( ~n720 & n1644 ) | ( n767 & n1644 ) ;
  assign n1646 = ( x232 & n724 ) | ( x232 & n968 ) | ( n724 & n968 ) ;
  assign n1651 = x126 & x240 ;
  assign n1652 = ~x80 & n1651 ;
  assign n1647 = n417 ^ x241 ^ x96 ;
  assign n1648 = n1647 ^ n889 ^ 1'b0 ;
  assign n1649 = n1460 | n1648 ;
  assign n1650 = n1649 ^ n1324 ^ x7 ;
  assign n1653 = n1652 ^ n1650 ^ 1'b0 ;
  assign n1654 = n1646 & ~n1653 ;
  assign n1658 = x106 & ~x135 ;
  assign n1655 = ( n410 & ~n1043 ) | ( n410 & n1629 ) | ( ~n1043 & n1629 ) ;
  assign n1656 = ~n1537 & n1655 ;
  assign n1657 = n1044 & ~n1656 ;
  assign n1659 = n1658 ^ n1657 ^ 1'b0 ;
  assign n1660 = n1144 & ~n1315 ;
  assign n1661 = n499 ^ x47 ^ 1'b0 ;
  assign n1662 = n1656 | n1661 ;
  assign n1663 = n1056 & n1451 ;
  assign n1664 = n1068 & n1625 ;
  assign n1665 = n1664 ^ n1102 ^ x83 ;
  assign n1666 = ( n676 & n689 ) | ( n676 & ~n1004 ) | ( n689 & ~n1004 ) ;
  assign n1667 = ( n639 & ~n1665 ) | ( n639 & n1666 ) | ( ~n1665 & n1666 ) ;
  assign n1668 = n892 & ~n1209 ;
  assign n1669 = n671 & n1668 ;
  assign n1670 = x128 & n293 ;
  assign n1671 = n1670 ^ x199 ^ 1'b0 ;
  assign n1672 = n1671 ^ n540 ^ 1'b0 ;
  assign n1673 = ( n1650 & n1669 ) | ( n1650 & ~n1672 ) | ( n1669 & ~n1672 ) ;
  assign n1674 = ( ~n1117 & n1132 ) | ( ~n1117 & n1301 ) | ( n1132 & n1301 ) ;
  assign n1675 = ~n474 & n977 ;
  assign n1676 = n1239 ^ n767 ^ 1'b0 ;
  assign n1677 = n987 ^ n593 ^ 1'b0 ;
  assign n1678 = ~n763 & n1677 ;
  assign n1679 = n1120 ^ x22 ^ 1'b0 ;
  assign n1680 = n1007 & ~n1679 ;
  assign n1683 = n1136 ^ n958 ^ n880 ;
  assign n1681 = n561 ^ n355 ^ x10 ;
  assign n1682 = ( ~n933 & n1570 ) | ( ~n933 & n1681 ) | ( n1570 & n1681 ) ;
  assign n1684 = n1683 ^ n1682 ^ 1'b0 ;
  assign n1685 = ( n548 & ~n1680 ) | ( n548 & n1684 ) | ( ~n1680 & n1684 ) ;
  assign n1686 = n1120 ^ n1063 ^ 1'b0 ;
  assign n1687 = n836 | n1686 ;
  assign n1688 = n299 & n955 ;
  assign n1691 = ( x24 & n408 ) | ( x24 & n461 ) | ( n408 & n461 ) ;
  assign n1689 = n329 & n1452 ;
  assign n1690 = n1689 ^ n598 ^ 1'b0 ;
  assign n1692 = n1691 ^ n1690 ^ n396 ;
  assign n1693 = n544 & n1692 ;
  assign n1694 = n1693 ^ n370 ^ 1'b0 ;
  assign n1695 = n1694 ^ n1448 ^ x187 ;
  assign n1696 = n1104 ^ x55 ^ 1'b0 ;
  assign n1697 = n1220 & ~n1696 ;
  assign n1698 = n1697 ^ n1589 ^ 1'b0 ;
  assign n1701 = ( x72 & ~x125 ) | ( x72 & n430 ) | ( ~x125 & n430 ) ;
  assign n1700 = ( ~n341 & n1430 ) | ( ~n341 & n1691 ) | ( n1430 & n1691 ) ;
  assign n1702 = n1701 ^ n1700 ^ 1'b0 ;
  assign n1703 = x220 & ~n1702 ;
  assign n1699 = n648 & ~n1235 ;
  assign n1704 = n1703 ^ n1699 ^ 1'b0 ;
  assign n1705 = n757 ^ n642 ^ n294 ;
  assign n1706 = ~x86 & n1705 ;
  assign n1707 = n1706 ^ x88 ^ 1'b0 ;
  assign n1708 = n335 & n1707 ;
  assign n1709 = ~x12 & n1708 ;
  assign n1710 = ( n434 & n1003 ) | ( n434 & ~n1077 ) | ( n1003 & ~n1077 ) ;
  assign n1712 = n473 ^ n443 ^ 1'b0 ;
  assign n1711 = x76 & ~n1098 ;
  assign n1713 = n1712 ^ n1711 ^ 1'b0 ;
  assign n1714 = n1713 ^ n1690 ^ n890 ;
  assign n1715 = ~n1206 & n1629 ;
  assign n1716 = ~n1714 & n1715 ;
  assign n1717 = n1716 ^ n952 ^ n825 ;
  assign n1718 = n1345 | n1717 ;
  assign n1719 = n1718 ^ n971 ^ 1'b0 ;
  assign n1720 = n1719 ^ n279 ^ x132 ;
  assign n1721 = n355 & n410 ;
  assign n1729 = n1555 ^ n1289 ^ 1'b0 ;
  assign n1723 = n1372 ^ n511 ^ n496 ;
  assign n1724 = n910 ^ n497 ^ 1'b0 ;
  assign n1725 = n550 | n1724 ;
  assign n1726 = n1723 | n1725 ;
  assign n1722 = n616 & ~n1130 ;
  assign n1727 = n1726 ^ n1722 ^ 1'b0 ;
  assign n1728 = x31 & n1727 ;
  assign n1730 = n1729 ^ n1728 ^ 1'b0 ;
  assign n1732 = ( x8 & ~x196 ) | ( x8 & n640 ) | ( ~x196 & n640 ) ;
  assign n1733 = ( x179 & n1531 ) | ( x179 & ~n1732 ) | ( n1531 & ~n1732 ) ;
  assign n1731 = x186 & ~n1717 ;
  assign n1734 = n1733 ^ n1731 ^ 1'b0 ;
  assign n1735 = ( ~n838 & n1676 ) | ( ~n838 & n1734 ) | ( n1676 & n1734 ) ;
  assign n1736 = n1330 ^ n325 ^ x18 ;
  assign n1737 = ~x182 & n1736 ;
  assign n1738 = ( n1469 & n1595 ) | ( n1469 & ~n1737 ) | ( n1595 & ~n1737 ) ;
  assign n1739 = n1205 ^ n1011 ^ 1'b0 ;
  assign n1740 = n1189 ^ x121 ^ x30 ;
  assign n1741 = n1740 ^ n1062 ^ 1'b0 ;
  assign n1742 = ( n1247 & n1488 ) | ( n1247 & ~n1741 ) | ( n1488 & ~n1741 ) ;
  assign n1743 = n929 ^ n656 ^ 1'b0 ;
  assign n1744 = n1743 ^ n654 ^ n417 ;
  assign n1745 = x232 ^ x209 ^ x198 ;
  assign n1746 = n1745 ^ n1690 ^ x177 ;
  assign n1747 = ~n662 & n1046 ;
  assign n1748 = n1747 ^ n338 ^ 1'b0 ;
  assign n1749 = n1748 ^ n1264 ^ x236 ;
  assign n1750 = ( n410 & n1746 ) | ( n410 & ~n1749 ) | ( n1746 & ~n1749 ) ;
  assign n1751 = n1750 ^ n1588 ^ 1'b0 ;
  assign n1752 = n1290 | n1751 ;
  assign n1753 = n352 & n1201 ;
  assign n1756 = n838 & ~n1268 ;
  assign n1757 = n1756 ^ n524 ^ 1'b0 ;
  assign n1754 = n1168 ^ x32 ^ 1'b0 ;
  assign n1755 = n313 & ~n1754 ;
  assign n1758 = n1757 ^ n1755 ^ 1'b0 ;
  assign n1759 = n634 ^ x80 ^ 1'b0 ;
  assign n1760 = n1759 ^ n290 ^ 1'b0 ;
  assign n1761 = n414 & ~n1760 ;
  assign n1767 = n431 & ~n990 ;
  assign n1768 = n1767 ^ n903 ^ 1'b0 ;
  assign n1762 = x148 & n1083 ;
  assign n1763 = ~n533 & n1762 ;
  assign n1764 = n1763 ^ n315 ^ 1'b0 ;
  assign n1765 = n730 | n1764 ;
  assign n1766 = n988 & ~n1765 ;
  assign n1769 = n1768 ^ n1766 ^ x192 ;
  assign n1770 = n1761 & ~n1769 ;
  assign n1771 = n1770 ^ x51 ^ 1'b0 ;
  assign n1772 = x76 & n1427 ;
  assign n1773 = ~n295 & n1772 ;
  assign n1774 = n1773 ^ n1148 ^ 1'b0 ;
  assign n1775 = n1289 & n1774 ;
  assign n1776 = ( n457 & n1158 ) | ( n457 & ~n1570 ) | ( n1158 & ~n1570 ) ;
  assign n1777 = n918 ^ n376 ^ 1'b0 ;
  assign n1778 = x59 & ~n1777 ;
  assign n1779 = x116 & ~n352 ;
  assign n1780 = ( n340 & n1745 ) | ( n340 & n1779 ) | ( n1745 & n1779 ) ;
  assign n1781 = n1780 ^ n1706 ^ 1'b0 ;
  assign n1782 = n1778 & ~n1781 ;
  assign n1783 = ( ~x145 & x158 ) | ( ~x145 & n313 ) | ( x158 & n313 ) ;
  assign n1784 = n1783 ^ n728 ^ 1'b0 ;
  assign n1785 = ( x208 & n554 ) | ( x208 & ~n1784 ) | ( n554 & ~n1784 ) ;
  assign n1786 = ( n623 & n1782 ) | ( n623 & n1785 ) | ( n1782 & n1785 ) ;
  assign n1787 = ~x232 & n269 ;
  assign n1788 = x30 & x237 ;
  assign n1789 = n1787 & n1788 ;
  assign n1790 = n724 ^ x124 ^ x32 ;
  assign n1792 = ~n647 & n699 ;
  assign n1793 = n1792 ^ x54 ^ 1'b0 ;
  assign n1791 = n469 ^ x159 ^ 1'b0 ;
  assign n1794 = n1793 ^ n1791 ^ 1'b0 ;
  assign n1795 = ~n1375 & n1794 ;
  assign n1796 = ( ~x35 & n1790 ) | ( ~x35 & n1795 ) | ( n1790 & n1795 ) ;
  assign n1798 = x111 & ~n516 ;
  assign n1799 = n1798 ^ n1014 ^ x123 ;
  assign n1797 = x252 & ~n798 ;
  assign n1800 = n1799 ^ n1797 ^ 1'b0 ;
  assign n1801 = x156 | n402 ;
  assign n1802 = n1801 ^ n1638 ^ n1630 ;
  assign n1806 = x153 & ~n357 ;
  assign n1805 = x37 & n261 ;
  assign n1803 = x39 & ~n724 ;
  assign n1804 = n1803 ^ x8 ^ 1'b0 ;
  assign n1807 = n1806 ^ n1805 ^ n1804 ;
  assign n1809 = x27 & n1173 ;
  assign n1810 = n1809 ^ n1447 ^ 1'b0 ;
  assign n1811 = ( x211 & ~n937 ) | ( x211 & n1810 ) | ( ~n937 & n1810 ) ;
  assign n1812 = n1406 | n1811 ;
  assign n1808 = n873 & n1775 ;
  assign n1813 = n1812 ^ n1808 ^ 1'b0 ;
  assign n1826 = n343 ^ x180 ^ x80 ;
  assign n1827 = n1826 ^ n1658 ^ n560 ;
  assign n1816 = x65 & n341 ;
  assign n1817 = ~n1535 & n1816 ;
  assign n1818 = n1817 ^ n597 ^ 1'b0 ;
  assign n1814 = n1270 ^ n280 ^ 1'b0 ;
  assign n1815 = x33 & ~n1814 ;
  assign n1819 = n1818 ^ n1815 ^ 1'b0 ;
  assign n1820 = x125 & n397 ;
  assign n1821 = n1820 ^ x56 ^ 1'b0 ;
  assign n1822 = n1821 ^ n1365 ^ n761 ;
  assign n1823 = n656 & ~n1353 ;
  assign n1824 = ( n1819 & ~n1822 ) | ( n1819 & n1823 ) | ( ~n1822 & n1823 ) ;
  assign n1825 = n829 & n1824 ;
  assign n1828 = n1827 ^ n1825 ^ 1'b0 ;
  assign n1836 = n1225 ^ n910 ^ x136 ;
  assign n1837 = n1836 ^ n1643 ^ n1102 ;
  assign n1829 = n877 ^ n397 ^ 1'b0 ;
  assign n1830 = x245 & ~n1829 ;
  assign n1831 = ~n982 & n1830 ;
  assign n1832 = n1831 ^ n1114 ^ 1'b0 ;
  assign n1833 = x188 & ~n1832 ;
  assign n1834 = n602 & n1833 ;
  assign n1835 = n1239 | n1834 ;
  assign n1838 = n1837 ^ n1835 ^ 1'b0 ;
  assign n1839 = ( x12 & x140 ) | ( x12 & ~x228 ) | ( x140 & ~x228 ) ;
  assign n1840 = n1839 ^ n1346 ^ n829 ;
  assign n1841 = n1478 ^ n791 ^ x173 ;
  assign n1842 = n1365 & n1841 ;
  assign n1843 = n1842 ^ n594 ^ 1'b0 ;
  assign n1844 = ( ~x72 & x91 ) | ( ~x72 & n1205 ) | ( x91 & n1205 ) ;
  assign n1845 = x25 & n1844 ;
  assign n1847 = x135 & n759 ;
  assign n1848 = n1847 ^ x158 ^ 1'b0 ;
  assign n1849 = n1848 ^ n490 ^ 1'b0 ;
  assign n1850 = n462 | n1849 ;
  assign n1851 = n1850 ^ n734 ^ x157 ;
  assign n1846 = n1644 ^ n796 ^ n780 ;
  assign n1852 = n1851 ^ n1846 ^ n1608 ;
  assign n1853 = n1277 ^ n669 ^ n590 ;
  assign n1854 = ( ~x148 & n450 ) | ( ~x148 & n711 ) | ( n450 & n711 ) ;
  assign n1855 = n1854 ^ x253 ^ x118 ;
  assign n1856 = n1352 & ~n1855 ;
  assign n1857 = n1853 & n1856 ;
  assign n1860 = ~n261 & n1188 ;
  assign n1861 = n1860 ^ x127 ^ 1'b0 ;
  assign n1862 = n1289 & ~n1861 ;
  assign n1863 = n1862 ^ n595 ^ 1'b0 ;
  assign n1858 = x218 ^ x39 ^ 1'b0 ;
  assign n1859 = n1858 ^ n1356 ^ n637 ;
  assign n1864 = n1863 ^ n1859 ^ n1791 ;
  assign n1865 = n290 & ~n1864 ;
  assign n1866 = n1865 ^ n1104 ^ 1'b0 ;
  assign n1872 = n264 & n568 ;
  assign n1873 = ~n885 & n1872 ;
  assign n1870 = n518 & ~n960 ;
  assign n1867 = n910 ^ n524 ^ 1'b0 ;
  assign n1868 = ( x30 & n847 ) | ( x30 & n1470 ) | ( n847 & n1470 ) ;
  assign n1869 = n1867 & ~n1868 ;
  assign n1871 = n1870 ^ n1869 ^ 1'b0 ;
  assign n1874 = n1873 ^ n1871 ^ n367 ;
  assign n1876 = n1640 ^ n1075 ^ 1'b0 ;
  assign n1875 = ( x67 & n287 ) | ( x67 & ~n895 ) | ( n287 & ~n895 ) ;
  assign n1877 = n1876 ^ n1875 ^ x244 ;
  assign n1878 = ~n504 & n1864 ;
  assign n1879 = n1878 ^ n1198 ^ n763 ;
  assign n1880 = n1879 ^ n470 ^ 1'b0 ;
  assign n1881 = ~n1517 & n1880 ;
  assign n1882 = n1360 & n1733 ;
  assign n1883 = ( n879 & ~n1854 ) | ( n879 & n1882 ) | ( ~n1854 & n1882 ) ;
  assign n1884 = n1535 ^ n1135 ^ n773 ;
  assign n1885 = n350 | n1571 ;
  assign n1886 = n1766 & n1885 ;
  assign n1888 = ( x21 & ~x219 ) | ( x21 & n330 ) | ( ~x219 & n330 ) ;
  assign n1887 = n499 & n1672 ;
  assign n1889 = n1888 ^ n1887 ^ n1744 ;
  assign n1890 = n831 & ~n1087 ;
  assign n1891 = ~n682 & n1890 ;
  assign n1892 = x146 & n816 ;
  assign n1893 = ~x211 & n1892 ;
  assign n1894 = ( x228 & ~n919 ) | ( x228 & n1893 ) | ( ~n919 & n1893 ) ;
  assign n1895 = n766 & n1007 ;
  assign n1896 = ~x28 & n1895 ;
  assign n1897 = ( n318 & n444 ) | ( n318 & n1703 ) | ( n444 & n1703 ) ;
  assign n1898 = ( n1324 & n1896 ) | ( n1324 & ~n1897 ) | ( n1896 & ~n1897 ) ;
  assign n1899 = n1091 ^ x228 ^ 1'b0 ;
  assign n1900 = ~n812 & n1899 ;
  assign n1901 = n1900 ^ n1247 ^ x159 ;
  assign n1903 = n1442 ^ x207 ^ 1'b0 ;
  assign n1902 = ( n428 & n744 ) | ( n428 & n840 ) | ( n744 & n840 ) ;
  assign n1904 = n1903 ^ n1902 ^ x74 ;
  assign n1905 = x92 & ~n814 ;
  assign n1906 = n1905 ^ n982 ^ 1'b0 ;
  assign n1907 = ( n257 & n1732 ) | ( n257 & ~n1906 ) | ( n1732 & ~n1906 ) ;
  assign n1908 = n1907 ^ n1701 ^ 1'b0 ;
  assign n1909 = n1908 ^ n1581 ^ x45 ;
  assign n1912 = ~n616 & n910 ;
  assign n1913 = n1912 ^ n732 ^ x17 ;
  assign n1914 = n368 & n1682 ;
  assign n1915 = n1914 ^ n564 ^ 1'b0 ;
  assign n1916 = ( n737 & n1913 ) | ( n737 & n1915 ) | ( n1913 & n1915 ) ;
  assign n1911 = n577 | n1795 ;
  assign n1910 = n1422 ^ x56 ^ 1'b0 ;
  assign n1917 = n1916 ^ n1911 ^ n1910 ;
  assign n1918 = n671 | n1206 ;
  assign n1919 = n1314 & ~n1918 ;
  assign n1920 = ( n444 & n598 ) | ( n444 & n1919 ) | ( n598 & n1919 ) ;
  assign n1921 = n1920 ^ n1589 ^ 1'b0 ;
  assign n1931 = n1001 ^ n787 ^ 1'b0 ;
  assign n1932 = n1173 & n1931 ;
  assign n1927 = n941 ^ x198 ^ 1'b0 ;
  assign n1928 = ~n971 & n1927 ;
  assign n1929 = n508 & n1928 ;
  assign n1930 = ~x191 & n1929 ;
  assign n1923 = x232 & ~n511 ;
  assign n1922 = n419 & ~n657 ;
  assign n1924 = n1923 ^ n1922 ^ n1231 ;
  assign n1925 = ~n1851 & n1924 ;
  assign n1926 = n384 & n1925 ;
  assign n1933 = n1932 ^ n1930 ^ n1926 ;
  assign n1934 = n916 & n1078 ;
  assign n1935 = n1934 ^ n1075 ^ 1'b0 ;
  assign n1936 = ( n291 & ~n438 ) | ( n291 & n996 ) | ( ~n438 & n996 ) ;
  assign n1937 = x100 & ~n1488 ;
  assign n1938 = n1937 ^ n340 ^ 1'b0 ;
  assign n1939 = ~x55 & n1254 ;
  assign n1940 = n1939 ^ x229 ^ 1'b0 ;
  assign n1941 = n1938 & n1940 ;
  assign n1942 = ~n1527 & n1941 ;
  assign n1943 = n1936 & n1942 ;
  assign n1944 = x87 & ~n1091 ;
  assign n1945 = ( x212 & n1604 ) | ( x212 & ~n1944 ) | ( n1604 & ~n1944 ) ;
  assign n1946 = n881 & ~n1945 ;
  assign n1947 = n259 & n1946 ;
  assign n1948 = ~n1460 & n1784 ;
  assign n1949 = n506 ^ x225 ^ 1'b0 ;
  assign n1950 = n1948 & ~n1949 ;
  assign n1951 = n336 & n1102 ;
  assign n1952 = n1951 ^ n358 ^ 1'b0 ;
  assign n1953 = ( x94 & ~n645 ) | ( x94 & n1590 ) | ( ~n645 & n1590 ) ;
  assign n1954 = n1161 ^ n410 ^ 1'b0 ;
  assign n1955 = n1954 ^ n1853 ^ 1'b0 ;
  assign n1956 = n1953 & ~n1955 ;
  assign n1957 = ~n585 & n1346 ;
  assign n1958 = ( n1380 & ~n1605 ) | ( n1380 & n1957 ) | ( ~n1605 & n1957 ) ;
  assign n1959 = n1482 ^ n799 ^ x97 ;
  assign n1960 = x209 ^ x27 ^ 1'b0 ;
  assign n1961 = x240 & n1960 ;
  assign n1962 = x202 & n1961 ;
  assign n1963 = ~x56 & n1962 ;
  assign n1964 = ( x137 & n1125 ) | ( x137 & ~n1963 ) | ( n1125 & ~n1963 ) ;
  assign n1969 = n576 ^ n408 ^ 1'b0 ;
  assign n1970 = ~n857 & n1969 ;
  assign n1971 = ~x41 & n1970 ;
  assign n1965 = x211 & n1042 ;
  assign n1966 = n1240 & n1965 ;
  assign n1967 = n1966 ^ n1047 ^ 1'b0 ;
  assign n1968 = n739 & n1967 ;
  assign n1972 = n1971 ^ n1968 ^ 1'b0 ;
  assign n1973 = n378 & ~n1972 ;
  assign n1974 = n334 & n459 ;
  assign n1976 = x237 & n327 ;
  assign n1977 = n1976 ^ n417 ^ 1'b0 ;
  assign n1975 = n475 & n1436 ;
  assign n1978 = n1977 ^ n1975 ^ n1075 ;
  assign n1979 = n944 ^ n738 ^ n284 ;
  assign n1980 = n709 & n1979 ;
  assign n1981 = n1978 & n1980 ;
  assign n1984 = n673 ^ n654 ^ x164 ;
  assign n1982 = n1047 ^ x212 ^ 1'b0 ;
  assign n1983 = n680 | n1982 ;
  assign n1985 = n1984 ^ n1983 ^ n926 ;
  assign n1986 = n495 ^ n361 ^ x151 ;
  assign n1987 = ~n1356 & n1986 ;
  assign n1988 = ~n1782 & n1987 ;
  assign n1993 = ~n445 & n656 ;
  assign n1994 = n1993 ^ n443 ^ 1'b0 ;
  assign n1992 = n692 | n1331 ;
  assign n1995 = n1994 ^ n1992 ^ 1'b0 ;
  assign n1989 = n595 ^ n382 ^ n325 ;
  assign n1990 = n1003 & n1989 ;
  assign n1991 = ~n1761 & n1990 ;
  assign n1996 = n1995 ^ n1991 ^ 1'b0 ;
  assign n1997 = n614 & ~n1996 ;
  assign n1998 = ( n1985 & n1988 ) | ( n1985 & ~n1997 ) | ( n1988 & ~n1997 ) ;
  assign n1999 = n408 & ~n1742 ;
  assign n2000 = n1363 & n1999 ;
  assign n2001 = ( n488 & ~n576 ) | ( n488 & n617 ) | ( ~n576 & n617 ) ;
  assign n2002 = n493 ^ x180 ^ 1'b0 ;
  assign n2003 = n2001 | n2002 ;
  assign n2004 = n2003 ^ n1799 ^ n428 ;
  assign n2005 = n853 & n2004 ;
  assign n2006 = n2005 ^ n548 ^ 1'b0 ;
  assign n2007 = n1452 ^ n530 ^ x185 ;
  assign n2008 = x0 & x218 ;
  assign n2009 = ( n845 & n929 ) | ( n845 & n2008 ) | ( n929 & n2008 ) ;
  assign n2010 = n1533 ^ n1001 ^ 1'b0 ;
  assign n2011 = n533 & ~n2010 ;
  assign n2012 = x220 ^ x38 ^ 1'b0 ;
  assign n2013 = x228 & n2012 ;
  assign n2014 = ( n370 & n874 ) | ( n370 & n2013 ) | ( n874 & n2013 ) ;
  assign n2015 = n2011 & ~n2014 ;
  assign n2016 = n284 & n2015 ;
  assign n2017 = n500 ^ n259 ^ x216 ;
  assign n2018 = x152 & n1746 ;
  assign n2019 = ~n1228 & n2018 ;
  assign n2020 = n2017 | n2019 ;
  assign n2023 = n1430 ^ x76 ^ 1'b0 ;
  assign n2024 = ~n587 & n2023 ;
  assign n2025 = x71 & n2024 ;
  assign n2026 = ~n724 & n2025 ;
  assign n2027 = n2026 ^ n984 ^ 1'b0 ;
  assign n2021 = n1093 ^ n269 ^ x204 ;
  assign n2022 = ( n1120 & n1391 ) | ( n1120 & n2021 ) | ( n1391 & n2021 ) ;
  assign n2028 = n2027 ^ n2022 ^ n724 ;
  assign n2029 = ( x33 & n429 ) | ( x33 & n537 ) | ( n429 & n537 ) ;
  assign n2030 = n2029 ^ n1924 ^ n1264 ;
  assign n2031 = n1030 ^ n320 ^ x72 ;
  assign n2032 = n2031 ^ x54 ^ 1'b0 ;
  assign n2033 = n1006 ^ n737 ^ n470 ;
  assign n2034 = n2033 ^ n1761 ^ 1'b0 ;
  assign n2035 = n436 & n2034 ;
  assign n2036 = x211 & n2035 ;
  assign n2037 = n2032 & n2036 ;
  assign n2038 = n2037 ^ x109 ^ 1'b0 ;
  assign n2039 = ~x117 & n551 ;
  assign n2040 = ~n284 & n518 ;
  assign n2041 = ( n1362 & ~n2039 ) | ( n1362 & n2040 ) | ( ~n2039 & n2040 ) ;
  assign n2042 = n306 & n711 ;
  assign n2043 = n2042 ^ n1759 ^ n1236 ;
  assign n2044 = n879 & ~n2043 ;
  assign n2045 = n2044 ^ n1725 ^ 1'b0 ;
  assign n2046 = n1757 ^ n750 ^ 1'b0 ;
  assign n2047 = n2045 & n2046 ;
  assign n2048 = x245 & n998 ;
  assign n2049 = n1535 ^ n1044 ^ 1'b0 ;
  assign n2050 = n987 | n1397 ;
  assign n2051 = ( ~n379 & n1411 ) | ( ~n379 & n2050 ) | ( n1411 & n2050 ) ;
  assign n2052 = n2051 ^ n626 ^ x167 ;
  assign n2054 = n1483 & n1493 ;
  assign n2055 = n2026 & n2054 ;
  assign n2053 = ~n331 & n1043 ;
  assign n2056 = n2055 ^ n2053 ^ 1'b0 ;
  assign n2057 = n1299 ^ n1189 ^ n299 ;
  assign n2058 = n1787 ^ n1411 ^ 1'b0 ;
  assign n2059 = x141 & n2058 ;
  assign n2060 = n1502 & n2059 ;
  assign n2061 = n2057 & n2060 ;
  assign n2062 = ( ~n814 & n1095 ) | ( ~n814 & n2061 ) | ( n1095 & n2061 ) ;
  assign n2063 = n1418 | n1845 ;
  assign n2065 = x63 & ~n790 ;
  assign n2066 = ~n464 & n2065 ;
  assign n2064 = ( x11 & ~n1229 ) | ( x11 & n2013 ) | ( ~n1229 & n2013 ) ;
  assign n2067 = n2066 ^ n2064 ^ 1'b0 ;
  assign n2068 = n1813 & n2067 ;
  assign n2069 = n1277 & n2068 ;
  assign n2070 = n2069 ^ n1375 ^ 1'b0 ;
  assign n2076 = ( ~x29 & n574 ) | ( ~x29 & n738 ) | ( n574 & n738 ) ;
  assign n2077 = n1284 ^ n877 ^ n551 ;
  assign n2078 = n2077 ^ n1810 ^ 1'b0 ;
  assign n2079 = n1423 | n2078 ;
  assign n2080 = n2076 | n2079 ;
  assign n2081 = n2080 ^ n1743 ^ 1'b0 ;
  assign n2071 = n802 ^ n396 ^ x176 ;
  assign n2072 = n1080 ^ n907 ^ 1'b0 ;
  assign n2073 = ~n692 & n2072 ;
  assign n2074 = ( n424 & n2071 ) | ( n424 & n2073 ) | ( n2071 & n2073 ) ;
  assign n2075 = n2074 ^ n1641 ^ 1'b0 ;
  assign n2082 = n2081 ^ n2075 ^ 1'b0 ;
  assign n2084 = n633 ^ x227 ^ 1'b0 ;
  assign n2083 = ( ~x114 & n426 ) | ( ~x114 & n1179 ) | ( n426 & n1179 ) ;
  assign n2085 = n2084 ^ n2083 ^ n1011 ;
  assign n2089 = n294 & ~n337 ;
  assign n2090 = x194 & ~n1104 ;
  assign n2091 = n2089 & n2090 ;
  assign n2092 = n2091 ^ x178 ^ 1'b0 ;
  assign n2087 = x138 & n663 ;
  assign n2088 = n604 & n2087 ;
  assign n2093 = n2092 ^ n2088 ^ 1'b0 ;
  assign n2086 = x74 & n584 ;
  assign n2094 = n2093 ^ n2086 ^ n2050 ;
  assign n2095 = n1807 ^ n341 ^ 1'b0 ;
  assign n2096 = ~n1752 & n2095 ;
  assign n2099 = x44 & n1300 ;
  assign n2100 = ~x128 & n2099 ;
  assign n2097 = ( x184 & n1059 ) | ( x184 & ~n1805 ) | ( n1059 & ~n1805 ) ;
  assign n2098 = x137 & n2097 ;
  assign n2101 = n2100 ^ n2098 ^ 1'b0 ;
  assign n2102 = n2101 ^ x166 ^ 1'b0 ;
  assign n2103 = n1146 & n2102 ;
  assign n2104 = n2103 ^ n1823 ^ 1'b0 ;
  assign n2105 = x196 | n1850 ;
  assign n2106 = n1644 ^ n572 ^ n416 ;
  assign n2107 = n573 ^ x64 ^ x7 ;
  assign n2108 = ~x207 & n2107 ;
  assign n2109 = ~n679 & n2108 ;
  assign n2110 = ( ~n867 & n918 ) | ( ~n867 & n2109 ) | ( n918 & n2109 ) ;
  assign n2111 = x149 & n492 ;
  assign n2112 = ~x119 & n2111 ;
  assign n2113 = n748 ^ n634 ^ 1'b0 ;
  assign n2114 = n1040 ^ n706 ^ 1'b0 ;
  assign n2115 = ~n2113 & n2114 ;
  assign n2116 = n1130 & n2115 ;
  assign n2117 = ( n1273 & n2112 ) | ( n1273 & n2116 ) | ( n2112 & n2116 ) ;
  assign n2118 = n516 & n595 ;
  assign n2119 = n2118 ^ n1805 ^ 1'b0 ;
  assign n2120 = n543 ^ x199 ^ 1'b0 ;
  assign n2121 = n2119 & ~n2120 ;
  assign n2122 = n905 | n1484 ;
  assign n2123 = ~n2121 & n2122 ;
  assign n2124 = ( n1851 & ~n2117 ) | ( n1851 & n2123 ) | ( ~n2117 & n2123 ) ;
  assign n2125 = n2089 ^ n449 ^ x3 ;
  assign n2126 = n438 & ~n2125 ;
  assign n2127 = ( n963 & n1743 ) | ( n963 & n2126 ) | ( n1743 & n2126 ) ;
  assign n2128 = ( ~n340 & n1315 ) | ( ~n340 & n1864 ) | ( n1315 & n1864 ) ;
  assign n2129 = n2032 & n2128 ;
  assign n2130 = n2127 & n2129 ;
  assign n2131 = n1375 ^ n284 ^ 1'b0 ;
  assign n2138 = x91 & ~n692 ;
  assign n2132 = n1134 ^ n287 ^ 1'b0 ;
  assign n2133 = n1858 ^ x116 ^ 1'b0 ;
  assign n2134 = n2132 | n2133 ;
  assign n2135 = n2134 ^ n1272 ^ x113 ;
  assign n2136 = n313 | n2135 ;
  assign n2137 = ~n1570 & n2136 ;
  assign n2139 = n2138 ^ n2137 ^ 1'b0 ;
  assign n2140 = n2139 ^ n1083 ^ 1'b0 ;
  assign n2141 = n1219 & ~n1630 ;
  assign n2142 = ~n1799 & n2141 ;
  assign n2154 = n1161 ^ n699 ^ n272 ;
  assign n2152 = ( n341 & n1012 ) | ( n341 & ~n1087 ) | ( n1012 & ~n1087 ) ;
  assign n2147 = ~n372 & n417 ;
  assign n2148 = n2147 ^ n780 ^ 1'b0 ;
  assign n2149 = n2148 ^ n679 ^ n572 ;
  assign n2150 = n1975 & n2149 ;
  assign n2151 = ~n541 & n2150 ;
  assign n2153 = n2152 ^ n2151 ^ 1'b0 ;
  assign n2143 = n1493 ^ n1059 ^ n841 ;
  assign n2144 = n1548 ^ n443 ^ 1'b0 ;
  assign n2145 = n372 | n2144 ;
  assign n2146 = ( ~x42 & n2143 ) | ( ~x42 & n2145 ) | ( n2143 & n2145 ) ;
  assign n2155 = n2154 ^ n2153 ^ n2146 ;
  assign n2156 = ~n332 & n434 ;
  assign n2157 = n2156 ^ n1617 ^ n1532 ;
  assign n2158 = n2157 ^ x20 ^ 1'b0 ;
  assign n2160 = n1487 & ~n2125 ;
  assign n2159 = ~n287 & n880 ;
  assign n2161 = n2160 ^ n2159 ^ 1'b0 ;
  assign n2162 = n1713 ^ n434 ^ 1'b0 ;
  assign n2163 = n2161 | n2162 ;
  assign n2164 = ( n408 & ~n1612 ) | ( n408 & n1832 ) | ( ~n1612 & n1832 ) ;
  assign n2165 = n1401 ^ x7 ^ 1'b0 ;
  assign n2166 = n373 & ~n2165 ;
  assign n2167 = n1685 & n2166 ;
  assign n2168 = ( n987 & n1161 ) | ( n987 & n1625 ) | ( n1161 & n1625 ) ;
  assign n2169 = n325 & n367 ;
  assign n2170 = ( ~n1541 & n2168 ) | ( ~n1541 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2172 = n668 & n809 ;
  assign n2173 = n2172 ^ n1258 ^ 1'b0 ;
  assign n2171 = n1641 ^ n999 ^ x233 ;
  assign n2174 = n2173 ^ n2171 ^ 1'b0 ;
  assign n2175 = n1714 & n2174 ;
  assign n2176 = x79 & n1101 ;
  assign n2177 = n2050 & n2176 ;
  assign n2178 = n695 ^ n626 ^ x229 ;
  assign n2183 = n1111 ^ n871 ^ 1'b0 ;
  assign n2184 = n1680 & ~n2183 ;
  assign n2179 = n468 & n1006 ;
  assign n2180 = ( x212 & n370 ) | ( x212 & ~n2179 ) | ( n370 & ~n2179 ) ;
  assign n2181 = n1598 ^ n992 ^ 1'b0 ;
  assign n2182 = n2180 & n2181 ;
  assign n2185 = n2184 ^ n2182 ^ 1'b0 ;
  assign n2186 = n707 & n2185 ;
  assign n2187 = n1832 ^ n306 ^ 1'b0 ;
  assign n2188 = n2187 ^ n504 ^ 1'b0 ;
  assign n2189 = n1052 & n2188 ;
  assign n2190 = n2189 ^ n1562 ^ 1'b0 ;
  assign n2191 = n2186 & ~n2190 ;
  assign n2192 = ( n971 & n2178 ) | ( n971 & n2191 ) | ( n2178 & n2191 ) ;
  assign n2193 = n741 & ~n1535 ;
  assign n2194 = n2193 ^ n1857 ^ 1'b0 ;
  assign n2195 = ( n333 & n785 ) | ( n333 & ~n1474 ) | ( n785 & ~n1474 ) ;
  assign n2196 = x151 & n2195 ;
  assign n2197 = ~n2175 & n2196 ;
  assign n2198 = n673 ^ x250 ^ 1'b0 ;
  assign n2199 = n1358 & ~n2198 ;
  assign n2200 = n2199 ^ x81 ^ 1'b0 ;
  assign n2201 = n1629 & n2200 ;
  assign n2202 = n1051 & ~n1280 ;
  assign n2203 = n2202 ^ x69 ^ 1'b0 ;
  assign n2204 = n2203 ^ n2073 ^ 1'b0 ;
  assign n2205 = n1029 | n2204 ;
  assign n2206 = n1852 ^ n1729 ^ n944 ;
  assign n2207 = x9 & ~n2206 ;
  assign n2208 = ~n682 & n2207 ;
  assign n2209 = n1057 ^ n309 ^ 1'b0 ;
  assign n2210 = ~n1074 & n2209 ;
  assign n2211 = n2210 ^ n941 ^ n706 ;
  assign n2212 = x45 & n580 ;
  assign n2213 = n2212 ^ n1134 ^ 1'b0 ;
  assign n2214 = n514 | n2213 ;
  assign n2215 = n2214 ^ n787 ^ 1'b0 ;
  assign n2216 = ( n558 & ~n1117 ) | ( n558 & n1455 ) | ( ~n1117 & n1455 ) ;
  assign n2217 = n2216 ^ n1133 ^ 1'b0 ;
  assign n2218 = n2217 ^ n1567 ^ n1211 ;
  assign n2220 = n647 ^ x109 ^ 1'b0 ;
  assign n2219 = x197 & ~n963 ;
  assign n2221 = n2220 ^ n2219 ^ 1'b0 ;
  assign n2222 = x203 & n1333 ;
  assign n2223 = ~n1244 & n2222 ;
  assign n2224 = n1622 & ~n2223 ;
  assign n2225 = n2221 & n2224 ;
  assign n2226 = ( n2215 & n2218 ) | ( n2215 & n2225 ) | ( n2218 & n2225 ) ;
  assign n2227 = n330 ^ x209 ^ x126 ;
  assign n2228 = n2227 ^ n378 ^ 1'b0 ;
  assign n2229 = n428 & n2228 ;
  assign n2230 = ~n322 & n2229 ;
  assign n2231 = ( n1372 & n1593 ) | ( n1372 & n2230 ) | ( n1593 & n2230 ) ;
  assign n2232 = n1721 & n2231 ;
  assign n2233 = n1305 ^ n372 ^ x159 ;
  assign n2246 = n1563 ^ n1263 ^ n457 ;
  assign n2234 = ( x230 & n355 ) | ( x230 & n770 ) | ( n355 & n770 ) ;
  assign n2235 = n872 & ~n1460 ;
  assign n2236 = ~x217 & n2235 ;
  assign n2237 = n2236 ^ n1187 ^ 1'b0 ;
  assign n2238 = ~n2027 & n2237 ;
  assign n2239 = n871 & n2238 ;
  assign n2240 = n2239 ^ x211 ^ 1'b0 ;
  assign n2241 = n769 ^ n533 ^ n338 ;
  assign n2242 = n1526 ^ x52 ^ 1'b0 ;
  assign n2243 = ~n2241 & n2242 ;
  assign n2244 = ( ~n2234 & n2240 ) | ( ~n2234 & n2243 ) | ( n2240 & n2243 ) ;
  assign n2245 = n1067 & ~n2244 ;
  assign n2247 = n2246 ^ n2245 ^ 1'b0 ;
  assign n2248 = ~n289 & n368 ;
  assign n2249 = n2248 ^ n1887 ^ 1'b0 ;
  assign n2250 = n598 & ~n870 ;
  assign n2251 = n2250 ^ n326 ^ 1'b0 ;
  assign n2252 = ( n405 & ~n618 ) | ( n405 & n877 ) | ( ~n618 & n877 ) ;
  assign n2253 = n2251 & ~n2252 ;
  assign n2254 = n1183 & n2253 ;
  assign n2255 = n322 | n1539 ;
  assign n2257 = n703 & n1545 ;
  assign n2258 = n2257 ^ n695 ^ 1'b0 ;
  assign n2256 = n1791 ^ n910 ^ x205 ;
  assign n2259 = n2258 ^ n2256 ^ 1'b0 ;
  assign n2260 = x17 & ~n2259 ;
  assign n2261 = n2255 | n2260 ;
  assign n2262 = n1592 ^ n642 ^ n259 ;
  assign n2263 = n2014 | n2262 ;
  assign n2264 = n1075 & ~n1130 ;
  assign n2265 = n447 & n2264 ;
  assign n2266 = n2265 ^ x209 ^ 1'b0 ;
  assign n2267 = n581 | n2266 ;
  assign n2268 = n1791 ^ n1726 ^ n1353 ;
  assign n2269 = x111 & ~n901 ;
  assign n2270 = n2269 ^ n1128 ^ 1'b0 ;
  assign n2271 = n2270 ^ n1280 ^ 1'b0 ;
  assign n2272 = n1712 & ~n2271 ;
  assign n2273 = n2272 ^ n552 ^ x9 ;
  assign n2274 = ( n493 & ~n969 ) | ( n493 & n2250 ) | ( ~n969 & n2250 ) ;
  assign n2275 = n2274 ^ n1903 ^ 1'b0 ;
  assign n2276 = x70 & n2275 ;
  assign n2277 = ( n262 & n709 ) | ( n262 & ~n1004 ) | ( n709 & ~n1004 ) ;
  assign n2278 = x53 & x185 ;
  assign n2279 = n2278 ^ x131 ^ 1'b0 ;
  assign n2280 = n2279 ^ x106 ^ 1'b0 ;
  assign n2281 = ( ~n706 & n2277 ) | ( ~n706 & n2280 ) | ( n2277 & n2280 ) ;
  assign n2282 = n2022 ^ n1769 ^ n452 ;
  assign n2283 = ( n446 & n533 ) | ( n446 & n1894 ) | ( n533 & n1894 ) ;
  assign n2284 = n1122 ^ n1009 ^ 1'b0 ;
  assign n2285 = n1477 ^ n1040 ^ 1'b0 ;
  assign n2286 = n2284 & n2285 ;
  assign n2292 = x252 & ~n1787 ;
  assign n2293 = n2292 ^ n1057 ^ 1'b0 ;
  assign n2289 = n744 ^ x14 ^ 1'b0 ;
  assign n2290 = n2289 ^ n2227 ^ x116 ;
  assign n2287 = n1309 ^ n1130 ^ n868 ;
  assign n2288 = n1949 & n2287 ;
  assign n2291 = n2290 ^ n2288 ^ 1'b0 ;
  assign n2294 = n2293 ^ n2291 ^ 1'b0 ;
  assign n2295 = n2286 & ~n2294 ;
  assign n2296 = n1093 ^ n702 ^ 1'b0 ;
  assign n2297 = ( x40 & n1280 ) | ( x40 & ~n2296 ) | ( n1280 & ~n2296 ) ;
  assign n2298 = n578 ^ x25 ^ 1'b0 ;
  assign n2299 = ~n322 & n2298 ;
  assign n2300 = n2299 ^ x254 ^ 1'b0 ;
  assign n2301 = ~n1659 & n2300 ;
  assign n2302 = ~n2297 & n2301 ;
  assign n2303 = n346 & n2302 ;
  assign n2304 = ~n812 & n1564 ;
  assign n2305 = n430 & n2304 ;
  assign n2306 = n2305 ^ n1061 ^ 1'b0 ;
  assign n2307 = n2306 ^ x49 ^ 1'b0 ;
  assign n2308 = n1665 | n2307 ;
  assign n2309 = n1526 ^ n1315 ^ 1'b0 ;
  assign n2310 = ~n1261 & n2309 ;
  assign n2312 = n455 ^ n431 ^ 1'b0 ;
  assign n2313 = ~n843 & n2312 ;
  assign n2311 = n348 & ~n1029 ;
  assign n2314 = n2313 ^ n2311 ^ 1'b0 ;
  assign n2315 = ~x54 & x110 ;
  assign n2316 = n1801 & ~n2315 ;
  assign n2317 = n2314 & n2316 ;
  assign n2318 = n1120 | n1594 ;
  assign n2319 = n2318 ^ n410 ^ 1'b0 ;
  assign n2320 = n2319 ^ n1179 ^ 1'b0 ;
  assign n2321 = x196 & ~n2320 ;
  assign n2322 = ( n831 & n2317 ) | ( n831 & ~n2321 ) | ( n2317 & ~n2321 ) ;
  assign n2323 = x212 ^ x190 ^ 1'b0 ;
  assign n2324 = n745 & n2323 ;
  assign n2325 = n2324 ^ n1732 ^ x198 ;
  assign n2326 = n2325 ^ n684 ^ 1'b0 ;
  assign n2327 = x190 & n2326 ;
  assign n2328 = n2327 ^ x150 ^ 1'b0 ;
  assign n2329 = x132 | n445 ;
  assign n2330 = ( n2293 & ~n2328 ) | ( n2293 & n2329 ) | ( ~n2328 & n2329 ) ;
  assign n2331 = n1250 ^ n343 ^ 1'b0 ;
  assign n2332 = x242 & n2331 ;
  assign n2333 = ( x204 & n416 ) | ( x204 & ~n753 ) | ( n416 & ~n753 ) ;
  assign n2334 = x42 & ~n609 ;
  assign n2335 = n2334 ^ x200 ^ 1'b0 ;
  assign n2336 = n2335 ^ n941 ^ n306 ;
  assign n2337 = ( n960 & n2333 ) | ( n960 & n2336 ) | ( n2333 & n2336 ) ;
  assign n2338 = ( ~x186 & n2332 ) | ( ~x186 & n2337 ) | ( n2332 & n2337 ) ;
  assign n2339 = n1428 ^ n1117 ^ 1'b0 ;
  assign n2340 = n748 ^ n462 ^ x155 ;
  assign n2341 = x81 & n2340 ;
  assign n2342 = x123 & ~n542 ;
  assign n2343 = n2342 ^ n642 ^ 1'b0 ;
  assign n2344 = n1380 ^ n1367 ^ n1018 ;
  assign n2345 = n2344 ^ x196 ^ 1'b0 ;
  assign n2346 = n2343 & ~n2345 ;
  assign n2347 = ~n2341 & n2346 ;
  assign n2348 = n256 & n2261 ;
  assign n2349 = n2347 & n2348 ;
  assign n2354 = n1390 ^ n602 ^ n287 ;
  assign n2351 = n256 ^ x235 ^ x208 ;
  assign n2352 = n1367 ^ x8 ^ 1'b0 ;
  assign n2353 = ~n2351 & n2352 ;
  assign n2355 = n2354 ^ n2353 ^ n730 ;
  assign n2350 = n2333 & ~n2349 ;
  assign n2356 = n2355 ^ n2350 ^ 1'b0 ;
  assign n2357 = ( ~x58 & n977 ) | ( ~x58 & n1625 ) | ( n977 & n1625 ) ;
  assign n2358 = ~n305 & n1956 ;
  assign n2359 = n2357 & n2358 ;
  assign n2360 = x213 & n295 ;
  assign n2361 = n877 & n2360 ;
  assign n2362 = n2361 ^ n1289 ^ 1'b0 ;
  assign n2363 = n773 & n2362 ;
  assign n2364 = n2363 ^ n831 ^ 1'b0 ;
  assign n2365 = x219 & ~x246 ;
  assign n2367 = ( ~x20 & n280 ) | ( ~x20 & n281 ) | ( n280 & n281 ) ;
  assign n2368 = ( x22 & x168 ) | ( x22 & n2367 ) | ( x168 & n2367 ) ;
  assign n2369 = n2368 ^ n1411 ^ x212 ;
  assign n2366 = n1074 | n1844 ;
  assign n2370 = n2369 ^ n2366 ^ 1'b0 ;
  assign n2371 = n2365 & n2370 ;
  assign n2372 = n2371 ^ n678 ^ 1'b0 ;
  assign n2373 = x14 & ~n473 ;
  assign n2374 = n386 & n2373 ;
  assign n2375 = n2374 ^ n317 ^ 1'b0 ;
  assign n2376 = n1873 | n2375 ;
  assign n2377 = n2376 ^ n358 ^ 1'b0 ;
  assign n2378 = x248 & ~n1477 ;
  assign n2379 = n2377 & n2378 ;
  assign n2380 = ( x24 & n1864 ) | ( x24 & ~n2089 ) | ( n1864 & ~n2089 ) ;
  assign n2381 = n491 & ~n702 ;
  assign n2382 = n2381 ^ n868 ^ 1'b0 ;
  assign n2383 = ~n331 & n2382 ;
  assign n2384 = n2383 ^ n2333 ^ x153 ;
  assign n2385 = x69 & ~n625 ;
  assign n2386 = n2385 ^ n669 ^ 1'b0 ;
  assign n2387 = n313 & ~n726 ;
  assign n2388 = n1863 & n2387 ;
  assign n2389 = n2138 & ~n2186 ;
  assign n2390 = ( n849 & n1328 ) | ( n849 & ~n2019 ) | ( n1328 & ~n2019 ) ;
  assign n2398 = ( n644 & n671 ) | ( n644 & ~n683 ) | ( n671 & ~n683 ) ;
  assign n2399 = ( n1994 & ~n2220 ) | ( n1994 & n2398 ) | ( ~n2220 & n2398 ) ;
  assign n2392 = n486 ^ n430 ^ 1'b0 ;
  assign n2393 = n289 | n2392 ;
  assign n2394 = n2393 ^ n526 ^ n403 ;
  assign n2395 = ( n374 & ~n474 ) | ( n374 & n2394 ) | ( ~n474 & n2394 ) ;
  assign n2396 = x192 & ~n1148 ;
  assign n2397 = ~n2395 & n2396 ;
  assign n2391 = n2341 ^ n1317 ^ x139 ;
  assign n2400 = n2399 ^ n2397 ^ n2391 ;
  assign n2401 = n2230 & n2400 ;
  assign n2402 = n1474 & ~n1745 ;
  assign n2403 = n2402 ^ n1977 ^ 1'b0 ;
  assign n2404 = x128 & n400 ;
  assign n2405 = n2404 ^ n1391 ^ 1'b0 ;
  assign n2406 = n608 ^ n314 ^ x93 ;
  assign n2407 = ( n1846 & ~n2405 ) | ( n1846 & n2406 ) | ( ~n2405 & n2406 ) ;
  assign n2408 = n2407 ^ x37 ^ 1'b0 ;
  assign n2409 = ~n2403 & n2408 ;
  assign n2410 = x179 ^ x143 ^ x105 ;
  assign n2411 = ( x28 & n623 ) | ( x28 & n999 ) | ( n623 & n999 ) ;
  assign n2412 = ( ~n1081 & n1192 ) | ( ~n1081 & n2411 ) | ( n1192 & n2411 ) ;
  assign n2413 = ( n464 & ~n690 ) | ( n464 & n1150 ) | ( ~n690 & n1150 ) ;
  assign n2414 = ~n537 & n2413 ;
  assign n2415 = ( n2410 & n2412 ) | ( n2410 & n2414 ) | ( n2412 & n2414 ) ;
  assign n2416 = n282 & n2220 ;
  assign n2417 = ~n1181 & n2416 ;
  assign n2418 = n2149 ^ x145 ^ 1'b0 ;
  assign n2419 = ~n1590 & n2418 ;
  assign n2420 = x203 & ~n2167 ;
  assign n2421 = n2420 ^ n1725 ^ 1'b0 ;
  assign n2422 = ~x235 & n2013 ;
  assign n2423 = ( x124 & n497 ) | ( x124 & ~n2422 ) | ( n497 & ~n2422 ) ;
  assign n2424 = n2423 ^ x91 ^ 1'b0 ;
  assign n2425 = n1461 & n2424 ;
  assign n2426 = n1944 ^ n1390 ^ 1'b0 ;
  assign n2427 = n2425 & ~n2426 ;
  assign n2428 = n337 & n1963 ;
  assign n2429 = n2428 ^ n1478 ^ 1'b0 ;
  assign n2430 = n915 & ~n2429 ;
  assign n2439 = ~n261 & n605 ;
  assign n2440 = n2439 ^ n1493 ^ 1'b0 ;
  assign n2441 = ( ~x54 & n941 ) | ( ~x54 & n956 ) | ( n941 & n956 ) ;
  assign n2442 = n2121 ^ n633 ^ x171 ;
  assign n2443 = x224 | n2442 ;
  assign n2444 = ( n2440 & ~n2441 ) | ( n2440 & n2443 ) | ( ~n2441 & n2443 ) ;
  assign n2431 = x86 & n749 ;
  assign n2432 = n2431 ^ n584 ^ 1'b0 ;
  assign n2433 = x113 & ~n2432 ;
  assign n2434 = n2433 ^ n1491 ^ 1'b0 ;
  assign n2435 = ~n2089 & n2434 ;
  assign n2436 = n2435 ^ n1133 ^ 1'b0 ;
  assign n2437 = n421 & n633 ;
  assign n2438 = ( x176 & n2436 ) | ( x176 & ~n2437 ) | ( n2436 & ~n2437 ) ;
  assign n2445 = n2444 ^ n2438 ^ 1'b0 ;
  assign n2446 = n2096 ^ n637 ^ 1'b0 ;
  assign n2447 = n262 | n2446 ;
  assign n2448 = n871 ^ x130 ^ 1'b0 ;
  assign n2449 = n2132 ^ n625 ^ x218 ;
  assign n2450 = ( x180 & n521 ) | ( x180 & n2449 ) | ( n521 & n2449 ) ;
  assign n2451 = ( ~x238 & n715 ) | ( ~x238 & n1841 ) | ( n715 & n1841 ) ;
  assign n2452 = ~n1656 & n1783 ;
  assign n2453 = n2452 ^ x197 ^ 1'b0 ;
  assign n2454 = n2453 ^ n617 ^ 1'b0 ;
  assign n2455 = ~n2451 & n2454 ;
  assign n2456 = ( n1538 & n2450 ) | ( n1538 & n2455 ) | ( n2450 & n2455 ) ;
  assign n2458 = n1086 ^ n469 ^ 1'b0 ;
  assign n2457 = n1046 & ~n1703 ;
  assign n2459 = n2458 ^ n2457 ^ 1'b0 ;
  assign n2460 = x101 & ~n2459 ;
  assign n2461 = ( x201 & n483 ) | ( x201 & n726 ) | ( n483 & n726 ) ;
  assign n2462 = n1202 | n2432 ;
  assign n2463 = n2462 ^ n547 ^ 1'b0 ;
  assign n2464 = n2463 ^ n1855 ^ n358 ;
  assign n2465 = n2464 ^ n1061 ^ 1'b0 ;
  assign n2466 = n2113 ^ n1409 ^ 1'b0 ;
  assign n2467 = ( n1314 & ~n2465 ) | ( n1314 & n2466 ) | ( ~n2465 & n2466 ) ;
  assign n2468 = n2467 ^ n1320 ^ 1'b0 ;
  assign n2469 = ( n799 & ~n2461 ) | ( n799 & n2468 ) | ( ~n2461 & n2468 ) ;
  assign n2475 = x16 | n1070 ;
  assign n2470 = n493 ^ x24 ^ 1'b0 ;
  assign n2471 = n1924 ^ n1616 ^ 1'b0 ;
  assign n2472 = n373 & n2471 ;
  assign n2473 = ~n2470 & n2472 ;
  assign n2474 = n1647 & n2473 ;
  assign n2476 = n2475 ^ n2474 ^ 1'b0 ;
  assign n2477 = ( n572 & n587 ) | ( n572 & ~n1284 ) | ( n587 & ~n1284 ) ;
  assign n2478 = n2477 ^ n1101 ^ n889 ;
  assign n2479 = n2478 ^ n1594 ^ 1'b0 ;
  assign n2480 = x185 & ~n1652 ;
  assign n2481 = n2480 ^ n1579 ^ 1'b0 ;
  assign n2483 = x39 & x131 ;
  assign n2484 = ~x191 & n2483 ;
  assign n2482 = ( x54 & ~x164 ) | ( x54 & n1455 ) | ( ~x164 & n1455 ) ;
  assign n2485 = n2484 ^ n2482 ^ 1'b0 ;
  assign n2486 = n2485 ^ n1385 ^ 1'b0 ;
  assign n2487 = n2486 ^ n1597 ^ 1'b0 ;
  assign n2488 = n1780 | n2487 ;
  assign n2489 = n1049 | n1179 ;
  assign n2490 = n2489 ^ n663 ^ 1'b0 ;
  assign n2491 = x140 & n1906 ;
  assign n2492 = n2361 & n2491 ;
  assign n2493 = n2490 & ~n2492 ;
  assign n2494 = n2488 & n2493 ;
  assign n2495 = ( ~n556 & n1372 ) | ( ~n556 & n1844 ) | ( n1372 & n1844 ) ;
  assign n2496 = n2495 ^ n1017 ^ 1'b0 ;
  assign n2497 = n470 | n2496 ;
  assign n2498 = n1799 & n2497 ;
  assign n2499 = ( ~n386 & n1482 ) | ( ~n386 & n1978 ) | ( n1482 & n1978 ) ;
  assign n2500 = x172 & n2499 ;
  assign n2501 = n576 ^ n396 ^ 1'b0 ;
  assign n2502 = n2501 ^ n1543 ^ n593 ;
  assign n2503 = ( x87 & n441 ) | ( x87 & n488 ) | ( n441 & n488 ) ;
  assign n2504 = ( ~n1573 & n1583 ) | ( ~n1573 & n2503 ) | ( n1583 & n2503 ) ;
  assign n2505 = n2504 ^ n1729 ^ 1'b0 ;
  assign n2506 = ~n398 & n2505 ;
  assign n2507 = n980 ^ n731 ^ n474 ;
  assign n2508 = ~n408 & n2507 ;
  assign n2509 = n1132 & n1939 ;
  assign n2510 = n1260 ^ x247 ^ 1'b0 ;
  assign n2511 = n1201 ^ n1121 ^ 1'b0 ;
  assign n2512 = n2510 & ~n2511 ;
  assign n2513 = n1430 ^ n663 ^ x246 ;
  assign n2514 = n2513 ^ n1369 ^ n1083 ;
  assign n2515 = ~n1716 & n2514 ;
  assign n2516 = n1599 & n2008 ;
  assign n2517 = ~x208 & n2516 ;
  assign n2518 = n1017 | n1442 ;
  assign n2519 = n1745 ^ n732 ^ n609 ;
  assign n2520 = n1874 & n2519 ;
  assign n2526 = n756 & ~n1501 ;
  assign n2527 = n2526 ^ n793 ^ 1'b0 ;
  assign n2528 = ( ~n607 & n642 ) | ( ~n607 & n2527 ) | ( n642 & n2527 ) ;
  assign n2529 = ~n822 & n2528 ;
  assign n2523 = n299 ^ x114 ^ 1'b0 ;
  assign n2524 = x187 | n2523 ;
  assign n2521 = ~n362 & n918 ;
  assign n2522 = ~x14 & n2521 ;
  assign n2525 = n2524 ^ n2522 ^ 1'b0 ;
  assign n2530 = n2529 ^ n2525 ^ 1'b0 ;
  assign n2531 = ( x75 & n269 ) | ( x75 & n722 ) | ( n269 & n722 ) ;
  assign n2533 = ( x69 & n623 ) | ( x69 & ~n1102 ) | ( n623 & ~n1102 ) ;
  assign n2532 = x8 | n1624 ;
  assign n2534 = n2533 ^ n2532 ^ n779 ;
  assign n2535 = n2531 & ~n2534 ;
  assign n2536 = ~n1451 & n2535 ;
  assign n2553 = n720 & ~n1396 ;
  assign n2554 = x41 & ~n2553 ;
  assign n2537 = n2513 ^ n884 ^ 1'b0 ;
  assign n2538 = x122 & n2537 ;
  assign n2539 = ~n1725 & n2538 ;
  assign n2540 = ~n2289 & n2539 ;
  assign n2541 = n2540 ^ n2407 ^ x87 ;
  assign n2542 = ( n380 & n763 ) | ( n380 & n2541 ) | ( n763 & n2541 ) ;
  assign n2549 = ~x109 & n1434 ;
  assign n2550 = ( n595 & n905 ) | ( n595 & n2549 ) | ( n905 & n2549 ) ;
  assign n2547 = n325 ^ x97 ^ 1'b0 ;
  assign n2543 = x43 & ~n1977 ;
  assign n2544 = n2543 ^ n404 ^ 1'b0 ;
  assign n2545 = n572 & ~n1689 ;
  assign n2546 = ~n2544 & n2545 ;
  assign n2548 = n2547 ^ n2546 ^ 1'b0 ;
  assign n2551 = n2550 ^ n2548 ^ n354 ;
  assign n2552 = ~n2542 & n2551 ;
  assign n2555 = n2554 ^ n2552 ^ 1'b0 ;
  assign n2556 = n1661 & ~n2555 ;
  assign n2557 = ~n428 & n2556 ;
  assign n2560 = n843 ^ x200 ^ 1'b0 ;
  assign n2558 = n2234 ^ n1372 ^ n524 ;
  assign n2559 = n2558 ^ n391 ^ 1'b0 ;
  assign n2561 = n2560 ^ n2559 ^ n580 ;
  assign n2562 = n1415 ^ n1328 ^ 1'b0 ;
  assign n2563 = x211 & ~n564 ;
  assign n2564 = n2116 ^ n1450 ^ 1'b0 ;
  assign n2565 = ( n698 & n2563 ) | ( n698 & n2564 ) | ( n2563 & n2564 ) ;
  assign n2574 = n1358 ^ n1209 ^ x87 ;
  assign n2566 = ( n520 & n554 ) | ( n520 & n768 ) | ( n554 & n768 ) ;
  assign n2567 = ( x187 & ~x222 ) | ( x187 & n2566 ) | ( ~x222 & n2566 ) ;
  assign n2568 = n1048 | n2440 ;
  assign n2569 = n2568 ^ x235 ^ 1'b0 ;
  assign n2570 = ~n795 & n2569 ;
  assign n2571 = n2570 ^ n843 ^ 1'b0 ;
  assign n2572 = ~n2567 & n2571 ;
  assign n2573 = n2572 ^ x86 ^ 1'b0 ;
  assign n2575 = n2574 ^ n2573 ^ n1243 ;
  assign n2576 = ( n514 & n633 ) | ( n514 & n2261 ) | ( n633 & n2261 ) ;
  assign n2577 = n1226 ^ x85 ^ 1'b0 ;
  assign n2578 = n1616 & ~n2577 ;
  assign n2579 = n2578 ^ n1631 ^ 1'b0 ;
  assign n2580 = n1336 & n2579 ;
  assign n2581 = n813 & n1372 ;
  assign n2582 = ~n2580 & n2581 ;
  assign n2583 = ( ~n1117 & n1605 ) | ( ~n1117 & n1782 ) | ( n1605 & n1782 ) ;
  assign n2584 = n2583 ^ n1006 ^ n886 ;
  assign n2585 = n443 | n2584 ;
  assign n2586 = ~x222 & n872 ;
  assign n2587 = n516 & n1461 ;
  assign n2588 = n2587 ^ x3 ^ 1'b0 ;
  assign n2589 = n2588 ^ n843 ^ 1'b0 ;
  assign n2590 = x4 & n2589 ;
  assign n2591 = n2586 & n2590 ;
  assign n2592 = ~n521 & n2591 ;
  assign n2593 = ( n348 & n1499 ) | ( n348 & n2592 ) | ( n1499 & n2592 ) ;
  assign n2594 = n2593 ^ n2006 ^ n1603 ;
  assign n2596 = x10 & x40 ;
  assign n2595 = n1733 ^ n499 ^ 1'b0 ;
  assign n2597 = n2596 ^ n2595 ^ n1687 ;
  assign n2598 = ~n1211 & n1913 ;
  assign n2599 = ~n1484 & n2598 ;
  assign n2600 = n1859 | n2599 ;
  assign n2601 = ( ~n1252 & n1802 ) | ( ~n1252 & n2600 ) | ( n1802 & n2600 ) ;
  assign n2602 = n2296 ^ n1666 ^ n584 ;
  assign n2603 = n284 ^ x170 ^ 1'b0 ;
  assign n2604 = n1605 & ~n2603 ;
  assign n2605 = n2215 ^ n773 ^ 1'b0 ;
  assign n2606 = x98 & n2605 ;
  assign n2607 = n2606 ^ n1462 ^ 1'b0 ;
  assign n2608 = ( n299 & n1219 ) | ( n299 & n1932 ) | ( n1219 & n1932 ) ;
  assign n2609 = ~n1397 & n2608 ;
  assign n2610 = ~n1804 & n2609 ;
  assign n2611 = ( n2604 & ~n2607 ) | ( n2604 & n2610 ) | ( ~n2607 & n2610 ) ;
  assign n2612 = x3 & ~n787 ;
  assign n2613 = ~n2354 & n2612 ;
  assign n2614 = n1080 ^ n807 ^ x39 ;
  assign n2615 = ( n363 & n584 ) | ( n363 & ~n1148 ) | ( n584 & ~n1148 ) ;
  assign n2616 = n1352 ^ x114 ^ 1'b0 ;
  assign n2617 = n2203 ^ n1188 ^ 1'b0 ;
  assign n2618 = n2407 & ~n2617 ;
  assign n2619 = ~x106 & n2618 ;
  assign n2620 = n532 & ~n2619 ;
  assign n2621 = n1050 | n1658 ;
  assign n2622 = x186 & ~n2621 ;
  assign n2623 = n2622 ^ n810 ^ 1'b0 ;
  assign n2624 = n2623 ^ n1873 ^ n576 ;
  assign n2629 = n1526 ^ n406 ^ 1'b0 ;
  assign n2630 = ( x35 & ~x56 ) | ( x35 & n2629 ) | ( ~x56 & n2629 ) ;
  assign n2625 = n482 & n1454 ;
  assign n2626 = n2625 ^ n1537 ^ 1'b0 ;
  assign n2627 = n579 & ~n1241 ;
  assign n2628 = ~n2626 & n2627 ;
  assign n2631 = n2630 ^ n2628 ^ n1191 ;
  assign n2632 = x140 & x212 ;
  assign n2633 = ~n2398 & n2632 ;
  assign n2634 = n2633 ^ n1380 ^ n656 ;
  assign n2635 = n455 & ~n769 ;
  assign n2636 = n1885 & ~n2635 ;
  assign n2637 = n2636 ^ n1650 ^ 1'b0 ;
  assign n2638 = n2450 ^ n1796 ^ n1483 ;
  assign n2639 = ~n662 & n2638 ;
  assign n2640 = ~n1176 & n1903 ;
  assign n2641 = n2640 ^ n2472 ^ 1'b0 ;
  assign n2642 = n640 & ~n2641 ;
  assign n2643 = n1338 ^ n1174 ^ 1'b0 ;
  assign n2644 = n2643 ^ n608 ^ 1'b0 ;
  assign n2645 = ~n1027 & n2644 ;
  assign n2646 = n2645 ^ n1030 ^ 1'b0 ;
  assign n2648 = n379 | n1701 ;
  assign n2649 = n1783 | n2648 ;
  assign n2647 = ( ~x132 & n1635 ) | ( ~x132 & n1816 ) | ( n1635 & n1816 ) ;
  assign n2650 = n2649 ^ n2647 ^ 1'b0 ;
  assign n2651 = n544 & n2650 ;
  assign n2652 = ~n502 & n644 ;
  assign n2653 = ~n1503 & n2652 ;
  assign n2654 = ~x63 & n1629 ;
  assign n2655 = n2653 | n2654 ;
  assign n2657 = n2507 ^ n871 ^ n618 ;
  assign n2658 = n1142 & ~n2657 ;
  assign n2659 = n2658 ^ n1787 ^ 1'b0 ;
  assign n2660 = n1736 & n2659 ;
  assign n2661 = n2660 ^ n1323 ^ 1'b0 ;
  assign n2656 = ~n2071 & n2441 ;
  assign n2662 = n2661 ^ n2656 ^ 1'b0 ;
  assign n2663 = n2638 ^ n2028 ^ 1'b0 ;
  assign n2664 = x140 & ~n1520 ;
  assign n2665 = n2664 ^ n1251 ^ 1'b0 ;
  assign n2666 = ( ~n1009 & n1176 ) | ( ~n1009 & n2665 ) | ( n1176 & n2665 ) ;
  assign n2667 = n1403 ^ n406 ^ 1'b0 ;
  assign n2668 = n645 ^ n318 ^ 1'b0 ;
  assign n2669 = n2668 ^ n1806 ^ 1'b0 ;
  assign n2670 = x87 | n2669 ;
  assign n2671 = n2670 ^ n366 ^ 1'b0 ;
  assign n2672 = ~n2667 & n2671 ;
  assign n2673 = n1380 & n2280 ;
  assign n2674 = ~n1231 & n1812 ;
  assign n2675 = n2674 ^ n730 ^ 1'b0 ;
  assign n2676 = n1267 ^ x125 ^ 1'b0 ;
  assign n2677 = ( n1136 & ~n1353 ) | ( n1136 & n2335 ) | ( ~n1353 & n2335 ) ;
  assign n2678 = n783 | n2677 ;
  assign n2679 = n2678 ^ n1378 ^ 1'b0 ;
  assign n2680 = n1674 ^ x15 ^ 1'b0 ;
  assign n2681 = n2680 ^ n1919 ^ 1'b0 ;
  assign n2682 = n545 & n2681 ;
  assign n2683 = n2682 ^ n1154 ^ n373 ;
  assign n2685 = n2017 ^ n1155 ^ n330 ;
  assign n2686 = ( n893 & n1644 ) | ( n893 & ~n2685 ) | ( n1644 & ~n2685 ) ;
  assign n2687 = ( n532 & n614 ) | ( n532 & ~n2686 ) | ( n614 & ~n2686 ) ;
  assign n2684 = ~x162 & n1381 ;
  assign n2688 = n2687 ^ n2684 ^ 1'b0 ;
  assign n2689 = n1067 ^ n560 ^ n262 ;
  assign n2690 = n1811 & ~n2689 ;
  assign n2691 = ~n391 & n2690 ;
  assign n2692 = ~x232 & n479 ;
  assign n2693 = n2692 ^ x37 ^ x23 ;
  assign n2694 = ~n1014 & n1511 ;
  assign n2695 = n1934 & ~n2694 ;
  assign n2696 = ( x84 & x152 ) | ( x84 & ~n733 ) | ( x152 & ~n733 ) ;
  assign n2697 = n1861 ^ n993 ^ x92 ;
  assign n2698 = n2696 & n2697 ;
  assign n2699 = n1438 & ~n2698 ;
  assign n2700 = n751 ^ n448 ^ n362 ;
  assign n2701 = ( ~x202 & n595 ) | ( ~x202 & n1454 ) | ( n595 & n1454 ) ;
  assign n2702 = ( x190 & n2700 ) | ( x190 & ~n2701 ) | ( n2700 & ~n2701 ) ;
  assign n2703 = ~n1092 & n2702 ;
  assign n2704 = ~n973 & n2703 ;
  assign n2705 = n921 ^ n816 ^ x0 ;
  assign n2706 = n352 | n1848 ;
  assign n2707 = n2706 ^ n272 ^ 1'b0 ;
  assign n2708 = n2333 & ~n2707 ;
  assign n2709 = n2708 ^ n1816 ^ 1'b0 ;
  assign n2710 = ( x4 & n2705 ) | ( x4 & n2709 ) | ( n2705 & n2709 ) ;
  assign n2711 = ( ~n1460 & n1542 ) | ( ~n1460 & n2710 ) | ( n1542 & n2710 ) ;
  assign n2712 = ( n1158 & ~n2170 ) | ( n1158 & n2711 ) | ( ~n2170 & n2711 ) ;
  assign n2713 = x99 & x143 ;
  assign n2714 = ~n999 & n2713 ;
  assign n2715 = n1156 & ~n2714 ;
  assign n2716 = n2715 ^ x3 ^ 1'b0 ;
  assign n2717 = x178 & n345 ;
  assign n2718 = ~n511 & n2717 ;
  assign n2719 = n2425 | n2718 ;
  assign n2720 = n2206 ^ n813 ^ 1'b0 ;
  assign n2721 = n2720 ^ n1461 ^ 1'b0 ;
  assign n2722 = ( x36 & ~x165 ) | ( x36 & n575 ) | ( ~x165 & n575 ) ;
  assign n2723 = n1391 ^ n590 ^ n326 ;
  assign n2724 = ( n1114 & ~n2705 ) | ( n1114 & n2723 ) | ( ~n2705 & n2723 ) ;
  assign n2725 = ( n1961 & n2125 ) | ( n1961 & n2724 ) | ( n2125 & n2724 ) ;
  assign n2726 = ( n403 & n2425 ) | ( n403 & ~n2725 ) | ( n2425 & ~n2725 ) ;
  assign n2727 = n875 & ~n1810 ;
  assign n2728 = n2727 ^ x27 ^ 1'b0 ;
  assign n2729 = n673 | n2728 ;
  assign n2730 = n2729 ^ n282 ^ 1'b0 ;
  assign n2731 = n2354 ^ n2068 ^ 1'b0 ;
  assign n2732 = n2731 ^ n436 ^ 1'b0 ;
  assign n2733 = ( x160 & ~x193 ) | ( x160 & n1506 ) | ( ~x193 & n1506 ) ;
  assign n2734 = n290 & n578 ;
  assign n2735 = n1351 & n2734 ;
  assign n2736 = x146 & ~n1222 ;
  assign n2737 = ~x114 & n2736 ;
  assign n2738 = ( x171 & n835 ) | ( x171 & n1374 ) | ( n835 & n1374 ) ;
  assign n2739 = n2738 ^ n1971 ^ n1590 ;
  assign n2740 = x127 & ~n1290 ;
  assign n2741 = ( n2737 & n2739 ) | ( n2737 & ~n2740 ) | ( n2739 & ~n2740 ) ;
  assign n2742 = x126 & ~n1611 ;
  assign n2743 = n2742 ^ n1939 ^ 1'b0 ;
  assign n2744 = n404 & ~n2743 ;
  assign n2745 = ( n822 & ~n1512 ) | ( n822 & n1793 ) | ( ~n1512 & n1793 ) ;
  assign n2746 = ( x2 & ~n552 ) | ( x2 & n621 ) | ( ~n552 & n621 ) ;
  assign n2747 = n2746 ^ n2645 ^ n491 ;
  assign n2748 = n2747 ^ n1006 ^ n774 ;
  assign n2749 = x155 & n916 ;
  assign n2750 = ( x102 & n793 ) | ( x102 & n1338 ) | ( n793 & n1338 ) ;
  assign n2751 = n2221 ^ n724 ^ 1'b0 ;
  assign n2752 = n2750 & ~n2751 ;
  assign n2753 = ( n2448 & n2749 ) | ( n2448 & ~n2752 ) | ( n2749 & ~n2752 ) ;
  assign n2754 = n1664 ^ n949 ^ n806 ;
  assign n2755 = n2754 ^ n733 ^ x129 ;
  assign n2758 = n353 & n1098 ;
  assign n2759 = ( n2145 & ~n2178 ) | ( n2145 & n2758 ) | ( ~n2178 & n2758 ) ;
  assign n2756 = x209 & ~n1187 ;
  assign n2757 = n2756 ^ x190 ^ 1'b0 ;
  assign n2760 = n2759 ^ n2757 ^ 1'b0 ;
  assign n2764 = n886 ^ n791 ^ 1'b0 ;
  assign n2763 = n1135 ^ n944 ^ x188 ;
  assign n2765 = n2764 ^ n2763 ^ n2039 ;
  assign n2761 = n1736 ^ n1552 ^ x238 ;
  assign n2762 = n2330 & ~n2761 ;
  assign n2766 = n2765 ^ n2762 ^ 1'b0 ;
  assign n2767 = ( ~x228 & n346 ) | ( ~x228 & n832 ) | ( n346 & n832 ) ;
  assign n2768 = n2767 ^ n1952 ^ x21 ;
  assign n2769 = n1398 ^ n355 ^ x174 ;
  assign n2770 = n1601 ^ n776 ^ n597 ;
  assign n2771 = ( n352 & ~n2769 ) | ( n352 & n2770 ) | ( ~n2769 & n2770 ) ;
  assign n2772 = n2156 ^ n1861 ^ 1'b0 ;
  assign n2773 = n1117 & n2772 ;
  assign n2774 = ( n1384 & n1919 ) | ( n1384 & n2773 ) | ( n1919 & n2773 ) ;
  assign n2775 = x143 & n2774 ;
  assign n2776 = n826 ^ n274 ^ 1'b0 ;
  assign n2777 = x73 & ~n2776 ;
  assign n2778 = ( n1116 & n1743 ) | ( n1116 & n2777 ) | ( n1743 & n2777 ) ;
  assign n2779 = n2778 ^ n1035 ^ n733 ;
  assign n2780 = ( n1838 & ~n2191 ) | ( n1838 & n2779 ) | ( ~n2191 & n2779 ) ;
  assign n2781 = n1327 & ~n2780 ;
  assign n2782 = ( x159 & ~n534 ) | ( x159 & n2781 ) | ( ~n534 & n2781 ) ;
  assign n2783 = ~n718 & n2367 ;
  assign n2784 = n2783 ^ n687 ^ 1'b0 ;
  assign n2785 = x20 & n2784 ;
  assign n2786 = n2785 ^ n2696 ^ 1'b0 ;
  assign n2787 = n1409 ^ x236 ^ 1'b0 ;
  assign n2788 = n322 | n2787 ;
  assign n2789 = n2788 ^ n706 ^ n578 ;
  assign n2790 = n2789 ^ n2203 ^ x139 ;
  assign n2791 = ( n1656 & n2786 ) | ( n1656 & n2790 ) | ( n2786 & n2790 ) ;
  assign n2792 = n1132 ^ n1044 ^ n542 ;
  assign n2793 = n2792 ^ x137 ^ 1'b0 ;
  assign n2794 = ( n887 & ~n2791 ) | ( n887 & n2793 ) | ( ~n2791 & n2793 ) ;
  assign n2795 = ( ~x202 & n1280 ) | ( ~x202 & n2369 ) | ( n1280 & n2369 ) ;
  assign n2796 = n1320 ^ n446 ^ x240 ;
  assign n2797 = n666 ^ x254 ^ 1'b0 ;
  assign n2798 = ~n2796 & n2797 ;
  assign n2799 = ~n2795 & n2798 ;
  assign n2800 = ~n800 & n2799 ;
  assign n2801 = n1830 & n1854 ;
  assign n2802 = n2801 ^ n343 ^ 1'b0 ;
  assign n2803 = n2802 ^ n2503 ^ 1'b0 ;
  assign n2804 = x11 & n2803 ;
  assign n2805 = ~n790 & n2804 ;
  assign n2806 = n618 ^ x201 ^ 1'b0 ;
  assign n2807 = n2399 & n2806 ;
  assign n2808 = n1906 ^ n1563 ^ 1'b0 ;
  assign n2810 = n855 ^ n297 ^ 1'b0 ;
  assign n2811 = ~n722 & n2810 ;
  assign n2809 = n516 & ~n1985 ;
  assign n2812 = n2811 ^ n2809 ^ 1'b0 ;
  assign n2813 = n1475 | n2812 ;
  assign n2814 = x191 | n2813 ;
  assign n2815 = n949 & ~n2761 ;
  assign n2816 = n1274 | n1446 ;
  assign n2817 = ~n2631 & n2816 ;
  assign n2818 = ~n1944 & n2817 ;
  assign n2819 = ~x14 & n426 ;
  assign n2820 = n1391 ^ n1043 ^ 1'b0 ;
  assign n2821 = ~n2819 & n2820 ;
  assign n2822 = x37 & ~n2821 ;
  assign n2823 = n432 ^ n393 ^ x218 ;
  assign n2824 = ( x44 & n449 ) | ( x44 & ~n2823 ) | ( n449 & ~n2823 ) ;
  assign n2831 = x156 & n841 ;
  assign n2832 = ~n551 & n2831 ;
  assign n2827 = n277 & n654 ;
  assign n2828 = n2827 ^ n1896 ^ 1'b0 ;
  assign n2829 = n851 & n1197 ;
  assign n2830 = ~n2828 & n2829 ;
  assign n2833 = n2832 ^ n2830 ^ n1006 ;
  assign n2825 = ( ~n473 & n1183 ) | ( ~n473 & n1469 ) | ( n1183 & n1469 ) ;
  assign n2826 = n2117 | n2825 ;
  assign n2834 = n2833 ^ n2826 ^ 1'b0 ;
  assign n2835 = n1687 | n1759 ;
  assign n2836 = n2506 ^ n2117 ^ 1'b0 ;
  assign n2837 = n2778 ^ n2529 ^ 1'b0 ;
  assign n2838 = n1555 | n2837 ;
  assign n2842 = x7 & ~x106 ;
  assign n2843 = ~x8 & n2842 ;
  assign n2844 = ~x153 & n365 ;
  assign n2845 = ~n1127 & n2844 ;
  assign n2846 = n2843 & n2845 ;
  assign n2839 = n2277 ^ n464 ^ x38 ;
  assign n2840 = n2839 ^ n2151 ^ 1'b0 ;
  assign n2841 = n2840 ^ n1787 ^ n1334 ;
  assign n2847 = n2846 ^ n2841 ^ n1660 ;
  assign n2848 = n2796 ^ n2215 ^ 1'b0 ;
  assign n2849 = ~n2847 & n2848 ;
  assign n2850 = n1108 ^ n695 ^ x226 ;
  assign n2851 = ~n2145 & n2850 ;
  assign n2852 = n2409 ^ n1708 ^ 1'b0 ;
  assign n2853 = n2851 & n2852 ;
  assign n2854 = n2853 ^ x96 ^ 1'b0 ;
  assign n2857 = n1478 ^ n789 ^ 1'b0 ;
  assign n2858 = n1986 | n2857 ;
  assign n2859 = n1088 ^ x115 ^ 1'b0 ;
  assign n2860 = n2859 ^ n1917 ^ n1290 ;
  assign n2861 = ( n756 & n2858 ) | ( n756 & n2860 ) | ( n2858 & n2860 ) ;
  assign n2855 = n585 ^ n291 ^ 1'b0 ;
  assign n2856 = n2297 | n2855 ;
  assign n2862 = n2861 ^ n2856 ^ n971 ;
  assign n2863 = x147 & ~n305 ;
  assign n2864 = n2863 ^ x50 ^ 1'b0 ;
  assign n2865 = x250 & ~n2864 ;
  assign n2866 = n2211 & n2865 ;
  assign n2867 = ~n1545 & n2866 ;
  assign n2868 = n1801 ^ n506 ^ 1'b0 ;
  assign n2869 = n2868 ^ n1562 ^ 1'b0 ;
  assign n2870 = n2492 ^ n619 ^ 1'b0 ;
  assign n2871 = n735 & n1475 ;
  assign n2872 = n720 & n1866 ;
  assign n2874 = n1418 | n2134 ;
  assign n2875 = x124 | n2874 ;
  assign n2876 = n930 & ~n1397 ;
  assign n2877 = x240 & n2876 ;
  assign n2878 = n2875 & ~n2877 ;
  assign n2879 = n2495 ^ n1112 ^ 1'b0 ;
  assign n2880 = n2878 | n2879 ;
  assign n2881 = x248 & ~n949 ;
  assign n2882 = n2031 ^ n820 ^ 1'b0 ;
  assign n2883 = n1482 & ~n2882 ;
  assign n2884 = ( n1468 & ~n2881 ) | ( n1468 & n2883 ) | ( ~n2881 & n2883 ) ;
  assign n2885 = n1075 & ~n2884 ;
  assign n2886 = n2880 & n2885 ;
  assign n2873 = ~n925 & n1377 ;
  assign n2887 = n2886 ^ n2873 ^ 1'b0 ;
  assign n2888 = n544 & ~n1123 ;
  assign n2889 = n2888 ^ x254 ^ 1'b0 ;
  assign n2890 = n2422 ^ n1301 ^ n515 ;
  assign n2891 = n2890 ^ n1973 ^ 1'b0 ;
  assign n2892 = x91 & n2891 ;
  assign n2895 = ~n758 & n2654 ;
  assign n2896 = n877 & n2895 ;
  assign n2893 = n1805 ^ n1012 ^ 1'b0 ;
  assign n2894 = ~n1440 & n2893 ;
  assign n2897 = n2896 ^ n2894 ^ n1016 ;
  assign n2898 = n665 & n1632 ;
  assign n2899 = n2898 ^ n515 ^ 1'b0 ;
  assign n2900 = n1608 | n2899 ;
  assign n2901 = n1591 | n2900 ;
  assign n2902 = n1458 & n2340 ;
  assign n2903 = ~n1194 & n2902 ;
  assign n2905 = n921 ^ n528 ^ x0 ;
  assign n2906 = ( n1362 & n2305 ) | ( n1362 & n2905 ) | ( n2305 & n2905 ) ;
  assign n2904 = n1220 ^ x92 ^ 1'b0 ;
  assign n2907 = n2906 ^ n2904 ^ 1'b0 ;
  assign n2908 = ~n2903 & n2907 ;
  assign n2912 = n907 | n2689 ;
  assign n2913 = n2912 ^ n297 ^ x0 ;
  assign n2914 = n2913 ^ n1963 ^ n327 ;
  assign n2915 = n2714 | n2914 ;
  assign n2916 = n2915 ^ n1941 ^ 1'b0 ;
  assign n2909 = n949 ^ n464 ^ x184 ;
  assign n2910 = x142 & n1133 ;
  assign n2911 = n2909 & n2910 ;
  assign n2917 = n2916 ^ n2911 ^ n2148 ;
  assign n2918 = n1547 ^ n1340 ^ 1'b0 ;
  assign n2919 = n2918 ^ n687 ^ x239 ;
  assign n2920 = n2578 ^ n2286 ^ 1'b0 ;
  assign n2921 = ~n997 & n2920 ;
  assign n2925 = ( ~x0 & x44 ) | ( ~x0 & x92 ) | ( x44 & x92 ) ;
  assign n2926 = n2925 ^ x250 ^ 1'b0 ;
  assign n2927 = n1198 & n2926 ;
  assign n2922 = x82 & ~n608 ;
  assign n2923 = n2922 ^ n1493 ^ 1'b0 ;
  assign n2924 = ( n1220 & n1997 ) | ( n1220 & n2923 ) | ( n1997 & n2923 ) ;
  assign n2928 = n2927 ^ n2924 ^ 1'b0 ;
  assign n2929 = n2154 & ~n2928 ;
  assign n2932 = x160 & n2031 ;
  assign n2933 = n2932 ^ n1374 ^ 1'b0 ;
  assign n2934 = n2933 ^ n1001 ^ 1'b0 ;
  assign n2930 = ~n1236 & n1864 ;
  assign n2931 = n338 | n2930 ;
  assign n2935 = n2934 ^ n2931 ^ n1569 ;
  assign n2936 = n2749 ^ n1900 ^ n1300 ;
  assign n2937 = n2936 ^ n2033 ^ n700 ;
  assign n2944 = n916 ^ x172 ^ x57 ;
  assign n2938 = x59 & n809 ;
  assign n2939 = n2938 ^ n1876 ^ 1'b0 ;
  assign n2940 = n421 | n1590 ;
  assign n2941 = n2940 ^ n1526 ^ 1'b0 ;
  assign n2942 = n2941 ^ n604 ^ 1'b0 ;
  assign n2943 = ~n2939 & n2942 ;
  assign n2945 = n2944 ^ n2943 ^ n1180 ;
  assign n2946 = ~n1133 & n2945 ;
  assign n2947 = n586 ^ n348 ^ 1'b0 ;
  assign n2948 = ( x132 & n376 ) | ( x132 & ~n1228 ) | ( n376 & ~n1228 ) ;
  assign n2949 = n1554 | n2948 ;
  assign n2950 = ~n1433 & n1545 ;
  assign n2951 = n1897 ^ n1150 ^ 1'b0 ;
  assign n2952 = n2178 | n2951 ;
  assign n2953 = n406 ^ x210 ^ 1'b0 ;
  assign n2954 = x107 & n2953 ;
  assign n2955 = ~n973 & n1062 ;
  assign n2956 = ~x75 & n2955 ;
  assign n2957 = ( n2952 & n2954 ) | ( n2952 & ~n2956 ) | ( n2954 & ~n2956 ) ;
  assign n2958 = ( ~n1360 & n2952 ) | ( ~n1360 & n2957 ) | ( n2952 & n2957 ) ;
  assign n2959 = n787 | n1861 ;
  assign n2960 = n2633 & ~n2959 ;
  assign n2961 = ( n891 & n2778 ) | ( n891 & n2960 ) | ( n2778 & n2960 ) ;
  assign n2962 = n2961 ^ n1128 ^ 1'b0 ;
  assign n2963 = ~n2958 & n2962 ;
  assign n2964 = n2950 & n2963 ;
  assign n2965 = ~x19 & n2964 ;
  assign n2966 = n2434 ^ n756 ^ x56 ;
  assign n2967 = n1901 & ~n2966 ;
  assign n2968 = ~x74 & n605 ;
  assign n2969 = n1778 ^ n956 ^ 1'b0 ;
  assign n2970 = ~n2968 & n2969 ;
  assign n2971 = n2970 ^ n783 ^ x98 ;
  assign n2972 = n2523 ^ n1535 ^ 1'b0 ;
  assign n2974 = x45 & n1634 ;
  assign n2973 = n533 & ~n1393 ;
  assign n2975 = n2974 ^ n2973 ^ 1'b0 ;
  assign n2976 = n883 ^ n734 ^ 1'b0 ;
  assign n2977 = n528 & n2976 ;
  assign n2978 = ( n936 & ~n1552 ) | ( n936 & n2700 ) | ( ~n1552 & n2700 ) ;
  assign n2982 = n1562 ^ n1137 ^ 1'b0 ;
  assign n2979 = n2495 ^ n1154 ^ 1'b0 ;
  assign n2980 = ~n1092 & n2979 ;
  assign n2981 = n2980 ^ n2186 ^ 1'b0 ;
  assign n2983 = n2982 ^ n2981 ^ 1'b0 ;
  assign n2984 = n1617 | n2305 ;
  assign n2985 = n2984 ^ n2236 ^ 1'b0 ;
  assign n2986 = x31 & ~n2519 ;
  assign n2987 = n868 & n1783 ;
  assign n2988 = x105 & n1430 ;
  assign n2989 = n2988 ^ n657 ^ 1'b0 ;
  assign n2990 = n1664 ^ n523 ^ 1'b0 ;
  assign n2991 = n2989 & n2990 ;
  assign n2992 = n2991 ^ n2970 ^ 1'b0 ;
  assign n2993 = x44 & n2992 ;
  assign n2994 = n2783 ^ n2134 ^ 1'b0 ;
  assign n2995 = n2994 ^ n961 ^ 1'b0 ;
  assign n2996 = n1560 | n2995 ;
  assign n2997 = n633 | n2996 ;
  assign n2998 = n748 & n2490 ;
  assign n2999 = ( x10 & ~n757 ) | ( x10 & n2998 ) | ( ~n757 & n2998 ) ;
  assign n3000 = n2999 ^ n2322 ^ n1478 ;
  assign n3001 = n3000 ^ n2398 ^ 1'b0 ;
  assign n3002 = x22 & ~n747 ;
  assign n3003 = ( ~n912 & n2593 ) | ( ~n912 & n3002 ) | ( n2593 & n3002 ) ;
  assign n3004 = n469 | n2296 ;
  assign n3005 = n2707 ^ n2065 ^ 1'b0 ;
  assign n3006 = n1629 & ~n3005 ;
  assign n3007 = n3006 ^ n1586 ^ 1'b0 ;
  assign n3008 = n421 | n3007 ;
  assign n3009 = n2051 | n3008 ;
  assign n3010 = n3009 ^ n618 ^ x96 ;
  assign n3011 = n941 & n2527 ;
  assign n3012 = n907 & n3011 ;
  assign n3013 = n652 & n2215 ;
  assign n3015 = n536 & ~n2406 ;
  assign n3014 = x179 & ~n1608 ;
  assign n3016 = n3015 ^ n3014 ^ 1'b0 ;
  assign n3020 = n389 & n2313 ;
  assign n3021 = n3020 ^ x73 ^ 1'b0 ;
  assign n3017 = n1380 ^ n956 ^ 1'b0 ;
  assign n3018 = ~n1723 & n3017 ;
  assign n3019 = n3018 ^ x45 ^ 1'b0 ;
  assign n3022 = n3021 ^ n3019 ^ n2654 ;
  assign n3023 = ( n1344 & n1506 ) | ( n1344 & ~n2489 ) | ( n1506 & ~n2489 ) ;
  assign n3024 = n771 & ~n937 ;
  assign n3025 = n3024 ^ n598 ^ 1'b0 ;
  assign n3026 = ~n894 & n3025 ;
  assign n3027 = ~n2662 & n3026 ;
  assign n3030 = n1245 ^ n485 ^ n341 ;
  assign n3028 = n662 ^ x231 ^ 1'b0 ;
  assign n3029 = n1006 | n3028 ;
  assign n3031 = n3030 ^ n3029 ^ 1'b0 ;
  assign n3032 = ( n547 & ~n695 ) | ( n547 & n2059 ) | ( ~n695 & n2059 ) ;
  assign n3033 = n3032 ^ n1465 ^ x10 ;
  assign n3034 = n1983 ^ x33 ^ 1'b0 ;
  assign n3035 = ( n293 & n370 ) | ( n293 & ~n3034 ) | ( n370 & ~n3034 ) ;
  assign n3036 = n2007 ^ x30 ^ 1'b0 ;
  assign n3037 = n3035 & n3036 ;
  assign n3038 = n680 | n1212 ;
  assign n3039 = ( x32 & x80 ) | ( x32 & ~x230 ) | ( x80 & ~x230 ) ;
  assign n3040 = ( x44 & n787 ) | ( x44 & ~n1250 ) | ( n787 & ~n1250 ) ;
  assign n3041 = ( ~n855 & n1411 ) | ( ~n855 & n3040 ) | ( n1411 & n3040 ) ;
  assign n3042 = x91 & ~n648 ;
  assign n3043 = n1726 ^ n1245 ^ 1'b0 ;
  assign n3044 = n3043 ^ x232 ^ 1'b0 ;
  assign n3045 = n3042 | n3044 ;
  assign n3046 = n863 & ~n3045 ;
  assign n3047 = n404 & ~n1066 ;
  assign n3048 = ~x14 & n3047 ;
  assign n3049 = ( ~n279 & n1054 ) | ( ~n279 & n3048 ) | ( n1054 & n3048 ) ;
  assign n3050 = ( ~n532 & n1299 ) | ( ~n532 & n1748 ) | ( n1299 & n1748 ) ;
  assign n3051 = n3049 & ~n3050 ;
  assign n3052 = n3046 & n3051 ;
  assign n3053 = n2047 & ~n3052 ;
  assign n3054 = n3053 ^ n376 ^ 1'b0 ;
  assign n3055 = ( n3039 & n3041 ) | ( n3039 & n3054 ) | ( n3041 & n3054 ) ;
  assign n3057 = x116 ^ x24 ^ 1'b0 ;
  assign n3058 = n285 & n3057 ;
  assign n3056 = n2645 ^ n2251 ^ x10 ;
  assign n3059 = n3058 ^ n3056 ^ n2791 ;
  assign n3060 = n2179 ^ n1710 ^ 1'b0 ;
  assign n3061 = ( n629 & n1077 ) | ( n629 & n2374 ) | ( n1077 & n2374 ) ;
  assign n3062 = ~n352 & n2573 ;
  assign n3063 = ( ~n326 & n3061 ) | ( ~n326 & n3062 ) | ( n3061 & n3062 ) ;
  assign n3064 = x159 & n516 ;
  assign n3065 = ~n879 & n3064 ;
  assign n3066 = n3065 ^ n1812 ^ 1'b0 ;
  assign n3067 = x118 ^ x4 ^ 1'b0 ;
  assign n3068 = n3067 ^ n626 ^ 1'b0 ;
  assign n3069 = ~n3066 & n3068 ;
  assign n3070 = ( n728 & n1489 ) | ( n728 & n3029 ) | ( n1489 & n3029 ) ;
  assign n3073 = n1264 ^ n1081 ^ 1'b0 ;
  assign n3074 = n3073 ^ n1851 ^ x107 ;
  assign n3071 = ~x149 & n1194 ;
  assign n3072 = x132 | n3071 ;
  assign n3075 = n3074 ^ n3072 ^ x5 ;
  assign n3076 = x142 & x186 ;
  assign n3077 = n3076 ^ x206 ^ 1'b0 ;
  assign n3078 = x241 & ~n687 ;
  assign n3079 = n2215 & n3078 ;
  assign n3080 = n3079 ^ n1261 ^ x118 ;
  assign n3081 = n3080 ^ n1672 ^ 1'b0 ;
  assign n3082 = n256 & ~n3081 ;
  assign n3083 = n3082 ^ n2701 ^ x214 ;
  assign n3084 = n1346 | n2689 ;
  assign n3085 = n2950 | n3084 ;
  assign n3088 = n636 ^ n632 ^ x207 ;
  assign n3086 = x126 & ~n1337 ;
  assign n3087 = n3086 ^ n1276 ^ 1'b0 ;
  assign n3089 = n3088 ^ n3087 ^ 1'b0 ;
  assign n3090 = n409 | n1028 ;
  assign n3091 = x253 | n3090 ;
  assign n3092 = n553 | n692 ;
  assign n3093 = n629 | n3092 ;
  assign n3094 = n757 ^ n631 ^ n317 ;
  assign n3095 = ( x66 & x246 ) | ( x66 & n990 ) | ( x246 & n990 ) ;
  assign n3096 = n3095 ^ n2414 ^ n558 ;
  assign n3097 = n826 ^ n452 ^ 1'b0 ;
  assign n3098 = n454 & ~n3097 ;
  assign n3099 = ~x158 & n3098 ;
  assign n3100 = x106 | n3099 ;
  assign n3101 = ( ~n392 & n995 ) | ( ~n392 & n1011 ) | ( n995 & n1011 ) ;
  assign n3102 = n3101 ^ n1667 ^ 1'b0 ;
  assign n3103 = n764 | n3102 ;
  assign n3105 = n2489 ^ n1988 ^ x241 ;
  assign n3104 = ( ~x138 & x242 ) | ( ~x138 & n633 ) | ( x242 & n633 ) ;
  assign n3106 = n3105 ^ n3104 ^ n2267 ;
  assign n3107 = n3006 ^ n2104 ^ 1'b0 ;
  assign n3108 = ~n432 & n1539 ;
  assign n3109 = n3108 ^ n639 ^ 1'b0 ;
  assign n3110 = n3109 ^ x250 ^ 1'b0 ;
  assign n3111 = n2039 ^ n1560 ^ n363 ;
  assign n3112 = ( n1132 & n1598 ) | ( n1132 & n2524 ) | ( n1598 & n2524 ) ;
  assign n3113 = ( ~n1503 & n3111 ) | ( ~n1503 & n3112 ) | ( n3111 & n3112 ) ;
  assign n3114 = n825 ^ n510 ^ n430 ;
  assign n3115 = ( ~x34 & x221 ) | ( ~x34 & x254 ) | ( x221 & x254 ) ;
  assign n3116 = ( n687 & ~n1163 ) | ( n687 & n3115 ) | ( ~n1163 & n3115 ) ;
  assign n3117 = n2549 ^ n871 ^ x66 ;
  assign n3118 = ( n1409 & ~n3116 ) | ( n1409 & n3117 ) | ( ~n3116 & n3117 ) ;
  assign n3119 = n2467 | n3118 ;
  assign n3120 = n3114 | n3119 ;
  assign n3121 = x101 ^ x14 ^ 1'b0 ;
  assign n3122 = ( ~n734 & n1488 ) | ( ~n734 & n1873 ) | ( n1488 & n1873 ) ;
  assign n3123 = ( ~n892 & n918 ) | ( ~n892 & n2686 ) | ( n918 & n2686 ) ;
  assign n3124 = n868 ^ x112 ^ 1'b0 ;
  assign n3125 = n1717 | n3124 ;
  assign n3126 = n3125 ^ n1789 ^ 1'b0 ;
  assign n3127 = ( n821 & n3123 ) | ( n821 & ~n3126 ) | ( n3123 & ~n3126 ) ;
  assign n3128 = n436 & n3127 ;
  assign n3129 = n3128 ^ n2374 ^ 1'b0 ;
  assign n3130 = n3129 ^ n890 ^ 1'b0 ;
  assign n3131 = ~n2960 & n3130 ;
  assign n3132 = x65 & n3131 ;
  assign n3133 = n3122 & n3132 ;
  assign n3134 = n1142 ^ n720 ^ 1'b0 ;
  assign n3135 = x43 & ~n3134 ;
  assign n3136 = ~x73 & n315 ;
  assign n3137 = n2596 | n3008 ;
  assign n3138 = n3137 ^ x216 ^ 1'b0 ;
  assign n3139 = n2324 ^ n616 ^ 1'b0 ;
  assign n3140 = x15 & n3139 ;
  assign n3141 = n3140 ^ n2160 ^ n1406 ;
  assign n3142 = n3141 ^ n1963 ^ 1'b0 ;
  assign n3143 = n561 & ~n2477 ;
  assign n3144 = n3143 ^ n1460 ^ 1'b0 ;
  assign n3145 = n1873 ^ n715 ^ n461 ;
  assign n3146 = ( n990 & n3144 ) | ( n990 & n3145 ) | ( n3144 & n3145 ) ;
  assign n3147 = n2629 ^ n1134 ^ x6 ;
  assign n3156 = n2305 ^ n1723 ^ n1178 ;
  assign n3153 = n452 | n2051 ;
  assign n3154 = n3153 ^ n1053 ^ 1'b0 ;
  assign n3148 = n1961 ^ n1516 ^ x227 ;
  assign n3149 = ( ~x114 & n835 ) | ( ~x114 & n3148 ) | ( n835 & n3148 ) ;
  assign n3150 = n761 ^ n665 ^ 1'b0 ;
  assign n3151 = ~n3149 & n3150 ;
  assign n3152 = ~n2596 & n3151 ;
  assign n3155 = n3154 ^ n3152 ^ 1'b0 ;
  assign n3157 = n3156 ^ n3155 ^ n2361 ;
  assign n3158 = ~n1152 & n3157 ;
  assign n3159 = n1826 & n3158 ;
  assign n3160 = x243 & ~n949 ;
  assign n3161 = ( n763 & n2507 ) | ( n763 & ~n3160 ) | ( n2507 & ~n3160 ) ;
  assign n3162 = ( ~n614 & n1787 ) | ( ~n614 & n2299 ) | ( n1787 & n2299 ) ;
  assign n3163 = n3162 ^ n2489 ^ n1181 ;
  assign n3164 = n436 & n3163 ;
  assign n3165 = n1857 & n3164 ;
  assign n3166 = n966 ^ n652 ^ x34 ;
  assign n3168 = n2057 ^ n532 ^ 1'b0 ;
  assign n3167 = ( x236 & n1922 ) | ( x236 & ~n2077 ) | ( n1922 & ~n2077 ) ;
  assign n3169 = n3168 ^ n3167 ^ n1913 ;
  assign n3170 = ( n3165 & n3166 ) | ( n3165 & n3169 ) | ( n3166 & n3169 ) ;
  assign n3171 = n566 & n2893 ;
  assign n3172 = ( n644 & n1247 ) | ( n644 & n1360 ) | ( n1247 & n1360 ) ;
  assign n3173 = n3172 ^ x56 ^ 1'b0 ;
  assign n3174 = ( x106 & ~n1181 ) | ( x106 & n2073 ) | ( ~n1181 & n2073 ) ;
  assign n3175 = ( n818 & n2398 ) | ( n818 & n3174 ) | ( n2398 & n3174 ) ;
  assign n3176 = n3175 ^ n2343 ^ 1'b0 ;
  assign n3177 = ~n1388 & n3176 ;
  assign n3191 = x96 & n504 ;
  assign n3192 = n1736 ^ n552 ^ 1'b0 ;
  assign n3193 = n3191 & n3192 ;
  assign n3194 = n742 ^ x248 ^ 1'b0 ;
  assign n3195 = n3193 & n3194 ;
  assign n3187 = n1768 ^ n1075 ^ n722 ;
  assign n3188 = n3187 ^ n400 ^ 1'b0 ;
  assign n3189 = n2569 & ~n3188 ;
  assign n3190 = ( x114 & n1816 ) | ( x114 & ~n3189 ) | ( n1816 & ~n3189 ) ;
  assign n3178 = n2550 ^ n1745 ^ 1'b0 ;
  assign n3179 = n879 ^ n699 ^ 1'b0 ;
  assign n3180 = n428 & n3179 ;
  assign n3181 = n901 | n2221 ;
  assign n3182 = n3181 ^ x31 ^ 1'b0 ;
  assign n3183 = n3180 & n3182 ;
  assign n3184 = ~n1672 & n3183 ;
  assign n3185 = n3184 ^ n835 ^ 1'b0 ;
  assign n3186 = n3178 & n3185 ;
  assign n3196 = n3195 ^ n3190 ^ n3186 ;
  assign n3197 = ( n989 & n1499 ) | ( n989 & n3196 ) | ( n1499 & n3196 ) ;
  assign n3199 = ~n1080 & n2324 ;
  assign n3200 = n3199 ^ n2941 ^ 1'b0 ;
  assign n3201 = n2230 & ~n3200 ;
  assign n3202 = n3201 ^ x128 ^ 1'b0 ;
  assign n3203 = ( x42 & n1554 ) | ( x42 & n3202 ) | ( n1554 & n3202 ) ;
  assign n3198 = n1888 ^ n995 ^ 1'b0 ;
  assign n3204 = n3203 ^ n3198 ^ n2478 ;
  assign n3205 = n1658 & ~n2157 ;
  assign n3206 = ( x224 & ~n761 ) | ( x224 & n2024 ) | ( ~n761 & n2024 ) ;
  assign n3207 = x231 & n3206 ;
  assign n3208 = n1362 & n3207 ;
  assign n3209 = n3205 | n3208 ;
  assign n3210 = n930 ^ x206 ^ 1'b0 ;
  assign n3211 = n327 & n523 ;
  assign n3212 = n789 & n3211 ;
  assign n3215 = n326 ^ x241 ^ 1'b0 ;
  assign n3216 = n808 & n3215 ;
  assign n3217 = n983 & n3182 ;
  assign n3218 = ~n3216 & n3217 ;
  assign n3213 = n374 & n1984 ;
  assign n3214 = n1851 & n3213 ;
  assign n3219 = n3218 ^ n3214 ^ x92 ;
  assign n3220 = n637 & ~n1721 ;
  assign n3221 = n2136 ^ n656 ^ 1'b0 ;
  assign n3222 = ~n3220 & n3221 ;
  assign n3223 = n3222 ^ n2749 ^ 1'b0 ;
  assign n3224 = n2045 & ~n2367 ;
  assign n3225 = n3224 ^ n1950 ^ 1'b0 ;
  assign n3226 = n1564 ^ n830 ^ n809 ;
  assign n3227 = ( n2686 & ~n3085 ) | ( n2686 & n3226 ) | ( ~n3085 & n3226 ) ;
  assign n3228 = n2148 ^ x53 ^ x47 ;
  assign n3229 = n3228 ^ n2643 ^ 1'b0 ;
  assign n3230 = ( ~n698 & n1569 ) | ( ~n698 & n3229 ) | ( n1569 & n3229 ) ;
  assign n3231 = ~n512 & n1548 ;
  assign n3232 = n1790 ^ n1746 ^ 1'b0 ;
  assign n3233 = x130 ^ x90 ^ x30 ;
  assign n3234 = ( x45 & n665 ) | ( x45 & n2258 ) | ( n665 & n2258 ) ;
  assign n3235 = ( ~n1854 & n3233 ) | ( ~n1854 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3236 = n477 & ~n951 ;
  assign n3237 = n3236 ^ n1671 ^ 1'b0 ;
  assign n3238 = n3237 ^ n331 ^ 1'b0 ;
  assign n3239 = n2573 ^ n1154 ^ n733 ;
  assign n3240 = n1502 | n2112 ;
  assign n3241 = n3240 ^ n1336 ^ 1'b0 ;
  assign n3242 = n3239 & ~n3241 ;
  assign n3243 = n3242 ^ n958 ^ 1'b0 ;
  assign n3244 = n2103 & ~n2722 ;
  assign n3245 = ~n952 & n3244 ;
  assign n3246 = ( n634 & ~n2630 ) | ( n634 & n2710 ) | ( ~n2630 & n2710 ) ;
  assign n3251 = n1045 & n1761 ;
  assign n3249 = ( ~n408 & n735 ) | ( ~n408 & n2368 ) | ( n735 & n2368 ) ;
  assign n3247 = ( n676 & ~n1745 ) | ( n676 & n1844 ) | ( ~n1745 & n1844 ) ;
  assign n3248 = n281 & n3247 ;
  assign n3250 = n3249 ^ n3248 ^ n1035 ;
  assign n3252 = n3251 ^ n3250 ^ 1'b0 ;
  assign n3253 = x119 & ~n3252 ;
  assign n3254 = n625 | n1469 ;
  assign n3255 = n1827 ^ n1140 ^ 1'b0 ;
  assign n3256 = n337 & n3255 ;
  assign n3257 = ( n1118 & ~n3254 ) | ( n1118 & n3256 ) | ( ~n3254 & n3256 ) ;
  assign n3261 = n707 ^ n335 ^ n331 ;
  assign n3258 = n1353 ^ n551 ^ x25 ;
  assign n3259 = n3258 ^ n1098 ^ 1'b0 ;
  assign n3260 = x5 & n3259 ;
  assign n3262 = n3261 ^ n3260 ^ 1'b0 ;
  assign n3269 = n2531 ^ n307 ^ 1'b0 ;
  assign n3270 = n1761 ^ n1245 ^ 1'b0 ;
  assign n3271 = n2289 & n3270 ;
  assign n3272 = n3271 ^ n796 ^ 1'b0 ;
  assign n3273 = ( ~n984 & n3269 ) | ( ~n984 & n3272 ) | ( n3269 & n3272 ) ;
  assign n3263 = n350 | n1283 ;
  assign n3264 = n2388 & ~n3263 ;
  assign n3265 = n3264 ^ n2143 ^ 1'b0 ;
  assign n3266 = n2314 | n3265 ;
  assign n3267 = x217 & ~n3266 ;
  assign n3268 = n3267 ^ n2206 ^ 1'b0 ;
  assign n3274 = n3273 ^ n3268 ^ 1'b0 ;
  assign n3275 = n1658 ^ n1101 ^ x59 ;
  assign n3276 = ( ~n544 & n2083 ) | ( ~n544 & n3275 ) | ( n2083 & n3275 ) ;
  assign n3277 = n3276 ^ n2296 ^ 1'b0 ;
  assign n3278 = n1632 & ~n3277 ;
  assign n3279 = n853 ^ n360 ^ x96 ;
  assign n3280 = n3279 ^ n2793 ^ 1'b0 ;
  assign n3281 = n1524 & ~n1986 ;
  assign n3282 = x41 & n307 ;
  assign n3283 = n3282 ^ n1610 ^ 1'b0 ;
  assign n3284 = n2447 | n2550 ;
  assign n3285 = n3283 | n3284 ;
  assign n3286 = ~n3281 & n3285 ;
  assign n3287 = x206 & n348 ;
  assign n3288 = ~x127 & n3287 ;
  assign n3289 = n3288 ^ n980 ^ x26 ;
  assign n3290 = n1721 & n3289 ;
  assign n3291 = x61 & n459 ;
  assign n3292 = n1014 & n3291 ;
  assign n3293 = n3292 ^ x157 ^ 1'b0 ;
  assign n3294 = n886 & ~n3293 ;
  assign n3295 = n951 ^ n492 ^ 1'b0 ;
  assign n3296 = n1053 | n3295 ;
  assign n3297 = n1111 & ~n3274 ;
  assign n3298 = ( n2597 & n3296 ) | ( n2597 & n3297 ) | ( n3296 & n3297 ) ;
  assign n3299 = ( ~x188 & n2056 ) | ( ~x188 & n2113 ) | ( n2056 & n2113 ) ;
  assign n3300 = n1732 ^ x29 ^ 1'b0 ;
  assign n3301 = n1136 & n3300 ;
  assign n3302 = n1425 ^ n807 ^ 1'b0 ;
  assign n3303 = ( n524 & n1362 ) | ( n524 & ~n3302 ) | ( n1362 & ~n3302 ) ;
  assign n3304 = n355 & ~n583 ;
  assign n3305 = n976 & n3304 ;
  assign n3306 = ~n3303 & n3305 ;
  assign n3307 = ( n533 & n722 ) | ( n533 & n1048 ) | ( n722 & n1048 ) ;
  assign n3308 = x3 & ~n3307 ;
  assign n3309 = n2405 & n3308 ;
  assign n3310 = x86 | n1039 ;
  assign n3311 = ( x179 & ~n285 ) | ( x179 & n3310 ) | ( ~n285 & n3310 ) ;
  assign n3312 = n3311 ^ n1140 ^ n905 ;
  assign n3313 = ~n3309 & n3312 ;
  assign n3314 = n526 ^ n380 ^ 1'b0 ;
  assign n3315 = n2532 & ~n2927 ;
  assign n3316 = ( ~n951 & n2629 ) | ( ~n951 & n3024 ) | ( n2629 & n3024 ) ;
  assign n3317 = n678 & n1112 ;
  assign n3318 = n3317 ^ n3034 ^ n2425 ;
  assign n3319 = ( ~n1369 & n3316 ) | ( ~n1369 & n3318 ) | ( n3316 & n3318 ) ;
  assign n3320 = ( ~n1420 & n2297 ) | ( ~n1420 & n3319 ) | ( n2297 & n3319 ) ;
  assign n3321 = x51 & n1877 ;
  assign n3322 = n1669 & n2668 ;
  assign n3323 = n1896 & ~n3322 ;
  assign n3324 = n322 | n3323 ;
  assign n3326 = ( x177 & n602 ) | ( x177 & n618 ) | ( n602 & n618 ) ;
  assign n3325 = n2262 ^ n521 ^ 1'b0 ;
  assign n3327 = n3326 ^ n3325 ^ x114 ;
  assign n3328 = n1433 & ~n3327 ;
  assign n3336 = n753 ^ x209 ^ x174 ;
  assign n3337 = ( n1062 & ~n2031 ) | ( n1062 & n3336 ) | ( ~n2031 & n3336 ) ;
  assign n3330 = x230 | n2461 ;
  assign n3331 = n3330 ^ n2153 ^ n1837 ;
  assign n3332 = n3065 ^ n1497 ^ 1'b0 ;
  assign n3333 = n2583 & n3332 ;
  assign n3334 = n3331 & n3333 ;
  assign n3329 = n372 | n3101 ;
  assign n3335 = n3334 ^ n3329 ^ 1'b0 ;
  assign n3338 = n3337 ^ n3335 ^ n2871 ;
  assign n3339 = n2901 | n3338 ;
  assign n3340 = n1826 ^ n1229 ^ n609 ;
  assign n3341 = ( n988 & n1290 ) | ( n988 & ~n2290 ) | ( n1290 & ~n2290 ) ;
  assign n3342 = n3341 ^ n316 ^ 1'b0 ;
  assign n3343 = n1204 & n3342 ;
  assign n3344 = n3071 | n3341 ;
  assign n3345 = n3343 | n3344 ;
  assign n3346 = n3340 & n3345 ;
  assign n3355 = n3061 ^ n2168 ^ 1'b0 ;
  assign n3356 = ~n3029 & n3355 ;
  assign n3357 = ~n1643 & n3356 ;
  assign n3358 = n3357 ^ n404 ^ 1'b0 ;
  assign n3351 = n1461 ^ n1258 ^ 1'b0 ;
  assign n3352 = x26 & x242 ;
  assign n3353 = ~n3351 & n3352 ;
  assign n3354 = ~n3202 & n3353 ;
  assign n3359 = n3358 ^ n3354 ^ 1'b0 ;
  assign n3347 = ( x229 & ~n329 ) | ( x229 & n1299 ) | ( ~n329 & n1299 ) ;
  assign n3348 = n3347 ^ n1793 ^ 1'b0 ;
  assign n3349 = n3348 ^ n2301 ^ 1'b0 ;
  assign n3350 = ~n1249 & n3349 ;
  assign n3360 = n3359 ^ n3350 ^ 1'b0 ;
  assign n3361 = ~n376 & n3360 ;
  assign n3362 = ( ~x183 & n1783 ) | ( ~x183 & n2299 ) | ( n1783 & n2299 ) ;
  assign n3363 = n3362 ^ x116 ^ 1'b0 ;
  assign n3364 = n3363 ^ n1430 ^ 1'b0 ;
  assign n3365 = ( n771 & n2121 ) | ( n771 & n2451 ) | ( n2121 & n2451 ) ;
  assign n3366 = n1798 ^ x132 ^ x56 ;
  assign n3367 = n3365 | n3366 ;
  assign n3368 = n3367 ^ n1746 ^ 1'b0 ;
  assign n3369 = n847 & n1109 ;
  assign n3370 = n3369 ^ n1568 ^ 1'b0 ;
  assign n3371 = n1201 & ~n3370 ;
  assign n3372 = x194 & ~n2696 ;
  assign n3373 = ~n1611 & n3372 ;
  assign n3374 = n536 & n3373 ;
  assign n3375 = n3374 ^ n1264 ^ 1'b0 ;
  assign n3376 = n933 ^ x129 ^ 1'b0 ;
  assign n3377 = ( ~x252 & n1639 ) | ( ~x252 & n3376 ) | ( n1639 & n3376 ) ;
  assign n3378 = ( n2036 & n2542 ) | ( n2036 & ~n3377 ) | ( n2542 & ~n3377 ) ;
  assign n3379 = n1771 | n2909 ;
  assign n3380 = n3379 ^ n1697 ^ 1'b0 ;
  assign n3381 = ~n3331 & n3380 ;
  assign n3382 = n1102 | n1738 ;
  assign n3383 = n3382 ^ n617 ^ x10 ;
  assign n3384 = n3383 ^ n1912 ^ n1146 ;
  assign n3385 = n3384 ^ n2947 ^ n540 ;
  assign n3386 = n2966 ^ n2755 ^ 1'b0 ;
  assign n3387 = n1837 & n3386 ;
  assign n3388 = n1354 & n1753 ;
  assign n3389 = n3388 ^ n768 ^ 1'b0 ;
  assign n3390 = n3389 ^ n444 ^ 1'b0 ;
  assign n3391 = ( ~n3269 & n3387 ) | ( ~n3269 & n3390 ) | ( n3387 & n3390 ) ;
  assign n3392 = ~x106 & n1503 ;
  assign n3393 = n1269 & n1614 ;
  assign n3394 = n1957 & ~n3393 ;
  assign n3395 = n3394 ^ n1352 ^ 1'b0 ;
  assign n3396 = n3395 ^ n2952 ^ 1'b0 ;
  assign n3397 = n1355 | n3396 ;
  assign n3398 = x193 & n1142 ;
  assign n3399 = ~n1392 & n3398 ;
  assign n3400 = n378 & ~n3399 ;
  assign n3401 = n3400 ^ n929 ^ 1'b0 ;
  assign n3402 = ( x12 & n3118 ) | ( x12 & ~n3401 ) | ( n3118 & ~n3401 ) ;
  assign n3403 = n1307 & ~n1457 ;
  assign n3404 = ~n1292 & n3403 ;
  assign n3405 = ~n1029 & n1088 ;
  assign n3406 = ~x180 & n3405 ;
  assign n3407 = n3406 ^ n1346 ^ 1'b0 ;
  assign n3408 = n3407 ^ n2109 ^ 1'b0 ;
  assign n3409 = n3404 | n3408 ;
  assign n3410 = n1311 | n2280 ;
  assign n3411 = n3044 ^ n1591 ^ x218 ;
  assign n3412 = n3411 ^ x50 ^ 1'b0 ;
  assign n3413 = x117 & n3412 ;
  assign n3414 = n3413 ^ n521 ^ 1'b0 ;
  assign n3415 = ~n3410 & n3414 ;
  assign n3416 = ( ~n435 & n1156 ) | ( ~n435 & n1280 ) | ( n1156 & n1280 ) ;
  assign n3417 = n1026 & n3416 ;
  assign n3418 = x185 & n3417 ;
  assign n3419 = n3418 ^ n2279 ^ n1586 ;
  assign n3420 = x61 & ~n1026 ;
  assign n3421 = n313 & ~n2935 ;
  assign n3422 = n3420 & n3421 ;
  assign n3428 = ~x186 & n3302 ;
  assign n3429 = n2710 & n3428 ;
  assign n3430 = ( n434 & n1249 ) | ( n434 & ~n3429 ) | ( n1249 & ~n3429 ) ;
  assign n3425 = ( n597 & n2440 ) | ( n597 & ~n2907 ) | ( n2440 & ~n2907 ) ;
  assign n3426 = n2315 ^ n1735 ^ 1'b0 ;
  assign n3427 = n3425 | n3426 ;
  assign n3423 = n338 & ~n1864 ;
  assign n3424 = n2208 & n3423 ;
  assign n3431 = n3430 ^ n3427 ^ n3424 ;
  assign n3432 = ( n1276 & ~n2836 ) | ( n1276 & n3431 ) | ( ~n2836 & n3431 ) ;
  assign n3433 = ~x213 & n956 ;
  assign n3434 = n3433 ^ n3099 ^ 1'b0 ;
  assign n3435 = ( n276 & ~n410 ) | ( n276 & n1173 ) | ( ~n410 & n1173 ) ;
  assign n3436 = ~n1037 & n1571 ;
  assign n3437 = ~n929 & n1875 ;
  assign n3438 = ( n1296 & n3436 ) | ( n1296 & ~n3437 ) | ( n3436 & ~n3437 ) ;
  assign n3439 = ~n3435 & n3438 ;
  assign n3440 = ~n3434 & n3439 ;
  assign n3441 = n3074 ^ x155 ^ 1'b0 ;
  assign n3442 = ~n684 & n1709 ;
  assign n3454 = n2179 ^ n892 ^ 1'b0 ;
  assign n3455 = n718 | n3454 ;
  assign n3456 = ( n1469 & n2001 ) | ( n1469 & ~n3455 ) | ( n2001 & ~n3455 ) ;
  assign n3447 = n1016 | n1848 ;
  assign n3448 = n3447 ^ n1338 ^ 1'b0 ;
  assign n3449 = n3448 ^ n1357 ^ n791 ;
  assign n3450 = n1173 ^ n357 ^ 1'b0 ;
  assign n3451 = n2856 | n3450 ;
  assign n3452 = n3451 ^ n2354 ^ 1'b0 ;
  assign n3453 = n3449 & n3452 ;
  assign n3443 = ~n977 & n1646 ;
  assign n3444 = ~n875 & n3443 ;
  assign n3445 = n3444 ^ n886 ^ 1'b0 ;
  assign n3446 = n1811 & ~n3445 ;
  assign n3457 = n3456 ^ n3453 ^ n3446 ;
  assign n3458 = n1848 ^ n893 ^ 1'b0 ;
  assign n3459 = n1127 | n3458 ;
  assign n3460 = n3459 ^ n1072 ^ x35 ;
  assign n3461 = ~n1268 & n2450 ;
  assign n3462 = n3461 ^ n1504 ^ 1'b0 ;
  assign n3463 = n3163 ^ n2414 ^ n1333 ;
  assign n3464 = n264 & n3463 ;
  assign n3465 = n3462 & n3464 ;
  assign n3466 = n1943 ^ n1783 ^ n1493 ;
  assign n3467 = n2065 ^ n1603 ^ n1077 ;
  assign n3468 = n2289 ^ x251 ^ x174 ;
  assign n3469 = n3468 ^ n2972 ^ x97 ;
  assign n3470 = n1268 | n3469 ;
  assign n3471 = n3467 & ~n3470 ;
  assign n3472 = x177 & ~n3115 ;
  assign n3473 = n1474 | n3472 ;
  assign n3474 = n3473 ^ n495 ^ 1'b0 ;
  assign n3475 = n3474 ^ n2981 ^ 1'b0 ;
  assign n3476 = n880 ^ x227 ^ 1'b0 ;
  assign n3477 = n3436 & ~n3476 ;
  assign n3478 = n806 & n3477 ;
  assign n3479 = x80 & ~n3478 ;
  assign n3480 = n2654 ^ n2247 ^ n1198 ;
  assign n3481 = n2943 & n3480 ;
  assign n3484 = n2507 ^ n256 ^ 1'b0 ;
  assign n3485 = n2289 & ~n3484 ;
  assign n3482 = n1359 ^ n483 ^ 1'b0 ;
  assign n3483 = n3482 ^ n2616 ^ n1903 ;
  assign n3486 = n3485 ^ n3483 ^ 1'b0 ;
  assign n3487 = x118 & n3486 ;
  assign n3488 = n1543 ^ n1345 ^ 1'b0 ;
  assign n3489 = n2393 ^ n689 ^ 1'b0 ;
  assign n3490 = ~n3488 & n3489 ;
  assign n3491 = n2329 ^ n2042 ^ n272 ;
  assign n3492 = n1050 | n3491 ;
  assign n3493 = ( n388 & n804 ) | ( n388 & ~n1608 ) | ( n804 & ~n1608 ) ;
  assign n3494 = n2156 | n2906 ;
  assign n3495 = n3494 ^ n1690 ^ 1'b0 ;
  assign n3496 = ( n3492 & ~n3493 ) | ( n3492 & n3495 ) | ( ~n3493 & n3495 ) ;
  assign n3497 = n2682 ^ n1810 ^ 1'b0 ;
  assign n3498 = n1850 | n3497 ;
  assign n3499 = ( x98 & n1231 ) | ( x98 & n1375 ) | ( n1231 & n1375 ) ;
  assign n3500 = ( x250 & n365 ) | ( x250 & n3499 ) | ( n365 & n3499 ) ;
  assign n3501 = n3500 ^ n1418 ^ n633 ;
  assign n3502 = n2457 ^ x23 ^ 1'b0 ;
  assign n3503 = ( n417 & n1738 ) | ( n417 & ~n3502 ) | ( n1738 & ~n3502 ) ;
  assign n3504 = ( n3498 & n3501 ) | ( n3498 & n3503 ) | ( n3501 & n3503 ) ;
  assign n3505 = x68 & ~n1898 ;
  assign n3506 = n3505 ^ n2321 ^ 1'b0 ;
  assign n3508 = n1522 ^ n1183 ^ n595 ;
  assign n3507 = ( x210 & ~n767 ) | ( x210 & n867 ) | ( ~n767 & n867 ) ;
  assign n3509 = n3508 ^ n3507 ^ 1'b0 ;
  assign n3510 = n3509 ^ n2518 ^ 1'b0 ;
  assign n3511 = n1127 ^ n1026 ^ x180 ;
  assign n3512 = n3511 ^ n1442 ^ n726 ;
  assign n3513 = n2599 ^ n1543 ^ 1'b0 ;
  assign n3514 = ( x39 & ~n3488 ) | ( x39 & n3513 ) | ( ~n3488 & n3513 ) ;
  assign n3515 = n3514 ^ n1320 ^ 1'b0 ;
  assign n3516 = ( x185 & ~x190 ) | ( x185 & x195 ) | ( ~x190 & x195 ) ;
  assign n3517 = n3516 ^ n699 ^ 1'b0 ;
  assign n3518 = n3517 ^ n3371 ^ n2574 ;
  assign n3519 = ~n1464 & n2933 ;
  assign n3520 = n1164 & n3519 ;
  assign n3521 = n3520 ^ n3393 ^ n831 ;
  assign n3522 = n3321 ^ n2517 ^ 1'b0 ;
  assign n3523 = n1691 & ~n3522 ;
  assign n3524 = ( n1086 & n1109 ) | ( n1086 & n2545 ) | ( n1109 & n2545 ) ;
  assign n3525 = x115 & ~n350 ;
  assign n3526 = ( n457 & ~n2390 ) | ( n457 & n3525 ) | ( ~n2390 & n3525 ) ;
  assign n3527 = n3526 ^ x83 ^ 1'b0 ;
  assign n3528 = ( n341 & n3524 ) | ( n341 & n3527 ) | ( n3524 & n3527 ) ;
  assign n3529 = n1977 | n2089 ;
  assign n3530 = n2599 & ~n3529 ;
  assign n3531 = n3530 ^ n404 ^ 1'b0 ;
  assign n3532 = x245 & ~n3531 ;
  assign n3533 = n3532 ^ n3122 ^ 1'b0 ;
  assign n3534 = n1672 & ~n3533 ;
  assign n3535 = n3030 ^ n2819 ^ 1'b0 ;
  assign n3536 = n3535 ^ n2542 ^ x136 ;
  assign n3537 = n2925 ^ n1130 ^ x12 ;
  assign n3538 = ~n2267 & n3537 ;
  assign n3539 = n3538 ^ n1921 ^ 1'b0 ;
  assign n3540 = n3000 & ~n3539 ;
  assign n3541 = n3536 & n3540 ;
  assign n3542 = ( n1179 & n1473 ) | ( n1179 & n1589 ) | ( n1473 & n1589 ) ;
  assign n3543 = ~n2315 & n3542 ;
  assign n3545 = ( n482 & n657 ) | ( n482 & ~n763 ) | ( n657 & ~n763 ) ;
  assign n3544 = n313 & n2125 ;
  assign n3546 = n3545 ^ n3544 ^ 1'b0 ;
  assign n3547 = n3543 & ~n3546 ;
  assign n3548 = n827 & n3547 ;
  assign n3549 = n3548 ^ n2794 ^ 1'b0 ;
  assign n3550 = ( x199 & ~n367 ) | ( x199 & n2354 ) | ( ~n367 & n2354 ) ;
  assign n3551 = n3550 ^ n2998 ^ n2231 ;
  assign n3552 = x168 & n938 ;
  assign n3553 = n3552 ^ n3029 ^ 1'b0 ;
  assign n3554 = n631 & n3553 ;
  assign n3555 = n432 & n3554 ;
  assign n3556 = n3555 ^ n3337 ^ n921 ;
  assign n3557 = n3556 ^ n2256 ^ 1'b0 ;
  assign n3558 = n3557 ^ n3198 ^ 1'b0 ;
  assign n3559 = ~n3551 & n3558 ;
  assign n3560 = n2692 ^ n1080 ^ 1'b0 ;
  assign n3561 = ~n2745 & n3560 ;
  assign n3562 = ( ~n381 & n1352 ) | ( ~n381 & n2904 ) | ( n1352 & n2904 ) ;
  assign n3563 = ~n873 & n3562 ;
  assign n3564 = n2092 & ~n3563 ;
  assign n3565 = ~n523 & n3564 ;
  assign n3566 = n1672 ^ x253 ^ 1'b0 ;
  assign n3567 = n633 & ~n1433 ;
  assign n3568 = n3567 ^ n693 ^ 1'b0 ;
  assign n3569 = ( x88 & n1589 ) | ( x88 & ~n3568 ) | ( n1589 & ~n3568 ) ;
  assign n3570 = n2481 & n3569 ;
  assign n3571 = ~n3566 & n3570 ;
  assign n3572 = n1280 ^ n864 ^ n303 ;
  assign n3573 = n362 | n3572 ;
  assign n3574 = n2374 ^ n1567 ^ 1'b0 ;
  assign n3575 = n1252 & n3574 ;
  assign n3576 = ( n3208 & n3459 ) | ( n3208 & n3575 ) | ( n3459 & n3575 ) ;
  assign n3577 = n2324 ^ n1612 ^ x157 ;
  assign n3578 = ( ~n1808 & n3576 ) | ( ~n1808 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3579 = n739 | n750 ;
  assign n3580 = n1046 ^ x18 ^ 1'b0 ;
  assign n3582 = ~n1663 & n3249 ;
  assign n3583 = n3582 ^ n1610 ^ 1'b0 ;
  assign n3581 = n1910 & ~n3275 ;
  assign n3584 = n3583 ^ n3581 ^ 1'b0 ;
  assign n3585 = ( n1511 & n1919 ) | ( n1511 & n3283 ) | ( n1919 & n3283 ) ;
  assign n3588 = n1128 | n1501 ;
  assign n3589 = n3588 ^ n1442 ^ 1'b0 ;
  assign n3590 = ~n1125 & n2489 ;
  assign n3591 = n3589 & n3590 ;
  assign n3587 = n1415 ^ n1287 ^ n1108 ;
  assign n3586 = n1845 ^ n1231 ^ 1'b0 ;
  assign n3592 = n3591 ^ n3587 ^ n3586 ;
  assign n3595 = n420 | n996 ;
  assign n3596 = n3595 ^ n1493 ^ 1'b0 ;
  assign n3597 = n890 & n3596 ;
  assign n3598 = n3597 ^ n1585 ^ 1'b0 ;
  assign n3593 = n1839 ^ n1197 ^ 1'b0 ;
  assign n3594 = n2545 & n3593 ;
  assign n3599 = n3598 ^ n3594 ^ n814 ;
  assign n3600 = n1347 | n3599 ;
  assign n3601 = ( ~n1173 & n1347 ) | ( ~n1173 & n3600 ) | ( n1347 & n3600 ) ;
  assign n3602 = n2670 ^ n1415 ^ 1'b0 ;
  assign n3604 = n1646 ^ n1346 ^ 1'b0 ;
  assign n3603 = n1017 & ~n2388 ;
  assign n3605 = n3604 ^ n3603 ^ 1'b0 ;
  assign n3606 = x154 & n481 ;
  assign n3607 = ~n516 & n3606 ;
  assign n3608 = n1448 & ~n3607 ;
  assign n3609 = n3608 ^ n3170 ^ n1517 ;
  assign n3610 = n642 | n1123 ;
  assign n3611 = n266 | n3610 ;
  assign n3612 = n841 & n3611 ;
  assign n3613 = ~x106 & n3612 ;
  assign n3614 = n3613 ^ n2773 ^ 1'b0 ;
  assign n3615 = n3614 ^ n3242 ^ 1'b0 ;
  assign n3616 = ~n2151 & n3615 ;
  assign n3617 = n2695 ^ n1975 ^ n1051 ;
  assign n3618 = n604 & n1166 ;
  assign n3619 = n780 & n3618 ;
  assign n3620 = n3619 ^ n402 ^ 1'b0 ;
  assign n3621 = n2243 & n3620 ;
  assign n3623 = n3249 ^ n393 ^ 1'b0 ;
  assign n3622 = n2789 ^ n1017 ^ n389 ;
  assign n3624 = n3623 ^ n3622 ^ 1'b0 ;
  assign n3625 = n2432 | n3624 ;
  assign n3631 = n934 | n1525 ;
  assign n3632 = n379 & ~n3631 ;
  assign n3626 = n875 ^ x32 ^ 1'b0 ;
  assign n3627 = n3148 & n3626 ;
  assign n3628 = n3172 & n3627 ;
  assign n3629 = ~n3608 & n3628 ;
  assign n3630 = n3629 ^ n2865 ^ 1'b0 ;
  assign n3633 = n3632 ^ n3630 ^ n1571 ;
  assign n3636 = n2113 ^ n1582 ^ 1'b0 ;
  assign n3634 = n703 ^ x205 ^ 1'b0 ;
  assign n3635 = ~n1116 & n3634 ;
  assign n3637 = n3636 ^ n3635 ^ 1'b0 ;
  assign n3638 = n3637 ^ n280 ^ 1'b0 ;
  assign n3639 = ~n3080 & n3638 ;
  assign n3640 = n3404 | n3512 ;
  assign n3647 = ( n652 & ~n995 ) | ( n652 & n1309 ) | ( ~n995 & n1309 ) ;
  assign n3648 = n2049 & n3647 ;
  assign n3649 = n3648 ^ n947 ^ 1'b0 ;
  assign n3650 = n2213 | n3649 ;
  assign n3641 = ( ~n657 & n947 ) | ( ~n657 & n1780 ) | ( n947 & n1780 ) ;
  assign n3642 = n2293 ^ n550 ^ 1'b0 ;
  assign n3643 = n1109 & n3642 ;
  assign n3644 = n3643 ^ n1034 ^ 1'b0 ;
  assign n3645 = n3644 ^ n1222 ^ 1'b0 ;
  assign n3646 = ( n2733 & n3641 ) | ( n2733 & n3645 ) | ( n3641 & n3645 ) ;
  assign n3651 = n3650 ^ n3646 ^ x138 ;
  assign n3652 = n1485 ^ n665 ^ x201 ;
  assign n3653 = ( n421 & n1819 ) | ( n421 & n3652 ) | ( n1819 & n3652 ) ;
  assign n3655 = ( ~n1251 & n1697 ) | ( ~n1251 & n2246 ) | ( n1697 & n2246 ) ;
  assign n3654 = n1031 | n3232 ;
  assign n3656 = n3655 ^ n3654 ^ 1'b0 ;
  assign n3659 = n3218 ^ n1391 ^ n731 ;
  assign n3657 = x173 & ~n1346 ;
  assign n3658 = ~n644 & n3657 ;
  assign n3660 = n3659 ^ n3658 ^ 1'b0 ;
  assign n3661 = n2554 & ~n3660 ;
  assign n3662 = n1537 ^ n654 ^ 1'b0 ;
  assign n3663 = n1280 | n3662 ;
  assign n3664 = n3663 ^ n870 ^ n826 ;
  assign n3665 = n3650 ^ n2930 ^ 1'b0 ;
  assign n3666 = ( n744 & ~n3664 ) | ( n744 & n3665 ) | ( ~n3664 & n3665 ) ;
  assign n3667 = ~n462 & n2966 ;
  assign n3668 = ~n272 & n3667 ;
  assign n3669 = ( ~n1086 & n1520 ) | ( ~n1086 & n3589 ) | ( n1520 & n3589 ) ;
  assign n3670 = n1736 & ~n2482 ;
  assign n3671 = ( n1216 & n3669 ) | ( n1216 & n3670 ) | ( n3669 & n3670 ) ;
  assign n3672 = n3671 ^ n2985 ^ 1'b0 ;
  assign n3673 = n2540 ^ n310 ^ 1'b0 ;
  assign n3674 = n1037 & ~n2582 ;
  assign n3675 = n2467 & n3674 ;
  assign n3676 = n1418 & ~n3675 ;
  assign n3677 = n3459 ^ n1681 ^ n1359 ;
  assign n3678 = ( ~n1854 & n1961 ) | ( ~n1854 & n3677 ) | ( n1961 & n3677 ) ;
  assign n3679 = n3292 ^ n3080 ^ 1'b0 ;
  assign n3680 = ( n616 & ~n3678 ) | ( n616 & n3679 ) | ( ~n3678 & n3679 ) ;
  assign n3681 = n1366 & ~n1870 ;
  assign n3682 = n3681 ^ n724 ^ 1'b0 ;
  assign n3683 = n1331 & ~n2001 ;
  assign n3684 = ( n3542 & ~n3682 ) | ( n3542 & n3683 ) | ( ~n3682 & n3683 ) ;
  assign n3685 = n2029 ^ x79 ^ 1'b0 ;
  assign n3686 = n1848 | n2968 ;
  assign n3687 = n3686 ^ n956 ^ 1'b0 ;
  assign n3688 = n1912 & ~n3687 ;
  assign n3689 = ( n884 & n980 ) | ( n884 & ~n1488 ) | ( n980 & ~n1488 ) ;
  assign n3690 = ( ~x17 & n1799 ) | ( ~x17 & n2606 ) | ( n1799 & n2606 ) ;
  assign n3691 = ~n1205 & n3690 ;
  assign n3692 = n3073 & n3691 ;
  assign n3693 = n2414 & n3692 ;
  assign n3694 = ( n547 & n2213 ) | ( n547 & n3074 ) | ( n2213 & n3074 ) ;
  assign n3695 = n1812 ^ x165 ^ 1'b0 ;
  assign n3696 = x184 & n3695 ;
  assign n3697 = ( x250 & ~n1497 ) | ( x250 & n3696 ) | ( ~n1497 & n3696 ) ;
  assign n3698 = n1011 & ~n1630 ;
  assign n3699 = n3698 ^ n1848 ^ 1'b0 ;
  assign n3700 = n3466 & n3699 ;
  assign n3701 = ~n3697 & n3700 ;
  assign n3702 = n2881 ^ n1501 ^ x195 ;
  assign n3703 = n855 ^ n821 ^ 1'b0 ;
  assign n3704 = ( n703 & n3702 ) | ( n703 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3705 = ~n1496 & n3704 ;
  assign n3706 = n3705 ^ n1004 ^ 1'b0 ;
  assign n3710 = n857 | n1671 ;
  assign n3711 = n393 | n3710 ;
  assign n3707 = n3261 ^ n3074 ^ n1550 ;
  assign n3708 = n1095 | n1477 ;
  assign n3709 = n3707 & ~n3708 ;
  assign n3712 = n3711 ^ n3709 ^ n1250 ;
  assign n3713 = n3712 ^ n1010 ^ 1'b0 ;
  assign n3714 = n2738 ^ n1824 ^ 1'b0 ;
  assign n3715 = n2554 & ~n3714 ;
  assign n3716 = ~n1505 & n2686 ;
  assign n3717 = ( x133 & n1289 ) | ( x133 & n2876 ) | ( n1289 & n2876 ) ;
  assign n3718 = ( n943 & n1631 ) | ( n943 & ~n2881 ) | ( n1631 & ~n2881 ) ;
  assign n3719 = n3718 ^ n872 ^ x95 ;
  assign n3720 = ( n1827 & n2547 ) | ( n1827 & ~n3719 ) | ( n2547 & ~n3719 ) ;
  assign n3721 = n3717 & ~n3720 ;
  assign n3722 = n3269 ^ n779 ^ 1'b0 ;
  assign n3723 = n881 & n2234 ;
  assign n3724 = n706 & n3723 ;
  assign n3725 = n1958 & n3724 ;
  assign n3726 = n2795 ^ n870 ^ 1'b0 ;
  assign n3727 = n1254 & ~n3726 ;
  assign n3728 = n2051 ^ n2035 ^ n1303 ;
  assign n3729 = n3728 ^ n476 ^ 1'b0 ;
  assign n3730 = ~n457 & n3729 ;
  assign n3731 = n534 & n3730 ;
  assign n3732 = ~n3727 & n3731 ;
  assign n3733 = x154 & ~n3732 ;
  assign n3734 = ~n2824 & n3733 ;
  assign n3735 = n3734 ^ n3027 ^ n2887 ;
  assign n3736 = n3735 ^ n2908 ^ n534 ;
  assign n3737 = n1132 & n3736 ;
  assign n3738 = n910 & ~n3305 ;
  assign n3739 = ( x112 & n2508 ) | ( x112 & ~n2571 ) | ( n2508 & ~n2571 ) ;
  assign n3740 = n2057 ^ n1957 ^ x186 ;
  assign n3741 = n2126 | n3303 ;
  assign n3742 = n889 | n3741 ;
  assign n3743 = n3740 & n3742 ;
  assign n3744 = n3743 ^ n1077 ^ 1'b0 ;
  assign n3745 = ( x217 & n461 ) | ( x217 & n3099 ) | ( n461 & n3099 ) ;
  assign n3746 = n3745 ^ n999 ^ 1'b0 ;
  assign n3747 = n443 | n3746 ;
  assign n3748 = n3747 ^ n365 ^ 1'b0 ;
  assign n3749 = n2406 ^ n1541 ^ 1'b0 ;
  assign n3750 = n1057 & n3749 ;
  assign n3751 = n3750 ^ n2929 ^ 1'b0 ;
  assign n3754 = ( ~n310 & n1723 ) | ( ~n310 & n3115 ) | ( n1723 & n3115 ) ;
  assign n3752 = n2881 ^ n341 ^ 1'b0 ;
  assign n3753 = n3752 ^ n590 ^ n553 ;
  assign n3755 = n3754 ^ n3753 ^ 1'b0 ;
  assign n3756 = ~n3296 & n3755 ;
  assign n3757 = n3756 ^ n3645 ^ n2345 ;
  assign n3761 = ( n1377 & n2573 ) | ( n1377 & ~n3071 ) | ( n2573 & ~n3071 ) ;
  assign n3758 = ~n702 & n1559 ;
  assign n3759 = n3758 ^ n1687 ^ 1'b0 ;
  assign n3760 = ~n919 & n3759 ;
  assign n3762 = n3761 ^ n3760 ^ x134 ;
  assign n3763 = ( n673 & n3082 ) | ( n673 & n3762 ) | ( n3082 & n3762 ) ;
  assign n3764 = n3388 ^ n2525 ^ n2145 ;
  assign n3765 = n3764 ^ n1780 ^ n1296 ;
  assign n3766 = n1136 ^ x158 ^ 1'b0 ;
  assign n3767 = n3766 ^ n3254 ^ 1'b0 ;
  assign n3768 = n2529 ^ n684 ^ 1'b0 ;
  assign n3769 = n3653 & n3768 ;
  assign n3770 = n534 | n969 ;
  assign n3771 = n1201 & n3770 ;
  assign n3772 = n3359 ^ n2474 ^ 1'b0 ;
  assign n3773 = n2887 ^ n626 ^ 1'b0 ;
  assign n3774 = x229 & n3773 ;
  assign n3775 = ( x12 & x156 ) | ( x12 & n471 ) | ( x156 & n471 ) ;
  assign n3776 = n1314 | n3775 ;
  assign n3782 = x205 ^ x147 ^ 1'b0 ;
  assign n3777 = n1393 ^ n378 ^ 1'b0 ;
  assign n3778 = n2258 | n3777 ;
  assign n3779 = ~x238 & n3566 ;
  assign n3780 = n3111 | n3779 ;
  assign n3781 = n3778 & ~n3780 ;
  assign n3783 = n3782 ^ n3781 ^ n3675 ;
  assign n3784 = ~n711 & n2700 ;
  assign n3785 = n3750 ^ n946 ^ n314 ;
  assign n3786 = ( n3587 & n3636 ) | ( n3587 & n3785 ) | ( n3636 & n3785 ) ;
  assign n3787 = n432 & ~n3226 ;
  assign n3788 = n678 & n3787 ;
  assign n3789 = n2374 | n3788 ;
  assign n3790 = x217 | n3789 ;
  assign n3791 = n3790 ^ n668 ^ 1'b0 ;
  assign n3792 = n3791 ^ n2739 ^ 1'b0 ;
  assign n3793 = n541 & n633 ;
  assign n3794 = n3793 ^ n2001 ^ 1'b0 ;
  assign n3795 = ~n1420 & n2116 ;
  assign n3796 = n961 | n3795 ;
  assign n3797 = ( n1251 & ~n3794 ) | ( n1251 & n3796 ) | ( ~n3794 & n3796 ) ;
  assign n3798 = n1986 ^ n962 ^ 1'b0 ;
  assign n3799 = n763 ^ x216 ^ 1'b0 ;
  assign n3800 = n1431 | n3799 ;
  assign n3801 = n1437 & ~n3800 ;
  assign n3802 = ( x81 & n3339 ) | ( x81 & n3801 ) | ( n3339 & n3801 ) ;
  assign n3803 = ( ~x99 & n663 ) | ( ~x99 & n1454 ) | ( n663 & n1454 ) ;
  assign n3804 = ~n841 & n3803 ;
  assign n3805 = n3804 ^ n1639 ^ n388 ;
  assign n3806 = n1928 ^ n963 ^ 1'b0 ;
  assign n3807 = ~n2231 & n2604 ;
  assign n3808 = n3807 ^ n3549 ^ 1'b0 ;
  assign n3809 = n3806 | n3808 ;
  assign n3810 = n1392 & n3761 ;
  assign n3811 = ( n1568 & ~n2227 ) | ( n1568 & n3810 ) | ( ~n2227 & n3810 ) ;
  assign n3822 = n3097 ^ n3071 ^ 1'b0 ;
  assign n3823 = ~n3488 & n3822 ;
  assign n3813 = n2087 ^ n1545 ^ 1'b0 ;
  assign n3812 = n434 & n1026 ;
  assign n3814 = n3813 ^ n3812 ^ 1'b0 ;
  assign n3815 = n3080 | n3459 ;
  assign n3816 = n3815 ^ n1701 ^ 1'b0 ;
  assign n3817 = n3816 ^ n1352 ^ x4 ;
  assign n3818 = ( n294 & n2790 ) | ( n294 & ~n2832 ) | ( n2790 & ~n2832 ) ;
  assign n3819 = n3413 & n3818 ;
  assign n3820 = ~n3817 & n3819 ;
  assign n3821 = n3814 & n3820 ;
  assign n3824 = n3823 ^ n3821 ^ n2832 ;
  assign n3825 = ~n1733 & n3067 ;
  assign n3826 = ~n829 & n3825 ;
  assign n3827 = n2161 ^ n2043 ^ 1'b0 ;
  assign n3828 = ~n3826 & n3827 ;
  assign n3829 = n3828 ^ n1331 ^ x119 ;
  assign n3830 = n1743 ^ n388 ^ 1'b0 ;
  assign n3831 = ( n1430 & ~n1827 ) | ( n1430 & n3830 ) | ( ~n1827 & n3830 ) ;
  assign n3832 = ~n3065 & n3831 ;
  assign n3833 = n800 & ~n1370 ;
  assign n3834 = n3833 ^ n1517 ^ 1'b0 ;
  assign n3835 = n1078 & n3218 ;
  assign n3837 = ( x242 & n1710 ) | ( x242 & ~n2569 ) | ( n1710 & ~n2569 ) ;
  assign n3838 = n910 & n3837 ;
  assign n3839 = n3838 ^ n2074 ^ 1'b0 ;
  assign n3840 = n3839 ^ n3309 ^ 1'b0 ;
  assign n3836 = x51 & n3073 ;
  assign n3841 = n3840 ^ n3836 ^ 1'b0 ;
  assign n3842 = n3754 ^ n597 ^ 1'b0 ;
  assign n3843 = n1211 | n3842 ;
  assign n3844 = n3843 ^ n2126 ^ n541 ;
  assign n3845 = n926 | n1845 ;
  assign n3846 = ( ~n2247 & n2262 ) | ( ~n2247 & n3845 ) | ( n2262 & n3845 ) ;
  assign n3847 = ( n3577 & ~n3844 ) | ( n3577 & n3846 ) | ( ~n3844 & n3846 ) ;
  assign n3848 = x237 & n644 ;
  assign n3849 = n3848 ^ x59 ^ 1'b0 ;
  assign n3850 = n903 & ~n3849 ;
  assign n3851 = n2113 & n3850 ;
  assign n3852 = ~n521 & n3117 ;
  assign n3853 = n3852 ^ x154 ^ 1'b0 ;
  assign n3854 = n3851 | n3853 ;
  assign n3855 = n3196 | n3854 ;
  assign n3856 = ( ~n1392 & n2833 ) | ( ~n1392 & n3855 ) | ( n2833 & n3855 ) ;
  assign n3857 = n3856 ^ n3742 ^ n3696 ;
  assign n3858 = ( n1619 & n3510 ) | ( n1619 & n3857 ) | ( n3510 & n3857 ) ;
  assign n3859 = n3858 ^ n3162 ^ n943 ;
  assign n3860 = x210 | n3305 ;
  assign n3861 = n891 ^ x40 ^ 1'b0 ;
  assign n3862 = ( n989 & ~n3860 ) | ( n989 & n3861 ) | ( ~n3860 & n3861 ) ;
  assign n3863 = ( n1598 & n2676 ) | ( n1598 & n3862 ) | ( n2676 & n3862 ) ;
  assign n3866 = n1939 ^ n1385 ^ 1'b0 ;
  assign n3867 = n1662 & n3866 ;
  assign n3864 = n867 | n2692 ;
  assign n3865 = n2205 & ~n3864 ;
  assign n3868 = n3867 ^ n3865 ^ n1700 ;
  assign n3869 = n795 ^ n358 ^ 1'b0 ;
  assign n3870 = n1445 & ~n3869 ;
  assign n3871 = n1908 & n3870 ;
  assign n3872 = n259 & n3871 ;
  assign n3873 = ( n1571 & n1649 ) | ( n1571 & n2065 ) | ( n1649 & n2065 ) ;
  assign n3874 = ( x249 & n1692 ) | ( x249 & ~n3873 ) | ( n1692 & ~n3873 ) ;
  assign n3875 = n675 ^ x46 ^ 1'b0 ;
  assign n3876 = ~n3874 & n3875 ;
  assign n3877 = n2436 ^ n1385 ^ 1'b0 ;
  assign n3878 = n1810 | n3877 ;
  assign n3879 = n3641 | n3878 ;
  assign n3880 = n3879 ^ n566 ^ 1'b0 ;
  assign n3881 = n1658 ^ n1374 ^ n340 ;
  assign n3882 = n2766 ^ n2617 ^ 1'b0 ;
  assign n3883 = n3881 | n3882 ;
  assign n3884 = n3839 ^ n2094 ^ 1'b0 ;
  assign n3885 = n3883 | n3884 ;
  assign n3887 = ( n276 & n1793 ) | ( n276 & ~n3849 ) | ( n1793 & ~n3849 ) ;
  assign n3886 = x186 & n619 ;
  assign n3888 = n3887 ^ n3886 ^ 1'b0 ;
  assign n3889 = n1451 ^ n1444 ^ n832 ;
  assign n3890 = n2758 & n2881 ;
  assign n3891 = ~n3889 & n3890 ;
  assign n3892 = ( n737 & n3888 ) | ( n737 & n3891 ) | ( n3888 & n3891 ) ;
  assign n3893 = ~n814 & n1044 ;
  assign n3894 = n730 & n3893 ;
  assign n3895 = x136 & ~n3894 ;
  assign n3896 = n3641 & n3895 ;
  assign n3899 = ~n474 & n516 ;
  assign n3900 = ~n3678 & n3899 ;
  assign n3901 = n1321 | n3900 ;
  assign n3897 = n3803 ^ n2143 ^ x93 ;
  assign n3898 = n3897 ^ n1331 ^ n613 ;
  assign n3902 = n3901 ^ n3898 ^ n741 ;
  assign n3903 = ( n2561 & n3896 ) | ( n2561 & n3902 ) | ( n3896 & n3902 ) ;
  assign n3904 = x158 & ~n1878 ;
  assign n3905 = ~n1690 & n3904 ;
  assign n3906 = n2522 ^ n1661 ^ 1'b0 ;
  assign n3907 = n2168 & n3906 ;
  assign n3908 = n2731 | n3219 ;
  assign n3909 = n2151 & ~n3908 ;
  assign n3910 = n1269 & ~n1604 ;
  assign n3911 = ( n700 & ~n3633 ) | ( n700 & n3910 ) | ( ~n3633 & n3910 ) ;
  assign n3912 = n1220 & ~n2913 ;
  assign n3913 = n297 & n3912 ;
  assign n3914 = n2357 | n3913 ;
  assign n3915 = n3914 ^ n3334 ^ 1'b0 ;
  assign n3916 = n1328 & ~n1361 ;
  assign n3917 = n3916 ^ n840 ^ 1'b0 ;
  assign n3918 = n3917 ^ n2553 ^ 1'b0 ;
  assign n3919 = n3918 ^ n3542 ^ n883 ;
  assign n3920 = n3919 ^ n3705 ^ n1662 ;
  assign n3921 = ( ~n1105 & n3915 ) | ( ~n1105 & n3920 ) | ( n3915 & n3920 ) ;
  assign n3922 = n3677 ^ n1822 ^ 1'b0 ;
  assign n3923 = ~n3162 & n3922 ;
  assign n3928 = n1503 ^ n609 ^ 1'b0 ;
  assign n3924 = ( x26 & n780 ) | ( x26 & ~n2138 ) | ( n780 & ~n2138 ) ;
  assign n3925 = n796 & ~n1174 ;
  assign n3926 = n3925 ^ n1442 ^ 1'b0 ;
  assign n3927 = ( x45 & n3924 ) | ( x45 & n3926 ) | ( n3924 & n3926 ) ;
  assign n3929 = n3928 ^ n3927 ^ 1'b0 ;
  assign n3930 = n3923 & ~n3929 ;
  assign n3933 = n2685 ^ n2050 ^ n1771 ;
  assign n3931 = ( x178 & ~n1989 ) | ( x178 & n2049 ) | ( ~n1989 & n2049 ) ;
  assign n3932 = ~n3438 & n3931 ;
  assign n3934 = n3933 ^ n3932 ^ 1'b0 ;
  assign n3935 = n3930 & n3934 ;
  assign n3936 = n1977 ^ n570 ^ 1'b0 ;
  assign n3937 = ~n2405 & n3936 ;
  assign n3938 = ~n1502 & n3937 ;
  assign n3939 = n3938 ^ n585 ^ 1'b0 ;
  assign n3940 = n3557 & n3939 ;
  assign n3941 = n2394 ^ n1559 ^ n1430 ;
  assign n3942 = n3941 ^ x58 ^ 1'b0 ;
  assign n3943 = n3129 & ~n3942 ;
  assign n3944 = x24 & n1703 ;
  assign n3945 = n3944 ^ n1304 ^ 1'b0 ;
  assign n3946 = ~n2234 & n3945 ;
  assign n3947 = ( n919 & n2995 ) | ( n919 & n3701 ) | ( n2995 & n3701 ) ;
  assign n3949 = n2904 ^ n1472 ^ x237 ;
  assign n3950 = n3949 ^ n2247 ^ 1'b0 ;
  assign n3951 = n842 & ~n3950 ;
  assign n3948 = n736 & n2125 ;
  assign n3952 = n3951 ^ n3948 ^ 1'b0 ;
  assign n3955 = ( x209 & n1337 ) | ( x209 & n1405 ) | ( n1337 & n1405 ) ;
  assign n3953 = n1535 ^ n373 ^ 1'b0 ;
  assign n3954 = n3953 ^ n1367 ^ 1'b0 ;
  assign n3956 = n3955 ^ n3954 ^ 1'b0 ;
  assign n3957 = ~n3465 & n3956 ;
  assign n3958 = ( ~n2427 & n3952 ) | ( ~n2427 & n3957 ) | ( n3952 & n3957 ) ;
  assign n3959 = n1552 & n3310 ;
  assign n3960 = n3959 ^ n1034 ^ 1'b0 ;
  assign n3961 = n3960 ^ n3716 ^ 1'b0 ;
  assign n3962 = n3867 & ~n3961 ;
  assign n3963 = n2282 ^ n294 ^ 1'b0 ;
  assign n3964 = n3693 & n3963 ;
  assign n3965 = n1197 & ~n2655 ;
  assign n3966 = n2749 & n3863 ;
  assign n3967 = n3031 ^ n2121 ^ n2087 ;
  assign n3968 = ( x73 & ~x161 ) | ( x73 & n3967 ) | ( ~x161 & n3967 ) ;
  assign n3969 = n358 & n3839 ;
  assign n3970 = n3969 ^ x46 ^ 1'b0 ;
  assign n3971 = ~n1162 & n1902 ;
  assign n3972 = n3971 ^ n1384 ^ 1'b0 ;
  assign n3973 = ~n3970 & n3972 ;
  assign n3974 = ~n840 & n2689 ;
  assign n3975 = n3687 ^ n1380 ^ 1'b0 ;
  assign n3976 = n1473 ^ n362 ^ 1'b0 ;
  assign n3977 = n3975 & n3976 ;
  assign n3978 = x154 | n2677 ;
  assign n3979 = n3977 | n3978 ;
  assign n3980 = n1375 & n3115 ;
  assign n3981 = n835 | n1022 ;
  assign n3982 = n3981 ^ x41 ^ 1'b0 ;
  assign n3983 = ( n782 & n1868 ) | ( n782 & ~n1943 ) | ( n1868 & ~n1943 ) ;
  assign n3984 = n3691 & n3983 ;
  assign n3985 = n3984 ^ n1685 ^ 1'b0 ;
  assign n3986 = n3982 | n3985 ;
  assign n3987 = n695 & n1427 ;
  assign n3988 = n1108 | n1745 ;
  assign n3989 = n3988 ^ n1739 ^ 1'b0 ;
  assign n3990 = n3639 ^ n2481 ^ 1'b0 ;
  assign n3991 = n481 & n3990 ;
  assign n3992 = ( n1064 & ~n2363 ) | ( n1064 & n2501 ) | ( ~n2363 & n2501 ) ;
  assign n3993 = n3992 ^ n1671 ^ 1'b0 ;
  assign n3994 = n627 & n3993 ;
  assign n3995 = ( n676 & n1278 ) | ( n676 & ~n2474 ) | ( n1278 & ~n2474 ) ;
  assign n3996 = n491 & n3433 ;
  assign n3997 = ~n1074 & n3309 ;
  assign n3998 = ( n3070 & n3996 ) | ( n3070 & ~n3997 ) | ( n3996 & ~n3997 ) ;
  assign n3999 = n2194 & n3998 ;
  assign n4000 = n1261 | n3824 ;
  assign n4001 = n3989 | n4000 ;
  assign n4002 = n2723 ^ n1209 ^ 1'b0 ;
  assign n4003 = ( ~n2585 & n2746 ) | ( ~n2585 & n2841 ) | ( n2746 & n2841 ) ;
  assign n4004 = n4003 ^ n2623 ^ 1'b0 ;
  assign n4006 = ( ~x6 & x200 ) | ( ~x6 & n2305 ) | ( x200 & n2305 ) ;
  assign n4007 = n4006 ^ n2230 ^ n1557 ;
  assign n4005 = n2379 ^ n731 ^ 1'b0 ;
  assign n4008 = n4007 ^ n4005 ^ n1738 ;
  assign n4009 = n2573 & ~n2697 ;
  assign n4010 = n1423 | n1838 ;
  assign n4011 = n4010 ^ n3289 ^ n388 ;
  assign n4012 = ~n771 & n4011 ;
  assign n4013 = n968 & n4012 ;
  assign n4014 = ~x241 & n3550 ;
  assign n4015 = n2657 ^ n2076 ^ n957 ;
  assign n4016 = ( n3964 & n4014 ) | ( n3964 & ~n4015 ) | ( n4014 & ~n4015 ) ;
  assign n4017 = n1906 ^ n1300 ^ n947 ;
  assign n4018 = n1145 ^ n564 ^ 1'b0 ;
  assign n4019 = n1188 & ~n4018 ;
  assign n4020 = n1664 & n4019 ;
  assign n4021 = n2178 & n4020 ;
  assign n4022 = n4021 ^ n3101 ^ 1'b0 ;
  assign n4023 = ~n617 & n4022 ;
  assign n4024 = n4017 & n4023 ;
  assign n4025 = ~n3549 & n4024 ;
  assign n4026 = ( ~n905 & n1287 ) | ( ~n905 & n4025 ) | ( n1287 & n4025 ) ;
  assign n4027 = n3913 ^ n486 ^ 1'b0 ;
  assign n4028 = n2824 ^ n2100 ^ 1'b0 ;
  assign n4029 = x80 & ~n2061 ;
  assign n4030 = n1083 & ~n4029 ;
  assign n4031 = n1908 ^ n835 ^ 1'b0 ;
  assign n4032 = x106 | n4031 ;
  assign n4033 = ~n1405 & n2049 ;
  assign n4034 = n4033 ^ n3724 ^ 1'b0 ;
  assign n4039 = n317 & n3525 ;
  assign n4040 = n4039 ^ n1409 ^ 1'b0 ;
  assign n4035 = n2613 ^ n616 ^ 1'b0 ;
  assign n4036 = n1233 | n4035 ;
  assign n4037 = x5 | n4036 ;
  assign n4038 = n865 | n4037 ;
  assign n4041 = n4040 ^ n4038 ^ 1'b0 ;
  assign n4042 = n4034 & n4041 ;
  assign n4043 = n1024 | n3285 ;
  assign n4044 = n773 ^ n609 ^ x187 ;
  assign n4045 = n4044 ^ n1877 ^ 1'b0 ;
  assign n4046 = ( n1105 & ~n3389 ) | ( n1105 & n4045 ) | ( ~n3389 & n4045 ) ;
  assign n4047 = n2558 ^ n766 ^ 1'b0 ;
  assign n4048 = n634 ^ n367 ^ 1'b0 ;
  assign n4049 = n3281 ^ n2868 ^ n1191 ;
  assign n4050 = n4048 & n4049 ;
  assign n4051 = n4047 & n4050 ;
  assign n4052 = n3105 ^ n1472 ^ n497 ;
  assign n4053 = ( n2653 & ~n4051 ) | ( n2653 & n4052 ) | ( ~n4051 & n4052 ) ;
  assign n4054 = n1133 ^ n929 ^ n520 ;
  assign n4055 = ( x243 & n605 ) | ( x243 & ~n2336 ) | ( n605 & ~n2336 ) ;
  assign n4056 = n4054 & ~n4055 ;
  assign n4057 = n2148 ^ n783 ^ 1'b0 ;
  assign n4060 = ( ~x78 & n1545 ) | ( ~x78 & n1630 ) | ( n1545 & n1630 ) ;
  assign n4058 = n2785 ^ n1414 ^ 1'b0 ;
  assign n4059 = n1309 | n4058 ;
  assign n4061 = n4060 ^ n4059 ^ n3360 ;
  assign n4062 = ( ~x238 & n4057 ) | ( ~x238 & n4061 ) | ( n4057 & n4061 ) ;
  assign n4064 = n2724 ^ n2071 ^ n363 ;
  assign n4065 = n4064 ^ n755 ^ 1'b0 ;
  assign n4066 = n4065 ^ n1740 ^ n1650 ;
  assign n4063 = ~n1821 & n2740 ;
  assign n4067 = n4066 ^ n4063 ^ 1'b0 ;
  assign n4068 = n4067 ^ n2995 ^ n2867 ;
  assign n4069 = ( n2359 & ~n4062 ) | ( n2359 & n4068 ) | ( ~n4062 & n4068 ) ;
  assign n4070 = ( ~n476 & n827 ) | ( ~n476 & n943 ) | ( n827 & n943 ) ;
  assign n4071 = n4070 ^ n1501 ^ 1'b0 ;
  assign n4072 = ~x248 & n4071 ;
  assign n4073 = ~n3191 & n4072 ;
  assign n4077 = ( x47 & n374 ) | ( x47 & ~n2528 ) | ( n374 & ~n2528 ) ;
  assign n4075 = ~n826 & n2580 ;
  assign n4074 = n759 & ~n2325 ;
  assign n4076 = n4075 ^ n4074 ^ 1'b0 ;
  assign n4078 = n4077 ^ n4076 ^ 1'b0 ;
  assign n4079 = n4073 & n4078 ;
  assign n4080 = n3600 ^ n2421 ^ n988 ;
  assign n4081 = n1954 & n4080 ;
  assign n4082 = n1235 ^ n272 ^ 1'b0 ;
  assign n4083 = x218 & n4082 ;
  assign n4084 = n704 & ~n1963 ;
  assign n4085 = ~n4083 & n4084 ;
  assign n4086 = n4085 ^ n4047 ^ n1122 ;
  assign n4087 = ~n1861 & n3460 ;
  assign n4088 = n2854 ^ n1775 ^ 1'b0 ;
  assign n4089 = ( n1421 & ~n3209 ) | ( n1421 & n4088 ) | ( ~n3209 & n4088 ) ;
  assign n4090 = n1623 ^ n1009 ^ 1'b0 ;
  assign n4091 = n4090 ^ x144 ^ 1'b0 ;
  assign n4092 = n2595 ^ n2447 ^ 1'b0 ;
  assign n4093 = x252 & n4092 ;
  assign n4094 = ~n2534 & n4093 ;
  assign n4095 = n4091 & n4094 ;
  assign n4099 = n1179 & n1267 ;
  assign n4098 = n666 & ~n3759 ;
  assign n4096 = n602 | n730 ;
  assign n4097 = n2933 | n4096 ;
  assign n4100 = n4099 ^ n4098 ^ n4097 ;
  assign n4101 = n1134 & ~n3643 ;
  assign n4102 = ( ~n637 & n1525 ) | ( ~n637 & n4101 ) | ( n1525 & n4101 ) ;
  assign n4103 = n1098 | n3435 ;
  assign n4104 = n4103 ^ n901 ^ 1'b0 ;
  assign n4105 = n315 | n4104 ;
  assign n4106 = n4102 & n4105 ;
  assign n4107 = n2135 ^ n871 ^ 1'b0 ;
  assign n4108 = n4107 ^ n2419 ^ n1158 ;
  assign n4109 = n2398 ^ n1020 ^ n990 ;
  assign n4110 = n4109 ^ n3071 ^ 1'b0 ;
  assign n4111 = n3704 ^ n1353 ^ 1'b0 ;
  assign n4112 = n4110 & n4111 ;
  assign n4113 = n1308 & n3553 ;
  assign n4114 = n4112 & n4113 ;
  assign n4115 = n2329 ^ n370 ^ 1'b0 ;
  assign n4116 = n2442 | n4115 ;
  assign n4117 = n1645 & ~n2737 ;
  assign n4118 = n4117 ^ n1750 ^ n765 ;
  assign n4120 = n1991 | n3779 ;
  assign n4121 = n4120 ^ n2482 ^ 1'b0 ;
  assign n4119 = ( ~x173 & n2390 ) | ( ~x173 & n2423 ) | ( n2390 & n2423 ) ;
  assign n4122 = n4121 ^ n4119 ^ 1'b0 ;
  assign n4123 = n4118 | n4122 ;
  assign n4124 = n3874 ^ n1782 ^ 1'b0 ;
  assign n4125 = n1164 & n4124 ;
  assign n4126 = n2343 ^ n1655 ^ n966 ;
  assign n4127 = n4126 ^ n2229 ^ 1'b0 ;
  assign n4128 = n3495 & n4127 ;
  assign n4129 = n4128 ^ x129 ^ 1'b0 ;
  assign n4130 = n1563 ^ n1211 ^ 1'b0 ;
  assign n4131 = n1427 & n4130 ;
  assign n4132 = ~n1846 & n4131 ;
  assign n4133 = n595 & ~n4132 ;
  assign n4134 = n402 & n4133 ;
  assign n4135 = ~n2453 & n3310 ;
  assign n4136 = ~n1533 & n4135 ;
  assign n4137 = n4136 ^ n1372 ^ n629 ;
  assign n4138 = n3232 ^ n2607 ^ n868 ;
  assign n4141 = n590 | n2333 ;
  assign n4142 = n1054 ^ n562 ^ n447 ;
  assign n4143 = ( ~n480 & n2310 ) | ( ~n480 & n4142 ) | ( n2310 & n4142 ) ;
  assign n4144 = n4143 ^ n3641 ^ 1'b0 ;
  assign n4145 = n4144 ^ n3834 ^ 1'b0 ;
  assign n4146 = n4141 | n4145 ;
  assign n4139 = ( n256 & n3843 ) | ( n256 & ~n3906 ) | ( n3843 & ~n3906 ) ;
  assign n4140 = ~n2628 & n4139 ;
  assign n4147 = n4146 ^ n4140 ^ 1'b0 ;
  assign n4149 = n782 & ~n2488 ;
  assign n4150 = ~n2040 & n4149 ;
  assign n4148 = n2773 ^ n2282 ^ 1'b0 ;
  assign n4151 = n4150 ^ n4148 ^ x175 ;
  assign n4152 = n2646 ^ n2564 ^ 1'b0 ;
  assign n4153 = n2437 ^ n1292 ^ 1'b0 ;
  assign n4154 = ( n2103 & n4152 ) | ( n2103 & ~n4153 ) | ( n4152 & ~n4153 ) ;
  assign n4155 = ~n1979 & n3155 ;
  assign n4156 = n1585 & ~n2205 ;
  assign n4157 = ( ~n3858 & n4155 ) | ( ~n3858 & n4156 ) | ( n4155 & n4156 ) ;
  assign n4158 = n1814 & ~n2791 ;
  assign n4161 = n2315 ^ n2084 ^ 1'b0 ;
  assign n4162 = n1493 & n4161 ;
  assign n4163 = n771 ^ n695 ^ n558 ;
  assign n4164 = n4163 ^ x37 ^ 1'b0 ;
  assign n4165 = n4162 & n4164 ;
  assign n4159 = ~n1016 & n4127 ;
  assign n4160 = n4159 ^ n2050 ^ 1'b0 ;
  assign n4166 = n4165 ^ n4160 ^ n2972 ;
  assign n4167 = ( x191 & ~n1078 ) | ( x191 & n2021 ) | ( ~n1078 & n2021 ) ;
  assign n4168 = n4167 ^ n853 ^ 1'b0 ;
  assign n4169 = n3393 ^ n841 ^ n468 ;
  assign n4170 = ~n2021 & n2569 ;
  assign n4171 = n4170 ^ n1447 ^ 1'b0 ;
  assign n4172 = n977 | n4171 ;
  assign n4173 = n4169 & ~n4172 ;
  assign n4174 = n1236 ^ n1098 ^ 1'b0 ;
  assign n4175 = n1197 & n4174 ;
  assign n4176 = n2505 & n3337 ;
  assign n4177 = ~n4175 & n4176 ;
  assign n4178 = n4177 ^ n2558 ^ n444 ;
  assign n4179 = n4178 ^ n3974 ^ n3488 ;
  assign n4180 = n4173 | n4179 ;
  assign n4181 = n2308 ^ n2167 ^ 1'b0 ;
  assign n4182 = ~n2123 & n4181 ;
  assign n4183 = n4182 ^ n3673 ^ n2704 ;
  assign n4184 = ~n497 & n682 ;
  assign n4185 = n4184 ^ n1599 ^ 1'b0 ;
  assign n4186 = n4185 ^ n2796 ^ n1758 ;
  assign n4187 = ( ~n2410 & n2825 ) | ( ~n2410 & n3352 ) | ( n2825 & n3352 ) ;
  assign n4188 = ~n4186 & n4187 ;
  assign n4189 = n2305 & n4188 ;
  assign n4190 = x216 ^ x207 ^ x82 ;
  assign n4191 = n1578 ^ n1409 ^ 1'b0 ;
  assign n4192 = ~n1857 & n4191 ;
  assign n4193 = n3888 & n4192 ;
  assign n4194 = n1741 & n4193 ;
  assign n4195 = n3644 ^ n276 ^ 1'b0 ;
  assign n4196 = n1048 | n4195 ;
  assign n4197 = n759 & n3596 ;
  assign n4198 = ~n2472 & n4197 ;
  assign n4199 = n1674 & ~n4198 ;
  assign n4200 = n2724 & n4199 ;
  assign n4201 = n4196 & n4200 ;
  assign n4202 = n3716 ^ n880 ^ 1'b0 ;
  assign n4203 = n1632 ^ n1102 ^ 1'b0 ;
  assign n4204 = ~n1464 & n4203 ;
  assign n4205 = x141 & ~n274 ;
  assign n4206 = ~n2073 & n4205 ;
  assign n4207 = n4206 ^ n652 ^ 1'b0 ;
  assign n4208 = n4204 & ~n4207 ;
  assign n4209 = n4208 ^ n1690 ^ n1258 ;
  assign n4210 = x237 & n4209 ;
  assign n4211 = ~n4139 & n4210 ;
  assign n4212 = ~n1512 & n1964 ;
  assign n4216 = n940 ^ x170 ^ 1'b0 ;
  assign n4217 = ~n469 & n4216 ;
  assign n4213 = n656 & n1692 ;
  assign n4214 = n2333 & n4213 ;
  assign n4215 = x10 & ~n4214 ;
  assign n4218 = n4217 ^ n4215 ^ n1874 ;
  assign n4223 = n2562 ^ n2236 ^ 1'b0 ;
  assign n4222 = n477 & ~n2071 ;
  assign n4224 = n4223 ^ n4222 ^ 1'b0 ;
  assign n4225 = n3037 ^ n268 ^ 1'b0 ;
  assign n4226 = n4224 & ~n4225 ;
  assign n4219 = n526 ^ x214 ^ 1'b0 ;
  assign n4220 = n4219 ^ n3514 ^ n3031 ;
  assign n4221 = ~n2878 & n4220 ;
  assign n4227 = n4226 ^ n4221 ^ 1'b0 ;
  assign n4228 = ~n1592 & n1948 ;
  assign n4229 = ~n1084 & n4228 ;
  assign n4230 = n790 & n3372 ;
  assign n4231 = n4230 ^ n4066 ^ n1513 ;
  assign n4232 = ( n1813 & n4229 ) | ( n1813 & ~n4231 ) | ( n4229 & ~n4231 ) ;
  assign n4233 = n4232 ^ n526 ^ 1'b0 ;
  assign n4234 = ~n1857 & n4233 ;
  assign n4235 = ~n3268 & n4234 ;
  assign n4236 = n1229 & ~n4013 ;
  assign n4237 = ~n374 & n4236 ;
  assign n4238 = ( x2 & n3225 ) | ( x2 & n3759 ) | ( n3225 & n3759 ) ;
  assign n4239 = n767 ^ n564 ^ 1'b0 ;
  assign n4240 = n4239 ^ n3450 ^ n1819 ;
  assign n4241 = n4240 ^ n3120 ^ 1'b0 ;
  assign n4242 = n2130 ^ n1249 ^ 1'b0 ;
  assign n4243 = ( n982 & n1739 ) | ( n982 & ~n2201 ) | ( n1739 & ~n2201 ) ;
  assign n4244 = ~n1346 & n4243 ;
  assign n4245 = x52 & n3203 ;
  assign n4246 = ~n1782 & n4245 ;
  assign n4247 = ( n3200 & n4029 ) | ( n3200 & ~n4246 ) | ( n4029 & ~n4246 ) ;
  assign n4248 = n4247 ^ n2268 ^ 1'b0 ;
  assign n4249 = ( x151 & n1304 ) | ( x151 & n2663 ) | ( n1304 & n2663 ) ;
  assign n4250 = ( x16 & ~n2019 ) | ( x16 & n3472 ) | ( ~n2019 & n3472 ) ;
  assign n4251 = ( n2631 & ~n2918 ) | ( n2631 & n4250 ) | ( ~n2918 & n4250 ) ;
  assign n4252 = ~n548 & n4251 ;
  assign n4253 = ~n4249 & n4252 ;
  assign n4256 = n3281 ^ n1113 ^ n841 ;
  assign n4255 = n1225 & n2158 ;
  assign n4254 = n2641 ^ n1535 ^ 1'b0 ;
  assign n4257 = n4256 ^ n4255 ^ n4254 ;
  assign n4259 = n3557 ^ n3243 ^ 1'b0 ;
  assign n4258 = n3609 ^ n350 ^ 1'b0 ;
  assign n4260 = n4259 ^ n4258 ^ n1053 ;
  assign n4263 = n1061 ^ n871 ^ 1'b0 ;
  assign n4264 = x87 & ~n4263 ;
  assign n4262 = n944 & n2724 ;
  assign n4265 = n4264 ^ n4262 ^ 1'b0 ;
  assign n4261 = n898 ^ n734 ^ n290 ;
  assign n4266 = n4265 ^ n4261 ^ n4211 ;
  assign n4267 = ( n704 & ~n2372 ) | ( n704 & n3410 ) | ( ~n2372 & n3410 ) ;
  assign n4268 = ( n598 & ~n1010 ) | ( n598 & n4267 ) | ( ~n1010 & n4267 ) ;
  assign n4269 = n4090 | n4268 ;
  assign n4270 = n779 & ~n4269 ;
  assign n4271 = ( ~x181 & n346 ) | ( ~x181 & n1902 ) | ( n346 & n1902 ) ;
  assign n4272 = ~n1627 & n4271 ;
  assign n4273 = ~n1501 & n4272 ;
  assign n4274 = ~n2274 & n4273 ;
  assign n4275 = n4274 ^ n3160 ^ 1'b0 ;
  assign n4276 = n2693 & ~n4275 ;
  assign n4277 = x123 ^ x7 ^ 1'b0 ;
  assign n4278 = n4276 & n4277 ;
  assign n4279 = ( n709 & n1845 ) | ( n709 & n3168 ) | ( n1845 & n3168 ) ;
  assign n4280 = n2578 & ~n4279 ;
  assign n4281 = n4280 ^ n4185 ^ 1'b0 ;
  assign n4282 = ( x152 & n3353 ) | ( x152 & ~n4281 ) | ( n3353 & ~n4281 ) ;
  assign n4283 = n2191 & n4282 ;
  assign n4284 = n1876 ^ n1273 ^ 1'b0 ;
  assign n4285 = x157 & n3563 ;
  assign n4286 = ( ~n1199 & n1701 ) | ( ~n1199 & n2685 ) | ( n1701 & n2685 ) ;
  assign n4287 = ~n295 & n4286 ;
  assign n4288 = ( ~n3541 & n4285 ) | ( ~n3541 & n4287 ) | ( n4285 & n4287 ) ;
  assign n4289 = ( n853 & n960 ) | ( n853 & ~n2093 ) | ( n960 & ~n2093 ) ;
  assign n4290 = n2851 ^ n2490 ^ 1'b0 ;
  assign n4291 = n4289 & n4290 ;
  assign n4292 = ( n4284 & ~n4288 ) | ( n4284 & n4291 ) | ( ~n4288 & n4291 ) ;
  assign n4293 = n3210 ^ n1511 ^ 1'b0 ;
  assign n4294 = ~n2351 & n4293 ;
  assign n4297 = ~n713 & n1287 ;
  assign n4298 = n4297 ^ n1123 ^ 1'b0 ;
  assign n4295 = n374 & ~n1247 ;
  assign n4296 = ~n4217 & n4295 ;
  assign n4299 = n4298 ^ n4296 ^ 1'b0 ;
  assign n4300 = n2032 & ~n4299 ;
  assign n4301 = n2365 ^ n1919 ^ 1'b0 ;
  assign n4302 = ( x170 & x248 ) | ( x170 & ~n4301 ) | ( x248 & ~n4301 ) ;
  assign n4303 = n4302 ^ n3187 ^ 1'b0 ;
  assign n4304 = n2274 & ~n4303 ;
  assign n4310 = n1037 ^ n936 ^ n893 ;
  assign n4311 = ~n3530 & n4310 ;
  assign n4312 = n4311 ^ x60 ^ 1'b0 ;
  assign n4313 = n4312 ^ n1425 ^ 1'b0 ;
  assign n4305 = n3513 ^ n3073 ^ 1'b0 ;
  assign n4306 = n1883 | n4305 ;
  assign n4307 = n4306 ^ n2434 ^ 1'b0 ;
  assign n4308 = n4307 ^ n3830 ^ n739 ;
  assign n4309 = ( ~n2701 & n2982 ) | ( ~n2701 & n4308 ) | ( n2982 & n4308 ) ;
  assign n4314 = n4313 ^ n4309 ^ n2623 ;
  assign n4315 = ( n933 & n1766 ) | ( n933 & ~n2009 ) | ( n1766 & ~n2009 ) ;
  assign n4316 = n3781 ^ n1727 ^ n1252 ;
  assign n4317 = n4315 | n4316 ;
  assign n4318 = n4226 | n4317 ;
  assign n4319 = ( x48 & n1729 ) | ( x48 & n3488 ) | ( n1729 & n3488 ) ;
  assign n4320 = n4040 & ~n4319 ;
  assign n4321 = n3663 & n4320 ;
  assign n4322 = ( ~n907 & n919 ) | ( ~n907 & n2896 ) | ( n919 & n2896 ) ;
  assign n4323 = n4322 ^ n3656 ^ 1'b0 ;
  assign n4324 = x58 & ~n4323 ;
  assign n4325 = n4321 & n4324 ;
  assign n4327 = n700 | n3543 ;
  assign n4326 = x198 & ~n2142 ;
  assign n4328 = n4327 ^ n4326 ^ 1'b0 ;
  assign n4329 = n3782 ^ n1006 ^ 1'b0 ;
  assign n4330 = n1154 ^ n666 ^ 1'b0 ;
  assign n4331 = n466 & ~n4330 ;
  assign n4332 = ( ~n3353 & n4329 ) | ( ~n3353 & n4331 ) | ( n4329 & n4331 ) ;
  assign n4333 = n4328 | n4332 ;
  assign n4334 = n4333 ^ n400 ^ 1'b0 ;
  assign n4335 = n2950 & ~n3766 ;
  assign n4336 = n343 & n668 ;
  assign n4337 = n887 & n4336 ;
  assign n4338 = ~n1800 & n4337 ;
  assign n4339 = n619 & n2407 ;
  assign n4340 = ~x2 & n4339 ;
  assign n4341 = n4340 ^ n3508 ^ n1068 ;
  assign n4342 = n2365 ^ n830 ^ 1'b0 ;
  assign n4343 = ( n3317 & n4341 ) | ( n3317 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4344 = n4338 | n4343 ;
  assign n4345 = n4335 & ~n4344 ;
  assign n4346 = n1864 & n2892 ;
  assign n4347 = n309 & ~n2215 ;
  assign n4348 = ~n1585 & n4347 ;
  assign n4349 = ( n2163 & n4081 ) | ( n2163 & ~n4348 ) | ( n4081 & ~n4348 ) ;
  assign n4350 = n3559 ^ n2956 ^ n1279 ;
  assign n4351 = n3281 ^ n331 ^ 1'b0 ;
  assign n4352 = n3569 & n4351 ;
  assign n4353 = n4352 ^ n3632 ^ 1'b0 ;
  assign n4354 = n898 ^ x254 ^ 1'b0 ;
  assign n4355 = x63 & n4354 ;
  assign n4356 = n4355 ^ n446 ^ 1'b0 ;
  assign n4357 = ~n841 & n2630 ;
  assign n4358 = n1853 | n2903 ;
  assign n4359 = ( n1405 & n4357 ) | ( n1405 & ~n4358 ) | ( n4357 & ~n4358 ) ;
  assign n4360 = n608 ^ n471 ^ x82 ;
  assign n4363 = ( x175 & n1064 ) | ( x175 & n1545 ) | ( n1064 & n1545 ) ;
  assign n4361 = n2886 ^ n2853 ^ 1'b0 ;
  assign n4362 = ~n1501 & n4361 ;
  assign n4364 = n4363 ^ n4362 ^ 1'b0 ;
  assign n4365 = n4364 ^ n616 ^ 1'b0 ;
  assign n4366 = n1574 & ~n4365 ;
  assign n4368 = n367 & n1853 ;
  assign n4369 = n2041 ^ n656 ^ x10 ;
  assign n4370 = n277 & ~n733 ;
  assign n4371 = n4369 & n4370 ;
  assign n4372 = n4368 & ~n4371 ;
  assign n4373 = n4372 ^ n1800 ^ 1'b0 ;
  assign n4367 = n835 | n2673 ;
  assign n4374 = n4373 ^ n4367 ^ 1'b0 ;
  assign n4378 = ( ~n363 & n1506 ) | ( ~n363 & n2293 ) | ( n1506 & n2293 ) ;
  assign n4375 = ( ~n340 & n1468 ) | ( ~n340 & n2114 ) | ( n1468 & n2114 ) ;
  assign n4376 = n633 | n657 ;
  assign n4377 = n4375 & n4376 ;
  assign n4379 = n4378 ^ n4377 ^ 1'b0 ;
  assign n4380 = n2490 & n3785 ;
  assign n4381 = n1502 & n4380 ;
  assign n4387 = n318 | n1977 ;
  assign n4388 = n4387 ^ n3279 ^ 1'b0 ;
  assign n4382 = n2398 ^ n1422 ^ 1'b0 ;
  assign n4383 = ( x158 & ~n1380 ) | ( x158 & n4382 ) | ( ~n1380 & n4382 ) ;
  assign n4384 = x156 | n4383 ;
  assign n4385 = n4384 ^ n3233 ^ 1'b0 ;
  assign n4386 = n1864 | n4385 ;
  assign n4389 = n4388 ^ n4386 ^ x56 ;
  assign n4390 = ~n1474 & n3482 ;
  assign n4391 = ( n2021 & ~n3914 ) | ( n2021 & n4390 ) | ( ~n3914 & n4390 ) ;
  assign n4393 = n1128 | n3374 ;
  assign n4392 = ~n995 & n1018 ;
  assign n4394 = n4393 ^ n4392 ^ 1'b0 ;
  assign n4395 = n623 | n1923 ;
  assign n4396 = x3 | n4395 ;
  assign n4397 = n4396 ^ n1752 ^ 1'b0 ;
  assign n4398 = n1446 | n4397 ;
  assign n4400 = n1222 | n2145 ;
  assign n4401 = n4400 ^ n3992 ^ 1'b0 ;
  assign n4399 = n393 & ~n2255 ;
  assign n4402 = n4401 ^ n4399 ^ 1'b0 ;
  assign n4403 = n4402 ^ n1422 ^ 1'b0 ;
  assign n4404 = n4398 | n4403 ;
  assign n4405 = n3165 ^ n1732 ^ n722 ;
  assign n4406 = n1843 ^ x74 ^ 1'b0 ;
  assign n4407 = n397 & n4406 ;
  assign n4408 = n4407 ^ n2397 ^ 1'b0 ;
  assign n4409 = n4405 | n4408 ;
  assign n4423 = ( x48 & n1111 ) | ( x48 & ~n1543 ) | ( n1111 & ~n1543 ) ;
  assign n4410 = ( n1045 & n1176 ) | ( n1045 & n1251 ) | ( n1176 & n1251 ) ;
  assign n4411 = n4410 ^ x106 ^ 1'b0 ;
  assign n4412 = n1093 & ~n4411 ;
  assign n4413 = x61 | n1687 ;
  assign n4414 = n3754 ^ n2696 ^ n2626 ;
  assign n4415 = ~n1511 & n4414 ;
  assign n4416 = ~n343 & n4415 ;
  assign n4417 = n2340 ^ n1563 ^ n1497 ;
  assign n4418 = ~n4416 & n4417 ;
  assign n4419 = n4418 ^ n2402 ^ 1'b0 ;
  assign n4420 = n4413 & ~n4419 ;
  assign n4421 = n1357 & n4420 ;
  assign n4422 = n4412 & ~n4421 ;
  assign n4424 = n4423 ^ n4422 ^ 1'b0 ;
  assign n4425 = ( n332 & n637 ) | ( n332 & ~n3049 ) | ( n637 & ~n3049 ) ;
  assign n4426 = x71 & x208 ;
  assign n4427 = n4426 ^ n999 ^ 1'b0 ;
  assign n4428 = n1691 ^ x240 ^ 1'b0 ;
  assign n4429 = ~n284 & n4428 ;
  assign n4430 = n4429 ^ n1236 ^ 1'b0 ;
  assign n4431 = n4427 | n4430 ;
  assign n4432 = n4431 ^ n2428 ^ 1'b0 ;
  assign n4433 = ~n416 & n3510 ;
  assign n4434 = ( n2737 & ~n3780 ) | ( n2737 & n4126 ) | ( ~n3780 & n4126 ) ;
  assign n4435 = n2386 ^ n2140 ^ 1'b0 ;
  assign n4436 = n3182 & n3801 ;
  assign n4437 = n3457 ^ n2340 ^ n1331 ;
  assign n4438 = ( n1231 & n2287 ) | ( n1231 & n4437 ) | ( n2287 & n4437 ) ;
  assign n4439 = n335 & n4438 ;
  assign n4440 = ~n540 & n1864 ;
  assign n4441 = x82 ^ x31 ^ 1'b0 ;
  assign n4442 = ~n2982 & n4441 ;
  assign n4443 = x171 & n4053 ;
  assign n4444 = n2365 & ~n3928 ;
  assign n4445 = n4444 ^ n4011 ^ 1'b0 ;
  assign n4450 = n4044 ^ n2702 ^ n2107 ;
  assign n4446 = n808 | n4214 ;
  assign n4447 = n1330 ^ n1233 ^ 1'b0 ;
  assign n4448 = n2421 & ~n4447 ;
  assign n4449 = n4446 & n4448 ;
  assign n4451 = n4450 ^ n4449 ^ 1'b0 ;
  assign n4452 = n405 & ~n4451 ;
  assign n4453 = ( n1264 & n3126 ) | ( n1264 & ~n4452 ) | ( n3126 & ~n4452 ) ;
  assign n4454 = ( ~n1580 & n2982 ) | ( ~n1580 & n3037 ) | ( n2982 & n3037 ) ;
  assign n4455 = ~n570 & n1963 ;
  assign n4458 = n1564 ^ n1483 ^ 1'b0 ;
  assign n4459 = ~n532 & n4458 ;
  assign n4456 = n2773 & n2921 ;
  assign n4457 = n3046 & n4456 ;
  assign n4460 = n4459 ^ n4457 ^ 1'b0 ;
  assign n4464 = n1384 & n2132 ;
  assign n4465 = ~n1064 & n2306 ;
  assign n4466 = ( ~n1708 & n4464 ) | ( ~n1708 & n4465 ) | ( n4464 & n4465 ) ;
  assign n4461 = n1465 ^ x176 ^ x10 ;
  assign n4462 = n4461 ^ n2108 ^ n880 ;
  assign n4463 = n4462 ^ n960 ^ x158 ;
  assign n4467 = n4466 ^ n4463 ^ n3907 ;
  assign n4468 = n604 & n2531 ;
  assign n4469 = n4468 ^ n544 ^ 1'b0 ;
  assign n4470 = ( x65 & n820 ) | ( x65 & n2613 ) | ( n820 & n2613 ) ;
  assign n4471 = n4470 ^ n490 ^ 1'b0 ;
  assign n4472 = ( ~n4308 & n4469 ) | ( ~n4308 & n4471 ) | ( n4469 & n4471 ) ;
  assign n4473 = n1349 ^ n523 ^ 1'b0 ;
  assign n4474 = n4473 ^ n3952 ^ n637 ;
  assign n4475 = n1601 & n2326 ;
  assign n4476 = n1097 & n4475 ;
  assign n4480 = n3336 ^ n2112 ^ 1'b0 ;
  assign n4481 = ( ~x207 & n707 ) | ( ~x207 & n4480 ) | ( n707 & n4480 ) ;
  assign n4477 = n486 & n1108 ;
  assign n4478 = n1357 & n4477 ;
  assign n4479 = n272 | n4478 ;
  assign n4482 = n4481 ^ n4479 ^ n2782 ;
  assign n4483 = n3004 ^ n1105 ^ 1'b0 ;
  assign n4484 = ~n1045 & n4483 ;
  assign n4485 = n2475 ^ n1714 ^ 1'b0 ;
  assign n4486 = n1264 & n4485 ;
  assign n4487 = n428 ^ x15 ^ 1'b0 ;
  assign n4488 = n1521 & n4487 ;
  assign n4489 = ~n2461 & n4488 ;
  assign n4490 = ~n4486 & n4489 ;
  assign n4491 = ( n1197 & n1771 ) | ( n1197 & n1801 ) | ( n1771 & n1801 ) ;
  assign n4492 = n2395 & n4491 ;
  assign n4493 = n2460 & ~n4427 ;
  assign n4494 = n4493 ^ n1136 ^ 1'b0 ;
  assign n4500 = n867 | n1305 ;
  assign n4501 = n885 | n4500 ;
  assign n4502 = n4501 ^ n3750 ^ n294 ;
  assign n4503 = n4502 ^ n1397 ^ n796 ;
  assign n4504 = n2835 & n4375 ;
  assign n4505 = ( n1889 & ~n4503 ) | ( n1889 & n4504 ) | ( ~n4503 & n4504 ) ;
  assign n4496 = n2904 ^ n1206 ^ 1'b0 ;
  assign n4497 = ~n1158 & n4496 ;
  assign n4498 = ( ~n374 & n966 ) | ( ~n374 & n4497 ) | ( n966 & n4497 ) ;
  assign n4495 = x104 & n4139 ;
  assign n4499 = n4498 ^ n4495 ^ 1'b0 ;
  assign n4506 = n4505 ^ n4499 ^ n4488 ;
  assign n4507 = n2737 ^ n580 ^ 1'b0 ;
  assign n4508 = n4256 & n4507 ;
  assign n4509 = ~n4286 & n4508 ;
  assign n4510 = n4296 ^ n4061 ^ n1135 ;
  assign n4511 = n2395 & n2699 ;
  assign n4512 = n410 & n4511 ;
  assign n4513 = n575 | n4484 ;
  assign n4515 = n367 & n2168 ;
  assign n4516 = n4515 ^ n855 ^ 1'b0 ;
  assign n4514 = n2363 | n3365 ;
  assign n4517 = n4516 ^ n4514 ^ n3438 ;
  assign n4518 = ( ~n1184 & n1687 ) | ( ~n1184 & n2213 ) | ( n1687 & n2213 ) ;
  assign n4519 = n3266 | n4518 ;
  assign n4520 = n444 | n4519 ;
  assign n4521 = n321 & ~n4520 ;
  assign n4522 = n421 | n3975 ;
  assign n4523 = n2510 ^ n1721 ^ 1'b0 ;
  assign n4524 = x146 & ~n4523 ;
  assign n4525 = n4522 & n4524 ;
  assign n4526 = n4525 ^ n1580 ^ 1'b0 ;
  assign n4527 = ( n1074 & ~n2559 ) | ( n1074 & n3322 ) | ( ~n2559 & n3322 ) ;
  assign n4528 = n1444 & ~n3892 ;
  assign n4529 = ( n479 & n795 ) | ( n479 & ~n3193 ) | ( n795 & ~n3193 ) ;
  assign n4530 = ~n518 & n1588 ;
  assign n4531 = ( n645 & n769 ) | ( n645 & ~n4530 ) | ( n769 & ~n4530 ) ;
  assign n4532 = ( x242 & ~n4529 ) | ( x242 & n4531 ) | ( ~n4529 & n4531 ) ;
  assign n4533 = ~n547 & n600 ;
  assign n4534 = n1921 & n4533 ;
  assign n4535 = n4534 ^ n3260 ^ 1'b0 ;
  assign n4538 = ~n1274 & n1333 ;
  assign n4539 = n3928 | n4538 ;
  assign n4540 = n1140 & ~n4539 ;
  assign n4541 = n262 | n305 ;
  assign n4542 = n4540 & ~n4541 ;
  assign n4536 = n4351 ^ n4327 ^ n3928 ;
  assign n4537 = ( n643 & n2089 ) | ( n643 & n4536 ) | ( n2089 & n4536 ) ;
  assign n4543 = n4542 ^ n4537 ^ n4139 ;
  assign n4544 = ~n1923 & n2608 ;
  assign n4545 = n2390 & ~n2689 ;
  assign n4546 = ~n4544 & n4545 ;
  assign n4547 = ~n2153 & n3372 ;
  assign n4548 = ~n990 & n2604 ;
  assign n4549 = ( n483 & n1832 ) | ( n483 & ~n4548 ) | ( n1832 & ~n4548 ) ;
  assign n4550 = ( n2699 & ~n4547 ) | ( n2699 & n4549 ) | ( ~n4547 & n4549 ) ;
  assign n4551 = n4550 ^ n1639 ^ x45 ;
  assign n4556 = n1487 ^ n1142 ^ 1'b0 ;
  assign n4555 = n2422 ^ n1239 ^ 1'b0 ;
  assign n4557 = n4556 ^ n4555 ^ n1934 ;
  assign n4552 = n3627 ^ n2906 ^ n280 ;
  assign n4553 = n4552 ^ n2333 ^ n1123 ;
  assign n4554 = ( n2191 & n3043 ) | ( n2191 & ~n4553 ) | ( n3043 & ~n4553 ) ;
  assign n4558 = n4557 ^ n4554 ^ n4476 ;
  assign n4559 = n713 & ~n3467 ;
  assign n4560 = ( x250 & ~n2024 ) | ( x250 & n2451 ) | ( ~n2024 & n2451 ) ;
  assign n4561 = n1408 | n1594 ;
  assign n4562 = n3163 | n4561 ;
  assign n4563 = n650 & n2250 ;
  assign n4564 = n4563 ^ n4019 ^ 1'b0 ;
  assign n4565 = ( x19 & n413 ) | ( x19 & ~n4564 ) | ( n413 & ~n4564 ) ;
  assign n4566 = ~n738 & n4565 ;
  assign n4567 = n4566 ^ n1035 ^ n964 ;
  assign n4568 = n3829 & ~n4567 ;
  assign n4569 = n3562 ^ n2684 ^ 1'b0 ;
  assign n4570 = ~n2241 & n4569 ;
  assign n4571 = ( n1688 & ~n2518 ) | ( n1688 & n2778 ) | ( ~n2518 & n2778 ) ;
  assign n4572 = n4571 ^ n3323 ^ 1'b0 ;
  assign n4573 = n4570 & n4572 ;
  assign n4574 = n4573 ^ n2374 ^ n1586 ;
  assign n4575 = ( ~x22 & n1603 ) | ( ~x22 & n2369 ) | ( n1603 & n2369 ) ;
  assign n4576 = n4313 ^ n2187 ^ 1'b0 ;
  assign n4577 = n2785 & ~n4576 ;
  assign n4578 = n1001 ^ x106 ^ 1'b0 ;
  assign n4579 = x116 & n4578 ;
  assign n4580 = ~n2667 & n4579 ;
  assign n4581 = n1372 & n4580 ;
  assign n4582 = n3358 ^ n923 ^ 1'b0 ;
  assign n4583 = n1867 & ~n4575 ;
  assign n4584 = n1116 | n4583 ;
  assign n4585 = n1290 & ~n4584 ;
  assign n4586 = n2707 | n4585 ;
  assign n4587 = n4586 ^ n4554 ^ 1'b0 ;
  assign n4589 = x127 & ~n2828 ;
  assign n4590 = n1390 ^ n335 ^ 1'b0 ;
  assign n4591 = ( n1130 & n4589 ) | ( n1130 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4588 = n4151 ^ x4 ^ 1'b0 ;
  assign n4592 = n4591 ^ n4588 ^ n2840 ;
  assign n4593 = n1226 & n2785 ;
  assign n4594 = n4593 ^ n1202 ^ n317 ;
  assign n4595 = n4594 ^ n1531 ^ 1'b0 ;
  assign n4596 = n739 ^ n432 ^ 1'b0 ;
  assign n4597 = ( n2408 & ~n4382 ) | ( n2408 & n4596 ) | ( ~n4382 & n4596 ) ;
  assign n4598 = n4597 ^ n595 ^ 1'b0 ;
  assign n4599 = x199 & ~n424 ;
  assign n4600 = n4599 ^ n2004 ^ 1'b0 ;
  assign n4601 = n4600 ^ n3141 ^ n766 ;
  assign n4602 = n744 & n3434 ;
  assign n4603 = n4602 ^ n4394 ^ 1'b0 ;
  assign n4604 = n2208 ^ n1864 ^ 1'b0 ;
  assign n4605 = n4604 ^ n4016 ^ n925 ;
  assign n4606 = ( n1688 & ~n2031 ) | ( n1688 & n3748 ) | ( ~n2031 & n3748 ) ;
  assign n4607 = n2270 ^ n645 ^ n584 ;
  assign n4608 = n2333 ^ n820 ^ 1'b0 ;
  assign n4609 = x102 | n4608 ;
  assign n4610 = n4609 ^ n1562 ^ 1'b0 ;
  assign n4611 = n4607 & n4610 ;
  assign n4612 = ( n2210 & ~n4551 ) | ( n2210 & n4611 ) | ( ~n4551 & n4611 ) ;
  assign n4615 = ~n345 & n2380 ;
  assign n4616 = n1353 & n4615 ;
  assign n4617 = n1438 & n4616 ;
  assign n4613 = ( n370 & ~n1309 ) | ( n370 & n3033 ) | ( ~n1309 & n3033 ) ;
  assign n4614 = ~n3966 & n4613 ;
  assign n4618 = n4617 ^ n4614 ^ 1'b0 ;
  assign n4621 = ( n825 & ~n2151 ) | ( n825 & n2477 ) | ( ~n2151 & n2477 ) ;
  assign n4619 = n2364 ^ n2019 ^ n1285 ;
  assign n4620 = ( n503 & n2283 ) | ( n503 & n4619 ) | ( n2283 & n4619 ) ;
  assign n4622 = n4621 ^ n4620 ^ n2928 ;
  assign n4623 = n579 & ~n4186 ;
  assign n4624 = n4622 & n4623 ;
  assign n4625 = n763 | n4481 ;
  assign n4626 = n3393 & ~n4625 ;
  assign n4627 = ~n1334 & n3566 ;
  assign n4628 = n806 ^ x40 ^ 1'b0 ;
  assign n4629 = n389 & ~n4628 ;
  assign n4630 = n4629 ^ n3157 ^ n2616 ;
  assign n4631 = n3160 & ~n3949 ;
  assign n4632 = ~n1739 & n4631 ;
  assign n4633 = n2594 & ~n4502 ;
  assign n4634 = n4632 & n4633 ;
  assign n4635 = n4390 ^ n330 ^ 1'b0 ;
  assign n4636 = ( ~x24 & n1009 ) | ( ~x24 & n4635 ) | ( n1009 & n4635 ) ;
  assign n4637 = ( n1706 & ~n2273 ) | ( n1706 & n4636 ) | ( ~n2273 & n4636 ) ;
  assign n4638 = n354 & ~n914 ;
  assign n4639 = n1268 ^ n1117 ^ 1'b0 ;
  assign n4640 = n1352 & n4639 ;
  assign n4641 = n4638 & n4640 ;
  assign n4642 = ( n2479 & n4049 ) | ( n2479 & n4641 ) | ( n4049 & n4641 ) ;
  assign n4643 = ~n863 & n4394 ;
  assign n4644 = n4643 ^ n3427 ^ 1'b0 ;
  assign n4645 = n3960 ^ n771 ^ n765 ;
  assign n4646 = ( n1375 & n1526 ) | ( n1375 & n2236 ) | ( n1526 & n2236 ) ;
  assign n4647 = n4646 ^ n2613 ^ 1'b0 ;
  assign n4648 = n2803 & n4647 ;
  assign n4649 = n1736 & n2210 ;
  assign n4650 = n4649 ^ n3485 ^ 1'b0 ;
  assign n4651 = n4650 ^ x72 ^ 1'b0 ;
  assign n4652 = n346 | n4651 ;
  assign n4653 = ( n4645 & n4648 ) | ( n4645 & ~n4652 ) | ( n4648 & ~n4652 ) ;
  assign n4654 = ~n370 & n3145 ;
  assign n4655 = n4654 ^ n907 ^ 1'b0 ;
  assign n4656 = ~n3918 & n4655 ;
  assign n4657 = n3061 & n4656 ;
  assign n4658 = ~n3448 & n4657 ;
  assign n4659 = ( n1077 & ~n1759 ) | ( n1077 & n4658 ) | ( ~n1759 & n4658 ) ;
  assign n4660 = n2939 ^ n877 ^ x42 ;
  assign n4661 = n3921 ^ n2073 ^ 1'b0 ;
  assign n4662 = ~n2987 & n4661 ;
  assign n4672 = n450 ^ x202 ^ x66 ;
  assign n4673 = n4672 ^ n3650 ^ n2510 ;
  assign n4669 = n609 & n1169 ;
  assign n4668 = ~n680 & n4376 ;
  assign n4670 = n4669 ^ n4668 ^ 1'b0 ;
  assign n4671 = n4670 ^ x55 ^ 1'b0 ;
  assign n4674 = n4673 ^ n4671 ^ x151 ;
  assign n4663 = n2501 ^ n1199 ^ 1'b0 ;
  assign n4664 = ~n1148 & n4663 ;
  assign n4665 = n4664 ^ n547 ^ n482 ;
  assign n4666 = n4665 ^ n1725 ^ n261 ;
  assign n4667 = n4182 & ~n4666 ;
  assign n4675 = n4674 ^ n4667 ^ 1'b0 ;
  assign n4676 = x112 & ~n3363 ;
  assign n4677 = n4676 ^ n836 ^ 1'b0 ;
  assign n4678 = n4677 ^ x239 ^ 1'b0 ;
  assign n4679 = n1926 ^ n1422 ^ n447 ;
  assign n4680 = n4679 ^ n2825 ^ n1137 ;
  assign n4681 = ~n3273 & n4119 ;
  assign n4682 = n4681 ^ n2170 ^ 1'b0 ;
  assign n4683 = n2461 ^ n1070 ^ 1'b0 ;
  assign n4684 = n1315 & n4683 ;
  assign n4685 = n4684 ^ n482 ^ 1'b0 ;
  assign n4686 = ~n1725 & n4685 ;
  assign n4687 = n4686 ^ n1488 ^ 1'b0 ;
  assign n4688 = n1034 & ~n4687 ;
  assign n4689 = n3722 ^ n2260 ^ 1'b0 ;
  assign n4690 = ~x3 & x248 ;
  assign n4691 = ( ~x142 & x245 ) | ( ~x142 & n1159 ) | ( x245 & n1159 ) ;
  assign n4692 = ( n1593 & n2066 ) | ( n1593 & ~n3594 ) | ( n2066 & ~n3594 ) ;
  assign n4693 = n1776 | n4692 ;
  assign n4694 = n4691 & ~n4693 ;
  assign n4695 = n1187 & ~n3280 ;
  assign n4696 = n2711 & ~n4085 ;
  assign n4697 = n4696 ^ n3664 ^ 1'b0 ;
  assign n4698 = n1644 | n4697 ;
  assign n4699 = n452 ^ n348 ^ 1'b0 ;
  assign n4700 = n4382 | n4699 ;
  assign n4701 = n4700 ^ n1464 ^ 1'b0 ;
  assign n4702 = n515 & n980 ;
  assign n4703 = ~x65 & n4702 ;
  assign n4704 = ~n4382 & n4703 ;
  assign n4705 = ~n2414 & n4704 ;
  assign n4706 = ( ~n1047 & n1279 ) | ( ~n1047 & n4066 ) | ( n1279 & n4066 ) ;
  assign n4710 = n615 & ~n2195 ;
  assign n4711 = n3926 ^ n1251 ^ n1184 ;
  assign n4712 = n4711 ^ n1052 ^ 1'b0 ;
  assign n4713 = ( n3813 & n4710 ) | ( n3813 & ~n4712 ) | ( n4710 & ~n4712 ) ;
  assign n4707 = x19 & ~x41 ;
  assign n4708 = n2560 | n4707 ;
  assign n4709 = n2972 | n4708 ;
  assign n4714 = n4713 ^ n4709 ^ 1'b0 ;
  assign n4715 = n3814 ^ n2849 ^ n580 ;
  assign n4716 = n2868 & n4289 ;
  assign n4717 = n2665 & n4716 ;
  assign n4718 = n4717 ^ n2758 ^ 1'b0 ;
  assign n4719 = ( n2685 & n4440 ) | ( n2685 & n4718 ) | ( n4440 & n4718 ) ;
  assign n4720 = n2945 ^ n1411 ^ n938 ;
  assign n4721 = n1910 ^ x191 ^ x42 ;
  assign n4722 = n4720 & n4721 ;
  assign n4723 = n2333 & n4722 ;
  assign n4724 = n4723 ^ n4313 ^ n923 ;
  assign n4725 = n4724 ^ n632 ^ 1'b0 ;
  assign n4726 = n3679 ^ n2308 ^ 1'b0 ;
  assign n4727 = n859 | n2998 ;
  assign n4728 = n4727 ^ n4208 ^ n2000 ;
  assign n4729 = ~n1342 & n4728 ;
  assign n4730 = n4729 ^ x16 ^ 1'b0 ;
  assign n4731 = n1040 & ~n1567 ;
  assign n4732 = ~n1834 & n4731 ;
  assign n4733 = n4732 ^ n1882 ^ 1'b0 ;
  assign n4734 = n2531 ^ n923 ^ n587 ;
  assign n4735 = n4734 ^ n1029 ^ 1'b0 ;
  assign n4736 = n540 | n818 ;
  assign n4737 = n4736 ^ n1123 ^ 1'b0 ;
  assign n4738 = n4737 ^ n1732 ^ 1'b0 ;
  assign n4739 = n4738 ^ x130 ^ 1'b0 ;
  assign n4740 = ( n3502 & n3957 ) | ( n3502 & n4739 ) | ( n3957 & n4739 ) ;
  assign n4741 = n321 | n4480 ;
  assign n4742 = x172 & n4741 ;
  assign n4743 = n1538 & n4742 ;
  assign n4744 = n4743 ^ n2850 ^ 1'b0 ;
  assign n4745 = n4744 ^ n2818 ^ n2665 ;
  assign n4752 = n3029 ^ n822 ^ 1'b0 ;
  assign n4753 = n343 & ~n4752 ;
  assign n4748 = n3545 ^ n2210 ^ 1'b0 ;
  assign n4746 = n1474 | n3322 ;
  assign n4747 = n435 | n4746 ;
  assign n4749 = n4748 ^ n4747 ^ n4731 ;
  assign n4750 = n3855 | n4749 ;
  assign n4751 = n1409 & ~n4750 ;
  assign n4754 = n4753 ^ n4751 ^ 1'b0 ;
  assign n4755 = n1054 & n1436 ;
  assign n4756 = n4755 ^ n1031 ^ 1'b0 ;
  assign n4757 = n2978 & n4756 ;
  assign n4758 = n4757 ^ n2124 ^ n2029 ;
  assign n4759 = n1529 ^ n1513 ^ n468 ;
  assign n4760 = ( n3115 & n3449 ) | ( n3115 & ~n4759 ) | ( n3449 & ~n4759 ) ;
  assign n4761 = n1491 ^ n1243 ^ n510 ;
  assign n4762 = n4761 ^ n3395 ^ 1'b0 ;
  assign n4763 = n3205 & ~n3690 ;
  assign n4764 = n2011 ^ x207 ^ 1'b0 ;
  assign n4765 = n4763 & n4764 ;
  assign n4766 = n2415 ^ n2240 ^ 1'b0 ;
  assign n4767 = ( n2413 & ~n3154 ) | ( n2413 & n3814 ) | ( ~n3154 & n3814 ) ;
  assign n4768 = n4766 | n4767 ;
  assign n4769 = n2238 | n4768 ;
  assign n4770 = ( n2985 & ~n3190 ) | ( n2985 & n4601 ) | ( ~n3190 & n4601 ) ;
  assign n4771 = n1420 ^ n648 ^ n461 ;
  assign n4773 = n1554 ^ x82 ^ 1'b0 ;
  assign n4774 = n4773 ^ n3776 ^ n3026 ;
  assign n4772 = n4620 ^ n1881 ^ n502 ;
  assign n4775 = n4774 ^ n4772 ^ n1567 ;
  assign n4776 = n4175 ^ x159 ^ 1'b0 ;
  assign n4777 = n4776 ^ n343 ^ 1'b0 ;
  assign n4778 = n4388 & n4777 ;
  assign n4779 = n2956 & n4778 ;
  assign n4780 = n2068 & ~n3598 ;
  assign n4781 = ~n3116 & n4780 ;
  assign n4782 = ( ~x230 & n2055 ) | ( ~x230 & n4165 ) | ( n2055 & n4165 ) ;
  assign n4783 = n4782 ^ n4041 ^ n301 ;
  assign n4784 = ~n2985 & n3759 ;
  assign n4785 = ~n4110 & n4784 ;
  assign n4786 = ( n1821 & ~n4066 ) | ( n1821 & n4785 ) | ( ~n4066 & n4785 ) ;
  assign n4787 = n4783 | n4786 ;
  assign n4788 = n4113 ^ n3245 ^ n2084 ;
  assign n4789 = n4175 ^ n3839 ^ 1'b0 ;
  assign n4790 = n1351 & ~n3366 ;
  assign n4792 = n1233 ^ x205 ^ 1'b0 ;
  assign n4793 = n1477 | n4792 ;
  assign n4791 = x66 | n3176 ;
  assign n4794 = n4793 ^ n4791 ^ 1'b0 ;
  assign n4795 = n1851 | n2329 ;
  assign n4796 = n4794 & ~n4795 ;
  assign n4797 = n4796 ^ n3186 ^ n1270 ;
  assign n4798 = n807 ^ n644 ^ 1'b0 ;
  assign n4799 = n2878 | n4798 ;
  assign n4800 = n4799 ^ n1855 ^ n1776 ;
  assign n4801 = n4800 ^ n3121 ^ n1208 ;
  assign n4802 = n1844 ^ n1035 ^ 1'b0 ;
  assign n4803 = x21 & n4802 ;
  assign n4804 = n3168 & n4803 ;
  assign n4805 = n1579 & n4804 ;
  assign n4806 = n2367 ^ n2013 ^ x18 ;
  assign n4807 = ( n384 & n4805 ) | ( n384 & n4806 ) | ( n4805 & n4806 ) ;
  assign n4808 = n4807 ^ n3062 ^ n1083 ;
  assign n4809 = n4808 ^ n526 ^ 1'b0 ;
  assign n4810 = n1296 ^ n766 ^ n613 ;
  assign n4811 = ( n1730 & n2781 ) | ( n1730 & ~n4810 ) | ( n2781 & ~n4810 ) ;
  assign n4817 = n2504 & n2749 ;
  assign n4818 = n4398 & n4817 ;
  assign n4812 = n1206 ^ n1057 ^ x216 ;
  assign n4813 = n4812 ^ n1568 ^ n901 ;
  assign n4814 = n4813 ^ n1816 ^ 1'b0 ;
  assign n4815 = n865 & n4814 ;
  assign n4816 = n4815 ^ n1353 ^ 1'b0 ;
  assign n4819 = n4818 ^ n4816 ^ n2068 ;
  assign n4821 = ~n2470 & n3046 ;
  assign n4820 = n2296 ^ n2249 ^ 1'b0 ;
  assign n4822 = n4821 ^ n4820 ^ n4242 ;
  assign n4823 = n3524 ^ n1579 ^ n1246 ;
  assign n4824 = ~n361 & n4777 ;
  assign n4825 = n1582 & n4824 ;
  assign n4826 = ( n2796 & n3285 ) | ( n2796 & ~n4292 ) | ( n3285 & ~n4292 ) ;
  assign n4827 = n4826 ^ n2613 ^ 1'b0 ;
  assign n4828 = n4827 ^ n4167 ^ 1'b0 ;
  assign n4830 = ( n695 & n2116 ) | ( n695 & n2707 ) | ( n2116 & n2707 ) ;
  assign n4831 = n1074 | n4830 ;
  assign n4832 = n4831 ^ n3495 ^ 1'b0 ;
  assign n4833 = n4832 ^ n348 ^ 1'b0 ;
  assign n4829 = x170 & ~n1870 ;
  assign n4834 = n4833 ^ n4829 ^ 1'b0 ;
  assign n4835 = ( ~n885 & n3711 ) | ( ~n885 & n4163 ) | ( n3711 & n4163 ) ;
  assign n4836 = n3223 & n4835 ;
  assign n4837 = n4836 ^ n4769 ^ 1'b0 ;
  assign n4838 = n1438 & ~n3563 ;
  assign n4839 = n4838 ^ n698 ^ n376 ;
  assign n4840 = ( n483 & n2985 ) | ( n483 & ~n4839 ) | ( n2985 & ~n4839 ) ;
  assign n4841 = ( ~n534 & n2333 ) | ( ~n534 & n3411 ) | ( n2333 & n3411 ) ;
  assign n4842 = n2832 ^ n399 ^ 1'b0 ;
  assign n4843 = n4842 ^ n1087 ^ 1'b0 ;
  assign n4844 = n2226 | n4843 ;
  assign n4845 = n4844 ^ n3041 ^ n510 ;
  assign n4846 = ~n4841 & n4845 ;
  assign n4847 = n4840 & n4846 ;
  assign n4849 = n845 ^ x84 ^ 1'b0 ;
  assign n4850 = n4849 ^ n1083 ^ n929 ;
  assign n4848 = n3049 ^ n880 ^ 1'b0 ;
  assign n4851 = n4850 ^ n4848 ^ n4703 ;
  assign n4852 = n4851 ^ n3509 ^ n2138 ;
  assign n4855 = n830 ^ n671 ^ 1'b0 ;
  assign n4856 = x211 & ~n4855 ;
  assign n4853 = n1437 | n1742 ;
  assign n4854 = n673 & ~n4853 ;
  assign n4857 = n4856 ^ n4854 ^ n1878 ;
  assign n4858 = n1543 | n4857 ;
  assign n4859 = ( n3177 & ~n4852 ) | ( n3177 & n4858 ) | ( ~n4852 & n4858 ) ;
  assign n4860 = n2475 ^ n1345 ^ n381 ;
  assign n4861 = n2036 & ~n4315 ;
  assign n4862 = ~n2355 & n4861 ;
  assign n4863 = n4862 ^ n2498 ^ n1372 ;
  assign n4864 = n1933 ^ n1782 ^ n1264 ;
  assign n4865 = n4864 ^ n2241 ^ 1'b0 ;
  assign n4866 = n1576 ^ n1136 ^ n331 ;
  assign n4867 = n2241 ^ x42 ^ 1'b0 ;
  assign n4868 = n4866 & ~n4867 ;
  assign n4869 = n4300 ^ n2274 ^ 1'b0 ;
  assign n4873 = n1625 ^ n1051 ^ 1'b0 ;
  assign n4871 = ~n822 & n1427 ;
  assign n4870 = ( ~n1428 & n2517 ) | ( ~n1428 & n4143 ) | ( n2517 & n4143 ) ;
  assign n4872 = n4871 ^ n4870 ^ n2559 ;
  assign n4874 = n4873 ^ n4872 ^ n365 ;
  assign n4875 = n3200 ^ n2578 ^ x162 ;
  assign n4876 = n1074 & ~n1669 ;
  assign n4877 = n2502 & n4738 ;
  assign n4878 = n4877 ^ n1525 ^ n600 ;
  assign n4879 = n4878 ^ n1875 ^ n960 ;
  assign n4880 = n4876 | n4879 ;
  assign n4881 = n4875 | n4880 ;
  assign n4885 = x168 & n1958 ;
  assign n4886 = n4885 ^ n912 ^ 1'b0 ;
  assign n4887 = n4886 ^ n3638 ^ 1'b0 ;
  assign n4888 = n4785 | n4887 ;
  assign n4889 = n4888 ^ x203 ^ 1'b0 ;
  assign n4882 = n381 & n1173 ;
  assign n4883 = n1678 & n2068 ;
  assign n4884 = n4882 & n4883 ;
  assign n4890 = n4889 ^ n4884 ^ 1'b0 ;
  assign n4891 = n2697 | n4890 ;
  assign n4892 = n4881 | n4891 ;
  assign n4893 = n4189 ^ n3928 ^ n1194 ;
  assign n4894 = x154 | n487 ;
  assign n4895 = n4894 ^ x146 ^ 1'b0 ;
  assign n4896 = ( ~x82 & x236 ) | ( ~x82 & n4363 ) | ( x236 & n4363 ) ;
  assign n4897 = n804 & ~n4896 ;
  assign n4898 = ~n3571 & n4897 ;
  assign n4899 = n2778 & n4898 ;
  assign n4900 = ~n4557 & n4899 ;
  assign n4901 = x10 | n2436 ;
  assign n4902 = n1854 | n4901 ;
  assign n4903 = ~n2673 & n4902 ;
  assign n4904 = n4903 ^ n4435 ^ 1'b0 ;
  assign n4905 = n4904 ^ n2453 ^ 1'b0 ;
  assign n4906 = n2880 ^ n1953 ^ 1'b0 ;
  assign n4907 = n2844 & n4906 ;
  assign n4908 = n2749 ^ n1807 ^ 1'b0 ;
  assign n4909 = ~n2858 & n4908 ;
  assign n4910 = n4909 ^ n4497 ^ 1'b0 ;
  assign n4911 = ( n695 & n1803 ) | ( n695 & ~n2389 ) | ( n1803 & ~n2389 ) ;
  assign n4912 = n4911 ^ n3632 ^ n1264 ;
  assign n4913 = ~n585 & n659 ;
  assign n4914 = n4913 ^ n4165 ^ 1'b0 ;
  assign n4915 = n4914 ^ n1963 ^ 1'b0 ;
  assign n4916 = n4912 & n4915 ;
  assign n4922 = x4 | n810 ;
  assign n4923 = n4922 ^ n1303 ^ n348 ;
  assign n4920 = x175 & ~n625 ;
  assign n4921 = ~n3475 & n4920 ;
  assign n4918 = n2868 ^ n1169 ^ 1'b0 ;
  assign n4917 = n1294 | n2379 ;
  assign n4919 = n4918 ^ n4917 ^ n3316 ;
  assign n4924 = n4923 ^ n4921 ^ n4919 ;
  assign n4926 = ( n632 & n851 ) | ( n632 & ~n3168 ) | ( n851 & ~n3168 ) ;
  assign n4927 = n4810 & n4926 ;
  assign n4928 = n4927 ^ n325 ^ 1'b0 ;
  assign n4925 = ( n1465 & ~n2548 ) | ( n1465 & n3021 ) | ( ~n2548 & n3021 ) ;
  assign n4929 = n4928 ^ n4925 ^ n2583 ;
  assign n4930 = ( n1112 & n3526 ) | ( n1112 & ~n4929 ) | ( n3526 & ~n4929 ) ;
  assign n4931 = n1006 | n1342 ;
  assign n4932 = n1836 | n4931 ;
  assign n4933 = n4932 ^ n3326 ^ n736 ;
  assign n4934 = n4933 ^ n2432 ^ 1'b0 ;
  assign n4935 = ( ~x236 & n1135 ) | ( ~x236 & n1418 ) | ( n1135 & n1418 ) ;
  assign n4936 = n4935 ^ n1196 ^ 1'b0 ;
  assign n4937 = n2626 & ~n4936 ;
  assign n4938 = n4937 ^ n2339 ^ 1'b0 ;
  assign n4939 = n4934 & ~n4938 ;
  assign n4940 = n3865 | n4310 ;
  assign n4941 = n4940 ^ n725 ^ 1'b0 ;
  assign n4942 = n4941 ^ n1183 ^ 1'b0 ;
  assign n4945 = n3332 ^ n1468 ^ 1'b0 ;
  assign n4943 = n2646 ^ n899 ^ 1'b0 ;
  assign n4944 = ~n1903 & n4943 ;
  assign n4946 = n4945 ^ n4944 ^ n1487 ;
  assign n4947 = n4946 ^ n4674 ^ 1'b0 ;
  assign n4948 = n290 & ~n473 ;
  assign n4949 = n1362 & n4948 ;
  assign n4950 = n4949 ^ n1736 ^ x101 ;
  assign n4951 = n1691 ^ n578 ^ x133 ;
  assign n4952 = ( n1244 & ~n2583 ) | ( n1244 & n4951 ) | ( ~n2583 & n4951 ) ;
  assign n4953 = ~n2405 & n2944 ;
  assign n4954 = ~n4327 & n4953 ;
  assign n4955 = n3575 & ~n4954 ;
  assign n4956 = n4952 & n4955 ;
  assign n4958 = x191 & n3008 ;
  assign n4957 = n4005 ^ n1180 ^ 1'b0 ;
  assign n4959 = n4958 ^ n4957 ^ n3338 ;
  assign n4960 = n566 | n1350 ;
  assign n4961 = n4960 ^ x181 ^ 1'b0 ;
  assign n4962 = n4961 ^ n4622 ^ 1'b0 ;
  assign n4963 = ( n1437 & n2905 ) | ( n1437 & n4436 ) | ( n2905 & n4436 ) ;
  assign n4964 = n3156 ^ n1409 ^ 1'b0 ;
  assign n4965 = n1445 & ~n4964 ;
  assign n4973 = ~n1235 & n2520 ;
  assign n4966 = n1922 ^ n820 ^ n276 ;
  assign n4967 = n4966 ^ n4503 ^ n3532 ;
  assign n4968 = x74 ^ x61 ^ 1'b0 ;
  assign n4969 = x232 & ~n4968 ;
  assign n4970 = n4969 ^ n2213 ^ 1'b0 ;
  assign n4971 = n4970 ^ n4127 ^ n1579 ;
  assign n4972 = n4967 & n4971 ;
  assign n4974 = n4973 ^ n4972 ^ 1'b0 ;
  assign n4975 = n4974 ^ n543 ^ 1'b0 ;
  assign n4976 = n4918 & ~n4962 ;
  assign n4977 = n3715 ^ n980 ^ 1'b0 ;
  assign n4978 = ( n2744 & n4521 ) | ( n2744 & ~n4977 ) | ( n4521 & ~n4977 ) ;
  assign n4979 = ~n1040 & n4978 ;
  assign n4980 = x144 & n1024 ;
  assign n4981 = n2630 | n4854 ;
  assign n4982 = n4980 & ~n4981 ;
  assign n4983 = n4982 ^ n3999 ^ n2364 ;
  assign n4984 = n3888 ^ n1052 ^ 1'b0 ;
  assign n4985 = ~n2844 & n4984 ;
  assign n4986 = n4985 ^ n396 ^ 1'b0 ;
  assign n4987 = n3852 ^ n2370 ^ n1704 ;
  assign n4988 = n1583 & ~n4480 ;
  assign n4989 = ~x240 & n4988 ;
  assign n4990 = n406 & n3982 ;
  assign n4991 = ~x99 & n4990 ;
  assign n4992 = n1645 | n4991 ;
  assign n4993 = n4989 & ~n4992 ;
  assign n4994 = n4987 | n4993 ;
  assign n4995 = n4994 ^ n4862 ^ 1'b0 ;
  assign n4998 = n4866 ^ n1637 ^ n758 ;
  assign n4996 = ( ~n544 & n1656 ) | ( ~n544 & n4048 ) | ( n1656 & n4048 ) ;
  assign n4997 = ( n1059 & n1682 ) | ( n1059 & ~n4996 ) | ( n1682 & ~n4996 ) ;
  assign n4999 = n4998 ^ n4997 ^ n2980 ;
  assign n5000 = ( ~n4986 & n4995 ) | ( ~n4986 & n4999 ) | ( n4995 & n4999 ) ;
  assign n5001 = ~n684 & n2171 ;
  assign n5002 = ~n3172 & n5001 ;
  assign n5003 = n5002 ^ n2094 ^ 1'b0 ;
  assign n5004 = n5003 ^ n4815 ^ x139 ;
  assign n5005 = n1581 & ~n4937 ;
  assign n5006 = n3184 ^ n1393 ^ 1'b0 ;
  assign n5007 = n5006 ^ n1901 ^ n1280 ;
  assign n5008 = n5005 | n5007 ;
  assign n5009 = n1933 & ~n5008 ;
  assign n5010 = n3191 ^ n1081 ^ 1'b0 ;
  assign n5011 = n1746 & n5010 ;
  assign n5012 = n2878 ^ n2744 ^ 1'b0 ;
  assign n5013 = ( n2534 & n4162 ) | ( n2534 & n5012 ) | ( n4162 & n5012 ) ;
  assign n5014 = ( n1006 & n5011 ) | ( n1006 & n5013 ) | ( n5011 & n5013 ) ;
  assign n5015 = n3894 ^ n352 ^ x246 ;
  assign n5016 = ~n1108 & n5015 ;
  assign n5017 = n2547 | n2985 ;
  assign n5018 = n4345 ^ n1251 ^ 1'b0 ;
  assign n5019 = n5017 & ~n5018 ;
  assign n5020 = n2599 | n4655 ;
  assign n5024 = n1678 & ~n1934 ;
  assign n5025 = n971 & n5024 ;
  assign n5021 = x52 | n3968 ;
  assign n5022 = ~x237 & n5021 ;
  assign n5023 = n4208 & n5022 ;
  assign n5026 = n5025 ^ n5023 ^ 1'b0 ;
  assign n5027 = n1372 ^ n1239 ^ 1'b0 ;
  assign n5028 = n5027 ^ x88 ^ 1'b0 ;
  assign n5029 = n4072 & ~n5028 ;
  assign n5030 = ( n436 & ~n1042 ) | ( n436 & n4208 ) | ( ~n1042 & n4208 ) ;
  assign n5031 = ~n1789 & n3126 ;
  assign n5032 = n3587 & n5031 ;
  assign n5033 = x68 & ~n5032 ;
  assign n5034 = n3107 & n5033 ;
  assign n5035 = n5034 ^ n4032 ^ 1'b0 ;
  assign n5037 = n827 | n995 ;
  assign n5038 = ( n1802 & ~n3363 ) | ( n1802 & n5037 ) | ( ~n3363 & n5037 ) ;
  assign n5036 = ~n445 & n4091 ;
  assign n5039 = n5038 ^ n5036 ^ n4942 ;
  assign n5041 = ~n1211 & n1917 ;
  assign n5042 = n5041 ^ n2659 ^ 1'b0 ;
  assign n5043 = n1365 ^ n1183 ^ 1'b0 ;
  assign n5044 = ( x248 & n3830 ) | ( x248 & ~n5043 ) | ( n3830 & ~n5043 ) ;
  assign n5045 = n3038 & n5044 ;
  assign n5046 = n5042 & n5045 ;
  assign n5047 = n502 | n5046 ;
  assign n5048 = n5047 ^ n1197 ^ 1'b0 ;
  assign n5040 = n3931 ^ n2868 ^ n711 ;
  assign n5049 = n5048 ^ n5040 ^ n2354 ;
  assign n5050 = ( n362 & n2330 ) | ( n362 & n5049 ) | ( n2330 & n5049 ) ;
  assign n5051 = n293 & n3336 ;
  assign n5052 = ( n2575 & ~n2856 ) | ( n2575 & n3799 ) | ( ~n2856 & n3799 ) ;
  assign n5053 = n5052 ^ n1001 ^ 1'b0 ;
  assign n5063 = ( x34 & n4006 ) | ( x34 & n4034 ) | ( n4006 & n4034 ) ;
  assign n5054 = n3289 ^ n936 ^ n614 ;
  assign n5055 = ~x5 & n2070 ;
  assign n5056 = n5055 ^ n1836 ^ 1'b0 ;
  assign n5057 = ( n790 & ~n1044 ) | ( n790 & n5056 ) | ( ~n1044 & n5056 ) ;
  assign n5058 = n5057 ^ n2616 ^ 1'b0 ;
  assign n5059 = n4911 & ~n5058 ;
  assign n5060 = ( n2076 & ~n3378 ) | ( n2076 & n3795 ) | ( ~n3378 & n3795 ) ;
  assign n5061 = n5060 ^ n4864 ^ n291 ;
  assign n5062 = ( n5054 & n5059 ) | ( n5054 & n5061 ) | ( n5059 & n5061 ) ;
  assign n5064 = n5063 ^ n5062 ^ n4916 ;
  assign n5065 = n3220 & ~n3970 ;
  assign n5066 = ( ~n764 & n1635 ) | ( ~n764 & n2602 ) | ( n1635 & n2602 ) ;
  assign n5072 = n426 | n3065 ;
  assign n5073 = n5072 ^ n2383 ^ 1'b0 ;
  assign n5067 = n2140 & n3611 ;
  assign n5068 = n5067 ^ n3854 ^ 1'b0 ;
  assign n5069 = n5068 ^ n3105 ^ 1'b0 ;
  assign n5070 = ~n2347 & n5069 ;
  assign n5071 = n5070 ^ n3888 ^ n1118 ;
  assign n5074 = n5073 ^ n5071 ^ 1'b0 ;
  assign n5075 = n944 ^ x126 ^ 1'b0 ;
  assign n5076 = ( x182 & n1688 ) | ( x182 & n3205 ) | ( n1688 & n3205 ) ;
  assign n5077 = ~n1050 & n1600 ;
  assign n5078 = n1186 & n5077 ;
  assign n5079 = n5078 ^ n3500 ^ 1'b0 ;
  assign n5080 = n5076 & ~n5079 ;
  assign n5081 = n5075 & ~n5080 ;
  assign n5086 = ( n479 & n1053 ) | ( n479 & ~n1556 ) | ( n1053 & ~n1556 ) ;
  assign n5082 = n2437 | n3594 ;
  assign n5083 = n731 & ~n2819 ;
  assign n5084 = ~n4407 & n5083 ;
  assign n5085 = n5082 | n5084 ;
  assign n5087 = n5086 ^ n5085 ^ n4301 ;
  assign n5088 = n4790 ^ n1235 ^ x79 ;
  assign n5089 = x193 ^ x133 ^ 1'b0 ;
  assign n5090 = ( ~n1272 & n1830 ) | ( ~n1272 & n5089 ) | ( n1830 & n5089 ) ;
  assign n5091 = n3362 & ~n4912 ;
  assign n5092 = ( n926 & ~n1579 ) | ( n926 & n3643 ) | ( ~n1579 & n3643 ) ;
  assign n5093 = ( n1277 & n4401 ) | ( n1277 & n5092 ) | ( n4401 & n5092 ) ;
  assign n5094 = n5093 ^ n3604 ^ n1280 ;
  assign n5095 = x99 & ~n2844 ;
  assign n5096 = n5095 ^ x92 ^ 1'b0 ;
  assign n5097 = n511 & n2642 ;
  assign n5098 = n1217 ^ n397 ^ 1'b0 ;
  assign n5104 = n2707 ^ n1180 ^ 1'b0 ;
  assign n5099 = n459 & n626 ;
  assign n5100 = n5099 ^ n731 ^ 1'b0 ;
  assign n5101 = n3395 ^ n406 ^ 1'b0 ;
  assign n5102 = n1996 & n5101 ;
  assign n5103 = ~n5100 & n5102 ;
  assign n5105 = n5104 ^ n5103 ^ 1'b0 ;
  assign n5106 = n3732 | n5105 ;
  assign n5107 = n2985 | n5106 ;
  assign n5109 = ( n1352 & n1859 ) | ( n1352 & ~n2127 ) | ( n1859 & ~n2127 ) ;
  assign n5108 = n392 & ~n2630 ;
  assign n5110 = n5109 ^ n5108 ^ 1'b0 ;
  assign n5111 = n1672 ^ n413 ^ 1'b0 ;
  assign n5112 = n5111 ^ n2524 ^ 1'b0 ;
  assign n5113 = n4619 | n5112 ;
  assign n5114 = n5113 ^ n1508 ^ 1'b0 ;
  assign n5115 = n3561 ^ n3253 ^ x159 ;
  assign n5120 = ( ~n736 & n816 ) | ( ~n736 & n3682 ) | ( n816 & n3682 ) ;
  assign n5116 = n2824 ^ n2794 ^ n492 ;
  assign n5117 = ( n1883 & n3059 ) | ( n1883 & n5116 ) | ( n3059 & n5116 ) ;
  assign n5118 = n1634 | n5117 ;
  assign n5119 = n1403 & ~n5118 ;
  assign n5121 = n5120 ^ n5119 ^ 1'b0 ;
  assign n5122 = n2138 ^ n1260 ^ n1243 ;
  assign n5123 = ~n4335 & n5122 ;
  assign n5124 = n595 | n679 ;
  assign n5125 = n879 ^ n547 ^ 1'b0 ;
  assign n5126 = n5125 ^ n1705 ^ x172 ;
  assign n5127 = ~n5124 & n5126 ;
  assign n5132 = n272 & ~n2016 ;
  assign n5133 = n5132 ^ n1652 ^ n374 ;
  assign n5134 = ( n1478 & ~n1844 ) | ( n1478 & n5133 ) | ( ~n1844 & n5133 ) ;
  assign n5135 = n4677 & n5134 ;
  assign n5128 = n4748 ^ n969 ^ x214 ;
  assign n5129 = n2384 ^ n490 ^ n455 ;
  assign n5130 = n2145 & ~n5129 ;
  assign n5131 = n5128 & ~n5130 ;
  assign n5136 = n5135 ^ n5131 ^ 1'b0 ;
  assign n5137 = n730 ^ x242 ^ x221 ;
  assign n5138 = n361 & n3711 ;
  assign n5139 = n5137 & n5138 ;
  assign n5140 = ~n3923 & n5139 ;
  assign n5141 = n1517 ^ x140 ^ 1'b0 ;
  assign n5142 = n2665 | n5141 ;
  assign n5143 = n3468 & ~n5142 ;
  assign n5144 = n5143 ^ n3254 ^ 1'b0 ;
  assign n5145 = n1403 & ~n5144 ;
  assign n5146 = n5140 & n5145 ;
  assign n5147 = n5100 ^ n3106 ^ 1'b0 ;
  assign n5148 = n5146 | n5147 ;
  assign n5149 = n5148 ^ n821 ^ n542 ;
  assign n5150 = ( n551 & n3290 ) | ( n551 & n4779 ) | ( n3290 & n4779 ) ;
  assign n5151 = n3438 ^ n3402 ^ n299 ;
  assign n5152 = n4118 ^ n1294 ^ 1'b0 ;
  assign n5153 = ~n2555 & n5152 ;
  assign n5154 = n3310 ^ n1307 ^ n1097 ;
  assign n5155 = n5154 ^ n1289 ^ n379 ;
  assign n5156 = x100 & n5155 ;
  assign n5157 = ~n4077 & n5156 ;
  assign n5160 = n2112 ^ n2101 ^ 1'b0 ;
  assign n5161 = ~n430 & n3024 ;
  assign n5162 = n566 & n5161 ;
  assign n5163 = n5162 ^ n3285 ^ 1'b0 ;
  assign n5164 = n745 & ~n5163 ;
  assign n5165 = ( n3289 & n5160 ) | ( n3289 & n5164 ) | ( n5160 & n5164 ) ;
  assign n5158 = n4984 ^ n1783 ^ x27 ;
  assign n5159 = n1091 & ~n5158 ;
  assign n5166 = n5165 ^ n5159 ^ 1'b0 ;
  assign n5167 = ( x47 & n2878 ) | ( x47 & n4239 ) | ( n2878 & n4239 ) ;
  assign n5168 = ~n654 & n1003 ;
  assign n5169 = n1381 ^ n321 ^ x2 ;
  assign n5170 = x209 & ~n5169 ;
  assign n5171 = n2461 & n5170 ;
  assign n5172 = n5171 ^ n4926 ^ 1'b0 ;
  assign n5173 = ~n1026 & n1700 ;
  assign n5174 = n3651 ^ n2033 ^ 1'b0 ;
  assign n5175 = ~n2825 & n5174 ;
  assign n5176 = n4251 & ~n5175 ;
  assign n5177 = n1252 & n3233 ;
  assign n5178 = n4256 & ~n5177 ;
  assign n5179 = n5178 ^ n545 ^ 1'b0 ;
  assign n5180 = ~n1469 & n4055 ;
  assign n5181 = n1685 & n5180 ;
  assign n5182 = n1433 | n5181 ;
  assign n5183 = n2617 & ~n5182 ;
  assign n5187 = n3629 ^ n1776 ^ 1'b0 ;
  assign n5188 = n2384 & n5187 ;
  assign n5184 = n483 ^ n366 ^ x209 ;
  assign n5185 = n3604 & ~n4502 ;
  assign n5186 = n5184 | n5185 ;
  assign n5189 = n5188 ^ n5186 ^ 1'b0 ;
  assign n5190 = x215 & ~n420 ;
  assign n5191 = ~n5189 & n5190 ;
  assign n5192 = n3500 & ~n5191 ;
  assign n5193 = n3009 & n5192 ;
  assign n5194 = n5183 | n5193 ;
  assign n5195 = n5194 ^ n3393 ^ 1'b0 ;
  assign n5196 = n4965 ^ x1 ^ 1'b0 ;
  assign n5197 = ~n2769 & n3722 ;
  assign n5198 = n3326 & n3717 ;
  assign n5199 = n5197 & n5198 ;
  assign n5200 = n2689 | n4796 ;
  assign n5201 = n3514 | n5200 ;
  assign n5202 = n3087 & ~n5201 ;
  assign n5203 = n2544 | n4781 ;
  assign n5204 = n5203 ^ n5129 ^ 1'b0 ;
  assign n5205 = n290 & n5204 ;
  assign n5207 = n763 | n937 ;
  assign n5206 = x40 & ~n4710 ;
  assign n5208 = n5207 ^ n5206 ^ 1'b0 ;
  assign n5209 = n3427 ^ n2189 ^ 1'b0 ;
  assign n5210 = ~n706 & n1174 ;
  assign n5211 = n1876 & ~n5210 ;
  assign n5212 = n5209 & n5211 ;
  assign n5213 = n1635 ^ n378 ^ 1'b0 ;
  assign n5214 = n291 & n5213 ;
  assign n5215 = x248 & n1251 ;
  assign n5216 = n5215 ^ n2629 ^ 1'b0 ;
  assign n5217 = n5216 ^ n4144 ^ 1'b0 ;
  assign n5218 = ~n284 & n656 ;
  assign n5219 = ~n1667 & n5218 ;
  assign n5220 = n3227 ^ n1233 ^ 1'b0 ;
  assign n5221 = ~n5219 & n5220 ;
  assign n5222 = n5221 ^ n5204 ^ 1'b0 ;
  assign n5223 = n4306 ^ n4264 ^ n1591 ;
  assign n5224 = n693 | n3658 ;
  assign n5225 = n5223 & ~n5224 ;
  assign n5226 = ( ~n497 & n947 ) | ( ~n497 & n3061 ) | ( n947 & n3061 ) ;
  assign n5227 = n865 & n5226 ;
  assign n5228 = n5227 ^ x151 ^ 1'b0 ;
  assign n5229 = x7 & n4849 ;
  assign n5230 = n5229 ^ n4043 ^ 1'b0 ;
  assign n5231 = n5228 | n5230 ;
  assign n5232 = n523 & n979 ;
  assign n5233 = n1397 & n5232 ;
  assign n5234 = n366 ^ x159 ^ 1'b0 ;
  assign n5235 = ( n4346 & n5233 ) | ( n4346 & n5234 ) | ( n5233 & n5234 ) ;
  assign n5236 = n2725 ^ n1698 ^ n877 ;
  assign n5237 = n2700 & n3407 ;
  assign n5238 = n5237 ^ n3561 ^ 1'b0 ;
  assign n5239 = ( n2050 & n2558 ) | ( n2050 & n4503 ) | ( n2558 & n4503 ) ;
  assign n5240 = ( n4509 & ~n5238 ) | ( n4509 & n5239 ) | ( ~n5238 & n5239 ) ;
  assign n5241 = n3787 & ~n5240 ;
  assign n5242 = n5241 ^ n4310 ^ 1'b0 ;
  assign n5243 = n2114 & ~n5228 ;
  assign n5244 = n5243 ^ n3135 ^ 1'b0 ;
  assign n5245 = n947 | n1184 ;
  assign n5246 = n3583 | n5245 ;
  assign n5247 = ~n262 & n731 ;
  assign n5248 = ~x145 & n5247 ;
  assign n5249 = n5248 ^ n3227 ^ n693 ;
  assign n5250 = n5249 ^ n3154 ^ 1'b0 ;
  assign n5251 = n5044 ^ n294 ^ 1'b0 ;
  assign n5252 = n5251 ^ n4966 ^ n608 ;
  assign n5253 = n1254 ^ n1214 ^ n1149 ;
  assign n5254 = ( n2771 & ~n3296 ) | ( n2771 & n5253 ) | ( ~n3296 & n5253 ) ;
  assign n5255 = x165 & ~n2451 ;
  assign n5256 = ~n3964 & n5255 ;
  assign n5257 = n2438 ^ n2428 ^ 1'b0 ;
  assign n5258 = ~n947 & n1836 ;
  assign n5259 = ~n1003 & n5258 ;
  assign n5260 = n2662 & n3828 ;
  assign n5261 = n5259 & n5260 ;
  assign n5262 = n4376 ^ n3347 ^ x81 ;
  assign n5263 = n5262 ^ n3290 ^ 1'b0 ;
  assign n5264 = n2904 ^ n2513 ^ n1385 ;
  assign n5265 = x49 & ~n5264 ;
  assign n5266 = n4421 ^ n3133 ^ n887 ;
  assign n5267 = ~n2553 & n5266 ;
  assign n5268 = n5267 ^ n3517 ^ 1'b0 ;
  assign n5269 = n3607 ^ n2059 ^ 1'b0 ;
  assign n5270 = n639 | n5269 ;
  assign n5271 = n5270 ^ n3849 ^ n3553 ;
  assign n5272 = n5271 ^ n1097 ^ 1'b0 ;
  assign n5274 = n4307 ^ n750 ^ 1'b0 ;
  assign n5273 = n2210 & ~n3826 ;
  assign n5275 = n5274 ^ n5273 ^ 1'b0 ;
  assign n5276 = ~n615 & n4808 ;
  assign n5277 = n5276 ^ n4986 ^ n402 ;
  assign n5278 = n4162 & ~n4183 ;
  assign n5279 = ~n3678 & n5278 ;
  assign n5283 = ~n1035 & n1461 ;
  assign n5284 = n5283 ^ n335 ^ 1'b0 ;
  assign n5280 = ~n461 & n2408 ;
  assign n5281 = n3125 & n5280 ;
  assign n5282 = n1447 & ~n5281 ;
  assign n5285 = n5284 ^ n5282 ^ 1'b0 ;
  assign n5286 = n1114 & n5285 ;
  assign n5287 = ~n3509 & n4163 ;
  assign n5288 = n5287 ^ n4306 ^ 1'b0 ;
  assign n5289 = n4922 ^ n301 ^ 1'b0 ;
  assign n5290 = n2384 ^ n2184 ^ n1179 ;
  assign n5291 = n5290 ^ x230 ^ 1'b0 ;
  assign n5292 = n2783 ^ n1750 ^ n763 ;
  assign n5293 = n774 ^ n374 ^ 1'b0 ;
  assign n5294 = n5293 ^ n2893 ^ n779 ;
  assign n5295 = n5294 ^ n977 ^ 1'b0 ;
  assign n5296 = n5295 ^ n3575 ^ n2041 ;
  assign n5297 = n5292 & ~n5296 ;
  assign n5298 = ~n1676 & n5297 ;
  assign n5299 = ~n3666 & n4264 ;
  assign n5300 = n2022 ^ n568 ^ n476 ;
  assign n5303 = ( ~n578 & n1309 ) | ( ~n578 & n2574 ) | ( n1309 & n2574 ) ;
  assign n5304 = n5303 ^ n2558 ^ n1837 ;
  assign n5301 = n3070 ^ n1384 ^ 1'b0 ;
  assign n5302 = ~n2254 & n5301 ;
  assign n5305 = n5304 ^ n5302 ^ 1'b0 ;
  assign n5306 = ~n5300 & n5305 ;
  assign n5307 = n4443 ^ n3754 ^ n2763 ;
  assign n5308 = ( n5299 & ~n5306 ) | ( n5299 & n5307 ) | ( ~n5306 & n5307 ) ;
  assign n5309 = n2132 ^ n1284 ^ 1'b0 ;
  assign n5310 = ( n1196 & n2071 ) | ( n1196 & n5309 ) | ( n2071 & n5309 ) ;
  assign n5311 = n2869 ^ n1462 ^ n832 ;
  assign n5312 = ~n1118 & n1348 ;
  assign n5313 = n5311 & n5312 ;
  assign n5314 = n736 & n3163 ;
  assign n5315 = n5314 ^ n1712 ^ 1'b0 ;
  assign n5316 = ~n2108 & n5315 ;
  assign n5317 = n915 & ~n4028 ;
  assign n5318 = n5317 ^ n1299 ^ 1'b0 ;
  assign n5319 = n763 | n5318 ;
  assign n5320 = n1646 | n5319 ;
  assign n5321 = ~n430 & n536 ;
  assign n5324 = n904 & n3376 ;
  assign n5322 = ( n1550 & n2720 ) | ( n1550 & ~n3042 ) | ( n2720 & ~n3042 ) ;
  assign n5323 = ( n932 & n5295 ) | ( n932 & n5322 ) | ( n5295 & n5322 ) ;
  assign n5325 = n5324 ^ n5323 ^ x97 ;
  assign n5326 = ( ~n871 & n2997 ) | ( ~n871 & n5325 ) | ( n2997 & n5325 ) ;
  assign n5327 = ( x241 & n2395 ) | ( x241 & ~n3058 ) | ( n2395 & ~n3058 ) ;
  assign n5328 = ( n573 & n2798 ) | ( n573 & ~n5327 ) | ( n2798 & ~n5327 ) ;
  assign n5329 = ( n802 & n1250 ) | ( n802 & n3440 ) | ( n1250 & n3440 ) ;
  assign n5330 = n5329 ^ n4169 ^ 1'b0 ;
  assign n5331 = ~n5328 & n5330 ;
  assign n5332 = n1287 ^ n264 ^ 1'b0 ;
  assign n5333 = n426 | n5332 ;
  assign n5334 = n3858 | n3966 ;
  assign n5340 = n4646 ^ n936 ^ 1'b0 ;
  assign n5335 = n3289 & ~n3587 ;
  assign n5336 = ~x192 & n5335 ;
  assign n5337 = n5336 ^ n3174 ^ n1298 ;
  assign n5338 = ( ~n2655 & n4066 ) | ( ~n2655 & n5337 ) | ( n4066 & n5337 ) ;
  assign n5339 = n3323 & ~n5338 ;
  assign n5341 = n5340 ^ n5339 ^ 1'b0 ;
  assign n5342 = n1569 ^ n1240 ^ x192 ;
  assign n5343 = n5342 ^ n868 ^ n419 ;
  assign n5344 = n5343 ^ n5244 ^ n3156 ;
  assign n5360 = n1743 ^ n722 ^ n530 ;
  assign n5361 = n5360 ^ x144 ^ 1'b0 ;
  assign n5362 = n4609 | n5361 ;
  assign n5363 = n5362 ^ n1251 ^ n704 ;
  assign n5357 = ~n1665 & n3148 ;
  assign n5358 = ~n3292 & n5357 ;
  assign n5359 = n5358 ^ n5342 ^ 1'b0 ;
  assign n5355 = n2076 ^ n1814 ^ n1442 ;
  assign n5354 = n367 & n3352 ;
  assign n5356 = n5355 ^ n5354 ^ 1'b0 ;
  assign n5364 = n5363 ^ n5359 ^ n5356 ;
  assign n5351 = n1246 | n1470 ;
  assign n5352 = n5351 ^ n2297 ^ 1'b0 ;
  assign n5345 = n1180 | n4854 ;
  assign n5346 = n5345 ^ n1997 ^ 1'b0 ;
  assign n5347 = n5346 ^ n2319 ^ 1'b0 ;
  assign n5348 = n466 & n2923 ;
  assign n5349 = n5348 ^ n558 ^ 1'b0 ;
  assign n5350 = n5347 & ~n5349 ;
  assign n5353 = n5352 ^ n5350 ^ 1'b0 ;
  assign n5365 = n5364 ^ n5353 ^ n1917 ;
  assign n5366 = ~n382 & n4870 ;
  assign n5367 = n5366 ^ n1298 ^ 1'b0 ;
  assign n5368 = ( n1090 & n2155 ) | ( n1090 & n3766 ) | ( n2155 & n3766 ) ;
  assign n5371 = n1045 ^ x221 ^ x82 ;
  assign n5369 = n618 | n2867 ;
  assign n5370 = n5369 ^ n4600 ^ 1'b0 ;
  assign n5372 = n5371 ^ n5370 ^ 1'b0 ;
  assign n5373 = ( n1146 & ~n3260 ) | ( n1146 & n3901 ) | ( ~n3260 & n3901 ) ;
  assign n5374 = n5373 ^ n3070 ^ 1'b0 ;
  assign n5375 = n5288 & n5374 ;
  assign n5376 = n1467 & n5375 ;
  assign n5377 = n449 & n2590 ;
  assign n5378 = n1879 & n5377 ;
  assign n5379 = n1202 | n5378 ;
  assign n5380 = n4352 & ~n5379 ;
  assign n5381 = ( ~n326 & n4864 ) | ( ~n326 & n5380 ) | ( n4864 & n5380 ) ;
  assign n5382 = n2377 ^ n693 ^ 1'b0 ;
  assign n5383 = n3967 | n5382 ;
  assign n5385 = ( ~n554 & n961 ) | ( ~n554 & n2794 ) | ( n961 & n2794 ) ;
  assign n5384 = n1352 | n2805 ;
  assign n5386 = n5385 ^ n5384 ^ 1'b0 ;
  assign n5387 = x193 & ~n4404 ;
  assign n5388 = n2738 ^ n1018 ^ x221 ;
  assign n5389 = n2998 & ~n5388 ;
  assign n5390 = n5389 ^ n4371 ^ 1'b0 ;
  assign n5391 = x103 & n4670 ;
  assign n5392 = n2870 & n5391 ;
  assign n5393 = ( n1161 & n3841 ) | ( n1161 & n5392 ) | ( n3841 & n5392 ) ;
  assign n5394 = n1969 & ~n2649 ;
  assign n5395 = n1910 | n3237 ;
  assign n5396 = n5395 ^ n3885 ^ 1'b0 ;
  assign n5397 = n5394 | n5396 ;
  assign n5398 = x225 & n1517 ;
  assign n5399 = n2525 | n5398 ;
  assign n5400 = n3377 & n5038 ;
  assign n5401 = n5400 ^ n765 ^ 1'b0 ;
  assign n5402 = n5076 ^ n1953 ^ 1'b0 ;
  assign n5403 = n2854 ^ n857 ^ 1'b0 ;
  assign n5404 = n5403 ^ n3909 ^ 1'b0 ;
  assign n5405 = n1489 & n5404 ;
  assign n5406 = ( n5401 & n5402 ) | ( n5401 & ~n5405 ) | ( n5402 & ~n5405 ) ;
  assign n5407 = n2602 ^ n1701 ^ n566 ;
  assign n5408 = n5407 ^ n4919 ^ n3307 ;
  assign n5409 = n2225 ^ n2112 ^ n576 ;
  assign n5410 = n5409 ^ n908 ^ 1'b0 ;
  assign n5411 = n1627 | n5410 ;
  assign n5412 = n2201 & ~n5411 ;
  assign n5413 = ~x49 & n5412 ;
  assign n5414 = n2246 | n5413 ;
  assign n5415 = n5408 | n5414 ;
  assign n5421 = n1563 | n3254 ;
  assign n5422 = n1887 | n5421 ;
  assign n5416 = ( x12 & ~n1494 ) | ( x12 & n3065 ) | ( ~n1494 & n3065 ) ;
  assign n5417 = ~n1344 & n5416 ;
  assign n5418 = ~n2076 & n5417 ;
  assign n5419 = n5418 ^ n1525 ^ 1'b0 ;
  assign n5420 = n881 & n5419 ;
  assign n5423 = n5422 ^ n5420 ^ 1'b0 ;
  assign n5424 = x217 & n5423 ;
  assign n5425 = ~x77 & n1452 ;
  assign n5426 = n5425 ^ n1985 ^ 1'b0 ;
  assign n5427 = n5424 & n5426 ;
  assign n5428 = n3946 & n4429 ;
  assign n5431 = ~x253 & n3939 ;
  assign n5432 = ~x5 & n434 ;
  assign n5433 = n1355 & n5432 ;
  assign n5434 = n4978 | n5433 ;
  assign n5435 = n5431 & ~n5434 ;
  assign n5429 = n5343 ^ n597 ^ 1'b0 ;
  assign n5430 = n3999 & n5429 ;
  assign n5436 = n5435 ^ n5430 ^ n2512 ;
  assign n5437 = n2723 & ~n3162 ;
  assign n5438 = n5437 ^ n2527 ^ 1'b0 ;
  assign n5439 = ~n2666 & n3249 ;
  assign n5440 = x164 & n2965 ;
  assign n5441 = n5440 ^ n4294 ^ n747 ;
  assign n5442 = n5439 & n5441 ;
  assign n5444 = n2087 ^ n1099 ^ x236 ;
  assign n5445 = n338 & ~n5444 ;
  assign n5446 = n5445 ^ n2325 ^ n1418 ;
  assign n5443 = n1616 ^ x39 ^ 1'b0 ;
  assign n5447 = n5446 ^ n5443 ^ 1'b0 ;
  assign n5448 = ~n1385 & n5447 ;
  assign n5450 = n1268 ^ n749 ^ 1'b0 ;
  assign n5451 = n293 & ~n5450 ;
  assign n5449 = n1873 ^ n632 ^ 1'b0 ;
  assign n5452 = n5451 ^ n5449 ^ n3542 ;
  assign n5453 = ( n809 & n2093 ) | ( n809 & n5452 ) | ( n2093 & n5452 ) ;
  assign n5454 = n2116 | n2243 ;
  assign n5455 = n570 & n5454 ;
  assign n5456 = ( n1692 & n2519 ) | ( n1692 & n3928 ) | ( n2519 & n3928 ) ;
  assign n5457 = ( n1619 & ~n3376 ) | ( n1619 & n5456 ) | ( ~n3376 & n5456 ) ;
  assign n5458 = n5457 ^ n3442 ^ n3129 ;
  assign n5459 = ( n5453 & n5455 ) | ( n5453 & ~n5458 ) | ( n5455 & ~n5458 ) ;
  assign n5460 = n3790 ^ n3309 ^ n3135 ;
  assign n5461 = n695 | n1184 ;
  assign n5462 = ~n831 & n4286 ;
  assign n5463 = ~n5461 & n5462 ;
  assign n5464 = ( n864 & n2267 ) | ( n864 & ~n5463 ) | ( n2267 & ~n5463 ) ;
  assign n5465 = n5464 ^ n3275 ^ 1'b0 ;
  assign n5466 = n3831 & ~n5465 ;
  assign n5478 = n1252 & n1264 ;
  assign n5479 = n5478 ^ n547 ^ 1'b0 ;
  assign n5477 = x156 & n500 ;
  assign n5480 = n5479 ^ n5477 ^ 1'b0 ;
  assign n5472 = ~n2135 & n4126 ;
  assign n5473 = n5472 ^ n4565 ^ 1'b0 ;
  assign n5469 = n3126 & n3249 ;
  assign n5470 = n5469 ^ n3636 ^ 1'b0 ;
  assign n5471 = n5470 ^ n516 ^ 1'b0 ;
  assign n5474 = n5473 ^ n5471 ^ n3801 ;
  assign n5475 = n5474 ^ n1356 ^ 1'b0 ;
  assign n5476 = n402 | n5475 ;
  assign n5467 = n2243 & n3341 ;
  assign n5468 = n5467 ^ n3524 ^ n1813 ;
  assign n5481 = n5480 ^ n5476 ^ n5468 ;
  assign n5482 = n5466 & ~n5481 ;
  assign n5483 = n1743 & n5482 ;
  assign n5484 = ~n5460 & n5483 ;
  assign n5485 = n3392 ^ n573 ^ 1'b0 ;
  assign n5486 = ( n3063 & ~n5051 ) | ( n3063 & n5485 ) | ( ~n5051 & n5485 ) ;
  assign n5488 = n1948 ^ n1824 ^ 1'b0 ;
  assign n5487 = n544 & n838 ;
  assign n5489 = n5488 ^ n5487 ^ 1'b0 ;
  assign n5490 = n5489 ^ n301 ^ 1'b0 ;
  assign n5491 = ( n2114 & n2192 ) | ( n2114 & ~n2700 ) | ( n2192 & ~n2700 ) ;
  assign n5492 = n3349 ^ n2862 ^ 1'b0 ;
  assign n5493 = n3112 ^ n2382 ^ n799 ;
  assign n5494 = ~n5492 & n5493 ;
  assign n5495 = ~n4762 & n5494 ;
  assign n5496 = n5491 & n5495 ;
  assign n5497 = n3436 & n5212 ;
  assign n5498 = n4242 ^ n3804 ^ n2724 ;
  assign n5499 = ( n1986 & n2314 ) | ( n1986 & ~n4928 ) | ( n2314 & ~n4928 ) ;
  assign n5500 = n802 | n2070 ;
  assign n5501 = n1645 | n5500 ;
  assign n5502 = n5499 & ~n5501 ;
  assign n5503 = n1737 ^ n1405 ^ x249 ;
  assign n5504 = ( n262 & n508 ) | ( n262 & n5503 ) | ( n508 & n5503 ) ;
  assign n5505 = n5504 ^ n4947 ^ 1'b0 ;
  assign n5506 = n5502 | n5505 ;
  assign n5507 = ~n1105 & n1574 ;
  assign n5508 = n5506 & ~n5507 ;
  assign n5509 = n3126 ^ n1004 ^ 1'b0 ;
  assign n5510 = n4634 & n5509 ;
  assign n5511 = n1761 & ~n4337 ;
  assign n5512 = n5511 ^ n3594 ^ 1'b0 ;
  assign n5513 = ( n2716 & ~n2889 ) | ( n2716 & n5512 ) | ( ~n2889 & n5512 ) ;
  assign n5514 = ( n376 & ~n1184 ) | ( n376 & n1390 ) | ( ~n1184 & n1390 ) ;
  assign n5515 = x11 & ~n5514 ;
  assign n5516 = n5515 ^ n3117 ^ 1'b0 ;
  assign n5517 = n2191 | n5516 ;
  assign n5519 = ~x106 & n1099 ;
  assign n5520 = n2779 & n5519 ;
  assign n5521 = ~n2906 & n5520 ;
  assign n5522 = n5521 ^ x241 ^ 1'b0 ;
  assign n5523 = ( n866 & n2805 ) | ( n866 & ~n5522 ) | ( n2805 & ~n5522 ) ;
  assign n5518 = n4883 & n4967 ;
  assign n5524 = n5523 ^ n5518 ^ 1'b0 ;
  assign n5525 = n5073 ^ n2195 ^ 1'b0 ;
  assign n5526 = ~n1991 & n5525 ;
  assign n5527 = n1763 ^ x94 ^ 1'b0 ;
  assign n5528 = n2654 | n5527 ;
  assign n5529 = n5528 ^ n3110 ^ 1'b0 ;
  assign n5530 = ( ~n1395 & n4268 ) | ( ~n1395 & n5529 ) | ( n4268 & n5529 ) ;
  assign n5531 = n2291 & ~n2345 ;
  assign n5532 = n5531 ^ n5071 ^ n4282 ;
  assign n5533 = n5532 ^ n2659 ^ 1'b0 ;
  assign n5534 = n3197 ^ n1487 ^ 1'b0 ;
  assign n5535 = n1681 & ~n5534 ;
  assign n5536 = n5535 ^ n1995 ^ 1'b0 ;
  assign n5537 = n2241 | n2432 ;
  assign n5538 = n4726 & ~n5537 ;
  assign n5539 = n4147 ^ n2116 ^ n331 ;
  assign n5540 = n3101 ^ n2833 ^ 1'b0 ;
  assign n5541 = ( n1709 & ~n2819 ) | ( n1709 & n5540 ) | ( ~n2819 & n5540 ) ;
  assign n5542 = n3955 ^ n3029 ^ n1894 ;
  assign n5543 = n5542 ^ n4544 ^ 1'b0 ;
  assign n5544 = ~n5541 & n5543 ;
  assign n5545 = n553 & ~n2912 ;
  assign n5546 = n1897 & ~n5545 ;
  assign n5547 = n5546 ^ n1953 ^ 1'b0 ;
  assign n5548 = n1582 ^ n516 ^ 1'b0 ;
  assign n5549 = n5547 & ~n5548 ;
  assign n5550 = x218 & n5549 ;
  assign n5551 = n548 & n5550 ;
  assign n5552 = x132 & ~n1977 ;
  assign n5553 = n1649 & n5552 ;
  assign n5554 = n1327 | n3068 ;
  assign n5555 = ~n5553 & n5554 ;
  assign n5556 = ~n3384 & n5555 ;
  assign n5559 = ~n403 & n3711 ;
  assign n5558 = n1957 & ~n4968 ;
  assign n5560 = n5559 ^ n5558 ^ 1'b0 ;
  assign n5557 = n3518 ^ x139 ^ 1'b0 ;
  assign n5561 = n5560 ^ n5557 ^ 1'b0 ;
  assign n5562 = n1807 & ~n1893 ;
  assign n5563 = n5562 ^ n4638 ^ 1'b0 ;
  assign n5564 = ( n457 & n5561 ) | ( n457 & n5563 ) | ( n5561 & n5563 ) ;
  assign n5565 = x239 & n391 ;
  assign n5566 = n5565 ^ n3909 ^ 1'b0 ;
  assign n5567 = n3220 ^ n1283 ^ 1'b0 ;
  assign n5568 = n5567 ^ n2782 ^ x120 ;
  assign n5569 = n767 | n5568 ;
  assign n5570 = n1812 | n5569 ;
  assign n5571 = ( n3279 & n3548 ) | ( n3279 & ~n3658 ) | ( n3548 & ~n3658 ) ;
  assign n5572 = n5571 ^ n3141 ^ 1'b0 ;
  assign n5573 = n5388 & n5572 ;
  assign n5574 = n1027 & n1358 ;
  assign n5575 = n3311 ^ n813 ^ 1'b0 ;
  assign n5576 = ( n311 & n5574 ) | ( n311 & n5575 ) | ( n5574 & n5575 ) ;
  assign n5577 = ( x87 & n551 ) | ( x87 & n810 ) | ( n551 & n810 ) ;
  assign n5578 = n3024 & n5577 ;
  assign n5579 = n5576 & n5578 ;
  assign n5580 = n3767 ^ n1180 ^ 1'b0 ;
  assign n5581 = ~n3851 & n5580 ;
  assign n5582 = n2520 ^ n1353 ^ 1'b0 ;
  assign n5585 = n4502 ^ n2730 ^ n1675 ;
  assign n5583 = n4710 ^ n4010 ^ n1780 ;
  assign n5584 = n5583 ^ n2733 ^ x189 ;
  assign n5586 = n5585 ^ n5584 ^ 1'b0 ;
  assign n5587 = n2451 | n5586 ;
  assign n5588 = n4725 ^ n4093 ^ 1'b0 ;
  assign n5589 = n5587 | n5588 ;
  assign n5591 = ~n4219 & n4961 ;
  assign n5592 = ~n431 & n5591 ;
  assign n5590 = x65 & x79 ;
  assign n5593 = n5592 ^ n5590 ^ 1'b0 ;
  assign n5594 = n5577 ^ n3449 ^ 1'b0 ;
  assign n5595 = n5593 & ~n5594 ;
  assign n5596 = ( ~x40 & n600 ) | ( ~x40 & n3437 ) | ( n600 & n3437 ) ;
  assign n5597 = ( ~n1304 & n2676 ) | ( ~n1304 & n5596 ) | ( n2676 & n5596 ) ;
  assign n5598 = ( ~n1297 & n2074 ) | ( ~n1297 & n5597 ) | ( n2074 & n5597 ) ;
  assign n5603 = n733 | n1086 ;
  assign n5604 = n5603 ^ n1205 ^ 1'b0 ;
  assign n5602 = ~n1312 & n3021 ;
  assign n5605 = n5604 ^ n5602 ^ 1'b0 ;
  assign n5599 = ( ~n2924 & n2936 ) | ( ~n2924 & n4281 ) | ( n2936 & n4281 ) ;
  assign n5600 = n3383 | n3476 ;
  assign n5601 = n5599 | n5600 ;
  assign n5606 = n5605 ^ n5601 ^ 1'b0 ;
  assign n5607 = ~n5470 & n5606 ;
  assign n5608 = ( n3243 & n5183 ) | ( n3243 & ~n5233 ) | ( n5183 & ~n5233 ) ;
  assign n5609 = ~n634 & n2340 ;
  assign n5610 = n5609 ^ n3659 ^ 1'b0 ;
  assign n5611 = n2163 | n5610 ;
  assign n5612 = n5611 ^ n2213 ^ 1'b0 ;
  assign n5613 = n5612 ^ n1875 ^ 1'b0 ;
  assign n5614 = ~n3228 & n3569 ;
  assign n5615 = ~n2011 & n5614 ;
  assign n5617 = n2821 & ~n3585 ;
  assign n5618 = n1192 & n5617 ;
  assign n5616 = x66 & ~n2676 ;
  assign n5619 = n5618 ^ n5616 ^ 1'b0 ;
  assign n5620 = ( n4590 & n5615 ) | ( n4590 & ~n5619 ) | ( n5615 & ~n5619 ) ;
  assign n5621 = n352 | n3801 ;
  assign n5622 = n3550 | n5621 ;
  assign n5623 = n1768 ^ n676 ^ 1'b0 ;
  assign n5624 = n5622 & ~n5623 ;
  assign n5625 = n5624 ^ n3690 ^ n2407 ;
  assign n5626 = n5625 ^ n374 ^ 1'b0 ;
  assign n5627 = n3126 & n5626 ;
  assign n5628 = n2408 & n3937 ;
  assign n5629 = n5628 ^ n2422 ^ 1'b0 ;
  assign n5630 = n2638 ^ n883 ^ 1'b0 ;
  assign n5631 = n5629 & ~n5630 ;
  assign n5632 = x32 & n329 ;
  assign n5633 = n1827 & n5632 ;
  assign n5634 = ( n1912 & ~n3705 ) | ( n1912 & n5633 ) | ( ~n3705 & n5633 ) ;
  assign n5635 = ~n1985 & n3410 ;
  assign n5636 = ~n5634 & n5635 ;
  assign n5637 = ~n5136 & n5636 ;
  assign n5638 = x30 | n1617 ;
  assign n5639 = n5638 ^ n1764 ^ 1'b0 ;
  assign n5640 = n5639 ^ n4007 ^ n973 ;
  assign n5644 = ~n1372 & n1415 ;
  assign n5645 = n5644 ^ n2921 ^ 1'b0 ;
  assign n5641 = n2819 ^ n1482 ^ n568 ;
  assign n5642 = ( n633 & n2303 ) | ( n633 & n3583 ) | ( n2303 & n3583 ) ;
  assign n5643 = n5641 & n5642 ;
  assign n5646 = n5645 ^ n5643 ^ 1'b0 ;
  assign n5647 = n5646 ^ n1666 ^ 1'b0 ;
  assign n5648 = n2240 | n2983 ;
  assign n5649 = n926 & ~n5648 ;
  assign n5650 = n1357 & n2238 ;
  assign n5651 = ~n5649 & n5650 ;
  assign n5652 = n5651 ^ n4030 ^ 1'b0 ;
  assign n5653 = n3054 & n4310 ;
  assign n5661 = n4390 | n5185 ;
  assign n5662 = n5661 ^ n1532 ^ 1'b0 ;
  assign n5654 = n808 & ~n974 ;
  assign n5655 = ~n2103 & n5654 ;
  assign n5656 = n5655 ^ n1539 ^ n1050 ;
  assign n5657 = n2184 ^ n1684 ^ 1'b0 ;
  assign n5658 = n5657 ^ n4348 ^ n886 ;
  assign n5659 = n5658 ^ n511 ^ 1'b0 ;
  assign n5660 = ( n3229 & n5656 ) | ( n3229 & ~n5659 ) | ( n5656 & ~n5659 ) ;
  assign n5663 = n5662 ^ n5660 ^ n734 ;
  assign n5666 = n3206 & n5292 ;
  assign n5664 = n3193 & n4607 ;
  assign n5665 = n2365 & ~n5664 ;
  assign n5667 = n5666 ^ n5665 ^ 1'b0 ;
  assign n5668 = n3795 & n4079 ;
  assign n5669 = n4691 ^ n1688 ^ x221 ;
  assign n5670 = n5114 | n5669 ;
  assign n5671 = n5670 ^ n662 ^ 1'b0 ;
  assign n5672 = ~n1834 & n3930 ;
  assign n5673 = n1557 & n1804 ;
  assign n5674 = n5673 ^ n1873 ^ 1'b0 ;
  assign n5675 = n1634 & n5674 ;
  assign n5676 = ~n4445 & n5675 ;
  assign n5677 = n1709 & ~n4095 ;
  assign n5680 = n3184 & n4163 ;
  assign n5678 = n1614 ^ n1267 ^ 1'b0 ;
  assign n5679 = n5678 ^ n2529 ^ n2356 ;
  assign n5681 = n5680 ^ n5679 ^ n4841 ;
  assign n5682 = n1228 & n1400 ;
  assign n5683 = ( n756 & ~n4053 ) | ( n756 & n5143 ) | ( ~n4053 & n5143 ) ;
  assign n5684 = n5683 ^ n1811 ^ 1'b0 ;
  assign n5685 = n5682 & n5684 ;
  assign n5686 = n1624 & n5685 ;
  assign n5687 = ( n1037 & n2270 ) | ( n1037 & ~n2893 ) | ( n2270 & ~n2893 ) ;
  assign n5688 = n1344 & n5687 ;
  assign n5689 = n5688 ^ n4148 ^ n3286 ;
  assign n5690 = n392 & ~n2105 ;
  assign n5691 = ~n4744 & n5690 ;
  assign n5692 = n1878 ^ n886 ^ 1'b0 ;
  assign n5693 = n5619 & ~n5692 ;
  assign n5694 = n2781 ^ n524 ^ 1'b0 ;
  assign n5695 = ( x83 & n1149 ) | ( x83 & ~n2527 ) | ( n1149 & ~n2527 ) ;
  assign n5696 = n5695 ^ n684 ^ 1'b0 ;
  assign n5697 = x210 & n5696 ;
  assign n5698 = n5694 & n5697 ;
  assign n5699 = ~n1644 & n5698 ;
  assign n5700 = n4911 ^ n3032 ^ 1'b0 ;
  assign n5701 = n5699 | n5700 ;
  assign n5702 = x3 | n2633 ;
  assign n5703 = ~n1107 & n5702 ;
  assign n5704 = n1531 ^ x84 ^ 1'b0 ;
  assign n5705 = x230 & ~n485 ;
  assign n5706 = n5704 & n5705 ;
  assign n5707 = ( x25 & ~n4557 ) | ( x25 & n5706 ) | ( ~n4557 & n5706 ) ;
  assign n5708 = n870 & n1697 ;
  assign n5709 = n5708 ^ n297 ^ 1'b0 ;
  assign n5710 = n4190 ^ n2709 ^ n2564 ;
  assign n5711 = x195 & n2276 ;
  assign n5712 = n3273 & n5711 ;
  assign n5716 = ( x236 & ~n3524 ) | ( x236 & n3559 ) | ( ~n3524 & n3559 ) ;
  assign n5714 = ~n720 & n1059 ;
  assign n5713 = n307 & n5302 ;
  assign n5715 = n5714 ^ n5713 ^ 1'b0 ;
  assign n5717 = n5716 ^ n5715 ^ 1'b0 ;
  assign n5718 = ~n2002 & n5717 ;
  assign n5719 = n5718 ^ n262 ^ 1'b0 ;
  assign n5720 = ~n5712 & n5719 ;
  assign n5721 = n1986 & n2917 ;
  assign n5722 = n3690 & n5721 ;
  assign n5723 = ( ~n1741 & n3418 ) | ( ~n1741 & n3430 ) | ( n3418 & n3430 ) ;
  assign n5724 = n1678 ^ x181 ^ 1'b0 ;
  assign n5725 = n5451 | n5724 ;
  assign n5726 = n5725 ^ n1819 ^ n898 ;
  assign n5727 = n1922 ^ x89 ^ 1'b0 ;
  assign n5728 = x142 & ~n5727 ;
  assign n5729 = n5728 ^ n2218 ^ n814 ;
  assign n5730 = ~n366 & n5729 ;
  assign n5731 = n4910 & ~n5730 ;
  assign n5732 = x116 & ~n5731 ;
  assign n5733 = n3802 & n5732 ;
  assign n5734 = n3942 ^ n322 ^ 1'b0 ;
  assign n5735 = n1912 & ~n5734 ;
  assign n5736 = ( n1641 & ~n3196 ) | ( n1641 & n5138 ) | ( ~n3196 & n5138 ) ;
  assign n5739 = n5542 ^ n1812 ^ 1'b0 ;
  assign n5737 = n1883 ^ n1261 ^ 1'b0 ;
  assign n5738 = ~n4502 & n5737 ;
  assign n5740 = n5739 ^ n5738 ^ 1'b0 ;
  assign n5741 = ( ~n777 & n5736 ) | ( ~n777 & n5740 ) | ( n5736 & n5740 ) ;
  assign n5742 = n2858 | n4890 ;
  assign n5743 = n2432 & ~n5742 ;
  assign n5744 = n5743 ^ n2201 ^ n1187 ;
  assign n5745 = x45 & n4217 ;
  assign n5746 = n5745 ^ n731 ^ 1'b0 ;
  assign n5747 = x231 & n3699 ;
  assign n5748 = n5747 ^ x244 ^ 1'b0 ;
  assign n5749 = n3178 ^ n2917 ^ n1415 ;
  assign n5750 = n4447 & ~n5749 ;
  assign n5751 = ( n626 & n733 ) | ( n626 & n1356 ) | ( n733 & n1356 ) ;
  assign n5752 = n295 & n5751 ;
  assign n5753 = ~n4048 & n5752 ;
  assign n5754 = n802 | n5753 ;
  assign n5755 = ( n280 & n864 ) | ( n280 & n914 ) | ( n864 & n914 ) ;
  assign n5756 = n4844 ^ n2299 ^ 1'b0 ;
  assign n5757 = n5755 | n5756 ;
  assign n5758 = n2263 | n5446 ;
  assign n5759 = ( x169 & n1014 ) | ( x169 & n3780 ) | ( n1014 & n3780 ) ;
  assign n5760 = ( n2411 & ~n3744 ) | ( n2411 & n5409 ) | ( ~n3744 & n5409 ) ;
  assign n5761 = n1118 | n1312 ;
  assign n5762 = n4848 & ~n5761 ;
  assign n5763 = n2380 & n5762 ;
  assign n5764 = n1030 ^ n536 ^ 1'b0 ;
  assign n5765 = ~n2014 & n5764 ;
  assign n5766 = ~n2001 & n5433 ;
  assign n5767 = x86 ^ x72 ^ 1'b0 ;
  assign n5768 = ( n3050 & n5766 ) | ( n3050 & ~n5767 ) | ( n5766 & ~n5767 ) ;
  assign n5769 = n3231 & ~n5768 ;
  assign n5770 = ~n5765 & n5769 ;
  assign n5772 = n1029 | n4268 ;
  assign n5771 = n3004 & ~n3809 ;
  assign n5773 = n5772 ^ n5771 ^ 1'b0 ;
  assign n5774 = ( n1412 & ~n2258 ) | ( n1412 & n4646 ) | ( ~n2258 & n4646 ) ;
  assign n5775 = ( x88 & x162 ) | ( x88 & ~n1075 ) | ( x162 & ~n1075 ) ;
  assign n5776 = ~n5774 & n5775 ;
  assign n5777 = n5776 ^ n1779 ^ 1'b0 ;
  assign n5778 = n4136 | n5777 ;
  assign n5779 = n2319 & ~n5778 ;
  assign n5780 = n4873 & n5779 ;
  assign n5781 = ~n2518 & n2768 ;
  assign n5782 = n2604 & ~n5781 ;
  assign n5783 = ~x133 & n5782 ;
  assign n5784 = n1251 | n1547 ;
  assign n5785 = n5784 ^ n4744 ^ x101 ;
  assign n5786 = ~n2014 & n3063 ;
  assign n5787 = ~n4076 & n5786 ;
  assign n5788 = n2201 | n5787 ;
  assign n5789 = n756 | n5788 ;
  assign n5792 = ~n863 & n5765 ;
  assign n5793 = ~n2823 & n5792 ;
  assign n5794 = ( n3368 & n3645 ) | ( n3368 & n5793 ) | ( n3645 & n5793 ) ;
  assign n5790 = n2500 & n3652 ;
  assign n5791 = n1550 & n5790 ;
  assign n5795 = n5794 ^ n5791 ^ n5627 ;
  assign n5802 = n4850 ^ n3021 ^ n841 ;
  assign n5796 = n1902 ^ n1816 ^ n1381 ;
  assign n5797 = n5796 ^ n272 ^ x29 ;
  assign n5798 = n5797 ^ n4163 ^ 1'b0 ;
  assign n5799 = n4857 | n5798 ;
  assign n5800 = n5799 ^ n3791 ^ n1578 ;
  assign n5801 = n919 & ~n5800 ;
  assign n5803 = n5802 ^ n5801 ^ 1'b0 ;
  assign n5804 = ( n262 & ~n542 ) | ( n262 & n3937 ) | ( ~n542 & n3937 ) ;
  assign n5805 = ( n257 & ~n1776 ) | ( n257 & n3449 ) | ( ~n1776 & n3449 ) ;
  assign n5806 = n3472 ^ n554 ^ 1'b0 ;
  assign n5807 = n2701 & n5806 ;
  assign n5808 = n5807 ^ n3110 ^ 1'b0 ;
  assign n5809 = ~n982 & n5808 ;
  assign n5810 = n579 & n5809 ;
  assign n5811 = n1464 & n5810 ;
  assign n5812 = ~n396 & n2685 ;
  assign n5813 = n1362 & n5812 ;
  assign n5814 = n3602 ^ n800 ^ 1'b0 ;
  assign n5815 = ~n5813 & n5814 ;
  assign n5816 = n3563 | n5815 ;
  assign n5817 = n5195 ^ n2103 ^ x80 ;
  assign n5818 = n5817 ^ n1526 ^ 1'b0 ;
  assign n5819 = n1543 & n5818 ;
  assign n5820 = ( n1366 & ~n1672 ) | ( n1366 & n5373 ) | ( ~n1672 & n5373 ) ;
  assign n5821 = n5820 ^ n5445 ^ 1'b0 ;
  assign n5822 = ~n3264 & n5821 ;
  assign n5823 = ( n2769 & n5286 ) | ( n2769 & ~n5811 ) | ( n5286 & ~n5811 ) ;
  assign n5824 = n261 | n859 ;
  assign n5825 = n1342 & ~n5824 ;
  assign n5826 = n3830 & ~n5825 ;
  assign n5827 = ( n585 & n2576 ) | ( n585 & n5826 ) | ( n2576 & n5826 ) ;
  assign n5828 = ~n2700 & n3756 ;
  assign n5829 = n4126 ^ n3066 ^ 1'b0 ;
  assign n5830 = ~n5030 & n5829 ;
  assign n5831 = n5830 ^ n5593 ^ 1'b0 ;
  assign n5832 = n5828 | n5831 ;
  assign n5833 = n5832 ^ n4051 ^ 1'b0 ;
  assign n5834 = n5833 ^ n1199 ^ n1010 ;
  assign n5837 = n2465 ^ n409 ^ 1'b0 ;
  assign n5838 = n313 & ~n5837 ;
  assign n5835 = n1391 & n2558 ;
  assign n5836 = n1356 & n5835 ;
  assign n5839 = n5838 ^ n5836 ^ n1884 ;
  assign n5840 = ( n1543 & n2455 ) | ( n1543 & ~n2638 ) | ( n2455 & ~n2638 ) ;
  assign n5841 = ~n1231 & n5840 ;
  assign n5842 = n5841 ^ n3095 ^ 1'b0 ;
  assign n5843 = n1070 & ~n2461 ;
  assign n5847 = n2019 | n3399 ;
  assign n5848 = n5847 ^ n1383 ^ 1'b0 ;
  assign n5844 = n2175 | n5665 ;
  assign n5845 = n5844 ^ n1873 ^ 1'b0 ;
  assign n5846 = n4939 & ~n5845 ;
  assign n5849 = n5848 ^ n5846 ^ n2299 ;
  assign n5850 = n2474 | n2718 ;
  assign n5851 = n5850 ^ n2241 ^ 1'b0 ;
  assign n5852 = n4077 ^ n3705 ^ 1'b0 ;
  assign n5853 = n2229 & n5852 ;
  assign n5854 = ~n3406 & n5853 ;
  assign n5855 = n1663 & n5854 ;
  assign n5856 = n1052 & ~n5855 ;
  assign n5857 = n5856 ^ x141 ^ 1'b0 ;
  assign n5860 = ( n1680 & n3070 ) | ( n1680 & ~n4396 ) | ( n3070 & ~n4396 ) ;
  assign n5861 = n5860 ^ n3682 ^ 1'b0 ;
  assign n5862 = n1959 & ~n5861 ;
  assign n5858 = n4575 ^ n1482 ^ 1'b0 ;
  assign n5859 = n3994 & n5858 ;
  assign n5863 = n5862 ^ n5859 ^ 1'b0 ;
  assign n5864 = n3155 ^ n2363 ^ x153 ;
  assign n5865 = n5864 ^ n4479 ^ 1'b0 ;
  assign n5866 = n2268 & ~n5865 ;
  assign n5869 = n3945 ^ n2201 ^ 1'b0 ;
  assign n5870 = n5869 ^ n1616 ^ 1'b0 ;
  assign n5871 = n1838 & n5870 ;
  assign n5867 = x44 & ~n3541 ;
  assign n5868 = n5867 ^ n904 ^ 1'b0 ;
  assign n5872 = n5871 ^ n5868 ^ 1'b0 ;
  assign n5873 = ~n462 & n1247 ;
  assign n5874 = n2906 ^ n2599 ^ n843 ;
  assign n5875 = n5864 & n5874 ;
  assign n5876 = ~n2531 & n5875 ;
  assign n5877 = n2760 & ~n3943 ;
  assign n5878 = ( n1451 & n5383 ) | ( n1451 & ~n5877 ) | ( n5383 & ~n5877 ) ;
  assign n5879 = n4518 | n5878 ;
  assign n5880 = n2077 ^ n1123 ^ 1'b0 ;
  assign n5881 = n5050 & ~n5880 ;
  assign n5882 = n5881 ^ n1813 ^ 1'b0 ;
  assign n5883 = n5037 | n5882 ;
  assign n5884 = n3278 | n5883 ;
  assign n5885 = ( ~n2270 & n2692 ) | ( ~n2270 & n5102 ) | ( n2692 & n5102 ) ;
  assign n5886 = n5885 ^ x85 ^ 1'b0 ;
  assign n5887 = n5507 | n5886 ;
  assign n5888 = n2623 ^ n937 ^ 1'b0 ;
  assign n5889 = n1269 & ~n5888 ;
  assign n5890 = n2016 | n2297 ;
  assign n5891 = n5890 ^ n4518 ^ 1'b0 ;
  assign n5892 = n3696 & n5891 ;
  assign n5893 = n1080 | n5892 ;
  assign n5894 = n5893 ^ n1031 ^ 1'b0 ;
  assign n5895 = n5416 ^ n2524 ^ n2057 ;
  assign n5896 = n5895 ^ n1635 ^ 1'b0 ;
  assign n5897 = n3117 & n3310 ;
  assign n5898 = n5897 ^ n3035 ^ 1'b0 ;
  assign n5899 = ~n3176 & n5898 ;
  assign n5900 = n5899 ^ n636 ^ n268 ;
  assign n5901 = n4529 ^ n3167 ^ 1'b0 ;
  assign n5902 = ( n1801 & ~n2148 ) | ( n1801 & n2846 ) | ( ~n2148 & n2846 ) ;
  assign n5903 = n5902 ^ n2399 ^ 1'b0 ;
  assign n5904 = n1174 | n1764 ;
  assign n5905 = n5904 ^ n1501 ^ 1'b0 ;
  assign n5906 = n1056 | n3100 ;
  assign n5907 = n4265 & ~n5906 ;
  assign n5908 = n5905 | n5907 ;
  assign n5909 = n5908 ^ n2450 ^ 1'b0 ;
  assign n5914 = n1315 | n1737 ;
  assign n5915 = n5540 ^ n3037 ^ n2694 ;
  assign n5916 = n5914 | n5915 ;
  assign n5912 = ~n1720 & n3915 ;
  assign n5910 = n2324 & ~n2978 ;
  assign n5911 = n2041 & ~n5910 ;
  assign n5913 = n5912 ^ n5911 ^ 1'b0 ;
  assign n5917 = n5916 ^ n5913 ^ x143 ;
  assign n5918 = ( n289 & n1654 ) | ( n289 & ~n2091 ) | ( n1654 & ~n2091 ) ;
  assign n5920 = x150 & n2291 ;
  assign n5921 = ~x208 & n5920 ;
  assign n5922 = n5921 ^ x57 ^ 1'b0 ;
  assign n5923 = n4670 & ~n5922 ;
  assign n5919 = n4967 ^ n3953 ^ n352 ;
  assign n5924 = n5923 ^ n5919 ^ n2361 ;
  assign n5925 = n5918 & ~n5924 ;
  assign n5926 = ~n4073 & n5925 ;
  assign n5927 = n1979 ^ n1225 ^ 1'b0 ;
  assign n5928 = n5926 | n5927 ;
  assign n5929 = n3364 ^ n1093 ^ 1'b0 ;
  assign n5930 = ( x8 & n5928 ) | ( x8 & n5929 ) | ( n5928 & n5929 ) ;
  assign n5931 = n4443 ^ x55 ^ 1'b0 ;
  assign n5932 = n1877 | n5568 ;
  assign n5933 = n5932 ^ n1084 ^ 1'b0 ;
  assign n5934 = ~n1752 & n5494 ;
  assign n5935 = n5933 & n5934 ;
  assign n5936 = x88 & ~n3767 ;
  assign n5937 = n5936 ^ x230 ^ 1'b0 ;
  assign n5938 = n5937 ^ n5448 ^ n3689 ;
  assign n5939 = n3151 ^ x126 ^ 1'b0 ;
  assign n5940 = ~n1176 & n5939 ;
  assign n5941 = n1796 ^ n447 ^ 1'b0 ;
  assign n5942 = n5940 & n5941 ;
  assign n5943 = x10 & n3372 ;
  assign n5944 = n1467 & n5943 ;
  assign n5945 = n5944 ^ n699 ^ n335 ;
  assign n5946 = n5945 ^ x86 ^ 1'b0 ;
  assign n5948 = n3650 ^ n2569 ^ n1053 ;
  assign n5947 = n3306 ^ n3016 ^ 1'b0 ;
  assign n5949 = n5948 ^ n5947 ^ n1850 ;
  assign n5950 = n3251 ^ n1359 ^ x10 ;
  assign n5951 = x178 & ~n510 ;
  assign n5952 = n5951 ^ n2382 ^ 1'b0 ;
  assign n5953 = ~n671 & n5952 ;
  assign n5954 = n3844 ^ n2541 ^ n1729 ;
  assign n5955 = n2388 | n5954 ;
  assign n5956 = x242 | n5955 ;
  assign n5957 = n5953 & n5956 ;
  assign n5958 = ~x38 & n5957 ;
  assign n5959 = n4723 & n5613 ;
  assign n5960 = n2325 | n5959 ;
  assign n5961 = n2730 & ~n5960 ;
  assign n5967 = n1372 ^ x68 ^ 1'b0 ;
  assign n5968 = n3073 & n5967 ;
  assign n5969 = n5968 ^ n2029 ^ n330 ;
  assign n5966 = n2723 ^ n1265 ^ n745 ;
  assign n5962 = ( n2961 & n3549 ) | ( n2961 & n4229 ) | ( n3549 & n4229 ) ;
  assign n5963 = n553 | n5962 ;
  assign n5964 = n5963 ^ n2216 ^ 1'b0 ;
  assign n5965 = n5964 ^ x12 ^ 1'b0 ;
  assign n5970 = n5969 ^ n5966 ^ n5965 ;
  assign n5971 = n4641 ^ n1406 ^ x176 ;
  assign n5972 = n5948 ^ n2104 ^ n1039 ;
  assign n5973 = ~n2657 & n3276 ;
  assign n5974 = n5972 & ~n5973 ;
  assign n5975 = n1379 | n2606 ;
  assign n5976 = n5974 | n5975 ;
  assign n5977 = n1802 | n5976 ;
  assign n5978 = ( ~n1150 & n5971 ) | ( ~n1150 & n5977 ) | ( n5971 & n5977 ) ;
  assign n5979 = ( n764 & n1104 ) | ( n764 & ~n2707 ) | ( n1104 & ~n2707 ) ;
  assign n5980 = n1532 | n5979 ;
  assign n5981 = n492 & n5980 ;
  assign n5982 = n3520 ^ n455 ^ 1'b0 ;
  assign n5983 = n3432 & n4322 ;
  assign n5986 = n3778 | n4850 ;
  assign n5987 = x252 | n5986 ;
  assign n5984 = n1405 ^ n380 ^ n280 ;
  assign n5985 = n5329 | n5984 ;
  assign n5988 = n5987 ^ n5985 ^ 1'b0 ;
  assign n5989 = n841 | n5185 ;
  assign n5990 = n5575 ^ n3526 ^ 1'b0 ;
  assign n5991 = n5990 ^ n3587 ^ n1949 ;
  assign n5992 = ( ~n1080 & n1537 ) | ( ~n1080 & n3002 ) | ( n1537 & n3002 ) ;
  assign n5993 = ~n1074 & n5992 ;
  assign n5994 = n5993 ^ n757 ^ 1'b0 ;
  assign n5995 = n5994 ^ n3645 ^ n309 ;
  assign n5996 = n5995 ^ n2132 ^ n1735 ;
  assign n5997 = n2126 ^ n1763 ^ 1'b0 ;
  assign n5998 = n1352 & n5997 ;
  assign n6002 = ( n675 & ~n1598 ) | ( n675 & n4970 ) | ( ~n1598 & n4970 ) ;
  assign n5999 = n5226 ^ n1144 ^ 1'b0 ;
  assign n6000 = n1518 & n5999 ;
  assign n6001 = ( n1003 & n4229 ) | ( n1003 & n6000 ) | ( n4229 & n6000 ) ;
  assign n6003 = n6002 ^ n6001 ^ n5702 ;
  assign n6004 = n544 & n4450 ;
  assign n6005 = n6004 ^ n4407 ^ 1'b0 ;
  assign n6006 = ~n2918 & n4852 ;
  assign n6007 = ~n4099 & n6006 ;
  assign n6008 = n6005 & n6007 ;
  assign n6009 = n814 | n4476 ;
  assign n6010 = x20 & x52 ;
  assign n6011 = ~n459 & n6010 ;
  assign n6012 = n1068 | n2899 ;
  assign n6013 = n446 | n6012 ;
  assign n6015 = n1949 | n4703 ;
  assign n6016 = n1228 & n2030 ;
  assign n6017 = ~n6015 & n6016 ;
  assign n6014 = n4423 ^ n711 ^ n528 ;
  assign n6018 = n6017 ^ n6014 ^ n3690 ;
  assign n6019 = ( ~n6011 & n6013 ) | ( ~n6011 & n6018 ) | ( n6013 & n6018 ) ;
  assign n6028 = ( ~n1053 & n2397 ) | ( ~n1053 & n5007 ) | ( n2397 & n5007 ) ;
  assign n6020 = x179 & ~n3872 ;
  assign n6021 = n6020 ^ n445 ^ 1'b0 ;
  assign n6022 = n2858 ^ n814 ^ n345 ;
  assign n6023 = n4264 ^ n3050 ^ n357 ;
  assign n6024 = n6023 ^ n3556 ^ 1'b0 ;
  assign n6025 = ~n6022 & n6024 ;
  assign n6026 = n2530 & n6025 ;
  assign n6027 = ~n6021 & n6026 ;
  assign n6029 = n6028 ^ n6027 ^ 1'b0 ;
  assign n6030 = n4882 & ~n6029 ;
  assign n6031 = n2114 ^ n1851 ^ n905 ;
  assign n6032 = n6031 ^ n5398 ^ 1'b0 ;
  assign n6034 = n378 & ~n1717 ;
  assign n6035 = n6034 ^ n1233 ^ 1'b0 ;
  assign n6033 = n976 | n3663 ;
  assign n6036 = n6035 ^ n6033 ^ 1'b0 ;
  assign n6037 = x254 & ~n6036 ;
  assign n6038 = ( n4101 & n4968 ) | ( n4101 & n6037 ) | ( n4968 & n6037 ) ;
  assign n6040 = n5488 ^ n4363 ^ 1'b0 ;
  assign n6041 = n6040 ^ n3169 ^ n2811 ;
  assign n6039 = n1063 & ~n1409 ;
  assign n6042 = n6041 ^ n6039 ^ 1'b0 ;
  assign n6043 = n6042 ^ n3632 ^ 1'b0 ;
  assign n6044 = n5794 | n6043 ;
  assign n6045 = n739 & n2255 ;
  assign n6046 = n6045 ^ n1475 ^ x49 ;
  assign n6047 = ( n1412 & n3374 ) | ( n1412 & n6046 ) | ( n3374 & n6046 ) ;
  assign n6048 = n3027 ^ n1118 ^ 1'b0 ;
  assign n6049 = n6047 & n6048 ;
  assign n6050 = n2388 ^ n715 ^ 1'b0 ;
  assign n6051 = ~n6049 & n6050 ;
  assign n6052 = n473 | n2835 ;
  assign n6053 = n2608 | n6052 ;
  assign n6054 = n4087 & n6053 ;
  assign n6055 = ~n4093 & n6054 ;
  assign n6057 = n1503 & ~n1883 ;
  assign n6058 = n6057 ^ n5507 ^ 1'b0 ;
  assign n6056 = n3643 ^ n3232 ^ 1'b0 ;
  assign n6059 = n6058 ^ n6056 ^ 1'b0 ;
  assign n6060 = ~n4410 & n6059 ;
  assign n6062 = n1714 ^ x223 ^ 1'b0 ;
  assign n6063 = n1638 & n6062 ;
  assign n6061 = x202 & n5695 ;
  assign n6064 = n6063 ^ n6061 ^ n618 ;
  assign n6065 = n1267 | n6064 ;
  assign n6066 = n4639 | n6065 ;
  assign n6067 = n2400 & n2944 ;
  assign n6068 = n6067 ^ n3368 ^ 1'b0 ;
  assign n6072 = n2569 & ~n4600 ;
  assign n6073 = n6072 ^ n2785 ^ 1'b0 ;
  assign n6069 = ~n1810 & n4856 ;
  assign n6070 = n6069 ^ n2394 ^ 1'b0 ;
  assign n6071 = n6070 ^ x130 ^ 1'b0 ;
  assign n6074 = n6073 ^ n6071 ^ 1'b0 ;
  assign n6075 = ( ~n4284 & n5091 ) | ( ~n4284 & n6074 ) | ( n5091 & n6074 ) ;
  assign n6076 = n2930 ^ n1181 ^ n376 ;
  assign n6077 = n6076 ^ n3760 ^ n2380 ;
  assign n6078 = x6 & n2585 ;
  assign n6079 = n6078 ^ n4144 ^ 1'b0 ;
  assign n6080 = n6079 ^ n5094 ^ 1'b0 ;
  assign n6081 = n1099 & ~n6080 ;
  assign n6082 = n2287 & n5683 ;
  assign n6083 = n6082 ^ n2723 ^ n1036 ;
  assign n6084 = ~n554 & n3528 ;
  assign n6085 = ~x193 & n6084 ;
  assign n6086 = n1104 | n1701 ;
  assign n6087 = n881 | n6086 ;
  assign n6088 = n2548 ^ n2057 ^ x254 ;
  assign n6089 = n6088 ^ n4841 ^ n796 ;
  assign n6090 = n6087 & n6089 ;
  assign n6091 = ~n673 & n6090 ;
  assign n6092 = ( ~n782 & n1700 ) | ( ~n782 & n3568 ) | ( n1700 & n3568 ) ;
  assign n6093 = n2745 | n3924 ;
  assign n6094 = x20 | n6093 ;
  assign n6095 = n6092 & n6094 ;
  assign n6096 = n6095 ^ n5037 ^ 1'b0 ;
  assign n6097 = n5169 ^ n2982 ^ 1'b0 ;
  assign n6098 = n4478 ^ n4041 ^ n334 ;
  assign n6099 = n6097 & ~n6098 ;
  assign n6100 = ~n3004 & n6099 ;
  assign n6101 = ( x223 & n1027 ) | ( x223 & ~n3759 ) | ( n1027 & ~n3759 ) ;
  assign n6102 = n5506 | n6101 ;
  assign n6103 = n3141 & ~n6102 ;
  assign n6104 = n3724 | n6103 ;
  assign n6105 = n6100 & ~n6104 ;
  assign n6106 = n393 & ~n843 ;
  assign n6107 = ~n1877 & n6106 ;
  assign n6108 = ( n3640 & n4526 ) | ( n3640 & ~n6107 ) | ( n4526 & ~n6107 ) ;
  assign n6109 = ( n676 & n4567 ) | ( n676 & n5219 ) | ( n4567 & n5219 ) ;
  assign n6110 = n4766 | n6109 ;
  assign n6111 = n281 & ~n1284 ;
  assign n6112 = n6110 & ~n6111 ;
  assign n6113 = n1952 & n6112 ;
  assign n6114 = ( n1201 & n2449 ) | ( n1201 & n3340 ) | ( n2449 & n3340 ) ;
  assign n6115 = n2192 | n6114 ;
  assign n6116 = n352 | n6115 ;
  assign n6117 = n6116 ^ n5367 ^ 1'b0 ;
  assign n6118 = n575 ^ x117 ^ 1'b0 ;
  assign n6119 = n5102 & ~n6118 ;
  assign n6120 = n6119 ^ n3316 ^ 1'b0 ;
  assign n6121 = n6120 ^ n5331 ^ 1'b0 ;
  assign n6122 = n1277 & n5953 ;
  assign n6123 = n2134 & n6122 ;
  assign n6124 = n3821 ^ n879 ^ 1'b0 ;
  assign n6125 = n2492 & n6124 ;
  assign n6127 = n1260 ^ n832 ^ 1'b0 ;
  assign n6128 = n669 | n6127 ;
  assign n6126 = n2408 & n4883 ;
  assign n6129 = n6128 ^ n6126 ^ 1'b0 ;
  assign n6130 = ( n940 & n1051 ) | ( n940 & ~n6129 ) | ( n1051 & ~n6129 ) ;
  assign n6131 = ( n1244 & n4862 ) | ( n1244 & n6130 ) | ( n4862 & n6130 ) ;
  assign n6132 = n6131 ^ x160 ^ 1'b0 ;
  assign n6133 = ( x53 & ~n3983 ) | ( x53 & n5682 ) | ( ~n3983 & n5682 ) ;
  assign n6134 = n307 & n6133 ;
  assign n6135 = n3425 & n6134 ;
  assign n6136 = n2782 & ~n6135 ;
  assign n6137 = x102 & n1867 ;
  assign n6138 = n6137 ^ n1630 ^ 1'b0 ;
  assign n6141 = n1837 & n2336 ;
  assign n6142 = n6141 ^ n947 ^ 1'b0 ;
  assign n6143 = n6142 ^ n2194 ^ n2100 ;
  assign n6139 = n3144 ^ n2152 ^ n1408 ;
  assign n6140 = n6139 ^ n4405 ^ 1'b0 ;
  assign n6144 = n6143 ^ n6140 ^ 1'b0 ;
  assign n6145 = n6138 & ~n6144 ;
  assign n6146 = ( n6132 & n6136 ) | ( n6132 & ~n6145 ) | ( n6136 & ~n6145 ) ;
  assign n6147 = n1650 ^ n468 ^ 1'b0 ;
  assign n6148 = ~n1590 & n6147 ;
  assign n6149 = n3066 ^ n1697 ^ n360 ;
  assign n6150 = n6149 ^ n2864 ^ n1217 ;
  assign n6151 = n6148 & ~n6150 ;
  assign n6152 = ~n5363 & n6151 ;
  assign n6153 = n6152 ^ n6005 ^ n4710 ;
  assign n6154 = ~n3913 & n6153 ;
  assign n6155 = ~n2419 & n6154 ;
  assign n6156 = n3931 ^ n3754 ^ 1'b0 ;
  assign n6157 = n2613 | n3338 ;
  assign n6158 = n459 | n6157 ;
  assign n6159 = ~n3675 & n6158 ;
  assign n6168 = ( n1641 & n2399 ) | ( n1641 & ~n4672 ) | ( n2399 & ~n4672 ) ;
  assign n6169 = n5914 | n6168 ;
  assign n6160 = n4488 ^ n2711 ^ 1'b0 ;
  assign n6161 = n6160 ^ n4090 ^ 1'b0 ;
  assign n6162 = n3253 & ~n6161 ;
  assign n6163 = ( n1254 & n2280 ) | ( n1254 & ~n6162 ) | ( n2280 & ~n6162 ) ;
  assign n6164 = n4650 ^ n2737 ^ 1'b0 ;
  assign n6165 = ~n6163 & n6164 ;
  assign n6166 = n4404 & n6165 ;
  assign n6167 = x234 & ~n6166 ;
  assign n6170 = n6169 ^ n6167 ^ 1'b0 ;
  assign n6171 = n4798 ^ x251 ^ x196 ;
  assign n6172 = n1427 & n6171 ;
  assign n6173 = n6172 ^ n1658 ^ 1'b0 ;
  assign n6174 = n6173 ^ n4086 ^ n2836 ;
  assign n6175 = n6174 ^ n5492 ^ n2757 ;
  assign n6176 = ~x174 & n728 ;
  assign n6177 = n6176 ^ n5739 ^ 1'b0 ;
  assign n6178 = n6175 | n6177 ;
  assign n6179 = n3805 ^ n2649 ^ n1963 ;
  assign n6180 = ~n1910 & n2950 ;
  assign n6181 = n6180 ^ n2571 ^ 1'b0 ;
  assign n6182 = n6181 ^ n3388 ^ 1'b0 ;
  assign n6188 = ( ~n799 & n1564 ) | ( ~n799 & n1985 ) | ( n1564 & n1985 ) ;
  assign n6189 = ~n3985 & n6188 ;
  assign n6190 = n3754 & n6189 ;
  assign n6183 = n1054 & n1169 ;
  assign n6184 = n6183 ^ n1279 ^ 1'b0 ;
  assign n6185 = n6184 ^ n2583 ^ 1'b0 ;
  assign n6186 = n414 & ~n6185 ;
  assign n6187 = ~n4185 & n6186 ;
  assign n6191 = n6190 ^ n6187 ^ 1'b0 ;
  assign n6192 = ( x40 & ~n703 ) | ( x40 & n861 ) | ( ~n703 & n861 ) ;
  assign n6193 = n6192 ^ x243 ^ 1'b0 ;
  assign n6194 = ( n4638 & n5420 ) | ( n4638 & n6193 ) | ( n5420 & n6193 ) ;
  assign n6195 = n3851 ^ n2308 ^ 1'b0 ;
  assign n6196 = ~n6194 & n6195 ;
  assign n6197 = n873 ^ n305 ^ x180 ;
  assign n6198 = n3110 & ~n5574 ;
  assign n6199 = n6197 & n6198 ;
  assign n6200 = n2541 ^ n1001 ^ 1'b0 ;
  assign n6201 = n4839 & ~n6200 ;
  assign n6202 = n526 | n1800 ;
  assign n6203 = ( n2803 & ~n4560 ) | ( n2803 & n6202 ) | ( ~n4560 & n6202 ) ;
  assign n6204 = n6074 ^ n938 ^ 1'b0 ;
  assign n6205 = n6204 ^ n1966 ^ n1650 ;
  assign n6206 = n6205 ^ n5259 ^ n2241 ;
  assign n6207 = n6206 ^ n6038 ^ n5240 ;
  assign n6217 = n1637 ^ n1634 ^ 1'b0 ;
  assign n6218 = n3247 & n6217 ;
  assign n6215 = ( ~x117 & n305 ) | ( ~x117 & n1493 ) | ( n305 & n1493 ) ;
  assign n6216 = ( x140 & ~n938 ) | ( x140 & n6215 ) | ( ~n938 & n6215 ) ;
  assign n6219 = n6218 ^ n6216 ^ 1'b0 ;
  assign n6208 = n1362 | n1864 ;
  assign n6209 = n2798 | n6208 ;
  assign n6210 = n5624 & n6209 ;
  assign n6211 = ~n1264 & n6210 ;
  assign n6212 = n4402 & ~n4812 ;
  assign n6213 = ( n1623 & n5480 ) | ( n1623 & n6212 ) | ( n5480 & n6212 ) ;
  assign n6214 = n6211 | n6213 ;
  assign n6220 = n6219 ^ n6214 ^ 1'b0 ;
  assign n6221 = n1506 & n1599 ;
  assign n6222 = n6221 ^ n3569 ^ 1'b0 ;
  assign n6223 = n4121 | n6222 ;
  assign n6224 = n1735 | n6223 ;
  assign n6225 = n3242 ^ n2217 ^ n1454 ;
  assign n6226 = n6225 ^ n6149 ^ x31 ;
  assign n6227 = ( n3724 & n6224 ) | ( n3724 & n6226 ) | ( n6224 & n6226 ) ;
  assign n6228 = n4771 ^ n3830 ^ n1691 ;
  assign n6229 = ( n954 & n3121 ) | ( n954 & n3598 ) | ( n3121 & n3598 ) ;
  assign n6230 = n3310 & ~n6229 ;
  assign n6231 = n6230 ^ n925 ^ 1'b0 ;
  assign n6232 = ~n1898 & n6231 ;
  assign n6233 = n6232 ^ n2840 ^ 1'b0 ;
  assign n6234 = n1599 & ~n4390 ;
  assign n6235 = n3557 & n6234 ;
  assign n6236 = n3032 | n6235 ;
  assign n6237 = n1284 | n6236 ;
  assign n6238 = n1882 ^ n1627 ^ x240 ;
  assign n6239 = n4636 | n6238 ;
  assign n6240 = n995 & ~n6239 ;
  assign n6241 = n6240 ^ n1750 ^ x17 ;
  assign n6242 = n4923 ^ n4815 ^ n933 ;
  assign n6243 = n2461 | n5946 ;
  assign n6244 = n5393 & ~n6243 ;
  assign n6245 = ( n5013 & n5037 ) | ( n5013 & ~n6235 ) | ( n5037 & ~n6235 ) ;
  assign n6246 = x11 & n5054 ;
  assign n6247 = ( ~n3466 & n4296 ) | ( ~n3466 & n5202 ) | ( n4296 & n5202 ) ;
  assign n6248 = n6246 | n6247 ;
  assign n6249 = x44 | n6248 ;
  assign n6250 = n3771 ^ n1813 ^ n958 ;
  assign n6251 = n1304 ^ n1136 ^ n724 ;
  assign n6252 = n6251 ^ n5162 ^ n441 ;
  assign n6253 = ( n5052 & n5695 ) | ( n5052 & ~n6252 ) | ( n5695 & ~n6252 ) ;
  assign n6254 = ( ~n1084 & n1166 ) | ( ~n1084 & n3928 ) | ( n1166 & n3928 ) ;
  assign n6255 = n1118 | n6254 ;
  assign n6256 = n2714 & ~n6255 ;
  assign n6257 = n4980 ^ n2149 ^ 1'b0 ;
  assign n6258 = n1018 & ~n6257 ;
  assign n6259 = n6258 ^ n5054 ^ 1'b0 ;
  assign n6260 = n4310 | n6259 ;
  assign n6261 = n2299 & ~n6260 ;
  assign n6262 = n6256 & n6261 ;
  assign n6263 = x75 & n4429 ;
  assign n6264 = n6263 ^ n515 ^ 1'b0 ;
  assign n6265 = n6264 ^ n4678 ^ n3425 ;
  assign n6266 = n5277 ^ n4536 ^ n1855 ;
  assign n6267 = n3607 ^ n3459 ^ 1'b0 ;
  assign n6268 = n6267 ^ n2127 ^ 1'b0 ;
  assign n6269 = n2164 & ~n6268 ;
  assign n6270 = n1372 ^ n611 ^ x254 ;
  assign n6271 = n6269 & ~n6270 ;
  assign n6272 = n4841 ^ n1961 ^ n1188 ;
  assign n6273 = n6272 ^ n5848 ^ n4444 ;
  assign n6274 = n2741 ^ n2586 ^ n2305 ;
  assign n6275 = n4264 | n6274 ;
  assign n6276 = ~n3901 & n6275 ;
  assign n6286 = n2780 ^ n1433 ^ n665 ;
  assign n6287 = ~n5774 & n6286 ;
  assign n6278 = n943 ^ x196 ^ 1'b0 ;
  assign n6279 = n305 | n6278 ;
  assign n6280 = n6279 ^ n4966 ^ 1'b0 ;
  assign n6281 = n5056 | n6280 ;
  assign n6282 = n6281 ^ n2317 ^ n1859 ;
  assign n6283 = ( n1208 & n1689 ) | ( n1208 & n5467 ) | ( n1689 & n5467 ) ;
  assign n6284 = ~n3563 & n6283 ;
  assign n6285 = n6282 & n6284 ;
  assign n6277 = n4864 ^ n2754 ^ n388 ;
  assign n6288 = n6287 ^ n6285 ^ n6277 ;
  assign n6289 = n1042 & ~n2303 ;
  assign n6290 = n2142 & n6289 ;
  assign n6291 = n1616 & ~n6290 ;
  assign n6292 = n987 ^ n796 ^ 1'b0 ;
  assign n6293 = n2291 & n6292 ;
  assign n6294 = ~n3831 & n6293 ;
  assign n6295 = x83 & ~n4004 ;
  assign n6296 = ( ~n1205 & n1607 ) | ( ~n1205 & n2566 ) | ( n1607 & n2566 ) ;
  assign n6297 = n6296 ^ n4925 ^ 1'b0 ;
  assign n6298 = n4382 | n6297 ;
  assign n6299 = n5439 | n6298 ;
  assign n6300 = n5117 ^ n3452 ^ 1'b0 ;
  assign n6301 = n3343 & ~n6300 ;
  assign n6302 = n1421 & n4664 ;
  assign n6303 = n3954 & n6302 ;
  assign n6304 = ( n417 & ~n926 ) | ( n417 & n4107 ) | ( ~n926 & n4107 ) ;
  assign n6305 = ~n3861 & n6304 ;
  assign n6306 = n2151 & n6305 ;
  assign n6307 = ( n2790 & ~n6303 ) | ( n2790 & n6306 ) | ( ~n6303 & n6306 ) ;
  assign n6308 = n6197 ^ n5557 ^ n518 ;
  assign n6309 = n5328 | n5556 ;
  assign n6310 = n6309 ^ n4185 ^ 1'b0 ;
  assign n6311 = n5078 ^ n3337 ^ n1003 ;
  assign n6312 = n6311 ^ n473 ^ 1'b0 ;
  assign n6317 = ~n374 & n2679 ;
  assign n6313 = n1664 ^ n287 ^ 1'b0 ;
  assign n6314 = n6313 ^ n2402 ^ n496 ;
  assign n6315 = n6314 ^ n4790 ^ n669 ;
  assign n6316 = ( n1268 & n2921 ) | ( n1268 & ~n6315 ) | ( n2921 & ~n6315 ) ;
  assign n6318 = n6317 ^ n6316 ^ x82 ;
  assign n6319 = n2246 ^ n768 ^ n632 ;
  assign n6320 = ( n404 & n2450 ) | ( n404 & n3830 ) | ( n2450 & n3830 ) ;
  assign n6321 = n6320 ^ n4441 ^ n346 ;
  assign n6322 = n6321 ^ n5604 ^ 1'b0 ;
  assign n6323 = ( ~n903 & n4417 ) | ( ~n903 & n5125 ) | ( n4417 & n5125 ) ;
  assign n6324 = n4889 | n6323 ;
  assign n6325 = n6322 | n6324 ;
  assign n6326 = n4750 ^ n2765 ^ n1879 ;
  assign n6327 = n2478 & ~n2716 ;
  assign n6328 = n6327 ^ n918 ^ 1'b0 ;
  assign n6329 = n6326 | n6328 ;
  assign n6330 = n3455 ^ n3328 ^ n941 ;
  assign n6331 = ( n818 & n2818 ) | ( n818 & ~n3322 ) | ( n2818 & ~n3322 ) ;
  assign n6332 = n2262 & n5244 ;
  assign n6333 = n3499 ^ n1938 ^ n967 ;
  assign n6334 = n5664 ^ n2014 ^ 1'b0 ;
  assign n6335 = n6334 ^ n2199 ^ n1484 ;
  assign n6336 = ~n6333 & n6335 ;
  assign n6337 = ( ~n3973 & n6113 ) | ( ~n3973 & n6336 ) | ( n6113 & n6336 ) ;
  assign n6338 = ( n946 & n1802 ) | ( n946 & ~n4876 ) | ( n1802 & ~n4876 ) ;
  assign n6339 = n2599 ^ n2265 ^ x96 ;
  assign n6340 = ( ~x124 & n5002 ) | ( ~x124 & n6130 ) | ( n5002 & n6130 ) ;
  assign n6341 = n6340 ^ n2319 ^ 1'b0 ;
  assign n6342 = n6341 ^ n5604 ^ n3942 ;
  assign n6343 = ~n6339 & n6342 ;
  assign n6344 = ~n6338 & n6343 ;
  assign n6345 = n6235 ^ n5162 ^ 1'b0 ;
  assign n6346 = ~n2024 & n5092 ;
  assign n6347 = n6346 ^ n2083 ^ 1'b0 ;
  assign n6348 = n5695 ^ n4589 ^ n1388 ;
  assign n6349 = ~n6347 & n6348 ;
  assign n6350 = n4196 ^ n2168 ^ 1'b0 ;
  assign n6351 = n6349 & ~n6350 ;
  assign n6352 = n3030 ^ n532 ^ 1'b0 ;
  assign n6353 = ( n1318 & n2048 ) | ( n1318 & n6352 ) | ( n2048 & n6352 ) ;
  assign n6354 = n3790 & ~n5574 ;
  assign n6355 = n6354 ^ x168 ^ 1'b0 ;
  assign n6356 = n6355 ^ n796 ^ 1'b0 ;
  assign n6357 = n6074 & ~n6356 ;
  assign n6360 = n3555 ^ n1793 ^ n374 ;
  assign n6359 = n4710 ^ n581 ^ 1'b0 ;
  assign n6358 = n4968 ^ n4575 ^ x65 ;
  assign n6361 = n6360 ^ n6359 ^ n6358 ;
  assign n6362 = n3271 ^ n3061 ^ x3 ;
  assign n6363 = n1790 | n6362 ;
  assign n6364 = n5051 | n6363 ;
  assign n6365 = n6364 ^ n2626 ^ n1297 ;
  assign n6371 = x90 & n2719 ;
  assign n6372 = n2217 & n6371 ;
  assign n6373 = ( ~n602 & n4182 ) | ( ~n602 & n6372 ) | ( n4182 & n6372 ) ;
  assign n6368 = n311 | n1506 ;
  assign n6369 = n6368 ^ n3127 ^ n1600 ;
  assign n6366 = n3455 ^ n2206 ^ 1'b0 ;
  assign n6367 = x214 & n6366 ;
  assign n6370 = n6369 ^ n6367 ^ n5433 ;
  assign n6374 = n6373 ^ n6370 ^ n3322 ;
  assign n6375 = ( n1074 & ~n1232 ) | ( n1074 & n1512 ) | ( ~n1232 & n1512 ) ;
  assign n6376 = n2697 ^ n2250 ^ n2149 ;
  assign n6377 = n6376 ^ n3491 ^ 1'b0 ;
  assign n6378 = n2559 | n5056 ;
  assign n6379 = n6377 & ~n6378 ;
  assign n6380 = ( n1208 & n1559 ) | ( n1208 & n6379 ) | ( n1559 & n6379 ) ;
  assign n6381 = ~n6375 & n6380 ;
  assign n6382 = n616 ^ x81 ^ 1'b0 ;
  assign n6383 = n600 & n1011 ;
  assign n6384 = ~n6382 & n6383 ;
  assign n6385 = n6384 ^ n2286 ^ 1'b0 ;
  assign n6386 = n737 | n6385 ;
  assign n6387 = n5322 ^ n4945 ^ n1650 ;
  assign n6388 = n6387 ^ n1924 ^ 1'b0 ;
  assign n6389 = n2723 & n3206 ;
  assign n6390 = n6389 ^ n4070 ^ 1'b0 ;
  assign n6391 = n1344 | n6390 ;
  assign n6392 = n6391 ^ x46 ^ 1'b0 ;
  assign n6393 = n2919 | n6392 ;
  assign n6394 = n6393 ^ n2771 ^ 1'b0 ;
  assign n6395 = n2812 ^ n1219 ^ n591 ;
  assign n6396 = ( ~x60 & n1067 ) | ( ~x60 & n6395 ) | ( n1067 & n6395 ) ;
  assign n6397 = n6396 ^ n4204 ^ n744 ;
  assign n6398 = ~n419 & n2408 ;
  assign n6399 = x144 | n901 ;
  assign n6400 = n6399 ^ n5953 ^ 1'b0 ;
  assign n6401 = n2954 & n6400 ;
  assign n6402 = n4389 ^ n4296 ^ n2170 ;
  assign n6403 = n2860 & n5745 ;
  assign n6404 = n6403 ^ n534 ^ 1'b0 ;
  assign n6405 = n4199 & n6404 ;
  assign n6406 = ( n528 & ~n5535 ) | ( n528 & n6367 ) | ( ~n5535 & n6367 ) ;
  assign n6407 = ~n441 & n4673 ;
  assign n6408 = n6407 ^ n2893 ^ 1'b0 ;
  assign n6409 = ( n1390 & n1526 ) | ( n1390 & n6408 ) | ( n1526 & n6408 ) ;
  assign n6410 = n290 & ~n6409 ;
  assign n6411 = ~n6406 & n6410 ;
  assign n6412 = n1421 & n5461 ;
  assign n6413 = ~n2427 & n6412 ;
  assign n6414 = n3918 ^ n2525 ^ 1'b0 ;
  assign n6415 = ( n4437 & n6413 ) | ( n4437 & n6414 ) | ( n6413 & n6414 ) ;
  assign n6416 = n6242 & ~n6415 ;
  assign n6417 = n6416 ^ x216 ^ 1'b0 ;
  assign n6426 = n1047 | n4773 ;
  assign n6418 = n408 ^ x197 ^ 1'b0 ;
  assign n6419 = ~n1748 & n6418 ;
  assign n6420 = n2017 ^ n1359 ^ x178 ;
  assign n6421 = n1130 ^ n334 ^ 1'b0 ;
  assign n6422 = ~n6420 & n6421 ;
  assign n6423 = ~n393 & n6422 ;
  assign n6424 = n6419 & ~n6423 ;
  assign n6425 = n1331 & n6424 ;
  assign n6427 = n6426 ^ n6425 ^ 1'b0 ;
  assign n6428 = ~n424 & n6336 ;
  assign n6429 = n3727 ^ n1292 ^ 1'b0 ;
  assign n6430 = n556 & n6429 ;
  assign n6431 = n6430 ^ x53 ^ 1'b0 ;
  assign n6432 = n6431 ^ n5169 ^ n3361 ;
  assign n6433 = n2909 ^ n634 ^ n594 ;
  assign n6434 = ( ~x123 & n5342 ) | ( ~x123 & n6433 ) | ( n5342 & n6433 ) ;
  assign n6435 = x149 | n4014 ;
  assign n6436 = ~n3424 & n6435 ;
  assign n6437 = ~n3514 & n6436 ;
  assign n6438 = ( n1568 & n2525 ) | ( n1568 & ~n6421 ) | ( n2525 & ~n6421 ) ;
  assign n6439 = n5202 ^ n2759 ^ 1'b0 ;
  assign n6440 = n659 & n6439 ;
  assign n6441 = n5128 ^ n3101 ^ n2574 ;
  assign n6442 = n6441 ^ n5500 ^ 1'b0 ;
  assign n6443 = n6048 ^ n4945 ^ 1'b0 ;
  assign n6444 = n6442 & ~n6443 ;
  assign n6445 = n3448 ^ n1750 ^ n452 ;
  assign n6446 = x178 & n3508 ;
  assign n6447 = ~x16 & n6446 ;
  assign n6448 = n3187 | n6447 ;
  assign n6449 = n6448 ^ n1152 ^ 1'b0 ;
  assign n6450 = n870 & ~n6449 ;
  assign n6451 = n6445 & n6450 ;
  assign n6452 = n4703 ^ n574 ^ 1'b0 ;
  assign n6453 = n2767 | n6452 ;
  assign n6454 = n1450 & ~n6453 ;
  assign n6455 = n6451 & n6454 ;
  assign n6456 = n6219 ^ n3484 ^ n3285 ;
  assign n6457 = n1497 ^ n1472 ^ 1'b0 ;
  assign n6458 = n6457 ^ n2982 ^ 1'b0 ;
  assign n6459 = n6458 ^ n3276 ^ 1'b0 ;
  assign n6463 = ( ~n1966 & n2128 ) | ( ~n1966 & n4006 ) | ( n2128 & n4006 ) ;
  assign n6464 = ( n374 & n3469 ) | ( n374 & n6463 ) | ( n3469 & n6463 ) ;
  assign n6460 = ( x125 & n1732 ) | ( x125 & n1868 ) | ( n1732 & n1868 ) ;
  assign n6461 = n6460 ^ n1312 ^ 1'b0 ;
  assign n6462 = n4959 | n6461 ;
  assign n6465 = n6464 ^ n6462 ^ 1'b0 ;
  assign n6466 = n2934 ^ n1385 ^ 1'b0 ;
  assign n6467 = n6466 ^ n468 ^ 1'b0 ;
  assign n6468 = x246 & ~n6467 ;
  assign n6469 = n2597 ^ n471 ^ 1'b0 ;
  assign n6470 = n1372 & ~n6469 ;
  assign n6471 = n3316 & ~n3383 ;
  assign n6472 = ~n1907 & n6471 ;
  assign n6473 = n6470 | n6472 ;
  assign n6474 = n6473 ^ n841 ^ n421 ;
  assign n6478 = n1337 ^ n445 ^ x251 ;
  assign n6479 = n6478 ^ n2402 ^ n1806 ;
  assign n6480 = n4917 ^ n1501 ^ x231 ;
  assign n6481 = ( n1467 & n6479 ) | ( n1467 & ~n6480 ) | ( n6479 & ~n6480 ) ;
  assign n6475 = ( n560 & n1026 ) | ( n560 & n5451 ) | ( n1026 & n5451 ) ;
  assign n6476 = n6475 ^ n3417 ^ 1'b0 ;
  assign n6477 = n1900 & ~n6476 ;
  assign n6482 = n6481 ^ n6477 ^ 1'b0 ;
  assign n6483 = ( n6468 & n6474 ) | ( n6468 & n6482 ) | ( n6474 & n6482 ) ;
  assign n6484 = n5407 & ~n6483 ;
  assign n6500 = n666 & n2657 ;
  assign n6501 = ~n3365 & n4319 ;
  assign n6502 = ( x120 & n6500 ) | ( x120 & ~n6501 ) | ( n6500 & ~n6501 ) ;
  assign n6503 = ( x150 & n586 ) | ( x150 & n1338 ) | ( n586 & n1338 ) ;
  assign n6504 = n6503 ^ n2767 ^ 1'b0 ;
  assign n6505 = n6502 & ~n6504 ;
  assign n6496 = n2340 ^ n1590 ^ 1'b0 ;
  assign n6497 = x12 & ~n6496 ;
  assign n6498 = x90 & n6497 ;
  assign n6499 = n6323 & n6498 ;
  assign n6485 = n1390 ^ n1014 ^ 1'b0 ;
  assign n6486 = ~n5604 & n6485 ;
  assign n6487 = n368 & n2547 ;
  assign n6488 = n6487 ^ n995 ^ 1'b0 ;
  assign n6489 = n6488 ^ n619 ^ 1'b0 ;
  assign n6490 = n2531 & n6489 ;
  assign n6491 = n6490 ^ n6073 ^ 1'b0 ;
  assign n6492 = n4444 & ~n6491 ;
  assign n6493 = n6414 ^ n3514 ^ n3393 ;
  assign n6494 = n6492 & n6493 ;
  assign n6495 = ~n6486 & n6494 ;
  assign n6506 = n6505 ^ n6499 ^ n6495 ;
  assign n6507 = n1268 ^ n616 ^ n414 ;
  assign n6508 = ( x154 & ~n3756 ) | ( x154 & n6507 ) | ( ~n3756 & n6507 ) ;
  assign n6509 = n4341 ^ n3998 ^ n3136 ;
  assign n6510 = ( n1752 & n3033 ) | ( n1752 & ~n3816 ) | ( n3033 & ~n3816 ) ;
  assign n6511 = n1155 | n4337 ;
  assign n6512 = n6511 ^ n3032 ^ 1'b0 ;
  assign n6513 = n2460 & ~n3264 ;
  assign n6514 = n6512 & n6513 ;
  assign n6515 = ( ~n732 & n5899 ) | ( ~n732 & n6514 ) | ( n5899 & n6514 ) ;
  assign n6519 = n3984 & n4087 ;
  assign n6520 = n1784 & n6519 ;
  assign n6516 = n2052 ^ n518 ^ 1'b0 ;
  assign n6517 = n1958 & ~n6516 ;
  assign n6518 = n891 & n6517 ;
  assign n6521 = n6520 ^ n6518 ^ n5464 ;
  assign n6522 = x154 & n2362 ;
  assign n6523 = n6522 ^ n1506 ^ 1'b0 ;
  assign n6524 = ( ~n2782 & n4476 ) | ( ~n2782 & n6523 ) | ( n4476 & n6523 ) ;
  assign n6525 = ( ~n1826 & n3840 ) | ( ~n1826 & n5610 ) | ( n3840 & n5610 ) ;
  assign n6526 = ( n1973 & n5714 ) | ( n1973 & ~n6525 ) | ( n5714 & ~n6525 ) ;
  assign n6527 = ~n2877 & n6526 ;
  assign n6528 = n1107 & n1814 ;
  assign n6529 = n3627 ^ n2476 ^ n730 ;
  assign n6530 = n6529 ^ n5669 ^ n3297 ;
  assign n6531 = n6523 ^ n2814 ^ 1'b0 ;
  assign n6532 = x187 & ~n6531 ;
  assign n6533 = ~n1576 & n6532 ;
  assign n6534 = n1950 ^ n406 ^ 1'b0 ;
  assign n6535 = ~n2665 & n6534 ;
  assign n6536 = n6533 & n6535 ;
  assign n6537 = n2339 | n2495 ;
  assign n6538 = n6537 ^ n5853 ^ 1'b0 ;
  assign n6541 = ( x3 & ~x221 ) | ( x3 & n457 ) | ( ~x221 & n457 ) ;
  assign n6540 = n1009 & n4896 ;
  assign n6539 = n2482 ^ n1317 ^ 1'b0 ;
  assign n6542 = n6541 ^ n6540 ^ n6539 ;
  assign n6543 = n6503 ^ n2705 ^ 1'b0 ;
  assign n6544 = n5110 ^ x96 ^ 1'b0 ;
  assign n6545 = n2405 | n6544 ;
  assign n6546 = ~n4023 & n4967 ;
  assign n6547 = n4756 & ~n6546 ;
  assign n6548 = n6545 & n6547 ;
  assign n6551 = ( n3289 & n3844 ) | ( n3289 & n4436 ) | ( n3844 & n4436 ) ;
  assign n6552 = n6551 ^ n1592 ^ n1035 ;
  assign n6549 = n5746 ^ n4564 ^ 1'b0 ;
  assign n6550 = n4478 | n6549 ;
  assign n6553 = n6552 ^ n6550 ^ 1'b0 ;
  assign n6554 = n3467 & n4238 ;
  assign n6555 = n6554 ^ n5084 ^ n1610 ;
  assign n6563 = n2059 ^ x176 ^ 1'b0 ;
  assign n6564 = ( n808 & n3952 ) | ( n808 & ~n6563 ) | ( n3952 & ~n6563 ) ;
  assign n6556 = n1080 | n1317 ;
  assign n6557 = n6556 ^ n2765 ^ 1'b0 ;
  assign n6558 = ~n1228 & n3289 ;
  assign n6559 = ~x81 & n6558 ;
  assign n6560 = n6559 ^ n3532 ^ 1'b0 ;
  assign n6561 = n6557 & ~n6560 ;
  assign n6562 = n6561 ^ x201 ^ 1'b0 ;
  assign n6565 = n6564 ^ n6562 ^ 1'b0 ;
  assign n6566 = x168 & n1066 ;
  assign n6567 = ( x156 & ~n544 ) | ( x156 & n2126 ) | ( ~n544 & n2126 ) ;
  assign n6568 = n6566 | n6567 ;
  assign n6569 = x104 & n3237 ;
  assign n6570 = n6569 ^ n3673 ^ 1'b0 ;
  assign n6571 = n6570 ^ n5038 ^ 1'b0 ;
  assign n6572 = n1901 & n6571 ;
  assign n6573 = n1256 & n6572 ;
  assign n6574 = n6573 ^ n1051 ^ 1'b0 ;
  assign n6575 = ( n1137 & n3148 ) | ( n1137 & ~n5176 ) | ( n3148 & ~n5176 ) ;
  assign n6576 = ~n2847 & n6575 ;
  assign n6577 = n6576 ^ n3478 ^ 1'b0 ;
  assign n6578 = n3483 & ~n5204 ;
  assign n6579 = n6578 ^ n5933 ^ 1'b0 ;
  assign n6580 = ( n477 & n791 ) | ( n477 & n6333 ) | ( n791 & n6333 ) ;
  assign n6581 = n903 & ~n6580 ;
  assign n6582 = n6581 ^ n1953 ^ 1'b0 ;
  assign n6583 = n329 & n5844 ;
  assign n6584 = n6583 ^ n1758 ^ 1'b0 ;
  assign n6585 = n2668 ^ n2607 ^ 1'b0 ;
  assign n6586 = x188 & ~n6585 ;
  assign n6587 = x165 & n3162 ;
  assign n6588 = n6587 ^ n3543 ^ 1'b0 ;
  assign n6589 = n4889 & ~n6588 ;
  assign n6590 = n2576 & n6589 ;
  assign n6591 = ~n521 & n6590 ;
  assign n6592 = n6586 & ~n6591 ;
  assign n6593 = n6592 ^ n277 ^ 1'b0 ;
  assign n6594 = ( n6582 & n6584 ) | ( n6582 & ~n6593 ) | ( n6584 & ~n6593 ) ;
  assign n6595 = n2411 ^ n1844 ^ n1639 ;
  assign n6596 = ( x185 & n5944 ) | ( x185 & ~n6595 ) | ( n5944 & ~n6595 ) ;
  assign n6597 = n1357 & n2170 ;
  assign n6598 = ( n1072 & ~n1204 ) | ( n1072 & n5357 ) | ( ~n1204 & n5357 ) ;
  assign n6599 = n6597 & n6598 ;
  assign n6606 = n2560 ^ n849 ^ x142 ;
  assign n6605 = n1768 | n5972 ;
  assign n6607 = n6606 ^ n6605 ^ 1'b0 ;
  assign n6600 = ( ~x65 & n380 ) | ( ~x65 & n3247 ) | ( n380 & n3247 ) ;
  assign n6601 = n6600 ^ n1007 ^ 1'b0 ;
  assign n6602 = x32 & ~n6601 ;
  assign n6603 = n6602 ^ x243 ^ 1'b0 ;
  assign n6604 = ~n1754 & n6603 ;
  assign n6608 = n6607 ^ n6604 ^ n4090 ;
  assign n6609 = n4105 & ~n6608 ;
  assign n6610 = n2328 & n6609 ;
  assign n6611 = ( x163 & n625 ) | ( x163 & n1785 ) | ( n625 & n1785 ) ;
  assign n6612 = n4882 ^ n849 ^ 1'b0 ;
  assign n6613 = ( n3303 & n6611 ) | ( n3303 & ~n6612 ) | ( n6611 & ~n6612 ) ;
  assign n6614 = n5082 ^ n2465 ^ 1'b0 ;
  assign n6615 = ~n4183 & n6614 ;
  assign n6616 = n1438 | n1768 ;
  assign n6617 = n3478 & ~n6616 ;
  assign n6618 = ( n554 & n977 ) | ( n554 & ~n6617 ) | ( n977 & ~n6617 ) ;
  assign n6619 = n2781 | n6618 ;
  assign n6620 = ( n3491 & n4769 ) | ( n3491 & n5032 ) | ( n4769 & n5032 ) ;
  assign n6621 = n6620 ^ n3383 ^ 1'b0 ;
  assign n6624 = n1558 & ~n2011 ;
  assign n6623 = n5416 ^ n1605 ^ n785 ;
  assign n6622 = n5357 ^ n2243 ^ 1'b0 ;
  assign n6625 = n6624 ^ n6623 ^ n6622 ;
  assign n6626 = n6625 ^ n5571 ^ n5085 ;
  assign n6627 = n6626 ^ n3393 ^ 1'b0 ;
  assign n6636 = n3594 ^ n1297 ^ 1'b0 ;
  assign n6628 = n2476 ^ n2263 ^ n2106 ;
  assign n6629 = n1232 ^ n376 ^ x69 ;
  assign n6630 = ~n2145 & n6629 ;
  assign n6631 = n6630 ^ n534 ^ 1'b0 ;
  assign n6632 = n6628 & n6631 ;
  assign n6633 = ~n1873 & n6632 ;
  assign n6634 = n6633 ^ n5301 ^ 1'b0 ;
  assign n6635 = n4070 | n6634 ;
  assign n6637 = n6636 ^ n6635 ^ 1'b0 ;
  assign n6638 = x138 & n6530 ;
  assign n6639 = n5334 & n6638 ;
  assign n6640 = n3039 ^ n1961 ^ n720 ;
  assign n6641 = ( n1181 & n1944 ) | ( n1181 & ~n6640 ) | ( n1944 & ~n6640 ) ;
  assign n6642 = n6641 ^ n5285 ^ 1'b0 ;
  assign n6643 = n4705 ^ n4540 ^ n845 ;
  assign n6644 = n633 & ~n4965 ;
  assign n6645 = n6644 ^ n3964 ^ x127 ;
  assign n6646 = n2490 ^ n1916 ^ n1768 ;
  assign n6647 = x13 & n6646 ;
  assign n6656 = ~n2952 & n4148 ;
  assign n6657 = n6656 ^ n6556 ^ 1'b0 ;
  assign n6648 = n777 | n5918 ;
  assign n6649 = ( ~n616 & n2354 ) | ( ~n616 & n6648 ) | ( n2354 & n6648 ) ;
  assign n6650 = n1671 ^ n261 ^ 1'b0 ;
  assign n6651 = n1052 & n6650 ;
  assign n6652 = ~n6649 & n6651 ;
  assign n6653 = n6652 ^ n3534 ^ 1'b0 ;
  assign n6654 = ( n1098 & ~n4268 ) | ( n1098 & n6653 ) | ( ~n4268 & n6653 ) ;
  assign n6655 = n3675 | n6654 ;
  assign n6658 = n6657 ^ n6655 ^ 1'b0 ;
  assign n6659 = ~n6647 & n6658 ;
  assign n6660 = n2455 | n2958 ;
  assign n6661 = n6421 ^ x5 ^ 1'b0 ;
  assign n6662 = x180 & ~n6661 ;
  assign n6663 = ~n1821 & n6145 ;
  assign n6664 = ~n6662 & n6663 ;
  assign n6665 = n5656 ^ n3702 ^ n1656 ;
  assign n6666 = n6665 ^ n3120 ^ n1484 ;
  assign n6667 = n6666 ^ n1916 ^ 1'b0 ;
  assign n6668 = n2256 ^ n2186 ^ 1'b0 ;
  assign n6669 = n6667 & n6668 ;
  assign n6670 = ( n4211 & ~n5173 ) | ( n4211 & n5317 ) | ( ~n5173 & n5317 ) ;
  assign n6671 = n3292 ^ n2071 ^ n1250 ;
  assign n6672 = ( n2649 & n3129 ) | ( n2649 & ~n4072 ) | ( n3129 & ~n4072 ) ;
  assign n6673 = ( n3198 & ~n6671 ) | ( n3198 & n6672 ) | ( ~n6671 & n6672 ) ;
  assign n6674 = n6673 ^ n5510 ^ n2021 ;
  assign n6675 = n3111 | n6115 ;
  assign n6676 = x200 & ~n6675 ;
  assign n6677 = n6676 ^ n5502 ^ 1'b0 ;
  assign n6678 = ~n1641 & n4728 ;
  assign n6679 = n2432 & n6678 ;
  assign n6680 = n2330 ^ n2156 ^ 1'b0 ;
  assign n6681 = ( n3673 & n5233 ) | ( n3673 & ~n6680 ) | ( n5233 & ~n6680 ) ;
  assign n6685 = n3874 ^ n2680 ^ 1'b0 ;
  assign n6686 = n6685 ^ n3524 ^ n3364 ;
  assign n6682 = ( n350 & n1627 ) | ( n350 & n2143 ) | ( n1627 & n2143 ) ;
  assign n6683 = ~n2179 & n6682 ;
  assign n6684 = ~n1502 & n6683 ;
  assign n6687 = n6686 ^ n6684 ^ 1'b0 ;
  assign n6688 = n4049 & ~n4144 ;
  assign n6689 = n698 & n6688 ;
  assign n6690 = ( ~n550 & n1174 ) | ( ~n550 & n1192 ) | ( n1174 & n1192 ) ;
  assign n6691 = n6690 ^ n3055 ^ n2180 ;
  assign n6692 = n6691 ^ n4034 ^ 1'b0 ;
  assign n6693 = ( n4864 & n6689 ) | ( n4864 & ~n6692 ) | ( n6689 & ~n6692 ) ;
  assign n6694 = ~n4986 & n6693 ;
  assign n6695 = n5969 & ~n6694 ;
  assign n6696 = n6100 ^ n3513 ^ n3393 ;
  assign n6697 = x132 | n3592 ;
  assign n6698 = ( n3281 & n5524 ) | ( n3281 & n6697 ) | ( n5524 & n6697 ) ;
  assign n6699 = n3465 ^ n3237 ^ n1521 ;
  assign n6700 = n3748 ^ n406 ^ 1'b0 ;
  assign n6701 = n3792 & n6700 ;
  assign n6702 = ~n2728 & n6701 ;
  assign n6703 = n2267 & n6702 ;
  assign n6704 = n6699 & ~n6703 ;
  assign n6705 = n6704 ^ n2977 ^ 1'b0 ;
  assign n6706 = n6705 ^ n4490 ^ 1'b0 ;
  assign n6707 = n6706 ^ n5458 ^ n3286 ;
  assign n6708 = n5889 | n6055 ;
  assign n6709 = ~n2117 & n2811 ;
  assign n6710 = n1173 & n6709 ;
  assign n6711 = n4766 | n6710 ;
  assign n6712 = n1174 & ~n6711 ;
  assign n6713 = n3274 ^ n1308 ^ 1'b0 ;
  assign n6714 = n864 & ~n6713 ;
  assign n6715 = n3413 & n6714 ;
  assign n6716 = n6712 & n6715 ;
  assign n6717 = n1354 & ~n4171 ;
  assign n6718 = n3254 & n6717 ;
  assign n6719 = ( ~n680 & n2785 ) | ( ~n680 & n6718 ) | ( n2785 & n6718 ) ;
  assign n6720 = n6719 ^ n4620 ^ n1818 ;
  assign n6721 = n6720 ^ n2187 ^ n693 ;
  assign n6722 = n4150 ^ n3667 ^ n921 ;
  assign n6723 = ( n4762 & ~n6721 ) | ( n4762 & n6722 ) | ( ~n6721 & n6722 ) ;
  assign n6724 = n5520 ^ n2322 ^ 1'b0 ;
  assign n6725 = ~n2911 & n6724 ;
  assign n6726 = x161 & ~n2514 ;
  assign n6727 = n1517 & n6726 ;
  assign n6728 = n4753 & ~n6727 ;
  assign n6729 = ~n4556 & n6728 ;
  assign n6730 = n6729 ^ n6679 ^ n5932 ;
  assign n6731 = n4112 ^ n941 ^ 1'b0 ;
  assign n6732 = ~n416 & n6731 ;
  assign n6733 = n2752 ^ n2138 ^ 1'b0 ;
  assign n6734 = n6732 & ~n6733 ;
  assign n6735 = n6264 & n6734 ;
  assign n6736 = n4583 ^ n4185 ^ n1874 ;
  assign n6737 = n3166 ^ n2330 ^ n430 ;
  assign n6738 = n3960 ^ n3365 ^ 1'b0 ;
  assign n6739 = ~n6737 & n6738 ;
  assign n6740 = n2189 & n6739 ;
  assign n6741 = n5514 ^ n1538 ^ 1'b0 ;
  assign n6742 = n6740 & n6741 ;
  assign n6743 = n2642 ^ n2281 ^ 1'b0 ;
  assign n6744 = n5560 ^ n3351 ^ 1'b0 ;
  assign n6745 = n5109 | n6744 ;
  assign n6746 = n2600 & n2878 ;
  assign n6747 = ~n1883 & n4261 ;
  assign n6748 = n6747 ^ n1683 ^ 1'b0 ;
  assign n6749 = n6748 ^ n2441 ^ 1'b0 ;
  assign n6750 = n6746 | n6749 ;
  assign n6754 = ( ~n290 & n2402 ) | ( ~n290 & n5704 ) | ( n2402 & n5704 ) ;
  assign n6751 = n3024 & n3362 ;
  assign n6752 = n642 & n6751 ;
  assign n6753 = n6752 ^ n493 ^ 1'b0 ;
  assign n6755 = n6754 ^ n6753 ^ n2794 ;
  assign n6756 = n2113 ^ n518 ^ 1'b0 ;
  assign n6757 = n6755 & n6756 ;
  assign n6758 = n3548 & ~n6681 ;
  assign n6759 = n3366 ^ n2735 ^ 1'b0 ;
  assign n6760 = n4741 ^ n3943 ^ 1'b0 ;
  assign n6761 = n3228 | n6760 ;
  assign n6764 = n3352 ^ n2356 ^ 1'b0 ;
  assign n6762 = n773 ^ n720 ^ 1'b0 ;
  assign n6763 = n3898 & n6762 ;
  assign n6765 = n6764 ^ n6763 ^ n1189 ;
  assign n6766 = n6765 ^ n1634 ^ n1192 ;
  assign n6767 = n6766 ^ n3855 ^ n3602 ;
  assign n6769 = ~n891 & n1928 ;
  assign n6770 = ~n1710 & n6769 ;
  assign n6771 = ( n2512 & n3126 ) | ( n2512 & ~n4961 ) | ( n3126 & ~n4961 ) ;
  assign n6772 = x122 & ~n3607 ;
  assign n6773 = ~n6771 & n6772 ;
  assign n6774 = n6773 ^ n3754 ^ n2078 ;
  assign n6775 = n421 | n1511 ;
  assign n6776 = n2977 | n6775 ;
  assign n6777 = ( n2946 & n6774 ) | ( n2946 & n6776 ) | ( n6774 & n6776 ) ;
  assign n6778 = ( x96 & n1505 ) | ( x96 & n4163 ) | ( n1505 & n4163 ) ;
  assign n6779 = n6777 & n6778 ;
  assign n6780 = n6770 & n6779 ;
  assign n6768 = n676 & n4156 ;
  assign n6781 = n6780 ^ n6768 ^ 1'b0 ;
  assign n6782 = n2995 | n4594 ;
  assign n6783 = n5846 ^ n3556 ^ 1'b0 ;
  assign n6784 = n3155 & ~n6783 ;
  assign n6785 = n2203 ^ n2113 ^ n1444 ;
  assign n6786 = n6785 ^ n2100 ^ n716 ;
  assign n6787 = ( n2422 & ~n4970 ) | ( n2422 & n5138 ) | ( ~n4970 & n5138 ) ;
  assign n6788 = ( n2356 & n3645 ) | ( n2356 & n3792 ) | ( n3645 & n3792 ) ;
  assign n6789 = n6788 ^ n5557 ^ n3315 ;
  assign n6790 = n615 | n6789 ;
  assign n6791 = n6790 ^ n6752 ^ 1'b0 ;
  assign n6792 = ( n1372 & ~n5602 ) | ( n1372 & n6791 ) | ( ~n5602 & n6791 ) ;
  assign n6797 = n4540 ^ n3465 ^ n2927 ;
  assign n6793 = n995 ^ x251 ^ x150 ;
  assign n6794 = n5488 & ~n6793 ;
  assign n6795 = n5210 & n6794 ;
  assign n6796 = n6795 ^ n4732 ^ n2351 ;
  assign n6798 = n6797 ^ n6796 ^ n5517 ;
  assign n6799 = ( x180 & n2867 ) | ( x180 & n6798 ) | ( n2867 & n6798 ) ;
  assign n6800 = n2881 & ~n4359 ;
  assign n6801 = n3205 ^ n2974 ^ 1'b0 ;
  assign n6802 = ~n4183 & n6801 ;
  assign n6803 = n6802 ^ x162 ^ 1'b0 ;
  assign n6804 = ( n348 & n642 ) | ( n348 & ~n1555 ) | ( n642 & ~n1555 ) ;
  assign n6805 = n6804 ^ n3251 ^ 1'b0 ;
  assign n6806 = n6805 ^ n2022 ^ n1047 ;
  assign n6807 = n6486 ^ n5910 ^ 1'b0 ;
  assign n6808 = n6807 ^ n1676 ^ 1'b0 ;
  assign n6809 = ( x229 & ~n2519 ) | ( x229 & n4465 ) | ( ~n2519 & n4465 ) ;
  assign n6810 = n4427 | n6809 ;
  assign n6811 = n4427 & ~n6810 ;
  assign n6812 = ( n1390 & n1944 ) | ( n1390 & ~n2567 ) | ( n1944 & ~n2567 ) ;
  assign n6813 = n6503 ^ n3048 ^ 1'b0 ;
  assign n6814 = n1655 | n6813 ;
  assign n6815 = ( n1763 & n5128 ) | ( n1763 & ~n6814 ) | ( n5128 & ~n6814 ) ;
  assign n6816 = n533 & ~n1297 ;
  assign n6817 = n6816 ^ x180 ^ 1'b0 ;
  assign n6818 = n6815 & n6817 ;
  assign n6819 = n6812 & n6818 ;
  assign n6820 = ~n5524 & n6819 ;
  assign n6822 = n1128 | n1388 ;
  assign n6823 = n6822 ^ n1574 ^ 1'b0 ;
  assign n6821 = n2643 ^ x19 ^ 1'b0 ;
  assign n6824 = n6823 ^ n6821 ^ n2502 ;
  assign n6825 = ~n3198 & n5573 ;
  assign n6826 = ( n1318 & n1538 ) | ( n1318 & ~n2838 ) | ( n1538 & ~n2838 ) ;
  assign n6827 = n1196 & ~n5229 ;
  assign n6828 = ~n6826 & n6827 ;
  assign n6829 = n6828 ^ n1563 ^ n725 ;
  assign n6830 = n4567 ^ n3965 ^ 1'b0 ;
  assign n6831 = ~n4779 & n6830 ;
  assign n6832 = n4085 ^ n2149 ^ n1911 ;
  assign n6833 = n6832 ^ n6130 ^ n1188 ;
  assign n6835 = n5169 ^ n2361 ^ 1'b0 ;
  assign n6836 = n6835 ^ n3557 ^ 1'b0 ;
  assign n6837 = x125 & ~n6836 ;
  assign n6834 = n1192 & ~n1388 ;
  assign n6838 = n6837 ^ n6834 ^ 1'b0 ;
  assign n6839 = x227 & n3730 ;
  assign n6840 = n4310 & n6839 ;
  assign n6841 = n6840 ^ n3694 ^ 1'b0 ;
  assign n6848 = n1556 & n2530 ;
  assign n6842 = n2619 ^ n1818 ^ 1'b0 ;
  assign n6843 = ~n3667 & n6842 ;
  assign n6844 = n6843 ^ n2164 ^ 1'b0 ;
  assign n6845 = n6844 ^ n5364 ^ 1'b0 ;
  assign n6846 = n4605 & ~n6845 ;
  assign n6847 = ( n1958 & ~n3306 ) | ( n1958 & n6846 ) | ( ~n3306 & n6846 ) ;
  assign n6849 = n6848 ^ n6847 ^ n321 ;
  assign n6850 = ~n1894 & n5688 ;
  assign n6856 = n826 & ~n2499 ;
  assign n6851 = n3587 ^ n1743 ^ 1'b0 ;
  assign n6852 = ( n4429 & n5223 ) | ( n4429 & n6851 ) | ( n5223 & n6851 ) ;
  assign n6853 = n2741 ^ n2355 ^ x22 ;
  assign n6854 = n6853 ^ n1252 ^ n295 ;
  assign n6855 = n6852 & ~n6854 ;
  assign n6857 = n6856 ^ n6855 ^ 1'b0 ;
  assign n6858 = n6857 ^ n938 ^ 1'b0 ;
  assign n6859 = n1301 | n4465 ;
  assign n6861 = ~n1158 & n2343 ;
  assign n6862 = n6861 ^ n660 ^ 1'b0 ;
  assign n6863 = n6862 ^ n5008 ^ n4199 ;
  assign n6860 = n331 & ~n5051 ;
  assign n6864 = n6863 ^ n6860 ^ n5082 ;
  assign n6865 = ( ~n1184 & n6611 ) | ( ~n1184 & n6864 ) | ( n6611 & n6864 ) ;
  assign n6866 = n1944 & ~n3156 ;
  assign n6867 = n3324 & ~n6449 ;
  assign n6868 = ~n987 & n6867 ;
  assign n6869 = n6868 ^ n2136 ^ 1'b0 ;
  assign n6870 = ~n6866 & n6869 ;
  assign n6871 = ( ~n6859 & n6865 ) | ( ~n6859 & n6870 ) | ( n6865 & n6870 ) ;
  assign n6872 = n1619 & ~n4337 ;
  assign n6875 = n713 | n1806 ;
  assign n6876 = ( n1588 & ~n3062 ) | ( n1588 & n6875 ) | ( ~n3062 & n6875 ) ;
  assign n6873 = ( n895 & ~n1270 ) | ( n895 & n4692 ) | ( ~n1270 & n4692 ) ;
  assign n6874 = n3648 & n6873 ;
  assign n6877 = n6876 ^ n6874 ^ 1'b0 ;
  assign n6878 = n6843 & ~n6877 ;
  assign n6879 = ( ~n3231 & n6872 ) | ( ~n3231 & n6878 ) | ( n6872 & n6878 ) ;
  assign n6880 = ~n602 & n2152 ;
  assign n6881 = n6880 ^ n3717 ^ 1'b0 ;
  assign n6882 = n1072 & ~n3019 ;
  assign n6883 = n4785 & n6882 ;
  assign n6884 = ( n1050 & n2236 ) | ( n1050 & n3939 ) | ( n2236 & n3939 ) ;
  assign n6885 = n6884 ^ n3578 ^ 1'b0 ;
  assign n6886 = ~n5270 & n6885 ;
  assign n6887 = n3783 & ~n6886 ;
  assign n6888 = ~n3467 & n5295 ;
  assign n6889 = n6888 ^ n3518 ^ 1'b0 ;
  assign n6890 = n3680 & n6889 ;
  assign n6891 = n6887 & n6890 ;
  assign n6892 = n6883 | n6891 ;
  assign n6893 = n6881 & ~n6892 ;
  assign n6894 = n5751 ^ n2519 ^ 1'b0 ;
  assign n6895 = n2256 & n6894 ;
  assign n6896 = n735 & n2065 ;
  assign n6897 = n2743 & n6896 ;
  assign n6898 = ~n3281 & n3798 ;
  assign n6899 = n6897 & n6898 ;
  assign n6900 = n6899 ^ n1348 ^ 1'b0 ;
  assign n6901 = n6895 & n6900 ;
  assign n6902 = n6901 ^ n4902 ^ 1'b0 ;
  assign n6903 = ~n4589 & n6902 ;
  assign n6904 = n6313 ^ n1672 ^ 1'b0 ;
  assign n6905 = ( ~n417 & n4975 ) | ( ~n417 & n6904 ) | ( n4975 & n6904 ) ;
  assign n6906 = ~n1671 & n4186 ;
  assign n6907 = n5707 | n6906 ;
  assign n6908 = x49 & ~n6558 ;
  assign n6911 = n3799 ^ n2864 ^ 1'b0 ;
  assign n6909 = n2333 ^ n2132 ^ 1'b0 ;
  assign n6910 = n6909 ^ n6612 ^ n2030 ;
  assign n6912 = n6911 ^ n6910 ^ 1'b0 ;
  assign n6914 = ( n558 & ~n2588 ) | ( n558 & n2840 ) | ( ~n2588 & n2840 ) ;
  assign n6913 = ( x184 & n2503 ) | ( x184 & ~n3857 ) | ( n2503 & ~n3857 ) ;
  assign n6915 = n6914 ^ n6913 ^ 1'b0 ;
  assign n6917 = ( ~n669 & n1130 ) | ( ~n669 & n1652 ) | ( n1130 & n1652 ) ;
  assign n6916 = n722 | n764 ;
  assign n6918 = n6917 ^ n6916 ^ 1'b0 ;
  assign n6919 = ( x181 & ~n838 ) | ( x181 & n6918 ) | ( ~n838 & n6918 ) ;
  assign n6920 = n4459 & ~n5380 ;
  assign n6921 = ~n4302 & n6920 ;
  assign n6922 = x92 & ~n6921 ;
  assign n6923 = n4480 & n6922 ;
  assign n6924 = n6923 ^ n6434 ^ n4870 ;
  assign n6925 = n1998 | n6924 ;
  assign n6926 = ~n462 & n1140 ;
  assign n6927 = n6926 ^ x243 ^ 1'b0 ;
  assign n6928 = n768 | n6927 ;
  assign n6929 = n6928 ^ n6228 ^ 1'b0 ;
  assign n6930 = n5137 & n6929 ;
  assign n6931 = n2238 ^ n1505 ^ n1267 ;
  assign n6932 = n1458 & ~n4634 ;
  assign n6933 = n6931 & n6932 ;
  assign n6934 = n1622 ^ n1120 ^ 1'b0 ;
  assign n6935 = ( n1675 & ~n6317 ) | ( n1675 & n6934 ) | ( ~n6317 & n6934 ) ;
  assign n6936 = ( n4498 & ~n4558 ) | ( n4498 & n6935 ) | ( ~n4558 & n6935 ) ;
  assign n6937 = n6936 ^ n2106 ^ 1'b0 ;
  assign n6938 = n6492 ^ n3334 ^ 1'b0 ;
  assign n6939 = ( n1348 & ~n1840 ) | ( n1348 & n6938 ) | ( ~n1840 & n6938 ) ;
  assign n6940 = ( n1390 & ~n2746 ) | ( n1390 & n6939 ) | ( ~n2746 & n6939 ) ;
  assign n6941 = ( n271 & n1601 ) | ( n271 & ~n2299 ) | ( n1601 & ~n2299 ) ;
  assign n6942 = n5102 ^ n481 ^ n470 ;
  assign n6943 = ( n5281 & n6941 ) | ( n5281 & n6942 ) | ( n6941 & n6942 ) ;
  assign n6944 = n426 & n1165 ;
  assign n6945 = ~n2411 & n6944 ;
  assign n6946 = n6945 ^ x18 ^ 1'b0 ;
  assign n6947 = n2558 & ~n6946 ;
  assign n6948 = n2438 & ~n4455 ;
  assign n6949 = ~n6947 & n6948 ;
  assign n6950 = n1208 & ~n4970 ;
  assign n6951 = n3144 & n3805 ;
  assign n6952 = n6950 & n6951 ;
  assign n6953 = n3974 ^ n1068 ^ 1'b0 ;
  assign n6954 = n954 | n6953 ;
  assign n6955 = n2240 | n6310 ;
  assign n6956 = ( n4109 & n6164 ) | ( n4109 & n6955 ) | ( n6164 & n6955 ) ;
  assign n6957 = n272 | n2522 ;
  assign n6958 = n3170 & ~n6957 ;
  assign n6960 = ( ~n421 & n1202 ) | ( ~n421 & n2731 ) | ( n1202 & n2731 ) ;
  assign n6961 = n3406 | n6960 ;
  assign n6962 = n1533 | n6961 ;
  assign n6963 = n6962 ^ x224 ^ 1'b0 ;
  assign n6959 = n5169 ^ n4204 ^ x203 ;
  assign n6964 = n6963 ^ n6959 ^ n3195 ;
  assign n6965 = n855 & ~n6964 ;
  assign n6966 = n6958 & n6965 ;
  assign n6967 = n284 & n2580 ;
  assign n6968 = n3448 & ~n6967 ;
  assign n6969 = ~n4577 & n6968 ;
  assign n6970 = n6868 | n6969 ;
  assign n6971 = n2746 & ~n6970 ;
  assign n6972 = n6971 ^ n5637 ^ 1'b0 ;
  assign n6973 = ~n6966 & n6972 ;
  assign n6975 = n2434 & ~n6873 ;
  assign n6976 = n6975 ^ n6945 ^ 1'b0 ;
  assign n6974 = x220 & n2595 ;
  assign n6977 = n6976 ^ n6974 ^ n4910 ;
  assign n6978 = n4570 ^ n3223 ^ n2419 ;
  assign n6979 = n4889 & ~n5522 ;
  assign n6980 = n3483 & n6979 ;
  assign n6981 = n6980 ^ n1776 ^ 1'b0 ;
  assign n6982 = n3846 ^ n3010 ^ n1192 ;
  assign n6983 = ( x158 & ~n2448 ) | ( x158 & n6982 ) | ( ~n2448 & n6982 ) ;
  assign n6984 = n2272 & ~n5805 ;
  assign n6985 = n6274 ^ n3619 ^ n1194 ;
  assign n6986 = n5807 | n6985 ;
  assign n6987 = n4224 & n6986 ;
  assign n6988 = ~n4877 & n6987 ;
  assign n6989 = n4346 ^ n998 ^ 1'b0 ;
  assign n6993 = n1270 & n4908 ;
  assign n6994 = ~n3790 & n6993 ;
  assign n6990 = ( x198 & ~n1727 ) | ( x198 & n2774 ) | ( ~n1727 & n2774 ) ;
  assign n6991 = n6990 ^ n3702 ^ 1'b0 ;
  assign n6992 = n6991 ^ n3607 ^ n2052 ;
  assign n6995 = n6994 ^ n6992 ^ n6345 ;
  assign n6999 = ( ~x69 & n490 ) | ( ~x69 & n1437 ) | ( n490 & n1437 ) ;
  assign n7000 = ( ~n863 & n2793 ) | ( ~n863 & n6999 ) | ( n2793 & n6999 ) ;
  assign n6996 = n2289 ^ x182 ^ 1'b0 ;
  assign n6997 = n6996 ^ n1727 ^ 1'b0 ;
  assign n6998 = n1798 & ~n6997 ;
  assign n7001 = n7000 ^ n6998 ^ n1124 ;
  assign n7002 = ~n421 & n6056 ;
  assign n7003 = n7002 ^ n5234 ^ 1'b0 ;
  assign n7004 = ~n2564 & n4332 ;
  assign n7005 = n291 & n2950 ;
  assign n7006 = ~n1913 & n7005 ;
  assign n7007 = ~n3523 & n6720 ;
  assign n7008 = n7007 ^ n5392 ^ 1'b0 ;
  assign n7009 = ~n7006 & n7008 ;
  assign n7014 = n2967 ^ n2011 ^ n789 ;
  assign n7010 = n1070 ^ x246 ^ 1'b0 ;
  assign n7011 = n436 & ~n7010 ;
  assign n7012 = n7011 ^ n4997 ^ n2673 ;
  assign n7013 = ( ~n4030 & n6107 ) | ( ~n4030 & n7012 ) | ( n6107 & n7012 ) ;
  assign n7015 = n7014 ^ n7013 ^ 1'b0 ;
  assign n7016 = n7015 ^ x152 ^ 1'b0 ;
  assign n7017 = n5678 ^ n3484 ^ n1320 ;
  assign n7019 = x226 | n1297 ;
  assign n7020 = ~n3257 & n7019 ;
  assign n7018 = n5225 ^ n4644 ^ n1130 ;
  assign n7021 = n7020 ^ n7018 ^ x182 ;
  assign n7022 = n3488 ^ n2504 ^ 1'b0 ;
  assign n7023 = ~n6482 & n7022 ;
  assign n7024 = n5395 ^ n3623 ^ n585 ;
  assign n7025 = n5140 ^ n725 ^ 1'b0 ;
  assign n7026 = n5456 ^ n4796 ^ n3223 ;
  assign n7027 = n2398 ^ n2305 ^ 1'b0 ;
  assign n7028 = n7027 ^ n3744 ^ n409 ;
  assign n7029 = n6135 & n7028 ;
  assign n7030 = ( n1769 & ~n3135 ) | ( n1769 & n3157 ) | ( ~n3135 & n3157 ) ;
  assign n7031 = n1935 & ~n7030 ;
  assign n7032 = ~n1640 & n6233 ;
  assign n7033 = n2655 & n3874 ;
  assign n7034 = ~x49 & n7033 ;
  assign n7035 = n2357 | n5129 ;
  assign n7036 = n7034 & ~n7035 ;
  assign n7037 = n4014 | n7036 ;
  assign n7038 = n7037 ^ n6555 ^ 1'b0 ;
  assign n7039 = n6580 ^ n3831 ^ n3107 ;
  assign n7040 = n7038 & ~n7039 ;
  assign n7041 = n6831 ^ n4942 ^ 1'b0 ;
  assign n7042 = n2001 | n7041 ;
  assign n7046 = n4296 ^ n2523 ^ 1'b0 ;
  assign n7043 = n2586 ^ n1841 ^ x231 ;
  assign n7044 = n7043 ^ n3601 ^ n780 ;
  assign n7045 = n5384 & ~n7044 ;
  assign n7047 = n7046 ^ n7045 ^ 1'b0 ;
  assign n7048 = n4156 & ~n7047 ;
  assign n7050 = n4540 ^ n2770 ^ n2415 ;
  assign n7049 = n3500 ^ n1683 ^ x161 ;
  assign n7051 = n7050 ^ n7049 ^ n6492 ;
  assign n7052 = ( n4724 & n6525 ) | ( n4724 & ~n6580 ) | ( n6525 & ~n6580 ) ;
  assign n7059 = n551 & ~n1022 ;
  assign n7060 = n7059 ^ n1035 ^ 1'b0 ;
  assign n7061 = n7060 ^ n3745 ^ x154 ;
  assign n7053 = ( x3 & n3345 ) | ( x3 & n3546 ) | ( n3345 & n3546 ) ;
  assign n7054 = ~n2514 & n6441 ;
  assign n7055 = n2315 & n7054 ;
  assign n7056 = n1674 ^ n673 ^ 1'b0 ;
  assign n7057 = ~n7055 & n7056 ;
  assign n7058 = ( n4068 & n7053 ) | ( n4068 & ~n7057 ) | ( n7053 & ~n7057 ) ;
  assign n7062 = n7061 ^ n7058 ^ 1'b0 ;
  assign n7063 = n3763 ^ n1175 ^ 1'b0 ;
  assign n7066 = n6111 ^ n5322 ^ 1'b0 ;
  assign n7067 = n6320 & n7066 ;
  assign n7068 = ( n827 & ~n1425 ) | ( n827 & n6856 ) | ( ~n1425 & n6856 ) ;
  assign n7069 = ( n5146 & n7067 ) | ( n5146 & n7068 ) | ( n7067 & n7068 ) ;
  assign n7064 = n2997 ^ n2870 ^ n853 ;
  assign n7065 = n4939 & n7064 ;
  assign n7070 = n7069 ^ n7065 ^ 1'b0 ;
  assign n7071 = n7070 ^ n4825 ^ 1'b0 ;
  assign n7072 = n1034 & n2662 ;
  assign n7073 = n7072 ^ n6657 ^ 1'b0 ;
  assign n7074 = n6274 ^ n1861 ^ 1'b0 ;
  assign n7075 = ~n5877 & n7074 ;
  assign n7078 = n499 & ~n3607 ;
  assign n7079 = n7078 ^ n6999 ^ 1'b0 ;
  assign n7076 = n6087 ^ n4083 ^ n337 ;
  assign n7077 = n5622 & ~n7076 ;
  assign n7080 = n7079 ^ n7077 ^ 1'b0 ;
  assign n7081 = ~n2956 & n4446 ;
  assign n7083 = ~n329 & n1114 ;
  assign n7084 = n7083 ^ n2414 ^ n526 ;
  assign n7085 = n7084 ^ n6483 ^ 1'b0 ;
  assign n7082 = n1109 & n2865 ;
  assign n7086 = n7085 ^ n7082 ^ 1'b0 ;
  assign n7087 = n663 & ~n6015 ;
  assign n7088 = n1352 | n1846 ;
  assign n7089 = ( n2696 & n7087 ) | ( n2696 & ~n7088 ) | ( n7087 & ~n7088 ) ;
  assign n7090 = n7089 ^ n5849 ^ 1'b0 ;
  assign n7091 = n1461 & ~n7090 ;
  assign n7092 = n7091 ^ n2280 ^ 1'b0 ;
  assign n7095 = n1843 ^ n1118 ^ 1'b0 ;
  assign n7093 = ~n3546 & n6641 ;
  assign n7094 = n7093 ^ n1001 ^ 1'b0 ;
  assign n7096 = n7095 ^ n7094 ^ 1'b0 ;
  assign n7097 = n2748 ^ n910 ^ 1'b0 ;
  assign n7098 = n7097 ^ n3998 ^ n1447 ;
  assign n7099 = ( ~n3377 & n6338 ) | ( ~n3377 & n6766 ) | ( n6338 & n6766 ) ;
  assign n7100 = n5869 & ~n5905 ;
  assign n7101 = ~n6518 & n7100 ;
  assign n7102 = n966 & ~n2128 ;
  assign n7103 = n2754 & ~n7102 ;
  assign n7104 = ~n2745 & n5378 ;
  assign n7105 = n3049 & ~n4732 ;
  assign n7106 = n7104 & n7105 ;
  assign n7107 = ~n523 & n7106 ;
  assign n7108 = n4793 ^ n3160 ^ n2583 ;
  assign n7109 = ~n1150 & n7108 ;
  assign n7110 = n7109 ^ n2545 ^ 1'b0 ;
  assign n7111 = n5367 & ~n7110 ;
  assign n7112 = n5296 & n7111 ;
  assign n7114 = n3180 ^ n2629 ^ 1'b0 ;
  assign n7115 = n430 | n7114 ;
  assign n7113 = n2389 & ~n4345 ;
  assign n7116 = n7115 ^ n7113 ^ x147 ;
  assign n7117 = ( ~n5138 & n6015 ) | ( ~n5138 & n7116 ) | ( n6015 & n7116 ) ;
  assign n7118 = n4733 ^ n3750 ^ n348 ;
  assign n7119 = ~n5037 & n5720 ;
  assign n7121 = n1547 | n1909 ;
  assign n7120 = n4329 ^ n2001 ^ 1'b0 ;
  assign n7122 = n7121 ^ n7120 ^ 1'b0 ;
  assign n7123 = n6347 ^ n4609 ^ x77 ;
  assign n7124 = n2339 | n3613 ;
  assign n7125 = n7124 ^ n2134 ^ 1'b0 ;
  assign n7126 = n7125 ^ n1179 ^ 1'b0 ;
  assign n7127 = x215 & ~n4756 ;
  assign n7128 = n4639 & ~n7127 ;
  assign n7129 = ( n2785 & n7126 ) | ( n2785 & ~n7128 ) | ( n7126 & ~n7128 ) ;
  assign n7130 = n3717 & n5659 ;
  assign n7131 = n2479 | n5816 ;
  assign n7132 = ~n334 & n4547 ;
  assign n7133 = n7132 ^ n1986 ^ 1'b0 ;
  assign n7134 = n5775 ^ x156 ^ 1'b0 ;
  assign n7135 = n2981 ^ n2655 ^ 1'b0 ;
  assign n7136 = n7135 ^ n1437 ^ x251 ;
  assign n7138 = ~n3198 & n3292 ;
  assign n7139 = ~n2723 & n5560 ;
  assign n7140 = ( n1114 & ~n7138 ) | ( n1114 & n7139 ) | ( ~n7138 & n7139 ) ;
  assign n7137 = n1776 | n3177 ;
  assign n7141 = n7140 ^ n7137 ^ 1'b0 ;
  assign n7142 = ( n3679 & n5089 ) | ( n3679 & ~n7141 ) | ( n5089 & ~n7141 ) ;
  assign n7143 = n3691 ^ n894 ^ 1'b0 ;
  assign n7144 = n327 & ~n7143 ;
  assign n7145 = ~n2189 & n7144 ;
  assign n7146 = n7145 ^ n4811 ^ n2409 ;
  assign n7147 = n6501 | n7146 ;
  assign n7148 = n7147 ^ x44 ^ 1'b0 ;
  assign n7149 = ( n910 & n4215 ) | ( n910 & ~n5340 ) | ( n4215 & ~n5340 ) ;
  assign n7150 = n4473 | n4872 ;
  assign n7151 = n7150 ^ n4777 ^ 1'b0 ;
  assign n7154 = n2633 | n3535 ;
  assign n7152 = n5622 ^ n1791 ^ n1573 ;
  assign n7153 = n5492 | n7152 ;
  assign n7155 = n7154 ^ n7153 ^ 1'b0 ;
  assign n7156 = n7151 & ~n7155 ;
  assign n7158 = n2724 ^ n1768 ^ 1'b0 ;
  assign n7157 = n6941 ^ n830 ^ n473 ;
  assign n7159 = n7158 ^ n7157 ^ n2641 ;
  assign n7160 = n6495 | n6562 ;
  assign n7165 = n3157 ^ n1232 ^ n1030 ;
  assign n7162 = n1485 | n2592 ;
  assign n7163 = n2846 & ~n7162 ;
  assign n7164 = n7163 ^ n3862 ^ n2390 ;
  assign n7166 = n7165 ^ n7164 ^ n1011 ;
  assign n7161 = ( x6 & n2043 ) | ( x6 & n2353 ) | ( n2043 & n2353 ) ;
  assign n7167 = n7166 ^ n7161 ^ n4282 ;
  assign n7168 = n7160 & n7167 ;
  assign n7169 = n1861 ^ x169 ^ 1'b0 ;
  assign n7170 = n3422 ^ n2547 ^ n980 ;
  assign n7171 = n741 & n6304 ;
  assign n7172 = n7171 ^ n449 ^ 1'b0 ;
  assign n7173 = ( n7169 & n7170 ) | ( n7169 & n7172 ) | ( n7170 & n7172 ) ;
  assign n7174 = n7173 ^ n3138 ^ 1'b0 ;
  assign n7175 = n1214 & ~n5556 ;
  assign n7176 = n734 & n7175 ;
  assign n7177 = n2220 ^ n2036 ^ 1'b0 ;
  assign n7178 = ~n6322 & n7177 ;
  assign n7179 = n7178 ^ n2051 ^ 1'b0 ;
  assign n7180 = ~n5532 & n7179 ;
  assign n7181 = n4730 ^ n1616 ^ 1'b0 ;
  assign n7189 = ( n544 & ~n1108 ) | ( n544 & n4553 ) | ( ~n1108 & n4553 ) ;
  assign n7182 = n4705 ^ n2822 ^ 1'b0 ;
  assign n7183 = n7182 ^ n683 ^ 1'b0 ;
  assign n7184 = ( n3413 & n3787 ) | ( n3413 & ~n3818 ) | ( n3787 & ~n3818 ) ;
  assign n7185 = ( ~n1328 & n2782 ) | ( ~n1328 & n7184 ) | ( n2782 & n7184 ) ;
  assign n7186 = n7161 & ~n7185 ;
  assign n7187 = n7186 ^ n4355 ^ 1'b0 ;
  assign n7188 = n7183 | n7187 ;
  assign n7190 = n7189 ^ n7188 ^ 1'b0 ;
  assign n7191 = x228 & n1959 ;
  assign n7192 = ( n4427 & ~n5359 ) | ( n4427 & n7191 ) | ( ~n5359 & n7191 ) ;
  assign n7196 = n6640 ^ n2998 ^ n1665 ;
  assign n7197 = n566 | n5046 ;
  assign n7198 = n7196 | n7197 ;
  assign n7193 = n1051 | n2856 ;
  assign n7194 = n7193 ^ n2838 ^ 1'b0 ;
  assign n7195 = n7194 ^ n2520 ^ n1688 ;
  assign n7199 = n7198 ^ n7195 ^ n3059 ;
  assign n7200 = ( n736 & ~n2904 ) | ( n736 & n3563 ) | ( ~n2904 & n3563 ) ;
  assign n7201 = ( ~n1269 & n3377 ) | ( ~n1269 & n7200 ) | ( n3377 & n7200 ) ;
  assign n7202 = n7201 ^ n1024 ^ 1'b0 ;
  assign n7203 = n2905 & n7202 ;
  assign n7204 = ( n7192 & n7199 ) | ( n7192 & n7203 ) | ( n7199 & n7203 ) ;
  assign n7207 = n4255 ^ x101 ^ 1'b0 ;
  assign n7205 = ~n1080 & n1165 ;
  assign n7206 = n7205 ^ n1884 ^ 1'b0 ;
  assign n7208 = n7207 ^ n7206 ^ 1'b0 ;
  assign n7209 = ( n3105 & ~n4898 ) | ( n3105 & n7208 ) | ( ~n4898 & n7208 ) ;
  assign n7210 = n1735 & ~n1873 ;
  assign n7211 = n4743 ^ n2541 ^ x187 ;
  assign n7212 = n2944 ^ n1612 ^ x136 ;
  assign n7213 = n7211 & n7212 ;
  assign n7214 = n7210 & n7213 ;
  assign n7216 = n4464 ^ n3985 ^ n728 ;
  assign n7217 = n3520 | n7216 ;
  assign n7215 = ( x170 & n652 ) | ( x170 & n5228 ) | ( n652 & n5228 ) ;
  assign n7218 = n7217 ^ n7215 ^ n5556 ;
  assign n7219 = n2763 | n2987 ;
  assign n7220 = n7219 ^ n6201 ^ 1'b0 ;
  assign n7221 = n6848 ^ n698 ^ x207 ;
  assign n7222 = n7221 ^ n3968 ^ 1'b0 ;
  assign n7223 = ~n1861 & n3435 ;
  assign n7224 = n5804 ^ n1957 ^ 1'b0 ;
  assign n7225 = ~n1265 & n7224 ;
  assign n7226 = n2909 ^ n593 ^ 1'b0 ;
  assign n7227 = n7226 ^ n5226 ^ x18 ;
  assign n7228 = n3425 ^ n1619 ^ 1'b0 ;
  assign n7230 = ( n702 & n2126 ) | ( n702 & n5080 ) | ( n2126 & n5080 ) ;
  assign n7231 = n7230 ^ n581 ^ 1'b0 ;
  assign n7229 = ~n299 & n4436 ;
  assign n7232 = n7231 ^ n7229 ^ 1'b0 ;
  assign n7233 = ~n7228 & n7232 ;
  assign n7234 = ~n7227 & n7233 ;
  assign n7235 = n4739 ^ n820 ^ n751 ;
  assign n7236 = n3065 ^ n1012 ^ x212 ;
  assign n7237 = n7236 ^ n5002 ^ n1101 ;
  assign n7238 = n7237 ^ n3105 ^ 1'b0 ;
  assign n7239 = n3010 ^ n1496 ^ 1'b0 ;
  assign n7242 = x154 & n436 ;
  assign n7243 = n7242 ^ n3667 ^ 1'b0 ;
  assign n7244 = n7243 ^ n2696 ^ 1'b0 ;
  assign n7245 = ~n1183 & n7244 ;
  assign n7240 = n2469 ^ n2223 ^ x239 ;
  assign n7241 = n7240 ^ n2101 ^ n666 ;
  assign n7246 = n7245 ^ n7241 ^ n2745 ;
  assign n7247 = n7239 & n7246 ;
  assign n7248 = n7238 & n7247 ;
  assign n7249 = n3524 ^ n912 ^ 1'b0 ;
  assign n7250 = ( n2161 & ~n6447 ) | ( n2161 & n7249 ) | ( ~n6447 & n7249 ) ;
  assign n7253 = n1691 & n2391 ;
  assign n7254 = ~n1468 & n7253 ;
  assign n7255 = ( ~n1072 & n4041 ) | ( ~n1072 & n7254 ) | ( n4041 & n7254 ) ;
  assign n7251 = n2310 ^ n757 ^ 1'b0 ;
  assign n7252 = n6778 & n7251 ;
  assign n7256 = n7255 ^ n7252 ^ n2730 ;
  assign n7257 = ( n2792 & n3205 ) | ( n2792 & n3638 ) | ( n3205 & n3638 ) ;
  assign n7258 = n5500 ^ n3125 ^ 1'b0 ;
  assign n7259 = ~n5828 & n7258 ;
  assign n7260 = ~n5843 & n7259 ;
  assign n7261 = n2691 ^ n2390 ^ 1'b0 ;
  assign n7262 = n7261 ^ n3634 ^ 1'b0 ;
  assign n7263 = n2845 & ~n7262 ;
  assign n7264 = ( ~n779 & n2725 ) | ( ~n779 & n4841 ) | ( n2725 & n4841 ) ;
  assign n7265 = ~n5490 & n7264 ;
  assign n7266 = n2583 | n6938 ;
  assign n7267 = n936 & ~n4085 ;
  assign n7268 = n7267 ^ n417 ^ 1'b0 ;
  assign n7269 = ( n1140 & n1342 ) | ( n1140 & n7268 ) | ( n1342 & n7268 ) ;
  assign n7270 = n5265 ^ n4364 ^ n707 ;
  assign n7271 = ~n7269 & n7270 ;
  assign n7272 = n7271 ^ n3289 ^ 1'b0 ;
  assign n7273 = n3596 ^ n1676 ^ 1'b0 ;
  assign n7274 = ~n2912 & n7273 ;
  assign n7275 = n2712 & n7274 ;
  assign n7276 = n3826 & n7275 ;
  assign n7277 = n4051 ^ n3515 ^ 1'b0 ;
  assign n7278 = ~n7276 & n7277 ;
  assign n7279 = n2785 & ~n5197 ;
  assign n7280 = n7279 ^ n4671 ^ 1'b0 ;
  assign n7281 = ( n374 & n4410 ) | ( n374 & n6742 ) | ( n4410 & n6742 ) ;
  assign n7282 = ~n6035 & n6622 ;
  assign n7283 = ( n983 & n5513 ) | ( n983 & ~n7282 ) | ( n5513 & ~n7282 ) ;
  assign n7284 = n4137 ^ n2157 ^ 1'b0 ;
  assign n7285 = ~n7158 & n7284 ;
  assign n7286 = n7285 ^ n5669 ^ n5395 ;
  assign n7287 = ~n971 & n3736 ;
  assign n7288 = n7287 ^ n2465 ^ 1'b0 ;
  assign n7289 = n7288 ^ n1573 ^ n1300 ;
  assign n7290 = n7289 ^ n4318 ^ 1'b0 ;
  assign n7291 = ~n7286 & n7290 ;
  assign n7292 = ~n461 & n1179 ;
  assign n7293 = ~n2531 & n7292 ;
  assign n7294 = n7293 ^ n2410 ^ n2325 ;
  assign n7295 = ~n5130 & n7294 ;
  assign n7296 = ~n2670 & n7295 ;
  assign n7297 = ~n2536 & n3114 ;
  assign n7298 = n7297 ^ n3735 ^ 1'b0 ;
  assign n7299 = n2059 ^ n1226 ^ 1'b0 ;
  assign n7300 = n4338 | n7299 ;
  assign n7301 = ~n6607 & n7300 ;
  assign n7302 = ( n615 & ~n1961 ) | ( n615 & n7301 ) | ( ~n1961 & n7301 ) ;
  assign n7303 = n3071 | n5921 ;
  assign n7304 = n7303 ^ n707 ^ 1'b0 ;
  assign n7305 = ~n1209 & n2030 ;
  assign n7306 = ~n4756 & n7305 ;
  assign n7307 = n2481 & ~n7306 ;
  assign n7308 = ( n2760 & n4429 ) | ( n2760 & ~n7307 ) | ( n4429 & ~n7307 ) ;
  assign n7309 = n3858 & ~n7308 ;
  assign n7310 = ~n4882 & n7309 ;
  assign n7311 = n7310 ^ n4310 ^ n532 ;
  assign n7312 = ~n726 & n2443 ;
  assign n7313 = n7312 ^ n5317 ^ 1'b0 ;
  assign n7314 = n2064 ^ n919 ^ x248 ;
  assign n7315 = ( n480 & ~n1823 ) | ( n480 & n7314 ) | ( ~n1823 & n7314 ) ;
  assign n7316 = n450 & ~n874 ;
  assign n7317 = ~n2243 & n7316 ;
  assign n7318 = n7317 ^ n3865 ^ n3761 ;
  assign n7319 = x163 & n1623 ;
  assign n7320 = n7318 & n7319 ;
  assign n7321 = n7315 & n7320 ;
  assign n7322 = n7321 ^ n5025 ^ n3640 ;
  assign n7323 = ( n4009 & n4118 ) | ( n4009 & ~n6330 ) | ( n4118 & ~n6330 ) ;
  assign n7324 = n5304 ^ n2008 ^ 1'b0 ;
  assign n7325 = n4737 ^ n4217 ^ n997 ;
  assign n7326 = n5124 ^ n1640 ^ n756 ;
  assign n7327 = n7326 ^ n6478 ^ n5133 ;
  assign n7328 = n7310 | n7327 ;
  assign n7329 = n7325 & ~n7328 ;
  assign n7330 = n7329 ^ n5900 ^ 1'b0 ;
  assign n7331 = n7324 & ~n7330 ;
  assign n7332 = n4001 ^ x232 ^ 1'b0 ;
  assign n7333 = ( n1059 & n4100 ) | ( n1059 & n6819 ) | ( n4100 & n6819 ) ;
  assign n7334 = n7333 ^ n3336 ^ n2154 ;
  assign n7335 = n7332 & n7334 ;
  assign n7336 = n7335 ^ n6797 ^ 1'b0 ;
  assign n7337 = n4553 ^ n430 ^ 1'b0 ;
  assign n7338 = n5121 & n5697 ;
  assign n7339 = n7338 ^ n5575 ^ 1'b0 ;
  assign n7340 = n7337 & ~n7339 ;
  assign n7341 = n4850 & n7340 ;
  assign n7342 = n450 ^ x248 ^ 1'b0 ;
  assign n7343 = n2588 ^ n1400 ^ n1387 ;
  assign n7344 = ~n7342 & n7343 ;
  assign n7345 = n7344 ^ n5787 ^ 1'b0 ;
  assign n7346 = x105 & n633 ;
  assign n7347 = ~n3195 & n7346 ;
  assign n7348 = n2497 | n7347 ;
  assign n7349 = n2939 & ~n7348 ;
  assign n7350 = ~n693 & n6218 ;
  assign n7351 = n1188 & ~n7350 ;
  assign n7352 = ~n1545 & n7351 ;
  assign n7353 = ( n3196 & ~n4315 ) | ( n3196 & n6960 ) | ( ~n4315 & n6960 ) ;
  assign n7354 = n7352 | n7353 ;
  assign n7355 = ( ~x147 & n4488 ) | ( ~x147 & n5579 ) | ( n4488 & n5579 ) ;
  assign n7357 = ( n438 & ~n1468 ) | ( n438 & n3507 ) | ( ~n1468 & n3507 ) ;
  assign n7356 = n1219 & ~n4271 ;
  assign n7358 = n7357 ^ n7356 ^ n1981 ;
  assign n7359 = n4632 & n7358 ;
  assign n7360 = n3070 & ~n4459 ;
  assign n7361 = ( n1482 & ~n2765 ) | ( n1482 & n7360 ) | ( ~n2765 & n7360 ) ;
  assign n7362 = x36 & n2957 ;
  assign n7363 = n7362 ^ n1423 ^ 1'b0 ;
  assign n7365 = ~n2602 & n2893 ;
  assign n7366 = n7365 ^ n3006 ^ 1'b0 ;
  assign n7364 = n1132 & ~n3165 ;
  assign n7367 = n7366 ^ n7364 ^ 1'b0 ;
  assign n7368 = ~n3604 & n6097 ;
  assign n7369 = ~n3361 & n7368 ;
  assign n7370 = n7369 ^ n3409 ^ n2337 ;
  assign n7371 = ( n7363 & ~n7367 ) | ( n7363 & n7370 ) | ( ~n7367 & n7370 ) ;
  assign n7373 = n668 & ~n5386 ;
  assign n7372 = ( n947 & ~n2443 ) | ( n947 & n4763 ) | ( ~n2443 & n4763 ) ;
  assign n7374 = n7373 ^ n7372 ^ 1'b0 ;
  assign n7379 = n3859 & n6222 ;
  assign n7375 = ( ~n2173 & n4499 ) | ( ~n2173 & n6341 ) | ( n4499 & n6341 ) ;
  assign n7376 = n7152 & ~n7238 ;
  assign n7377 = n7376 ^ n706 ^ 1'b0 ;
  assign n7378 = ~n7375 & n7377 ;
  assign n7380 = n7379 ^ n7378 ^ 1'b0 ;
  assign n7381 = n7380 ^ n4109 ^ 1'b0 ;
  assign n7382 = n1175 & n7381 ;
  assign n7385 = n5987 & ~n6202 ;
  assign n7386 = n7385 ^ n5688 ^ 1'b0 ;
  assign n7387 = n4152 ^ n1521 ^ 1'b0 ;
  assign n7388 = n7386 & ~n7387 ;
  assign n7389 = n6421 & n7388 ;
  assign n7383 = n5408 ^ n1823 ^ n807 ;
  assign n7384 = ~n1834 & n7383 ;
  assign n7390 = n7389 ^ n7384 ^ 1'b0 ;
  assign n7391 = n3801 ^ n492 ^ x3 ;
  assign n7392 = n4827 & ~n7391 ;
  assign n7393 = x154 | n2154 ;
  assign n7394 = n7393 ^ n3881 ^ 1'b0 ;
  assign n7395 = n7394 ^ n3479 ^ 1'b0 ;
  assign n7396 = n5805 ^ n2070 ^ 1'b0 ;
  assign n7399 = n2881 ^ n1159 ^ n666 ;
  assign n7400 = ~n1403 & n7399 ;
  assign n7401 = n5418 & n7400 ;
  assign n7397 = n4478 ^ x142 ^ 1'b0 ;
  assign n7398 = n3328 | n7397 ;
  assign n7402 = n7401 ^ n7398 ^ n2377 ;
  assign n7403 = n5105 ^ n3750 ^ 1'b0 ;
  assign n7404 = n7403 ^ n4881 ^ n3331 ;
  assign n7405 = n7404 ^ n3746 ^ x3 ;
  assign n7406 = ~n2247 & n3832 ;
  assign n7407 = n4820 | n7406 ;
  assign n7408 = n7405 | n7407 ;
  assign n7409 = ~n2297 & n7143 ;
  assign n7410 = ( n2114 & n2934 ) | ( n2114 & ~n7401 ) | ( n2934 & ~n7401 ) ;
  assign n7411 = n7410 ^ n1574 ^ 1'b0 ;
  assign n7412 = n7411 ^ n1016 ^ n905 ;
  assign n7413 = ( ~n4267 & n4968 ) | ( ~n4267 & n5739 ) | ( n4968 & n5739 ) ;
  assign n7415 = n2923 ^ n1442 ^ n738 ;
  assign n7414 = n6541 ^ n3667 ^ n2306 ;
  assign n7416 = n7415 ^ n7414 ^ n5405 ;
  assign n7417 = ( n2310 & n7413 ) | ( n2310 & ~n7416 ) | ( n7413 & ~n7416 ) ;
  assign n7418 = n3783 & n6534 ;
  assign n7419 = n7418 ^ n5025 ^ 1'b0 ;
  assign n7420 = n6947 ^ n6549 ^ n297 ;
  assign n7421 = n3684 & ~n7420 ;
  assign n7422 = n3772 & ~n4796 ;
  assign n7423 = ~n4645 & n7422 ;
  assign n7424 = ~n2195 & n7423 ;
  assign n7425 = x28 & ~n7424 ;
  assign n7426 = n7425 ^ n5431 ^ 1'b0 ;
  assign n7427 = n1979 & ~n7426 ;
  assign n7428 = n3073 ^ n2153 ^ 1'b0 ;
  assign n7430 = n2260 & n3711 ;
  assign n7431 = ~n1385 & n7430 ;
  assign n7429 = n2596 ^ n334 ^ x63 ;
  assign n7432 = n7431 ^ n7429 ^ 1'b0 ;
  assign n7433 = n6696 & n7432 ;
  assign n7434 = n7433 ^ n5843 ^ 1'b0 ;
  assign n7435 = n2492 | n6105 ;
  assign n7436 = n7435 ^ n1662 ^ 1'b0 ;
  assign n7437 = n2495 ^ n1443 ^ x90 ;
  assign n7438 = n1658 ^ x162 ^ 1'b0 ;
  assign n7439 = n5080 & n7438 ;
  assign n7440 = ~n2175 & n2281 ;
  assign n7441 = n7440 ^ n6224 ^ n4723 ;
  assign n7442 = ( ~n7285 & n7439 ) | ( ~n7285 & n7441 ) | ( n7439 & n7441 ) ;
  assign n7443 = n7437 & ~n7442 ;
  assign n7444 = ~n4131 & n7443 ;
  assign n7445 = n1152 & n6628 ;
  assign n7446 = n2106 ^ n715 ^ n345 ;
  assign n7447 = n2336 ^ n1517 ^ 1'b0 ;
  assign n7448 = ( n838 & n4056 ) | ( n838 & n7447 ) | ( n4056 & n7447 ) ;
  assign n7449 = n6538 ^ n3716 ^ 1'b0 ;
  assign n7464 = ( n734 & ~n1720 ) | ( n734 & n2100 ) | ( ~n1720 & n2100 ) ;
  assign n7457 = n673 | n6197 ;
  assign n7458 = n7457 ^ n2495 ^ 1'b0 ;
  assign n7459 = ~n2074 & n3645 ;
  assign n7460 = n7458 & n7459 ;
  assign n7461 = ( n1484 & ~n1605 ) | ( n1484 & n7460 ) | ( ~n1605 & n7460 ) ;
  assign n7456 = n4150 | n4890 ;
  assign n7462 = n7461 ^ n7456 ^ 1'b0 ;
  assign n7454 = ( n1725 & n3752 ) | ( n1725 & n7326 ) | ( n3752 & n7326 ) ;
  assign n7455 = n7454 ^ n1087 ^ 1'b0 ;
  assign n7451 = n2033 & ~n2825 ;
  assign n7452 = ~n2527 & n7451 ;
  assign n7453 = n7452 ^ n1173 ^ 1'b0 ;
  assign n7463 = n7462 ^ n7455 ^ n7453 ;
  assign n7465 = n7464 ^ n7463 ^ n1511 ;
  assign n7450 = n1518 & ~n6934 ;
  assign n7466 = n7465 ^ n7450 ^ 1'b0 ;
  assign n7467 = n1276 & ~n2308 ;
  assign n7469 = n1730 & ~n4743 ;
  assign n7470 = n7469 ^ n2861 ^ 1'b0 ;
  assign n7471 = ~n2308 & n7470 ;
  assign n7468 = n1034 & n1559 ;
  assign n7472 = n7471 ^ n7468 ^ 1'b0 ;
  assign n7473 = ( n2466 & n7467 ) | ( n2466 & ~n7472 ) | ( n7467 & ~n7472 ) ;
  assign n7474 = ( n1072 & n1315 ) | ( n1072 & ~n1672 ) | ( n1315 & ~n1672 ) ;
  assign n7475 = ( n1754 & n3149 ) | ( n1754 & n7474 ) | ( n3149 & n7474 ) ;
  assign n7476 = n2950 & n3247 ;
  assign n7477 = n1383 | n7476 ;
  assign n7478 = n2522 & n6082 ;
  assign n7480 = x102 & ~n3356 ;
  assign n7479 = n7425 ^ n3262 ^ 1'b0 ;
  assign n7481 = n7480 ^ n7479 ^ n5086 ;
  assign n7486 = ~n982 & n1197 ;
  assign n7487 = n7486 ^ n1564 ^ 1'b0 ;
  assign n7482 = ( ~n2789 & n2864 ) | ( ~n2789 & n3813 ) | ( n2864 & n3813 ) ;
  assign n7483 = ~n587 & n7482 ;
  assign n7484 = n7483 ^ n2017 ^ 1'b0 ;
  assign n7485 = ( n2000 & n2351 ) | ( n2000 & ~n7484 ) | ( n2351 & ~n7484 ) ;
  assign n7488 = n7487 ^ n7485 ^ n6780 ;
  assign n7489 = n6486 ^ n5405 ^ n2782 ;
  assign n7490 = n1721 | n7489 ;
  assign n7491 = n3365 ^ n2835 ^ 1'b0 ;
  assign n7492 = n7491 ^ n2210 ^ n602 ;
  assign n7494 = n1957 ^ x148 ^ 1'b0 ;
  assign n7493 = ~n1211 & n1851 ;
  assign n7495 = n7494 ^ n7493 ^ n2588 ;
  assign n7496 = ( n1941 & n7492 ) | ( n1941 & ~n7495 ) | ( n7492 & ~n7495 ) ;
  assign n7497 = n5716 ^ n1639 ^ 1'b0 ;
  assign n7498 = n1588 & n7497 ;
  assign n7499 = n7113 ^ n5112 ^ 1'b0 ;
  assign n7500 = n2894 | n3746 ;
  assign n7501 = n3178 & ~n4712 ;
  assign n7502 = n3239 & ~n4190 ;
  assign n7503 = n7502 ^ n2699 ^ 1'b0 ;
  assign n7504 = ~n6555 & n6990 ;
  assign n7505 = n7504 ^ n3728 ^ 1'b0 ;
  assign n7506 = n5575 ^ n3048 ^ 1'b0 ;
  assign n7507 = n6695 | n7506 ;
  assign n7508 = n1645 & n7507 ;
  assign n7509 = n5457 ^ n3115 ^ n2297 ;
  assign n7510 = n1044 | n7509 ;
  assign n7517 = n1709 & n4076 ;
  assign n7518 = ( n2412 & n5270 ) | ( n2412 & ~n7517 ) | ( n5270 & ~n7517 ) ;
  assign n7519 = n7518 ^ n4155 ^ 1'b0 ;
  assign n7513 = n3737 ^ n2657 ^ n2610 ;
  assign n7511 = n1863 ^ n1418 ^ x210 ;
  assign n7512 = ~n1906 & n7511 ;
  assign n7514 = n7513 ^ n7512 ^ 1'b0 ;
  assign n7515 = n2536 | n4656 ;
  assign n7516 = n7514 & ~n7515 ;
  assign n7520 = n7519 ^ n7516 ^ 1'b0 ;
  assign n7521 = n4743 ^ n3702 ^ 1'b0 ;
  assign n7522 = ( n280 & n7076 ) | ( n280 & n7521 ) | ( n7076 & n7521 ) ;
  assign n7523 = n2781 & ~n7522 ;
  assign n7524 = n7523 ^ n6045 ^ n5851 ;
  assign n7525 = n5528 ^ x225 ^ 1'b0 ;
  assign n7526 = n6624 | n7525 ;
  assign n7527 = ( n2952 & n5430 ) | ( n2952 & ~n7526 ) | ( n5430 & ~n7526 ) ;
  assign n7528 = ( ~n728 & n5744 ) | ( ~n728 & n7527 ) | ( n5744 & n7527 ) ;
  assign n7529 = n2746 ^ n1667 ^ 1'b0 ;
  assign n7530 = x207 & n952 ;
  assign n7531 = ~n2753 & n7530 ;
  assign n7532 = n7529 | n7531 ;
  assign n7533 = n1205 & ~n7532 ;
  assign n7534 = ~n5425 & n7533 ;
  assign n7535 = n7534 ^ n2071 ^ n1525 ;
  assign n7538 = ( n1729 & n2148 ) | ( n1729 & n5675 ) | ( n2148 & n5675 ) ;
  assign n7536 = ~n1893 & n2466 ;
  assign n7537 = n7536 ^ n907 ^ 1'b0 ;
  assign n7539 = n7538 ^ n7537 ^ n495 ;
  assign n7540 = n7539 ^ n2456 ^ 1'b0 ;
  assign n7541 = n7535 & n7540 ;
  assign n7542 = ( n632 & n2730 ) | ( n632 & n3778 ) | ( n2730 & n3778 ) ;
  assign n7543 = n1415 & n5422 ;
  assign n7544 = ~n7542 & n7543 ;
  assign n7545 = ~n1438 & n2524 ;
  assign n7546 = n7545 ^ n481 ^ 1'b0 ;
  assign n7547 = n1733 | n7546 ;
  assign n7548 = ( x178 & ~n2702 ) | ( x178 & n3122 ) | ( ~n2702 & n3122 ) ;
  assign n7549 = n7548 ^ n1597 ^ 1'b0 ;
  assign n7550 = x32 & ~n2643 ;
  assign n7551 = ~n2981 & n7550 ;
  assign n7552 = n3022 | n6895 ;
  assign n7553 = ( x144 & ~n3001 ) | ( x144 & n7552 ) | ( ~n3001 & n7552 ) ;
  assign n7554 = n6602 ^ n695 ^ 1'b0 ;
  assign n7555 = n7554 ^ n5061 ^ 1'b0 ;
  assign n7556 = n4501 ^ n4425 ^ 1'b0 ;
  assign n7557 = n7555 | n7556 ;
  assign n7558 = n5729 ^ n3722 ^ n3044 ;
  assign n7559 = ( n2534 & n3740 ) | ( n2534 & ~n5529 ) | ( n3740 & ~n5529 ) ;
  assign n7560 = n7234 | n7559 ;
  assign n7561 = n7558 & ~n7560 ;
  assign n7566 = n4007 | n4220 ;
  assign n7567 = n3550 & ~n7566 ;
  assign n7568 = n1405 & n7567 ;
  assign n7569 = n7568 ^ n6282 ^ n3711 ;
  assign n7570 = n7569 ^ n891 ^ 1'b0 ;
  assign n7571 = ~n6891 & n7570 ;
  assign n7562 = n4016 | n6883 ;
  assign n7563 = n7562 ^ n543 ^ 1'b0 ;
  assign n7564 = n7563 ^ n3771 ^ n1421 ;
  assign n7565 = n7564 ^ n5849 ^ n4749 ;
  assign n7572 = n7571 ^ n7565 ^ n2965 ;
  assign n7573 = n4322 ^ n2191 ^ 1'b0 ;
  assign n7574 = n7573 ^ x81 ^ 1'b0 ;
  assign n7580 = n2685 ^ n2386 ^ 1'b0 ;
  assign n7581 = ~n3410 & n7580 ;
  assign n7582 = n7581 ^ n3385 ^ 1'b0 ;
  assign n7575 = x174 & n580 ;
  assign n7576 = n634 & n7575 ;
  assign n7577 = n6326 & n7576 ;
  assign n7578 = ( n2227 & ~n5639 ) | ( n2227 & n7577 ) | ( ~n5639 & n7577 ) ;
  assign n7579 = ( ~n3663 & n6562 ) | ( ~n3663 & n7578 ) | ( n6562 & n7578 ) ;
  assign n7583 = n7582 ^ n7579 ^ n5439 ;
  assign n7584 = n2170 ^ n1150 ^ x77 ;
  assign n7585 = n483 | n602 ;
  assign n7586 = n1805 & ~n7585 ;
  assign n7587 = n6529 ^ n1870 ^ 1'b0 ;
  assign n7588 = ~n7586 & n7587 ;
  assign n7589 = n7588 ^ n5126 ^ n534 ;
  assign n7590 = n2775 & n7589 ;
  assign n7591 = n6757 ^ n6296 ^ 1'b0 ;
  assign n7592 = n1994 & ~n7591 ;
  assign n7593 = n7389 ^ n2785 ^ 1'b0 ;
  assign n7600 = n4987 ^ n1168 ^ 1'b0 ;
  assign n7601 = n7474 ^ n3779 ^ 1'b0 ;
  assign n7602 = n7600 & ~n7601 ;
  assign n7603 = n7602 ^ n4328 ^ n1650 ;
  assign n7604 = ~x80 & n7603 ;
  assign n7594 = x38 & n291 ;
  assign n7595 = n1516 & n7594 ;
  assign n7596 = n5488 & n7595 ;
  assign n7597 = n7596 ^ n4469 ^ 1'b0 ;
  assign n7598 = n7597 ^ n3573 ^ 1'b0 ;
  assign n7599 = n4538 | n7598 ;
  assign n7605 = n7604 ^ n7599 ^ n2241 ;
  assign n7607 = ~n904 & n2412 ;
  assign n7608 = ~n1158 & n7607 ;
  assign n7609 = n7608 ^ n1434 ^ 1'b0 ;
  assign n7606 = n1708 & ~n6874 ;
  assign n7610 = n7609 ^ n7606 ^ 1'b0 ;
  assign n7611 = n2513 ^ n1489 ^ 1'b0 ;
  assign n7612 = n7611 ^ n1153 ^ n988 ;
  assign n7613 = n3151 ^ n1251 ^ n891 ;
  assign n7614 = ( ~n1354 & n2490 ) | ( ~n1354 & n7613 ) | ( n2490 & n7613 ) ;
  assign n7615 = n6011 ^ n2354 ^ 1'b0 ;
  assign n7616 = ( n7612 & ~n7614 ) | ( n7612 & n7615 ) | ( ~n7614 & n7615 ) ;
  assign n7617 = n1315 ^ n449 ^ x219 ;
  assign n7618 = n1153 & ~n7617 ;
  assign n7619 = n1832 & n7618 ;
  assign n7620 = n1894 | n7619 ;
  assign n7621 = n6423 & ~n7620 ;
  assign n7622 = n7621 ^ n7201 ^ n3471 ;
  assign n7624 = ~n1475 & n2341 ;
  assign n7625 = ~n4773 & n7624 ;
  assign n7623 = n1398 & n2408 ;
  assign n7626 = n7625 ^ n7623 ^ 1'b0 ;
  assign n7627 = n4321 ^ n3258 ^ 1'b0 ;
  assign n7628 = ( n2719 & n7626 ) | ( n2719 & ~n7627 ) | ( n7626 & ~n7627 ) ;
  assign n7629 = ~n1488 & n2778 ;
  assign n7630 = n7629 ^ n4201 ^ 1'b0 ;
  assign n7631 = n1334 ^ x109 ^ 1'b0 ;
  assign n7632 = n7630 & ~n7631 ;
  assign n7637 = ( n749 & ~n2659 ) | ( n749 & n3837 ) | ( ~n2659 & n3837 ) ;
  assign n7633 = n2838 ^ n2163 ^ 1'b0 ;
  assign n7634 = n2894 & ~n4102 ;
  assign n7635 = ( n6164 & ~n7633 ) | ( n6164 & n7634 ) | ( ~n7633 & n7634 ) ;
  assign n7636 = n7635 ^ n4730 ^ x160 ;
  assign n7638 = n7637 ^ n7636 ^ n5530 ;
  assign n7639 = ( ~n2397 & n7632 ) | ( ~n2397 & n7638 ) | ( n7632 & n7638 ) ;
  assign n7643 = n4555 ^ n1753 ^ 1'b0 ;
  assign n7640 = ~n1858 & n3361 ;
  assign n7641 = n7640 ^ n3573 ^ 1'b0 ;
  assign n7642 = n274 | n7641 ;
  assign n7644 = n7643 ^ n7642 ^ 1'b0 ;
  assign n7645 = ~n4296 & n7644 ;
  assign n7646 = n7645 ^ x56 ^ 1'b0 ;
  assign n7654 = n6421 ^ n4306 ^ 1'b0 ;
  assign n7655 = n3490 & ~n7654 ;
  assign n7651 = ( ~n761 & n890 ) | ( ~n761 & n7613 ) | ( n890 & n7613 ) ;
  assign n7652 = n4933 ^ n4741 ^ 1'b0 ;
  assign n7653 = n7651 & ~n7652 ;
  assign n7647 = n4429 ^ n2918 ^ 1'b0 ;
  assign n7648 = n7647 ^ n5480 ^ 1'b0 ;
  assign n7649 = ~n678 & n7648 ;
  assign n7650 = n7649 ^ n4627 ^ 1'b0 ;
  assign n7656 = n7655 ^ n7653 ^ n7650 ;
  assign n7662 = ~n3502 & n6884 ;
  assign n7657 = n2145 | n2673 ;
  assign n7658 = ( x34 & n3992 ) | ( x34 & ~n5441 ) | ( n3992 & ~n5441 ) ;
  assign n7659 = n1054 & ~n7658 ;
  assign n7660 = n3788 | n7659 ;
  assign n7661 = n7657 & ~n7660 ;
  assign n7663 = n7662 ^ n7661 ^ n3247 ;
  assign n7664 = ~n1346 & n2721 ;
  assign n7665 = ( x31 & n761 ) | ( x31 & n798 ) | ( n761 & n798 ) ;
  assign n7666 = n7664 & ~n7665 ;
  assign n7667 = ~n954 & n7666 ;
  assign n7668 = n7667 ^ n3058 ^ 1'b0 ;
  assign n7670 = n3472 ^ n979 ^ n261 ;
  assign n7671 = ( x179 & n3239 ) | ( x179 & n7670 ) | ( n3239 & n7670 ) ;
  assign n7669 = n2861 ^ n1957 ^ 1'b0 ;
  assign n7672 = n7671 ^ n7669 ^ x160 ;
  assign n7673 = x133 & n3830 ;
  assign n7674 = ( n2542 & n5168 ) | ( n2542 & ~n7673 ) | ( n5168 & ~n7673 ) ;
  assign n7675 = n4280 & n6488 ;
  assign n7676 = n7675 ^ n6639 ^ n4819 ;
  assign n7677 = ~n1764 & n3031 ;
  assign n7678 = ~n4261 & n7677 ;
  assign n7679 = ( ~n4028 & n4079 ) | ( ~n4028 & n7678 ) | ( n4079 & n7678 ) ;
  assign n7680 = n2887 & n4748 ;
  assign n7681 = ~n6124 & n7680 ;
  assign n7682 = ( n806 & n1684 ) | ( n806 & n2968 ) | ( n1684 & n2968 ) ;
  assign n7683 = ~n518 & n7682 ;
  assign n7684 = n3930 & n7683 ;
  assign n7685 = n7684 ^ n2047 ^ 1'b0 ;
  assign n7686 = n2325 ^ n352 ^ 1'b0 ;
  assign n7687 = ( x220 & ~n4720 ) | ( x220 & n7686 ) | ( ~n4720 & n7686 ) ;
  assign n7688 = n7687 ^ n2458 ^ n738 ;
  assign n7689 = n7688 ^ n1287 ^ 1'b0 ;
  assign n7690 = n7282 ^ n1474 ^ 1'b0 ;
  assign n7691 = n7689 | n7690 ;
  assign n7693 = n3967 ^ n1592 ^ n1483 ;
  assign n7692 = n6373 ^ n5809 ^ 1'b0 ;
  assign n7694 = n7693 ^ n7692 ^ n1181 ;
  assign n7695 = n6753 ^ x11 ^ 1'b0 ;
  assign n7696 = n2440 | n7695 ;
  assign n7697 = ( n5044 & ~n5855 ) | ( n5044 & n7696 ) | ( ~n5855 & n7696 ) ;
  assign n7701 = ( n365 & ~n1050 ) | ( n365 & n1936 ) | ( ~n1050 & n1936 ) ;
  assign n7702 = n7701 ^ n2382 ^ 1'b0 ;
  assign n7703 = n5823 | n7702 ;
  assign n7698 = ~n1095 & n2156 ;
  assign n7699 = n5166 | n7698 ;
  assign n7700 = n7671 | n7699 ;
  assign n7704 = n7703 ^ n7700 ^ 1'b0 ;
  assign n7705 = n7697 & ~n7704 ;
  assign n7706 = n3673 ^ n1297 ^ 1'b0 ;
  assign n7711 = n409 & ~n996 ;
  assign n7707 = n1697 ^ n901 ^ 1'b0 ;
  assign n7708 = n7707 ^ n1057 ^ n368 ;
  assign n7709 = ( n1350 & n1411 ) | ( n1350 & n7708 ) | ( n1411 & n7708 ) ;
  assign n7710 = ( n2036 & n6937 ) | ( n2036 & n7709 ) | ( n6937 & n7709 ) ;
  assign n7712 = n7711 ^ n7710 ^ 1'b0 ;
  assign n7713 = n4839 & ~n5087 ;
  assign n7714 = ( ~n4106 & n4121 ) | ( ~n4106 & n4609 ) | ( n4121 & n4609 ) ;
  assign n7715 = n7714 ^ n4656 ^ 1'b0 ;
  assign n7716 = n7713 & ~n7715 ;
  assign n7717 = n5246 & n7716 ;
  assign n7718 = n7717 ^ n2916 ^ 1'b0 ;
  assign n7719 = x184 & ~n1841 ;
  assign n7720 = n4010 & ~n7719 ;
  assign n7721 = ~n1571 & n7720 ;
  assign n7722 = n7721 ^ n1697 ^ 1'b0 ;
  assign n7724 = n1274 | n1361 ;
  assign n7723 = n287 | n7034 ;
  assign n7725 = n7724 ^ n7723 ^ 1'b0 ;
  assign n7726 = ( n2646 & ~n4879 ) | ( n2646 & n7725 ) | ( ~n4879 & n7725 ) ;
  assign n7727 = ( n399 & n7722 ) | ( n399 & ~n7726 ) | ( n7722 & ~n7726 ) ;
  assign n7728 = n1861 | n7420 ;
  assign n7729 = n7728 ^ n5966 ^ 1'b0 ;
  assign n7740 = n1656 ^ n677 ^ 1'b0 ;
  assign n7737 = n6872 ^ n6362 ^ 1'b0 ;
  assign n7738 = ~n2061 & n7737 ;
  assign n7739 = n5951 & n7738 ;
  assign n7741 = n7740 ^ n7739 ^ 1'b0 ;
  assign n7742 = n7741 ^ n1692 ^ n609 ;
  assign n7730 = n4731 ^ n2390 ^ 1'b0 ;
  assign n7731 = n1414 | n7730 ;
  assign n7732 = ( ~n475 & n3256 ) | ( ~n475 & n7731 ) | ( n3256 & n7731 ) ;
  assign n7733 = ( n609 & n1427 ) | ( n609 & n4973 ) | ( n1427 & n4973 ) ;
  assign n7734 = ~n7732 & n7733 ;
  assign n7735 = n541 & n757 ;
  assign n7736 = n7734 | n7735 ;
  assign n7743 = n7742 ^ n7736 ^ 1'b0 ;
  assign n7744 = ( ~x186 & n1186 ) | ( ~x186 & n2531 ) | ( n1186 & n2531 ) ;
  assign n7745 = n7744 ^ n2121 ^ 1'b0 ;
  assign n7746 = n5133 ^ n1591 ^ n946 ;
  assign n7753 = n1581 | n3027 ;
  assign n7751 = ( n3485 & ~n4064 ) | ( n3485 & n7314 ) | ( ~n4064 & n7314 ) ;
  assign n7752 = n7751 ^ n7744 ^ 1'b0 ;
  assign n7747 = n1347 & ~n2596 ;
  assign n7748 = n2654 & n7747 ;
  assign n7749 = n1374 | n7748 ;
  assign n7750 = n4144 & ~n7749 ;
  assign n7754 = n7753 ^ n7752 ^ n7750 ;
  assign n7755 = n4274 ^ n3218 ^ n1365 ;
  assign n7756 = n3722 ^ n1425 ^ n894 ;
  assign n7757 = ( ~n1434 & n7755 ) | ( ~n1434 & n7756 ) | ( n7755 & n7756 ) ;
  assign n7759 = ~x21 & n3286 ;
  assign n7760 = n1938 & ~n7759 ;
  assign n7761 = n7760 ^ n2368 ^ 1'b0 ;
  assign n7762 = n7761 ^ n2707 ^ 1'b0 ;
  assign n7758 = n4198 | n4255 ;
  assign n7763 = n7762 ^ n7758 ^ n5442 ;
  assign n7766 = ( n1274 & ~n4739 ) | ( n1274 & n6620 ) | ( ~n4739 & n6620 ) ;
  assign n7764 = n4325 ^ n2273 ^ n2039 ;
  assign n7765 = ~n2876 & n7764 ;
  assign n7767 = n7766 ^ n7765 ^ 1'b0 ;
  assign n7768 = n374 & ~n2573 ;
  assign n7769 = n7768 ^ n5056 ^ 1'b0 ;
  assign n7770 = n310 & ~n597 ;
  assign n7771 = ( ~n835 & n6011 ) | ( ~n835 & n7770 ) | ( n6011 & n7770 ) ;
  assign n7772 = n449 & ~n7771 ;
  assign n7773 = ~n7769 & n7772 ;
  assign n7774 = n3322 ^ x110 ^ 1'b0 ;
  assign n7775 = n7774 ^ n379 ^ 1'b0 ;
  assign n7776 = n4352 | n6312 ;
  assign n7777 = n1443 | n7776 ;
  assign n7778 = n2303 | n6940 ;
  assign n7779 = n7778 ^ n3275 ^ 1'b0 ;
  assign n7782 = n4919 ^ n2083 ^ 1'b0 ;
  assign n7783 = n7782 ^ n7422 ^ n4669 ;
  assign n7781 = ~n497 & n5625 ;
  assign n7784 = n7783 ^ n7781 ^ n6139 ;
  assign n7780 = n954 | n3176 ;
  assign n7785 = n7784 ^ n7780 ^ 1'b0 ;
  assign n7786 = n1812 & ~n5169 ;
  assign n7787 = ( n3526 & ~n4438 ) | ( n3526 & n7786 ) | ( ~n4438 & n7786 ) ;
  assign n7788 = ~n2160 & n7787 ;
  assign n7793 = n2345 | n4621 ;
  assign n7794 = n7793 ^ n5025 ^ 1'b0 ;
  assign n7789 = n3507 ^ n1125 ^ 1'b0 ;
  assign n7790 = x252 & ~n7789 ;
  assign n7791 = n2126 | n7790 ;
  assign n7792 = n7791 ^ n1274 ^ 1'b0 ;
  assign n7795 = n7794 ^ n7792 ^ x208 ;
  assign n7796 = n6705 ^ n969 ^ 1'b0 ;
  assign n7797 = n594 | n4355 ;
  assign n7798 = n7797 ^ n4782 ^ n2731 ;
  assign n7813 = n2051 ^ n692 ^ 1'b0 ;
  assign n7814 = ~n5932 & n7813 ;
  assign n7811 = n365 & ~n1556 ;
  assign n7812 = n2415 & n7811 ;
  assign n7799 = x155 & n5075 ;
  assign n7800 = ~n6061 & n7799 ;
  assign n7801 = n7626 & n7800 ;
  assign n7802 = ( n1344 & n1920 ) | ( n1344 & ~n7801 ) | ( n1920 & ~n7801 ) ;
  assign n7803 = ( n2238 & n3887 ) | ( n2238 & ~n6486 ) | ( n3887 & ~n6486 ) ;
  assign n7804 = n2975 | n7803 ;
  assign n7805 = n7804 ^ x144 ^ 1'b0 ;
  assign n7806 = n7805 ^ n6267 ^ n2825 ;
  assign n7807 = ~x210 & n1483 ;
  assign n7808 = ~n4417 & n7807 ;
  assign n7809 = n7806 & ~n7808 ;
  assign n7810 = ~n7802 & n7809 ;
  assign n7815 = n7814 ^ n7812 ^ n7810 ;
  assign n7816 = n6445 ^ n4167 ^ 1'b0 ;
  assign n7817 = ~n3233 & n7816 ;
  assign n7820 = ( n516 & n1337 ) | ( n516 & ~n1414 ) | ( n1337 & ~n1414 ) ;
  assign n7821 = ( n1264 & n2754 ) | ( n1264 & n7820 ) | ( n2754 & n7820 ) ;
  assign n7818 = n337 & n1956 ;
  assign n7819 = n7818 ^ n997 ^ 1'b0 ;
  assign n7822 = n7821 ^ n7819 ^ n4230 ;
  assign n7823 = ~n7817 & n7822 ;
  assign n7824 = n7823 ^ n3121 ^ n461 ;
  assign n7825 = n5025 ^ x54 ^ 1'b0 ;
  assign n7826 = n7824 | n7825 ;
  assign n7829 = ~n718 & n1948 ;
  assign n7830 = n2093 & n7829 ;
  assign n7827 = x52 & ~n480 ;
  assign n7828 = n3332 | n7827 ;
  assign n7831 = n7830 ^ n7828 ^ n853 ;
  assign n7834 = n3302 ^ n3289 ^ 1'b0 ;
  assign n7835 = n1106 ^ n759 ^ 1'b0 ;
  assign n7836 = n7834 | n7835 ;
  assign n7832 = n1452 ^ n709 ^ 1'b0 ;
  assign n7833 = n381 & n7832 ;
  assign n7837 = n7836 ^ n7833 ^ 1'b0 ;
  assign n7838 = n3067 & n4816 ;
  assign n7839 = n7814 & n7838 ;
  assign n7840 = n7839 ^ n6562 ^ 1'b0 ;
  assign n7841 = n2377 ^ n1684 ^ x242 ;
  assign n7842 = ( ~n1390 & n3043 ) | ( ~n1390 & n7841 ) | ( n3043 & n7841 ) ;
  assign n7843 = n7842 ^ n3411 ^ 1'b0 ;
  assign n7844 = n7843 ^ n6632 ^ 1'b0 ;
  assign n7845 = n6299 & ~n7844 ;
  assign n7846 = ~n3039 & n7845 ;
  assign n7847 = n5234 ^ n1599 ^ 1'b0 ;
  assign n7848 = ~n5032 & n7847 ;
  assign n7849 = n3546 ^ n907 ^ 1'b0 ;
  assign n7850 = n6173 & n7849 ;
  assign n7852 = ~n2463 & n4279 ;
  assign n7853 = n7852 ^ n350 ^ 1'b0 ;
  assign n7851 = n1093 & n3792 ;
  assign n7854 = n7853 ^ n7851 ^ 1'b0 ;
  assign n7855 = x82 & n406 ;
  assign n7856 = n7855 ^ n2909 ^ 1'b0 ;
  assign n7857 = n3104 & ~n7856 ;
  assign n7858 = n584 | n3050 ;
  assign n7859 = n7858 ^ n7566 ^ 1'b0 ;
  assign n7860 = n7859 ^ n3563 ^ n1525 ;
  assign n7861 = ~n6765 & n7860 ;
  assign n7862 = n7861 ^ n1219 ^ 1'b0 ;
  assign n7863 = x15 & ~n7862 ;
  assign n7864 = n7863 ^ n1059 ^ 1'b0 ;
  assign n7866 = n2520 ^ x230 ^ 1'b0 ;
  assign n7867 = n3715 & n7866 ;
  assign n7865 = n6886 ^ n1897 ^ n995 ;
  assign n7868 = n7867 ^ n7865 ^ 1'b0 ;
  assign n7869 = ~n1334 & n7868 ;
  assign n7870 = n2419 & ~n7786 ;
  assign n7871 = n7870 ^ n2987 ^ n431 ;
  assign n7872 = n855 & n881 ;
  assign n7873 = n7872 ^ n4257 ^ 1'b0 ;
  assign n7883 = n946 & ~n5128 ;
  assign n7876 = n1357 ^ x31 ^ 1'b0 ;
  assign n7877 = n2132 | n7876 ;
  assign n7875 = x158 & n3679 ;
  assign n7878 = n7877 ^ n7875 ^ 1'b0 ;
  assign n7879 = n5456 ^ n2494 ^ n2297 ;
  assign n7880 = n6632 ^ n6193 ^ n1014 ;
  assign n7881 = n7879 | n7880 ;
  assign n7882 = n7878 & n7881 ;
  assign n7874 = n4840 ^ n4224 ^ 1'b0 ;
  assign n7884 = n7883 ^ n7882 ^ n7874 ;
  assign n7885 = n6523 ^ n1324 ^ 1'b0 ;
  assign n7886 = n1569 | n7885 ;
  assign n7887 = n7886 ^ n4800 ^ n280 ;
  assign n7888 = n1255 ^ n281 ^ 1'b0 ;
  assign n7889 = ~n3678 & n7888 ;
  assign n7890 = ~n1956 & n5172 ;
  assign n7891 = n1511 | n4766 ;
  assign n7892 = n813 | n7891 ;
  assign n7893 = n7892 ^ n3727 ^ 1'b0 ;
  assign n7894 = ~n4134 & n7893 ;
  assign n7896 = n1057 & n2013 ;
  assign n7897 = n7896 ^ n314 ^ 1'b0 ;
  assign n7898 = ~n1603 & n7897 ;
  assign n7899 = n7898 ^ n2739 ^ 1'b0 ;
  assign n7900 = n753 | n7899 ;
  assign n7901 = n1742 ^ n1028 ^ 1'b0 ;
  assign n7902 = n295 & n7901 ;
  assign n7903 = ~n7900 & n7902 ;
  assign n7895 = n7342 ^ n821 ^ 1'b0 ;
  assign n7904 = n7903 ^ n7895 ^ 1'b0 ;
  assign n7905 = n2047 ^ n1656 ^ 1'b0 ;
  assign n7906 = n3703 ^ x143 ^ 1'b0 ;
  assign n7907 = n7905 | n7906 ;
  assign n7908 = ( n6225 & n7904 ) | ( n6225 & ~n7907 ) | ( n7904 & ~n7907 ) ;
  assign n7909 = n2399 & n7651 ;
  assign n7911 = n4302 ^ n1460 ^ 1'b0 ;
  assign n7910 = ( n2230 & n2340 ) | ( n2230 & ~n3298 ) | ( n2340 & ~n3298 ) ;
  assign n7912 = n7911 ^ n7910 ^ n2533 ;
  assign n7913 = n4530 ^ n2203 ^ n1882 ;
  assign n7914 = x121 | n1406 ;
  assign n7915 = n2134 | n7914 ;
  assign n7916 = n389 | n7915 ;
  assign n7917 = ( x118 & n1241 ) | ( x118 & ~n3548 ) | ( n1241 & ~n3548 ) ;
  assign n7918 = ( n7913 & n7916 ) | ( n7913 & ~n7917 ) | ( n7916 & ~n7917 ) ;
  assign n7919 = ( x125 & ~n1132 ) | ( x125 & n7918 ) | ( ~n1132 & n7918 ) ;
  assign n7920 = ( ~x55 & n3937 ) | ( ~x55 & n4997 ) | ( n3937 & n4997 ) ;
  assign n7921 = ~n3852 & n5169 ;
  assign n7922 = ( n1378 & n1791 ) | ( n1378 & ~n7921 ) | ( n1791 & ~n7921 ) ;
  assign n7923 = ~n905 & n7922 ;
  assign n7924 = n7923 ^ n3630 ^ 1'b0 ;
  assign n7925 = ( ~n3449 & n3932 ) | ( ~n3449 & n7924 ) | ( n3932 & n7924 ) ;
  assign n7926 = ~x246 & n5531 ;
  assign n7927 = n955 | n7926 ;
  assign n7928 = ( n925 & ~n2728 ) | ( n925 & n7927 ) | ( ~n2728 & n7927 ) ;
  assign n7929 = ( n2512 & ~n3717 ) | ( n2512 & n7928 ) | ( ~n3717 & n7928 ) ;
  assign n7930 = ( ~n1081 & n7925 ) | ( ~n1081 & n7929 ) | ( n7925 & n7929 ) ;
  assign n7931 = ~n3688 & n6139 ;
  assign n7932 = n7931 ^ n6390 ^ 1'b0 ;
  assign n7933 = ~n3814 & n6714 ;
  assign n7934 = n7933 ^ n6139 ^ 1'b0 ;
  assign n7936 = n2549 & ~n4386 ;
  assign n7935 = n511 & ~n1346 ;
  assign n7937 = n7936 ^ n7935 ^ n4383 ;
  assign n7938 = n7788 & ~n7937 ;
  assign n7939 = ~n6325 & n7938 ;
  assign n7942 = n2833 ^ n2178 ^ 1'b0 ;
  assign n7943 = n1443 & ~n7942 ;
  assign n7941 = n4025 ^ n3091 ^ n1265 ;
  assign n7940 = n1255 ^ n399 ^ 1'b0 ;
  assign n7944 = n7943 ^ n7941 ^ n7940 ;
  assign n7946 = n2778 ^ n1018 ^ 1'b0 ;
  assign n7947 = n1078 & n7946 ;
  assign n7948 = ~n4306 & n7947 ;
  assign n7949 = n7948 ^ n4933 ^ 1'b0 ;
  assign n7945 = n2411 & ~n3909 ;
  assign n7950 = n7949 ^ n7945 ^ 1'b0 ;
  assign n7951 = n7950 ^ n7617 ^ n4609 ;
  assign n7952 = n7951 ^ n2369 ^ x252 ;
  assign n7956 = n1004 | n1863 ;
  assign n7957 = n7956 ^ n2125 ^ 1'b0 ;
  assign n7958 = n7474 ^ n2377 ^ 1'b0 ;
  assign n7959 = n7957 & ~n7958 ;
  assign n7953 = n2265 | n4363 ;
  assign n7954 = n4329 | n7953 ;
  assign n7955 = n4113 | n7954 ;
  assign n7960 = n7959 ^ n7955 ^ 1'b0 ;
  assign n7961 = ~n3998 & n7960 ;
  assign n7968 = n7621 ^ n7217 ^ 1'b0 ;
  assign n7962 = n1460 & n2270 ;
  assign n7963 = n7962 ^ n4343 ^ n2624 ;
  assign n7964 = n3223 ^ n3013 ^ 1'b0 ;
  assign n7965 = n2109 | n7964 ;
  assign n7966 = n7965 ^ n2501 ^ n863 ;
  assign n7967 = ~n7963 & n7966 ;
  assign n7969 = n7968 ^ n7967 ^ 1'b0 ;
  assign n7970 = ( ~n597 & n3973 ) | ( ~n597 & n4724 ) | ( n3973 & n4724 ) ;
  assign n7971 = n607 & n7970 ;
  assign n7972 = n2510 ^ n1665 ^ x97 ;
  assign n7973 = ( n303 & n1417 ) | ( n303 & n7972 ) | ( n1417 & n7972 ) ;
  assign n7974 = n7422 & ~n7973 ;
  assign n7975 = n5482 ^ n2339 ^ 1'b0 ;
  assign n7976 = n4806 & ~n7975 ;
  assign n7977 = n1204 & ~n2379 ;
  assign n7978 = ~n7976 & n7977 ;
  assign n7983 = n1458 ^ n1452 ^ n1342 ;
  assign n7980 = n4556 ^ n1493 ^ 1'b0 ;
  assign n7979 = ~n1199 & n4199 ;
  assign n7981 = n7980 ^ n7979 ^ 1'b0 ;
  assign n7982 = n441 | n7981 ;
  assign n7984 = n7983 ^ n7982 ^ 1'b0 ;
  assign n7985 = n5097 & ~n7984 ;
  assign n7986 = n7985 ^ n1827 ^ 1'b0 ;
  assign n7987 = ( n7496 & ~n7978 ) | ( n7496 & n7986 ) | ( ~n7978 & n7986 ) ;
  assign n7988 = n2735 & ~n3032 ;
  assign n7989 = n7644 ^ n1589 ^ n963 ;
  assign n7990 = n1496 ^ n753 ^ n693 ;
  assign n7991 = n7990 ^ n7311 ^ 1'b0 ;
  assign n7992 = n7991 ^ n7650 ^ n2177 ;
  assign n7993 = ~n4055 & n5869 ;
  assign n7994 = ~n1118 & n2606 ;
  assign n7995 = ~n7993 & n7994 ;
  assign n7996 = ~n5622 & n7995 ;
  assign n7997 = n6313 & ~n7552 ;
  assign n7998 = n7996 & n7997 ;
  assign n7999 = n7998 ^ n466 ^ 1'b0 ;
  assign n8000 = n543 | n4267 ;
  assign n8001 = n756 ^ x10 ^ 1'b0 ;
  assign n8006 = n6222 ^ n880 ^ 1'b0 ;
  assign n8002 = ( x28 & ~x112 ) | ( x28 & n1448 ) | ( ~x112 & n1448 ) ;
  assign n8003 = n8002 ^ n1363 ^ 1'b0 ;
  assign n8004 = n4355 & ~n8003 ;
  assign n8005 = n7559 | n8004 ;
  assign n8007 = n8006 ^ n8005 ^ n1336 ;
  assign n8008 = ( n1380 & ~n5185 ) | ( n1380 & n7226 ) | ( ~n5185 & n7226 ) ;
  assign n8009 = n7806 & n8008 ;
  assign n8010 = n8009 ^ n4109 ^ 1'b0 ;
  assign n8011 = n6272 ^ n3332 ^ n2555 ;
  assign n8012 = n8011 ^ n5002 ^ 1'b0 ;
  assign n8013 = n5116 ^ n5097 ^ n3775 ;
  assign n8014 = ( ~n1660 & n5921 ) | ( ~n1660 & n7039 ) | ( n5921 & n7039 ) ;
  assign n8015 = ( n1950 & ~n5980 ) | ( n1950 & n8014 ) | ( ~n5980 & n8014 ) ;
  assign n8016 = n3374 ^ x70 ^ 1'b0 ;
  assign n8017 = n8016 ^ n3345 ^ 1'b0 ;
  assign n8018 = n6382 & ~n8017 ;
  assign n8019 = n5357 & ~n5992 ;
  assign n8020 = n8019 ^ n1727 ^ 1'b0 ;
  assign n8021 = n3332 ^ x155 ^ 1'b0 ;
  assign n8022 = ~n3576 & n8021 ;
  assign n8023 = n8022 ^ n1754 ^ n357 ;
  assign n8024 = n2332 | n6546 ;
  assign n8025 = n7332 ^ n3802 ^ 1'b0 ;
  assign n8026 = n2583 ^ n1720 ^ 1'b0 ;
  assign n8027 = n5796 | n8026 ;
  assign n8028 = n8027 ^ n6114 ^ 1'b0 ;
  assign n8029 = ~n3059 & n8028 ;
  assign n8030 = n3806 & n8029 ;
  assign n8031 = n8030 ^ n7294 ^ n7126 ;
  assign n8032 = n4038 ^ n3627 ^ 1'b0 ;
  assign n8033 = n8032 ^ n5492 ^ n4638 ;
  assign n8034 = ( n2145 & ~n6290 ) | ( n2145 & n8033 ) | ( ~n6290 & n8033 ) ;
  assign n8035 = n3599 | n8034 ;
  assign n8036 = n8031 | n8035 ;
  assign n8037 = n4552 ^ n2823 ^ 1'b0 ;
  assign n8038 = n1173 & ~n8037 ;
  assign n8039 = n8038 ^ n2337 ^ n934 ;
  assign n8040 = n3371 & n8039 ;
  assign n8041 = n8040 ^ n4204 ^ 1'b0 ;
  assign n8042 = n1907 | n8041 ;
  assign n8043 = n6316 ^ n2410 ^ 1'b0 ;
  assign n8044 = n8043 ^ n1418 ^ 1'b0 ;
  assign n8045 = n956 | n1348 ;
  assign n8046 = n8045 ^ n2004 ^ 1'b0 ;
  assign n8047 = ~n3012 & n8046 ;
  assign n8048 = n5150 ^ x253 ^ 1'b0 ;
  assign n8049 = n2931 & n8048 ;
  assign n8050 = ( n686 & n8047 ) | ( n686 & n8049 ) | ( n8047 & n8049 ) ;
  assign n8051 = n5500 ^ n769 ^ x197 ;
  assign n8055 = n6737 ^ n3861 ^ 1'b0 ;
  assign n8056 = n8055 ^ n715 ^ 1'b0 ;
  assign n8052 = x65 & ~n5160 ;
  assign n8053 = n8052 ^ n6060 ^ n5737 ;
  assign n8054 = n4278 & ~n8053 ;
  assign n8057 = n8056 ^ n8054 ^ 1'b0 ;
  assign n8058 = n3868 & n3984 ;
  assign n8059 = n2236 & n8058 ;
  assign n8060 = n8059 ^ n3292 ^ n1216 ;
  assign n8061 = n2602 ^ n838 ^ 1'b0 ;
  assign n8062 = n7060 & n8061 ;
  assign n8063 = n8062 ^ n2735 ^ 1'b0 ;
  assign n8064 = ( n3441 & n7862 ) | ( n3441 & n8063 ) | ( n7862 & n8063 ) ;
  assign n8065 = x120 & ~n883 ;
  assign n8066 = n8065 ^ n2428 ^ 1'b0 ;
  assign n8067 = ( n5408 & ~n5589 ) | ( n5408 & n6814 ) | ( ~n5589 & n6814 ) ;
  assign n8068 = n8066 & ~n8067 ;
  assign n8069 = n8068 ^ n3794 ^ 1'b0 ;
  assign n8070 = ( ~n870 & n2744 ) | ( ~n870 & n5266 ) | ( n2744 & n5266 ) ;
  assign n8071 = n5789 & n7634 ;
  assign n8072 = ~n8070 & n8071 ;
  assign n8073 = n6587 & ~n8072 ;
  assign n8074 = ~n1597 & n2211 ;
  assign n8075 = n7682 & n8074 ;
  assign n8076 = ( ~n2143 & n5716 ) | ( ~n2143 & n6317 ) | ( n5716 & n6317 ) ;
  assign n8077 = n8076 ^ n1161 ^ 1'b0 ;
  assign n8078 = ~n8075 & n8077 ;
  assign n8079 = n354 & n2398 ;
  assign n8080 = n2869 | n3878 ;
  assign n8081 = n7281 & ~n8080 ;
  assign n8082 = ~n8079 & n8081 ;
  assign n8083 = n7972 ^ n1455 ^ 1'b0 ;
  assign n8084 = ( ~n3141 & n4373 ) | ( ~n3141 & n8083 ) | ( n4373 & n8083 ) ;
  assign n8085 = ( x37 & ~n988 ) | ( x37 & n1879 ) | ( ~n988 & n1879 ) ;
  assign n8086 = n6140 ^ n4937 ^ 1'b0 ;
  assign n8087 = n444 & ~n8086 ;
  assign n8088 = n871 & n8087 ;
  assign n8089 = n1405 & n6382 ;
  assign n8090 = n681 & n8089 ;
  assign n8091 = n894 ^ n357 ^ 1'b0 ;
  assign n8092 = ( n2955 & n3500 ) | ( n2955 & n8091 ) | ( n3500 & n8091 ) ;
  assign n8093 = n5820 ^ n4474 ^ x252 ;
  assign n8094 = n4520 & ~n8093 ;
  assign n8095 = n8094 ^ n4337 ^ 1'b0 ;
  assign n8096 = n8092 & ~n8095 ;
  assign n8097 = n1183 & ~n4502 ;
  assign n8098 = n3032 ^ n2807 ^ n2466 ;
  assign n8099 = n3257 & n8098 ;
  assign n8100 = n8097 | n8099 ;
  assign n8101 = n6805 ^ n2246 ^ n1488 ;
  assign n8102 = ~n904 & n6662 ;
  assign n8103 = ~n5577 & n8102 ;
  assign n8104 = x203 | n8103 ;
  assign n8105 = n6708 ^ n4879 ^ n2688 ;
  assign n8106 = n1383 & n2860 ;
  assign n8107 = n2547 & ~n8106 ;
  assign n8108 = ~n1907 & n8107 ;
  assign n8109 = ~n4421 & n8108 ;
  assign n8110 = n3920 & ~n8109 ;
  assign n8111 = n2904 & n8110 ;
  assign n8112 = ~n3622 & n4533 ;
  assign n8113 = n1142 & ~n1361 ;
  assign n8114 = n279 & n8113 ;
  assign n8115 = n4212 | n8114 ;
  assign n8116 = n1017 | n8115 ;
  assign n8117 = n8116 ^ n1006 ^ 1'b0 ;
  assign n8118 = n3283 ^ x34 ^ 1'b0 ;
  assign n8119 = n482 & n8118 ;
  assign n8120 = n382 & ~n627 ;
  assign n8121 = x97 & n8120 ;
  assign n8122 = ~n8119 & n8121 ;
  assign n8123 = ( n335 & ~n864 ) | ( n335 & n1662 ) | ( ~n864 & n1662 ) ;
  assign n8124 = n8123 ^ n2036 ^ 1'b0 ;
  assign n8125 = n2261 | n6881 ;
  assign n8126 = n918 & n1063 ;
  assign n8127 = n6718 & n8126 ;
  assign n8128 = ( n3653 & n4394 ) | ( n3653 & n8127 ) | ( n4394 & n8127 ) ;
  assign n8129 = n6145 & n8128 ;
  assign n8130 = ~n8125 & n8129 ;
  assign n8131 = ( n8122 & n8124 ) | ( n8122 & n8130 ) | ( n8124 & n8130 ) ;
  assign n8132 = n5332 ^ n4109 ^ n2761 ;
  assign n8133 = ( ~n3417 & n7097 ) | ( ~n3417 & n8132 ) | ( n7097 & n8132 ) ;
  assign n8134 = n8133 ^ n3778 ^ 1'b0 ;
  assign n8135 = n8134 ^ n7375 ^ 1'b0 ;
  assign n8136 = n5276 | n8135 ;
  assign n8145 = n3796 ^ n886 ^ 1'b0 ;
  assign n8140 = x62 & ~n3942 ;
  assign n8137 = ( n881 & n1411 ) | ( n881 & n1525 ) | ( n1411 & n1525 ) ;
  assign n8138 = n1030 | n8137 ;
  assign n8139 = x240 | n8138 ;
  assign n8141 = n8140 ^ n8139 ^ 1'b0 ;
  assign n8142 = ~n642 & n8141 ;
  assign n8143 = n8142 ^ n5573 ^ 1'b0 ;
  assign n8144 = ~n6018 & n8143 ;
  assign n8146 = n8145 ^ n8144 ^ 1'b0 ;
  assign n8147 = n7274 ^ n5521 ^ n3239 ;
  assign n8148 = n8147 ^ n406 ^ 1'b0 ;
  assign n8149 = ( n2486 & ~n3621 ) | ( n2486 & n7138 ) | ( ~n3621 & n7138 ) ;
  assign n8150 = n8149 ^ n3653 ^ 1'b0 ;
  assign n8151 = x94 & ~n8150 ;
  assign n8152 = n8151 ^ n5779 ^ n2132 ;
  assign n8153 = ( n912 & ~n1427 ) | ( n912 & n3016 ) | ( ~n1427 & n3016 ) ;
  assign n8154 = n2655 | n8153 ;
  assign n8155 = n5238 ^ n3420 ^ 1'b0 ;
  assign n8156 = n3878 ^ n2970 ^ n1787 ;
  assign n8157 = n6456 | n8156 ;
  assign n8158 = n8155 | n8157 ;
  assign n8159 = n3316 ^ n2905 ^ 1'b0 ;
  assign n8160 = n4123 ^ n1634 ^ 1'b0 ;
  assign n8161 = ~n5105 & n8160 ;
  assign n8162 = x55 & n8161 ;
  assign n8163 = n8162 ^ n8154 ^ n1090 ;
  assign n8164 = x129 & n256 ;
  assign n8165 = n8164 ^ n1337 ^ 1'b0 ;
  assign n8166 = ~n7564 & n8165 ;
  assign n8167 = n2755 & n8166 ;
  assign n8168 = n3080 ^ n2157 ^ 1'b0 ;
  assign n8169 = n2758 & n8168 ;
  assign n8170 = n8169 ^ x97 ^ 1'b0 ;
  assign n8171 = n3056 & ~n6340 ;
  assign n8172 = x195 | n1118 ;
  assign n8173 = n3704 & ~n8172 ;
  assign n8174 = n8173 ^ n1396 ^ 1'b0 ;
  assign n8175 = ( n5128 & n5435 ) | ( n5128 & ~n5593 ) | ( n5435 & ~n5593 ) ;
  assign n8176 = ~n1277 & n6844 ;
  assign n8177 = ~n8175 & n8176 ;
  assign n8178 = ( ~n6053 & n7086 ) | ( ~n6053 & n7635 ) | ( n7086 & n7635 ) ;
  assign n8179 = n7895 ^ n4984 ^ 1'b0 ;
  assign n8180 = n5574 ^ n4704 ^ n3629 ;
  assign n8181 = n8180 ^ n6341 ^ 1'b0 ;
  assign n8182 = n8179 & n8181 ;
  assign n8183 = n6597 ^ n4658 ^ n291 ;
  assign n8184 = n8183 ^ n2838 ^ n2655 ;
  assign n8185 = n508 | n5574 ;
  assign n8186 = ( ~n2939 & n8184 ) | ( ~n2939 & n8185 ) | ( n8184 & n8185 ) ;
  assign n8187 = n7526 ^ n6285 ^ n6241 ;
  assign n8190 = n8132 ^ n1906 ^ 1'b0 ;
  assign n8188 = n6171 ^ n3803 ^ n684 ;
  assign n8189 = n5693 & n8188 ;
  assign n8191 = n8190 ^ n8189 ^ 1'b0 ;
  assign n8192 = n2805 & n8191 ;
  assign n8193 = n8192 ^ n1493 ^ 1'b0 ;
  assign n8194 = n4777 & ~n8193 ;
  assign n8195 = n8174 ^ n3760 ^ n2472 ;
  assign n8200 = n1586 ^ x99 ^ 1'b0 ;
  assign n8197 = n2773 ^ n1325 ^ 1'b0 ;
  assign n8198 = n2161 | n8197 ;
  assign n8199 = ( n617 & ~n1444 ) | ( n617 & n8198 ) | ( ~n1444 & n8198 ) ;
  assign n8196 = ( n274 & n2110 ) | ( n274 & n3417 ) | ( n2110 & n3417 ) ;
  assign n8201 = n8200 ^ n8199 ^ n8196 ;
  assign n8202 = n2056 & ~n3292 ;
  assign n8203 = n8202 ^ x81 ^ 1'b0 ;
  assign n8204 = n2645 ^ n1501 ^ 1'b0 ;
  assign n8205 = n8204 ^ n2718 ^ 1'b0 ;
  assign n8206 = ( n4292 & n8203 ) | ( n4292 & n8205 ) | ( n8203 & n8205 ) ;
  assign n8207 = n6649 ^ n5097 ^ 1'b0 ;
  assign n8208 = n8206 & ~n8207 ;
  assign n8209 = n1458 & ~n7121 ;
  assign n8210 = n2475 | n2767 ;
  assign n8211 = n8210 ^ n3075 ^ 1'b0 ;
  assign n8213 = n3987 & ~n6115 ;
  assign n8214 = n8213 ^ n3996 ^ 1'b0 ;
  assign n8212 = n3521 ^ n2768 ^ 1'b0 ;
  assign n8215 = n8214 ^ n8212 ^ 1'b0 ;
  assign n8216 = n1037 & n2989 ;
  assign n8217 = ~n4218 & n8216 ;
  assign n8225 = n2438 ^ n2112 ^ 1'b0 ;
  assign n8218 = n2621 ^ n2368 ^ n2201 ;
  assign n8219 = ( n3050 & n5456 ) | ( n3050 & ~n7533 ) | ( n5456 & ~n7533 ) ;
  assign n8220 = ( ~n2530 & n7515 ) | ( ~n2530 & n8219 ) | ( n7515 & n8219 ) ;
  assign n8221 = n4720 & ~n7900 ;
  assign n8222 = n2800 & n8221 ;
  assign n8223 = ( n8218 & ~n8220 ) | ( n8218 & n8222 ) | ( ~n8220 & n8222 ) ;
  assign n8224 = n4366 & ~n8223 ;
  assign n8226 = n8225 ^ n8224 ^ 1'b0 ;
  assign n8227 = ( ~x58 & n614 ) | ( ~x58 & n3324 ) | ( n614 & n3324 ) ;
  assign n8228 = n8227 ^ n6964 ^ 1'b0 ;
  assign n8229 = n1155 & ~n8228 ;
  assign n8230 = n8226 & ~n8229 ;
  assign n8231 = ( n477 & n3521 ) | ( n477 & n4926 ) | ( n3521 & n4926 ) ;
  assign n8232 = n7683 ^ n3110 ^ 1'b0 ;
  assign n8233 = n8231 & n8232 ;
  assign n8234 = n8233 ^ n4454 ^ n2444 ;
  assign n8235 = n3833 ^ n3361 ^ n2482 ;
  assign n8236 = n8235 ^ n7462 ^ n3781 ;
  assign n8237 = n8236 ^ n6071 ^ n5639 ;
  assign n8238 = n736 & n5531 ;
  assign n8239 = ~n5872 & n8238 ;
  assign n8240 = n7540 ^ n6909 ^ n2063 ;
  assign n8243 = n1787 ^ n1078 ^ x210 ;
  assign n8244 = n8243 ^ n7761 ^ n6512 ;
  assign n8241 = n4369 ^ n2135 ^ 1'b0 ;
  assign n8242 = n8241 ^ n1403 ^ 1'b0 ;
  assign n8245 = n8244 ^ n8242 ^ n4478 ;
  assign n8246 = ~n967 & n2860 ;
  assign n8247 = n8246 ^ n2213 ^ 1'b0 ;
  assign n8248 = x225 & n6188 ;
  assign n8249 = ~n8247 & n8248 ;
  assign n8250 = n8249 ^ n5210 ^ n2328 ;
  assign n8251 = n8250 ^ n1790 ^ 1'b0 ;
  assign n8252 = n5645 | n8251 ;
  assign n8253 = n8245 | n8252 ;
  assign n8254 = n4775 ^ n3832 ^ 1'b0 ;
  assign n8255 = n7243 ^ n2710 ^ 1'b0 ;
  assign n8256 = ~n2573 & n8255 ;
  assign n8257 = ( n997 & n8254 ) | ( n997 & ~n8256 ) | ( n8254 & ~n8256 ) ;
  assign n8258 = ( n487 & n5063 ) | ( n487 & ~n8177 ) | ( n5063 & ~n8177 ) ;
  assign n8262 = ~n1800 & n3781 ;
  assign n8260 = ~n1006 & n3858 ;
  assign n8261 = n8260 ^ n7464 ^ 1'b0 ;
  assign n8263 = n8262 ^ n8261 ^ n5073 ;
  assign n8259 = n6251 ^ n5706 ^ 1'b0 ;
  assign n8264 = n8263 ^ n8259 ^ 1'b0 ;
  assign n8265 = n3009 | n8264 ;
  assign n8266 = n3766 & ~n8265 ;
  assign n8267 = n8266 ^ n7113 ^ 1'b0 ;
  assign n8268 = n2614 ^ n1989 ^ n480 ;
  assign n8269 = n8268 ^ n2913 ^ 1'b0 ;
  assign n8270 = ( ~n4976 & n5216 ) | ( ~n4976 & n8269 ) | ( n5216 & n8269 ) ;
  assign n8271 = ( n558 & n2217 ) | ( n558 & ~n6369 ) | ( n2217 & ~n6369 ) ;
  assign n8272 = n8271 ^ n8177 ^ n6725 ;
  assign n8273 = n2383 ^ x249 ^ 1'b0 ;
  assign n8274 = n1476 | n8273 ;
  assign n8275 = n8274 ^ n3068 ^ 1'b0 ;
  assign n8276 = n8275 ^ n8200 ^ n3534 ;
  assign n8277 = n834 | n1148 ;
  assign n8278 = n8276 | n8277 ;
  assign n8279 = ( n1924 & n2716 ) | ( n1924 & ~n2783 ) | ( n2716 & ~n2783 ) ;
  assign n8280 = n4037 | n8279 ;
  assign n8281 = n7079 ^ n6545 ^ n686 ;
  assign n8282 = n2608 ^ n607 ^ 1'b0 ;
  assign n8283 = ~n6128 & n7013 ;
  assign n8284 = ~n6138 & n8283 ;
  assign n8285 = ( n3142 & n6991 ) | ( n3142 & n8284 ) | ( n6991 & n8284 ) ;
  assign n8286 = ~n8282 & n8285 ;
  assign n8287 = n8286 ^ x199 ^ 1'b0 ;
  assign n8288 = n3175 & ~n8287 ;
  assign n8289 = n1474 ^ n1011 ^ 1'b0 ;
  assign n8290 = n8289 ^ n2704 ^ n2052 ;
  assign n8291 = n8290 ^ n2834 ^ n1223 ;
  assign n8292 = ( n2792 & ~n5463 ) | ( n2792 & n8291 ) | ( ~n5463 & n8291 ) ;
  assign n8293 = n8292 ^ n5969 ^ 1'b0 ;
  assign n8294 = ( n5165 & n5253 ) | ( n5165 & ~n6935 ) | ( n5253 & ~n6935 ) ;
  assign n8295 = n4260 ^ n2400 ^ 1'b0 ;
  assign n8296 = n758 & n8295 ;
  assign n8297 = ~n2192 & n4911 ;
  assign n8298 = ( n5401 & ~n6290 ) | ( n5401 & n8297 ) | ( ~n6290 & n8297 ) ;
  assign n8299 = n7801 ^ n4504 ^ n544 ;
  assign n8300 = ~n7081 & n8299 ;
  assign n8301 = ~n8298 & n8300 ;
  assign n8302 = n3356 ^ n1726 ^ 1'b0 ;
  assign n8303 = n2745 | n8302 ;
  assign n8304 = n5610 | n8303 ;
  assign n8305 = n842 & n1816 ;
  assign n8306 = n8305 ^ n6746 ^ 1'b0 ;
  assign n8307 = n5503 ^ n3100 ^ 1'b0 ;
  assign n8308 = n8307 ^ n6082 ^ 1'b0 ;
  assign n8309 = n8306 & ~n8308 ;
  assign n8312 = n2206 ^ n1875 ^ x22 ;
  assign n8311 = n562 | n5425 ;
  assign n8313 = n8312 ^ n8311 ^ n5300 ;
  assign n8310 = ~n3430 & n3904 ;
  assign n8314 = n8313 ^ n8310 ^ 1'b0 ;
  assign n8315 = ~n835 & n7164 ;
  assign n8316 = n8315 ^ n7198 ^ 1'b0 ;
  assign n8317 = n2354 ^ n1166 ^ n884 ;
  assign n8318 = ( n838 & n895 ) | ( n838 & ~n6623 ) | ( n895 & ~n6623 ) ;
  assign n8319 = ( ~n6701 & n8317 ) | ( ~n6701 & n8318 ) | ( n8317 & n8318 ) ;
  assign n8320 = n2820 & n4998 ;
  assign n8322 = n5992 ^ n2461 ^ 1'b0 ;
  assign n8323 = n2704 | n8322 ;
  assign n8324 = x32 | n8323 ;
  assign n8321 = ( n2009 & ~n6754 ) | ( n2009 & n7392 ) | ( ~n6754 & n7392 ) ;
  assign n8325 = n8324 ^ n8321 ^ n7611 ;
  assign n8326 = n3279 & ~n4540 ;
  assign n8327 = n1881 & ~n8326 ;
  assign n8328 = ( x177 & n6249 ) | ( x177 & n8327 ) | ( n6249 & n8327 ) ;
  assign n8329 = ~n3219 & n3888 ;
  assign n8330 = n8329 ^ n5309 ^ 1'b0 ;
  assign n8331 = n8330 ^ n5000 ^ n969 ;
  assign n8332 = n713 | n8331 ;
  assign n8333 = ~n1365 & n2925 ;
  assign n8334 = n7015 ^ n816 ^ 1'b0 ;
  assign n8335 = ( ~n8140 & n8333 ) | ( ~n8140 & n8334 ) | ( n8333 & n8334 ) ;
  assign n8336 = ( n6707 & ~n7761 ) | ( n6707 & n8335 ) | ( ~n7761 & n8335 ) ;
  assign n8338 = x3 & n6225 ;
  assign n8339 = n8338 ^ n5680 ^ 1'b0 ;
  assign n8340 = n8339 ^ n6224 ^ 1'b0 ;
  assign n8337 = n5730 ^ n4501 ^ n3655 ;
  assign n8341 = n8340 ^ n8337 ^ n6222 ;
  assign n8342 = ~n2808 & n3126 ;
  assign n8343 = ~n3319 & n8342 ;
  assign n8344 = ~n2001 & n4856 ;
  assign n8345 = n5086 ^ n3296 ^ n3155 ;
  assign n8346 = n1859 & ~n4805 ;
  assign n8347 = n3983 ^ n3434 ^ 1'b0 ;
  assign n8348 = ~n8346 & n8347 ;
  assign n8349 = n7637 ^ n2445 ^ 1'b0 ;
  assign n8350 = n6101 | n8349 ;
  assign n8351 = n3753 | n5015 ;
  assign n8352 = n8351 ^ n3816 ^ 1'b0 ;
  assign n8353 = n4789 ^ n2821 ^ 1'b0 ;
  assign n8354 = n6435 & ~n8353 ;
  assign n8355 = ( n426 & n2519 ) | ( n426 & ~n8354 ) | ( n2519 & ~n8354 ) ;
  assign n8356 = n1969 & n4724 ;
  assign n8357 = ~n5086 & n8356 ;
  assign n8358 = n7783 | n8357 ;
  assign n8359 = n7142 ^ n5306 ^ n4556 ;
  assign n8360 = ~n5979 & n7972 ;
  assign n8361 = n8360 ^ n4758 ^ 1'b0 ;
  assign n8362 = ( x29 & n3754 ) | ( x29 & ~n8361 ) | ( n3754 & ~n8361 ) ;
  assign n8363 = n8362 ^ n1318 ^ 1'b0 ;
  assign n8364 = n5204 & ~n7522 ;
  assign n8365 = n8364 ^ n7283 ^ 1'b0 ;
  assign n8372 = n376 | n2659 ;
  assign n8373 = n8372 ^ n2464 ^ 1'b0 ;
  assign n8366 = n2177 | n7609 ;
  assign n8367 = n3042 | n8366 ;
  assign n8368 = n8367 ^ n7721 ^ n280 ;
  assign n8369 = n8368 ^ n2561 ^ 1'b0 ;
  assign n8370 = ( n3762 & ~n7485 ) | ( n3762 & n8369 ) | ( ~n7485 & n8369 ) ;
  assign n8371 = n7373 & n8370 ;
  assign n8374 = n8373 ^ n8371 ^ 1'b0 ;
  assign n8375 = n8374 ^ n4060 ^ n1854 ;
  assign n8376 = n7285 ^ n2738 ^ 1'b0 ;
  assign n8377 = ( n4169 & ~n4466 ) | ( n4169 & n8019 ) | ( ~n4466 & n8019 ) ;
  assign n8378 = n8227 & ~n8377 ;
  assign n8379 = n8378 ^ n1111 ^ 1'b0 ;
  assign n8380 = n8379 ^ n8122 ^ n6037 ;
  assign n8381 = n8380 ^ n488 ^ 1'b0 ;
  assign n8382 = n8156 ^ n2377 ^ 1'b0 ;
  assign n8383 = ( n1683 & n4544 ) | ( n1683 & n8382 ) | ( n4544 & n8382 ) ;
  assign n8384 = ~n5049 & n8383 ;
  assign n8385 = n2558 | n6525 ;
  assign n8386 = n4443 | n8385 ;
  assign n8387 = n8386 ^ n6937 ^ 1'b0 ;
  assign n8388 = n2374 ^ n1975 ^ 1'b0 ;
  assign n8389 = n5461 & ~n8388 ;
  assign n8390 = n8389 ^ n5658 ^ n1487 ;
  assign n8391 = ~n2934 & n3452 ;
  assign n8392 = n8391 ^ n1784 ^ 1'b0 ;
  assign n8393 = ( n1678 & n8390 ) | ( n1678 & ~n8392 ) | ( n8390 & ~n8392 ) ;
  assign n8394 = n3246 & n8393 ;
  assign n8395 = n4209 & ~n8172 ;
  assign n8396 = n6624 & n8395 ;
  assign n8397 = n8396 ^ n2807 ^ 1'b0 ;
  assign n8398 = ( n1623 & ~n4165 ) | ( n1623 & n6445 ) | ( ~n4165 & n6445 ) ;
  assign n8399 = n8397 & ~n8398 ;
  assign n8400 = n632 & ~n8399 ;
  assign n8401 = ~n758 & n8400 ;
  assign n8402 = ~n4163 & n5017 ;
  assign n8404 = n4958 ^ n1166 ^ 1'b0 ;
  assign n8405 = n4007 | n8404 ;
  assign n8406 = ~x22 & x184 ;
  assign n8407 = n3939 & n4897 ;
  assign n8408 = ~n6876 & n8407 ;
  assign n8409 = ( n3049 & n8406 ) | ( n3049 & n8408 ) | ( n8406 & n8408 ) ;
  assign n8410 = ( ~n6404 & n8405 ) | ( ~n6404 & n8409 ) | ( n8405 & n8409 ) ;
  assign n8403 = ( x93 & ~n578 ) | ( x93 & n3598 ) | ( ~n578 & n3598 ) ;
  assign n8411 = n8410 ^ n8403 ^ n6194 ;
  assign n8412 = ( n1721 & n5599 ) | ( n1721 & ~n8357 ) | ( n5599 & ~n8357 ) ;
  assign n8413 = n2031 & ~n2963 ;
  assign n8414 = ~n2663 & n6732 ;
  assign n8415 = n8414 ^ n5233 ^ 1'b0 ;
  assign n8416 = ~n3050 & n8415 ;
  assign n8417 = n5604 ^ n4335 ^ 1'b0 ;
  assign n8418 = n5687 & n8417 ;
  assign n8419 = ( ~x34 & n8416 ) | ( ~x34 & n8418 ) | ( n8416 & n8418 ) ;
  assign n8420 = ~n3607 & n8419 ;
  assign n8421 = ~n8413 & n8420 ;
  assign n8422 = n6131 & ~n7042 ;
  assign n8424 = ( x248 & ~n3254 ) | ( x248 & n6589 ) | ( ~n3254 & n6589 ) ;
  assign n8423 = ( n297 & n2322 ) | ( n297 & ~n2557 ) | ( n2322 & ~n2557 ) ;
  assign n8425 = n8424 ^ n8423 ^ 1'b0 ;
  assign n8426 = n6908 ^ n5054 ^ 1'b0 ;
  assign n8433 = n3696 ^ x25 ^ 1'b0 ;
  assign n8434 = n8433 ^ n5634 ^ 1'b0 ;
  assign n8435 = ~n3366 & n8434 ;
  assign n8428 = n7770 ^ n4611 ^ 1'b0 ;
  assign n8429 = n1995 & ~n8428 ;
  assign n8427 = n1438 & n2107 ;
  assign n8430 = n8429 ^ n8427 ^ n645 ;
  assign n8431 = n898 & ~n6901 ;
  assign n8432 = n8430 | n8431 ;
  assign n8436 = n8435 ^ n8432 ^ 1'b0 ;
  assign n8437 = n3175 ^ n963 ^ x120 ;
  assign n8438 = n8437 ^ n1284 ^ n832 ;
  assign n8439 = n5111 & ~n7261 ;
  assign n8440 = n8438 & n8439 ;
  assign n8441 = n8440 ^ n6564 ^ n1740 ;
  assign n8442 = n3465 ^ n258 ^ x188 ;
  assign n8443 = n7261 | n8442 ;
  assign n8444 = n7978 & ~n8443 ;
  assign n8445 = n3487 & ~n4692 ;
  assign n8446 = n1049 & n8445 ;
  assign n8447 = n4812 & n8446 ;
  assign n8448 = n8447 ^ n3117 ^ n1560 ;
  assign n8449 = ~n1688 & n5356 ;
  assign n8450 = ~n4364 & n6014 ;
  assign n8451 = ~n3967 & n4678 ;
  assign n8452 = ~n8450 & n8451 ;
  assign n8453 = n6553 & n6680 ;
  assign n8454 = n616 & ~n637 ;
  assign n8455 = n8454 ^ n3273 ^ 1'b0 ;
  assign n8456 = ( n3563 & n6511 ) | ( n3563 & ~n8455 ) | ( n6511 & ~n8455 ) ;
  assign n8457 = n8456 ^ x55 ^ 1'b0 ;
  assign n8458 = ( n8452 & n8453 ) | ( n8452 & ~n8457 ) | ( n8453 & ~n8457 ) ;
  assign n8459 = ~n3707 & n4719 ;
  assign n8460 = n8459 ^ n4112 ^ 1'b0 ;
  assign n8461 = n4143 | n8460 ;
  assign n8462 = n4781 ^ n4160 ^ n3720 ;
  assign n8463 = n4838 ^ n2041 ^ x39 ;
  assign n8464 = n8463 ^ n5682 ^ 1'b0 ;
  assign n8467 = n1840 & n4224 ;
  assign n8468 = ~n8011 & n8467 ;
  assign n8465 = ( n946 & n4701 ) | ( n946 & n7696 ) | ( n4701 & n7696 ) ;
  assign n8466 = n4312 | n8465 ;
  assign n8469 = n8468 ^ n8466 ^ 1'b0 ;
  assign n8470 = n4095 ^ n1256 ^ n1135 ;
  assign n8471 = n6184 ^ n2811 ^ 1'b0 ;
  assign n8472 = n3431 & ~n8471 ;
  assign n8473 = x7 & ~n7921 ;
  assign n8474 = ~n8472 & n8473 ;
  assign n8475 = ( ~n6060 & n8470 ) | ( ~n6060 & n8474 ) | ( n8470 & n8474 ) ;
  assign n8482 = n3750 ^ n1588 ^ 1'b0 ;
  assign n8483 = ( x227 & n6107 ) | ( x227 & n8482 ) | ( n6107 & n8482 ) ;
  assign n8476 = n2643 ^ n2562 ^ 1'b0 ;
  assign n8477 = n4970 & ~n8476 ;
  assign n8478 = n8165 ^ n789 ^ x104 ;
  assign n8479 = n8478 ^ n1120 ^ 1'b0 ;
  assign n8480 = n8477 & ~n8479 ;
  assign n8481 = ~n5791 & n8480 ;
  assign n8484 = n8483 ^ n8481 ^ 1'b0 ;
  assign n8485 = n5157 ^ n2017 ^ 1'b0 ;
  assign n8486 = n6359 & ~n8485 ;
  assign n8487 = n2793 & ~n3478 ;
  assign n8488 = n1467 ^ n1127 ^ n947 ;
  assign n8489 = n2834 & n8488 ;
  assign n8490 = ~n8487 & n8489 ;
  assign n8491 = n8257 ^ n6823 ^ 1'b0 ;
  assign n8492 = n813 & n8491 ;
  assign n8493 = n7165 ^ n3717 ^ n2781 ;
  assign n8494 = ( n952 & n2213 ) | ( n952 & ~n4298 ) | ( n2213 & ~n4298 ) ;
  assign n8495 = n8494 ^ n3038 ^ n675 ;
  assign n8496 = n8495 ^ n1464 ^ n929 ;
  assign n8497 = n5082 ^ x219 ^ 1'b0 ;
  assign n8498 = n4529 ^ n3472 ^ 1'b0 ;
  assign n8499 = n8498 ^ n500 ^ 1'b0 ;
  assign n8500 = n8497 & ~n8499 ;
  assign n8501 = n331 & ~n6335 ;
  assign n8502 = n5264 & n8501 ;
  assign n8503 = ( n3632 & n7282 ) | ( n3632 & ~n8502 ) | ( n7282 & ~n8502 ) ;
  assign n8504 = n8503 ^ n4032 ^ n2599 ;
  assign n8509 = n6176 ^ n5669 ^ 1'b0 ;
  assign n8505 = n3532 & n3727 ;
  assign n8506 = n8505 ^ n1926 ^ 1'b0 ;
  assign n8507 = n3594 & n8506 ;
  assign n8508 = n3327 & n8507 ;
  assign n8510 = n8509 ^ n8508 ^ n2158 ;
  assign n8511 = n8510 ^ n1405 ^ 1'b0 ;
  assign n8512 = n4331 & n8511 ;
  assign n8513 = ( n566 & n1461 ) | ( n566 & ~n1844 ) | ( n1461 & ~n1844 ) ;
  assign n8514 = ( ~x166 & n1625 ) | ( ~x166 & n8513 ) | ( n1625 & n8513 ) ;
  assign n8515 = n5958 ^ n636 ^ 1'b0 ;
  assign n8516 = n8515 ^ n7151 ^ 1'b0 ;
  assign n8517 = n8514 & n8516 ;
  assign n8518 = n6996 ^ n6076 ^ x102 ;
  assign n8519 = n4712 & n8518 ;
  assign n8520 = n7088 ^ n5238 ^ x54 ;
  assign n8521 = n764 & n8520 ;
  assign n8522 = n8521 ^ n1958 ^ 1'b0 ;
  assign n8523 = ~n1521 & n5420 ;
  assign n8524 = n2887 & ~n4837 ;
  assign n8525 = n3382 & n8524 ;
  assign n8526 = n6129 ^ n4803 ^ 1'b0 ;
  assign n8527 = ~n2721 & n8526 ;
  assign n8528 = n1888 ^ n1216 ^ 1'b0 ;
  assign n8529 = n758 | n8528 ;
  assign n8530 = ( n686 & n8527 ) | ( n686 & ~n8529 ) | ( n8527 & ~n8529 ) ;
  assign n8531 = ~n8525 & n8530 ;
  assign n8532 = ~n1861 & n2321 ;
  assign n8533 = n8532 ^ n1425 ^ 1'b0 ;
  assign n8534 = ~n2028 & n8533 ;
  assign n8535 = x50 | n8534 ;
  assign n8536 = ( n321 & n2175 ) | ( n321 & n5797 ) | ( n2175 & n5797 ) ;
  assign n8537 = n8536 ^ n3516 ^ n1372 ;
  assign n8538 = n8537 ^ n5418 ^ n2064 ;
  assign n8539 = ( n4997 & ~n5326 ) | ( n4997 & n8538 ) | ( ~n5326 & n8538 ) ;
  assign n8540 = n8539 ^ n3180 ^ n3083 ;
  assign n8541 = n5857 ^ n2325 ^ x131 ;
  assign n8544 = n7163 ^ n6460 ^ 1'b0 ;
  assign n8545 = x142 & ~n8544 ;
  assign n8543 = ~x183 & n1953 ;
  assign n8542 = ( n2999 & ~n4830 ) | ( n2999 & n8498 ) | ( ~n4830 & n8498 ) ;
  assign n8546 = n8545 ^ n8543 ^ n8542 ;
  assign n8549 = n2434 & n4770 ;
  assign n8547 = n1564 & ~n8290 ;
  assign n8548 = ~n5535 & n8547 ;
  assign n8550 = n8549 ^ n8548 ^ n1312 ;
  assign n8551 = n287 | n5226 ;
  assign n8552 = n2749 & n8551 ;
  assign n8553 = n4258 & n8552 ;
  assign n8554 = n8553 ^ n4518 ^ 1'b0 ;
  assign n8555 = n2807 & ~n6640 ;
  assign n8558 = ( x239 & n2280 ) | ( x239 & n5610 ) | ( n2280 & n5610 ) ;
  assign n8559 = n8558 ^ n7808 ^ 1'b0 ;
  assign n8556 = ( ~n331 & n818 ) | ( ~n331 & n5050 ) | ( n818 & n5050 ) ;
  assign n8557 = ( ~n2869 & n4620 ) | ( ~n2869 & n8556 ) | ( n4620 & n8556 ) ;
  assign n8560 = n8559 ^ n8557 ^ 1'b0 ;
  assign n8561 = ( ~n1136 & n8555 ) | ( ~n1136 & n8560 ) | ( n8555 & n8560 ) ;
  assign n8564 = ( x235 & ~n1342 ) | ( x235 & n1393 ) | ( ~n1342 & n1393 ) ;
  assign n8562 = n1353 ^ n806 ^ 1'b0 ;
  assign n8563 = x12 & n8562 ;
  assign n8565 = n8564 ^ n8563 ^ 1'b0 ;
  assign n8566 = n8244 ^ n5899 ^ 1'b0 ;
  assign n8567 = ( n919 & ~n3382 ) | ( n919 & n8566 ) | ( ~n3382 & n8566 ) ;
  assign n8568 = n8396 ^ n7561 ^ 1'b0 ;
  assign n8569 = n7064 ^ n1986 ^ x244 ;
  assign n8570 = n2880 | n8569 ;
  assign n8571 = n8570 ^ n5309 ^ 1'b0 ;
  assign n8572 = n1798 & ~n8571 ;
  assign n8573 = n8572 ^ n2858 ^ 1'b0 ;
  assign n8574 = n4132 ^ n2714 ^ n1739 ;
  assign n8576 = n6889 ^ n3271 ^ 1'b0 ;
  assign n8577 = n1438 & n8576 ;
  assign n8575 = ~x159 & n3096 ;
  assign n8578 = n8577 ^ n8575 ^ 1'b0 ;
  assign n8579 = n6462 ^ n4087 ^ 1'b0 ;
  assign n8580 = ( ~n7752 & n8578 ) | ( ~n7752 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8581 = n2684 ^ n2547 ^ 1'b0 ;
  assign n8582 = ( ~n2854 & n4190 ) | ( ~n2854 & n6486 ) | ( n4190 & n6486 ) ;
  assign n8583 = ~n933 & n1503 ;
  assign n8584 = ~x192 & n8583 ;
  assign n8585 = ( n1197 & n1828 ) | ( n1197 & n8584 ) | ( n1828 & n8584 ) ;
  assign n8586 = ( n4542 & ~n7613 ) | ( n4542 & n7852 ) | ( ~n7613 & n7852 ) ;
  assign n8587 = n7333 & ~n8586 ;
  assign n8588 = ~n8585 & n8587 ;
  assign n8589 = n8588 ^ n8335 ^ 1'b0 ;
  assign n8593 = n7236 ^ n2246 ^ 1'b0 ;
  assign n8591 = n5457 ^ n3655 ^ n3038 ;
  assign n8592 = n3639 & ~n8591 ;
  assign n8594 = n8593 ^ n8592 ^ 1'b0 ;
  assign n8590 = x77 & ~n4060 ;
  assign n8595 = n8594 ^ n8590 ^ 1'b0 ;
  assign n8596 = n3949 ^ n3512 ^ 1'b0 ;
  assign n8597 = n5097 & n8596 ;
  assign n8598 = n8597 ^ n1779 ^ 1'b0 ;
  assign n8599 = n4961 ^ n2035 ^ 1'b0 ;
  assign n8600 = n8187 ^ n5836 ^ n4102 ;
  assign n8601 = ( n4617 & n8599 ) | ( n4617 & n8600 ) | ( n8599 & n8600 ) ;
  assign n8602 = n3844 ^ x109 ^ 1'b0 ;
  assign n8603 = ~n7255 & n8602 ;
  assign n8604 = n2714 ^ n1297 ^ x2 ;
  assign n8605 = n2289 ^ n1650 ^ n1414 ;
  assign n8606 = n8605 ^ n7511 ^ n2985 ;
  assign n8607 = ( n3633 & n8604 ) | ( n3633 & n8606 ) | ( n8604 & n8606 ) ;
  assign n8608 = n8607 ^ n2406 ^ 1'b0 ;
  assign n8609 = ~n3298 & n7092 ;
  assign n8610 = n8608 & n8609 ;
  assign n8614 = n1784 | n2746 ;
  assign n8615 = n7422 | n8614 ;
  assign n8616 = n4816 & n8615 ;
  assign n8611 = n1855 | n5238 ;
  assign n8612 = n4444 | n8611 ;
  assign n8613 = n8612 ^ n3457 ^ n1703 ;
  assign n8617 = n8616 ^ n8613 ^ n4601 ;
  assign n8618 = n4970 ^ n2167 ^ 1'b0 ;
  assign n8619 = ( n1356 & n3578 ) | ( n1356 & ~n8618 ) | ( n3578 & ~n8618 ) ;
  assign n8620 = n1560 ^ n1488 ^ n677 ;
  assign n8621 = n1920 & ~n8620 ;
  assign n8626 = n2738 ^ n2458 ^ n1973 ;
  assign n8622 = n1913 & n7586 ;
  assign n8623 = n4501 ^ n269 ^ 1'b0 ;
  assign n8624 = ~n8622 & n8623 ;
  assign n8625 = ~n733 & n8624 ;
  assign n8627 = n8626 ^ n8625 ^ 1'b0 ;
  assign n8628 = n4533 & n8627 ;
  assign n8629 = ~n8621 & n8628 ;
  assign n8630 = n8629 ^ n7850 ^ 1'b0 ;
  assign n8631 = ( x46 & n8619 ) | ( x46 & n8630 ) | ( n8619 & n8630 ) ;
  assign n8632 = n7600 ^ n4801 ^ n2135 ;
  assign n8635 = n6035 ^ n3894 ^ n2009 ;
  assign n8633 = n402 | n3167 ;
  assign n8634 = n7357 | n8633 ;
  assign n8636 = n8635 ^ n8634 ^ 1'b0 ;
  assign n8637 = n2273 | n8636 ;
  assign n8638 = n2045 & n3019 ;
  assign n8639 = n8638 ^ n284 ^ 1'b0 ;
  assign n8640 = n8637 | n8639 ;
  assign n8641 = n8640 ^ n4577 ^ n2391 ;
  assign n8642 = ( n282 & ~n666 ) | ( n282 & n2293 ) | ( ~n666 & n2293 ) ;
  assign n8643 = n2027 ^ n1220 ^ 1'b0 ;
  assign n8644 = n3089 & ~n8643 ;
  assign n8645 = ( n6184 & n8642 ) | ( n6184 & n8644 ) | ( n8642 & n8644 ) ;
  assign n8646 = n5466 ^ n868 ^ n320 ;
  assign n8647 = n8645 | n8646 ;
  assign n8648 = n5189 ^ n4359 ^ n1697 ;
  assign n8649 = n7274 ^ n4912 ^ 1'b0 ;
  assign n8674 = x12 & n3785 ;
  assign n8675 = n8674 ^ n617 ^ 1'b0 ;
  assign n8676 = n3169 ^ n2063 ^ 1'b0 ;
  assign n8677 = n8675 & ~n8676 ;
  assign n8658 = n3388 ^ n2065 ^ n378 ;
  assign n8659 = n6375 ^ x112 ^ 1'b0 ;
  assign n8660 = n4006 ^ n2513 ^ n2287 ;
  assign n8661 = ~n272 & n4093 ;
  assign n8662 = ~n2655 & n8661 ;
  assign n8665 = n4935 | n5470 ;
  assign n8666 = n1591 & ~n8665 ;
  assign n8663 = n2881 ^ n2367 ^ 1'b0 ;
  assign n8664 = ~n2001 & n8663 ;
  assign n8667 = n8666 ^ n8664 ^ 1'b0 ;
  assign n8668 = n6136 | n6748 ;
  assign n8669 = n8667 | n8668 ;
  assign n8670 = ( n8660 & ~n8662 ) | ( n8660 & n8669 ) | ( ~n8662 & n8669 ) ;
  assign n8671 = ( n4707 & n8659 ) | ( n4707 & n8670 ) | ( n8659 & n8670 ) ;
  assign n8672 = n8658 | n8671 ;
  assign n8673 = n8672 ^ n2178 ^ 1'b0 ;
  assign n8650 = n5201 & ~n5516 ;
  assign n8651 = ~n374 & n8650 ;
  assign n8654 = ~n3133 & n8317 ;
  assign n8655 = n4332 & n8654 ;
  assign n8652 = ( n901 & n1430 ) | ( n901 & ~n1975 ) | ( n1430 & ~n1975 ) ;
  assign n8653 = n8652 ^ n4026 ^ 1'b0 ;
  assign n8656 = n8655 ^ n8653 ^ 1'b0 ;
  assign n8657 = ~n8651 & n8656 ;
  assign n8678 = n8677 ^ n8673 ^ n8657 ;
  assign n8679 = n637 | n834 ;
  assign n8680 = n6998 | n8679 ;
  assign n8684 = n1700 & ~n3318 ;
  assign n8685 = n4116 & n8684 ;
  assign n8681 = ~n2216 & n3844 ;
  assign n8682 = ~n4383 & n6517 ;
  assign n8683 = ~n8681 & n8682 ;
  assign n8686 = n8685 ^ n8683 ^ n7552 ;
  assign n8687 = x213 & n2957 ;
  assign n8688 = n8687 ^ n2765 ^ 1'b0 ;
  assign n8689 = ~x83 & x88 ;
  assign n8690 = n3184 | n8689 ;
  assign n8691 = n8688 | n8690 ;
  assign n8692 = n8691 ^ n7061 ^ n4463 ;
  assign n8693 = n1582 | n8692 ;
  assign n8694 = n8693 ^ n7619 ^ 1'b0 ;
  assign n8695 = ( n877 & n6311 ) | ( n877 & ~n8694 ) | ( n6311 & ~n8694 ) ;
  assign n8697 = n2573 & n6816 ;
  assign n8696 = n1961 & ~n6533 ;
  assign n8698 = n8697 ^ n8696 ^ 1'b0 ;
  assign n8699 = ( x134 & n3272 ) | ( x134 & n8698 ) | ( n3272 & n8698 ) ;
  assign n8700 = x6 & n7194 ;
  assign n8702 = ~n1396 & n5461 ;
  assign n8701 = n1184 & ~n4288 ;
  assign n8703 = n8702 ^ n8701 ^ n5680 ;
  assign n8704 = n8700 & n8703 ;
  assign n8705 = n7617 ^ n1578 ^ 1'b0 ;
  assign n8706 = n5492 ^ n4386 ^ 1'b0 ;
  assign n8707 = ( x215 & n1425 ) | ( x215 & ~n1573 ) | ( n1425 & ~n1573 ) ;
  assign n8708 = ( n804 & n2592 ) | ( n804 & n8707 ) | ( n2592 & n8707 ) ;
  assign n8709 = ( n3587 & ~n4949 ) | ( n3587 & n8708 ) | ( ~n4949 & n8708 ) ;
  assign n8710 = ( n5065 & n6438 ) | ( n5065 & ~n8709 ) | ( n6438 & ~n8709 ) ;
  assign n8711 = n6339 & ~n8710 ;
  assign n8712 = ( n7983 & n8706 ) | ( n7983 & ~n8711 ) | ( n8706 & ~n8711 ) ;
  assign n8713 = ( n8170 & ~n8705 ) | ( n8170 & n8712 ) | ( ~n8705 & n8712 ) ;
  assign n8714 = n1497 & n2441 ;
  assign n8715 = n8714 ^ n5797 ^ 1'b0 ;
  assign n8716 = ( n461 & ~n1175 ) | ( n461 & n8715 ) | ( ~n1175 & n8715 ) ;
  assign n8717 = n8716 ^ n4088 ^ n277 ;
  assign n8718 = ( n4152 & ~n6076 ) | ( n4152 & n8717 ) | ( ~n6076 & n8717 ) ;
  assign n8719 = n3509 ^ n1392 ^ 1'b0 ;
  assign n8720 = n5513 ^ n2408 ^ 1'b0 ;
  assign n8721 = n5964 | n8720 ;
  assign n8722 = ~n787 & n1447 ;
  assign n8723 = ~n1554 & n8722 ;
  assign n8724 = ( n1083 & ~n4730 ) | ( n1083 & n8723 ) | ( ~n4730 & n8723 ) ;
  assign n8725 = ( n2794 & ~n3968 ) | ( n2794 & n8579 ) | ( ~n3968 & n8579 ) ;
  assign n8728 = n1703 ^ n1383 ^ 1'b0 ;
  assign n8729 = n1671 | n8728 ;
  assign n8730 = ( ~n874 & n1975 ) | ( ~n874 & n8729 ) | ( n1975 & n8729 ) ;
  assign n8731 = ( n1655 & ~n4189 ) | ( n1655 & n8730 ) | ( ~n4189 & n8730 ) ;
  assign n8726 = n8103 ^ n3735 ^ n1226 ;
  assign n8727 = n8726 ^ n6554 ^ n4461 ;
  assign n8732 = n8731 ^ n8727 ^ n8384 ;
  assign n8733 = ( ~n1033 & n2737 ) | ( ~n1033 & n5372 ) | ( n2737 & n5372 ) ;
  assign n8742 = n6290 | n7734 ;
  assign n8743 = n8742 ^ n6887 ^ 1'b0 ;
  assign n8734 = ( x241 & n1786 ) | ( x241 & n4871 ) | ( n1786 & n4871 ) ;
  assign n8736 = n618 & ~n1818 ;
  assign n8737 = n8736 ^ n4609 ^ 1'b0 ;
  assign n8735 = n2308 ^ x160 ^ 1'b0 ;
  assign n8738 = n8737 ^ n8735 ^ 1'b0 ;
  assign n8739 = n7897 & ~n8738 ;
  assign n8740 = n8739 ^ n3501 ^ 1'b0 ;
  assign n8741 = ( n1719 & ~n8734 ) | ( n1719 & n8740 ) | ( ~n8734 & n8740 ) ;
  assign n8744 = n8743 ^ n8741 ^ 1'b0 ;
  assign n8745 = n4224 ^ n2326 ^ 1'b0 ;
  assign n8746 = n5322 ^ n2503 ^ 1'b0 ;
  assign n8747 = n2236 | n8746 ;
  assign n8748 = n2213 | n8747 ;
  assign n8749 = n8745 & ~n8748 ;
  assign n8754 = n355 & ~n1301 ;
  assign n8755 = n5169 | n5979 ;
  assign n8756 = n435 | n8755 ;
  assign n8757 = ( ~n2944 & n8754 ) | ( ~n2944 & n8756 ) | ( n8754 & n8756 ) ;
  assign n8750 = x167 & n908 ;
  assign n8751 = n1922 & n8750 ;
  assign n8752 = ( n2092 & n7327 ) | ( n2092 & n8751 ) | ( n7327 & n8751 ) ;
  assign n8753 = n2143 & ~n8752 ;
  assign n8758 = n8757 ^ n8753 ^ 1'b0 ;
  assign n8761 = x69 & ~n5592 ;
  assign n8762 = n8761 ^ n4165 ^ 1'b0 ;
  assign n8763 = n6843 | n8762 ;
  assign n8759 = n6856 & ~n7771 ;
  assign n8760 = ~n3144 & n8759 ;
  assign n8764 = n8763 ^ n8760 ^ n2217 ;
  assign n8765 = n4068 | n8764 ;
  assign n8766 = n8765 ^ n3487 ^ 1'b0 ;
  assign n8767 = n8766 ^ n4276 ^ 1'b0 ;
  assign n8768 = n473 & n1315 ;
  assign n8769 = ( ~n2440 & n6121 ) | ( ~n2440 & n8768 ) | ( n6121 & n8768 ) ;
  assign n8775 = x143 & ~n8644 ;
  assign n8770 = ~n336 & n2400 ;
  assign n8771 = ~n5953 & n7057 ;
  assign n8772 = n8770 & ~n8771 ;
  assign n8773 = n8772 ^ n3818 ^ 1'b0 ;
  assign n8774 = n5140 | n8773 ;
  assign n8776 = n8775 ^ n8774 ^ n683 ;
  assign n8777 = n7724 ^ n731 ^ 1'b0 ;
  assign n8778 = ( n6612 & n6669 ) | ( n6612 & n7085 ) | ( n6669 & n7085 ) ;
  assign n8779 = n5843 ^ n3337 ^ 1'b0 ;
  assign n8780 = ( ~n7658 & n8326 ) | ( ~n7658 & n8779 ) | ( n8326 & n8779 ) ;
  assign n8781 = ( n491 & n6977 ) | ( n491 & ~n7126 ) | ( n6977 & ~n7126 ) ;
  assign n8782 = n8563 ^ n1400 ^ 1'b0 ;
  assign n8783 = ~n3456 & n8782 ;
  assign n8784 = ~n8781 & n8783 ;
  assign n8785 = n8784 ^ n7030 ^ 1'b0 ;
  assign n8786 = n1588 ^ x248 ^ 1'b0 ;
  assign n8787 = ( x59 & n2904 ) | ( x59 & ~n8786 ) | ( n2904 & ~n8786 ) ;
  assign n8788 = n1267 | n2858 ;
  assign n8789 = n2963 | n8788 ;
  assign n8790 = n8789 ^ n3250 ^ n1852 ;
  assign n8791 = ( n1221 & ~n2167 ) | ( n1221 & n8790 ) | ( ~n2167 & n8790 ) ;
  assign n8792 = n6409 ^ n3960 ^ n3857 ;
  assign n8793 = ( x160 & n8731 ) | ( x160 & n8792 ) | ( n8731 & n8792 ) ;
  assign n8794 = n3799 | n3826 ;
  assign n8795 = n8794 ^ n3669 ^ 1'b0 ;
  assign n8796 = n8795 ^ n7410 ^ 1'b0 ;
  assign n8797 = x43 & ~n8796 ;
  assign n8800 = ( n2828 & ~n6771 ) | ( n2828 & n7230 ) | ( ~n6771 & n7230 ) ;
  assign n8798 = n8122 ^ n925 ^ 1'b0 ;
  assign n8799 = ~n4847 & n8798 ;
  assign n8801 = n8800 ^ n8799 ^ 1'b0 ;
  assign n8802 = ( n291 & n548 ) | ( n291 & n4805 ) | ( n548 & n4805 ) ;
  assign n8803 = ( ~n1246 & n1858 ) | ( ~n1246 & n8802 ) | ( n1858 & n8802 ) ;
  assign n8804 = n4208 | n8803 ;
  assign n8805 = n8804 ^ n3335 ^ 1'b0 ;
  assign n8806 = n431 & n4083 ;
  assign n8807 = n8806 ^ n6092 ^ 1'b0 ;
  assign n8808 = ( n5940 & ~n8805 ) | ( n5940 & n8807 ) | ( ~n8805 & n8807 ) ;
  assign n8809 = n2091 | n8808 ;
  assign n8810 = n2814 ^ n2009 ^ n1601 ;
  assign n8811 = n8509 ^ n6396 ^ n1601 ;
  assign n8812 = ~n3351 & n8811 ;
  assign n8813 = ~n8810 & n8812 ;
  assign n8814 = n8813 ^ n3305 ^ n1985 ;
  assign n8815 = n6115 & n8814 ;
  assign n8816 = n8815 ^ n6694 ^ 1'b0 ;
  assign n8817 = n1984 ^ n1508 ^ n1410 ;
  assign n8818 = ( n698 & ~n907 ) | ( n698 & n1527 ) | ( ~n907 & n1527 ) ;
  assign n8819 = n8818 ^ n2672 ^ n615 ;
  assign n8820 = n8819 ^ n1786 ^ 1'b0 ;
  assign n8821 = n8817 & n8820 ;
  assign n8822 = n889 & ~n4601 ;
  assign n8823 = n8821 | n8822 ;
  assign n8824 = n4680 ^ n3542 ^ 1'b0 ;
  assign n8825 = n3514 & n8824 ;
  assign n8826 = ( n1878 & n3611 ) | ( n1878 & n6580 ) | ( n3611 & n6580 ) ;
  assign n8827 = ~n700 & n3418 ;
  assign n8829 = n952 & ~n1331 ;
  assign n8830 = ~n1672 & n8829 ;
  assign n8828 = ( n1314 & ~n3330 ) | ( n1314 & n6541 ) | ( ~n3330 & n6541 ) ;
  assign n8831 = n8830 ^ n8828 ^ 1'b0 ;
  assign n8832 = ~n8827 & n8831 ;
  assign n8833 = ~n3196 & n5289 ;
  assign n8836 = n7637 ^ x219 ^ 1'b0 ;
  assign n8834 = n3759 ^ n3353 ^ 1'b0 ;
  assign n8835 = n637 & n8834 ;
  assign n8837 = n8836 ^ n8835 ^ 1'b0 ;
  assign n8838 = x171 & ~n8837 ;
  assign n8839 = n7208 ^ n4104 ^ 1'b0 ;
  assign n8840 = n8839 ^ n7087 ^ 1'b0 ;
  assign n8841 = n8840 ^ n5846 ^ n5763 ;
  assign n8842 = n8468 ^ n7413 ^ n7115 ;
  assign n8843 = n3878 ^ n3855 ^ n626 ;
  assign n8844 = n8843 ^ n4776 ^ n476 ;
  assign n8845 = ( n1007 & n3735 ) | ( n1007 & n5484 ) | ( n3735 & n5484 ) ;
  assign n8846 = n7494 ^ n4208 ^ 1'b0 ;
  assign n8847 = ~n8845 & n8846 ;
  assign n8848 = ~x19 & n4986 ;
  assign n8849 = ( n7013 & n7708 ) | ( n7013 & n8848 ) | ( n7708 & n8848 ) ;
  assign n8850 = n7698 ^ n6379 ^ n4499 ;
  assign n8851 = ( n580 & ~n4553 ) | ( n580 & n5610 ) | ( ~n4553 & n5610 ) ;
  assign n8852 = n1159 | n8851 ;
  assign n8853 = n8852 ^ n6295 ^ 1'b0 ;
  assign n8854 = x173 & n1034 ;
  assign n8855 = n3089 & ~n3905 ;
  assign n8856 = n8854 & n8855 ;
  assign n8857 = n6401 ^ n3823 ^ 1'b0 ;
  assign n8858 = n8857 ^ n4352 ^ n2036 ;
  assign n8859 = ~x72 & n938 ;
  assign n8860 = ~n357 & n8859 ;
  assign n8861 = ( n1912 & n2258 ) | ( n1912 & n8860 ) | ( n2258 & n8860 ) ;
  assign n8862 = ( x58 & ~n4904 ) | ( x58 & n8861 ) | ( ~n4904 & n8861 ) ;
  assign n8863 = n8011 ^ n5493 ^ 1'b0 ;
  assign n8864 = n2723 & n8863 ;
  assign n8865 = n1465 & ~n8864 ;
  assign n8866 = n6782 | n8111 ;
  assign n8867 = n595 & n605 ;
  assign n8868 = n8867 ^ n1092 ^ 1'b0 ;
  assign n8869 = n8868 ^ n5418 ^ n883 ;
  assign n8870 = n5155 ^ n5036 ^ n1943 ;
  assign n8871 = n1838 & n4147 ;
  assign n8872 = n8871 ^ n3100 ^ 1'b0 ;
  assign n8873 = ( n5383 & ~n5915 ) | ( n5383 & n8872 ) | ( ~n5915 & n8872 ) ;
  assign n8874 = ~n6921 & n8873 ;
  assign n8875 = n8874 ^ n3984 ^ 1'b0 ;
  assign n8876 = ~n7627 & n7782 ;
  assign n8877 = n8876 ^ n3833 ^ 1'b0 ;
  assign n8878 = ( n2097 & n3444 ) | ( n2097 & n5420 ) | ( n3444 & n5420 ) ;
  assign n8879 = ~n1981 & n2908 ;
  assign n8880 = ~n4864 & n8879 ;
  assign n8881 = ( n1438 & n8878 ) | ( n1438 & n8880 ) | ( n8878 & n8880 ) ;
  assign n8883 = n3868 ^ n1101 ^ n327 ;
  assign n8882 = n693 ^ x94 ^ 1'b0 ;
  assign n8884 = n8883 ^ n8882 ^ n4358 ;
  assign n8885 = ( n3374 & ~n3772 ) | ( n3374 & n5357 ) | ( ~n3772 & n5357 ) ;
  assign n8886 = n8885 ^ n499 ^ x150 ;
  assign n8887 = n4375 ^ n2867 ^ x248 ;
  assign n8888 = ( n654 & n1118 ) | ( n654 & ~n2280 ) | ( n1118 & ~n2280 ) ;
  assign n8889 = n8888 ^ x159 ^ 1'b0 ;
  assign n8890 = n8889 ^ n2287 ^ n1726 ;
  assign n8891 = n4316 ^ n1211 ^ 1'b0 ;
  assign n8892 = ~n8890 & n8891 ;
  assign n8893 = n2576 ^ n2402 ^ 1'b0 ;
  assign n8894 = ( ~x74 & n6706 ) | ( ~x74 & n8893 ) | ( n6706 & n8893 ) ;
  assign n8895 = ( n4723 & ~n6910 ) | ( n4723 & n8894 ) | ( ~n6910 & n8894 ) ;
  assign n8896 = n7818 ^ n1344 ^ n1018 ;
  assign n8897 = n3543 & n8896 ;
  assign n8898 = n8897 ^ n6064 ^ 1'b0 ;
  assign n8899 = x77 & n1408 ;
  assign n8900 = n7163 ^ n1320 ^ 1'b0 ;
  assign n8901 = ~n1428 & n8900 ;
  assign n8902 = n8901 ^ n3903 ^ x121 ;
  assign n8903 = ( n6148 & n6192 ) | ( n6148 & n8902 ) | ( n6192 & n8902 ) ;
  assign n8904 = ~n2403 & n8903 ;
  assign n8905 = ( n3378 & n6819 ) | ( n3378 & n8904 ) | ( n6819 & n8904 ) ;
  assign n8906 = ~n2936 & n8905 ;
  assign n8911 = n6190 ^ n4867 ^ n2394 ;
  assign n8908 = n3431 ^ n2750 ^ 1'b0 ;
  assign n8909 = n4113 ^ n2987 ^ 1'b0 ;
  assign n8910 = n8908 & ~n8909 ;
  assign n8912 = n8911 ^ n8910 ^ 1'b0 ;
  assign n8913 = ~n700 & n8912 ;
  assign n8914 = n7170 & n8913 ;
  assign n8915 = n1744 & n8914 ;
  assign n8907 = ( x11 & n611 ) | ( x11 & ~n2626 ) | ( n611 & ~n2626 ) ;
  assign n8916 = n8915 ^ n8907 ^ 1'b0 ;
  assign n8917 = ( ~n1106 & n1556 ) | ( ~n1106 & n2364 ) | ( n1556 & n2364 ) ;
  assign n8918 = n1122 ^ x126 ^ x122 ;
  assign n8919 = n1701 | n8918 ;
  assign n8920 = n8919 ^ n2620 ^ 1'b0 ;
  assign n8921 = ~n8917 & n8920 ;
  assign n8922 = ( n5803 & n7596 ) | ( n5803 & ~n8921 ) | ( n7596 & ~n8921 ) ;
  assign n8923 = n7711 ^ n7181 ^ n4758 ;
  assign n8924 = n8148 ^ n2386 ^ 1'b0 ;
  assign n8934 = n3557 ^ x231 ^ 1'b0 ;
  assign n8935 = n5191 | n8934 ;
  assign n8925 = n6721 ^ n5061 ^ 1'b0 ;
  assign n8926 = ~n3745 & n8925 ;
  assign n8927 = ~n961 & n8926 ;
  assign n8928 = n2158 & n7019 ;
  assign n8929 = n8928 ^ n2769 ^ 1'b0 ;
  assign n8930 = n8929 ^ n5612 ^ n2365 ;
  assign n8931 = n8930 ^ n4877 ^ 1'b0 ;
  assign n8932 = ~n7448 & n8931 ;
  assign n8933 = n8927 & n8932 ;
  assign n8936 = n8935 ^ n8933 ^ n7675 ;
  assign n8937 = n2260 & ~n2820 ;
  assign n8941 = n3168 ^ n3076 ^ 1'b0 ;
  assign n8938 = n2279 | n4206 ;
  assign n8939 = n3692 | n8938 ;
  assign n8940 = n8939 ^ n5480 ^ n3996 ;
  assign n8942 = n8941 ^ n8940 ^ 1'b0 ;
  assign n8943 = n8937 & n8942 ;
  assign n8949 = n4363 ^ n2365 ^ n1464 ;
  assign n8948 = n899 | n4255 ;
  assign n8950 = n8949 ^ n8948 ^ 1'b0 ;
  assign n8944 = ~n3673 & n8734 ;
  assign n8945 = n4876 & n8944 ;
  assign n8946 = n1821 ^ n1362 ^ n423 ;
  assign n8947 = n8945 & n8946 ;
  assign n8951 = n8950 ^ n8947 ^ n2746 ;
  assign n8952 = ( n1859 & ~n4533 ) | ( n1859 & n7688 ) | ( ~n4533 & n7688 ) ;
  assign n8953 = n8952 ^ n3133 ^ 1'b0 ;
  assign n8954 = n7836 ^ n5978 ^ 1'b0 ;
  assign n8955 = n5706 | n8954 ;
  assign n8956 = ( x71 & n8953 ) | ( x71 & n8955 ) | ( n8953 & n8955 ) ;
  assign n8961 = ~n1790 & n2905 ;
  assign n8962 = n8961 ^ n1051 ^ 1'b0 ;
  assign n8963 = n4104 ^ n821 ^ 1'b0 ;
  assign n8964 = n3455 | n8963 ;
  assign n8965 = n8964 ^ n4570 ^ n1988 ;
  assign n8966 = n3953 | n8965 ;
  assign n8967 = n3623 & ~n8966 ;
  assign n8968 = n5712 | n8967 ;
  assign n8969 = n8962 | n8968 ;
  assign n8957 = n8433 ^ n289 ^ 1'b0 ;
  assign n8958 = ~n2215 & n8957 ;
  assign n8959 = n8470 ^ n2790 ^ 1'b0 ;
  assign n8960 = ( n2647 & n8958 ) | ( n2647 & n8959 ) | ( n8958 & n8959 ) ;
  assign n8970 = n8969 ^ n8960 ^ n1218 ;
  assign n8971 = n6746 ^ n6503 ^ 1'b0 ;
  assign n8973 = ( n1244 & n1548 ) | ( n1244 & n2258 ) | ( n1548 & n2258 ) ;
  assign n8974 = n8973 ^ n2284 ^ 1'b0 ;
  assign n8975 = n8974 ^ n8929 ^ n294 ;
  assign n8972 = n7708 ^ n3528 ^ n2620 ;
  assign n8976 = n8975 ^ n8972 ^ n4368 ;
  assign n8977 = ( n2858 & n5364 ) | ( n2858 & ~n6754 ) | ( n5364 & ~n6754 ) ;
  assign n8978 = n6204 ^ n1884 ^ 1'b0 ;
  assign n8979 = n8978 ^ n7636 ^ 1'b0 ;
  assign n8980 = n8977 & ~n8979 ;
  assign n8981 = ( ~n2227 & n6267 ) | ( ~n2227 & n8980 ) | ( n6267 & n8980 ) ;
  assign n8982 = n2391 ^ n1635 ^ 1'b0 ;
  assign n8983 = n8982 ^ n8199 ^ n1964 ;
  assign n8984 = n2722 ^ n894 ^ 1'b0 ;
  assign n8985 = ( n1127 & ~n1150 ) | ( n1127 & n2822 ) | ( ~n1150 & n2822 ) ;
  assign n8986 = ( ~x111 & n8941 ) | ( ~x111 & n8985 ) | ( n8941 & n8985 ) ;
  assign n8987 = n8790 & ~n8986 ;
  assign n8988 = n2985 & n8987 ;
  assign n8989 = n3546 ^ n391 ^ 1'b0 ;
  assign n8990 = n2280 | n8989 ;
  assign n8994 = n5664 ^ n3101 ^ n1857 ;
  assign n8993 = ~x82 & n3110 ;
  assign n8995 = n8994 ^ n8993 ^ 1'b0 ;
  assign n8991 = ~n1442 & n2189 ;
  assign n8992 = n8991 ^ n2889 ^ 1'b0 ;
  assign n8996 = n8995 ^ n8992 ^ n5337 ;
  assign n8997 = ~n419 & n8996 ;
  assign n8998 = ~n5378 & n8997 ;
  assign n8999 = n8990 & n8998 ;
  assign n9000 = n1882 | n8999 ;
  assign n9001 = n9000 ^ n4137 ^ 1'b0 ;
  assign n9002 = n633 ^ n496 ^ 1'b0 ;
  assign n9003 = n5793 ^ n2629 ^ 1'b0 ;
  assign n9004 = n2145 & ~n9003 ;
  assign n9005 = ~n654 & n796 ;
  assign n9006 = n9005 ^ n3788 ^ 1'b0 ;
  assign n9007 = n9006 ^ n1776 ^ 1'b0 ;
  assign n9008 = n2865 & n9007 ;
  assign n9009 = n7613 ^ n5987 ^ n1845 ;
  assign n9010 = ( x224 & x238 ) | ( x224 & n1075 ) | ( x238 & n1075 ) ;
  assign n9011 = n9010 ^ n5726 ^ 1'b0 ;
  assign n9012 = n9009 & n9011 ;
  assign n9013 = n1986 & ~n6683 ;
  assign n9014 = n5855 | n9013 ;
  assign n9018 = n1192 ^ x66 ^ 1'b0 ;
  assign n9015 = ( n1721 & ~n2440 ) | ( n1721 & n3664 ) | ( ~n2440 & n3664 ) ;
  assign n9016 = n9015 ^ n1886 ^ 1'b0 ;
  assign n9017 = ~n3629 & n9016 ;
  assign n9019 = n9018 ^ n9017 ^ 1'b0 ;
  assign n9020 = ( n6694 & ~n7102 ) | ( n6694 & n9019 ) | ( ~n7102 & n9019 ) ;
  assign n9023 = ( n1428 & n2380 ) | ( n1428 & n4427 ) | ( n2380 & n4427 ) ;
  assign n9024 = ( n3264 & n8279 ) | ( n3264 & n9023 ) | ( n8279 & n9023 ) ;
  assign n9021 = n8396 ^ n7055 ^ n3315 ;
  assign n9022 = ~n4271 & n9021 ;
  assign n9025 = n9024 ^ n9022 ^ 1'b0 ;
  assign n9026 = n9025 ^ x78 ^ 1'b0 ;
  assign n9027 = ~n7740 & n9026 ;
  assign n9028 = n9027 ^ n3503 ^ 1'b0 ;
  assign n9029 = n4672 ^ n2993 ^ 1'b0 ;
  assign n9030 = ~n3985 & n9029 ;
  assign n9031 = n5703 ^ x74 ^ 1'b0 ;
  assign n9032 = n9030 & ~n9031 ;
  assign n9033 = ( n2638 & n7406 ) | ( n2638 & n7788 ) | ( n7406 & n7788 ) ;
  assign n9034 = n9033 ^ n8655 ^ 1'b0 ;
  assign n9035 = n5921 ^ n632 ^ 1'b0 ;
  assign n9036 = n7394 ^ n1576 ^ 1'b0 ;
  assign n9037 = n4343 | n9036 ;
  assign n9038 = n9037 ^ n5054 ^ 1'b0 ;
  assign n9039 = n9038 ^ n3429 ^ 1'b0 ;
  assign n9045 = n1261 ^ x65 ^ 1'b0 ;
  assign n9046 = n1149 | n9045 ;
  assign n9047 = ( x198 & ~n4253 ) | ( x198 & n9046 ) | ( ~n4253 & n9046 ) ;
  assign n9040 = ( n887 & n2705 ) | ( n887 & n6632 ) | ( n2705 & n6632 ) ;
  assign n9041 = n9040 ^ n6529 ^ n358 ;
  assign n9042 = ( n2374 & n6109 ) | ( n2374 & ~n7413 ) | ( n6109 & ~n7413 ) ;
  assign n9043 = n4588 | n9042 ;
  assign n9044 = n9041 & n9043 ;
  assign n9048 = n9047 ^ n9044 ^ n1913 ;
  assign n9049 = ( n3200 & n3310 ) | ( n3200 & n6061 ) | ( n3310 & n6061 ) ;
  assign n9050 = n9049 ^ n3906 ^ n3491 ;
  assign n9051 = n4596 | n9050 ;
  assign n9052 = n3569 | n9051 ;
  assign n9053 = n9052 ^ n6215 ^ 1'b0 ;
  assign n9054 = n6725 ^ n1400 ^ 1'b0 ;
  assign n9055 = x8 & n5715 ;
  assign n9056 = n7165 & n9055 ;
  assign n9057 = n9056 ^ n8964 ^ n8352 ;
  assign n9058 = n7494 ^ n6673 ^ n521 ;
  assign n9059 = n8913 | n9058 ;
  assign n9060 = ~n820 & n1745 ;
  assign n9061 = n9060 ^ n2833 ^ n1083 ;
  assign n9062 = n6358 & n6526 ;
  assign n9063 = n9062 ^ n7522 ^ 1'b0 ;
  assign n9064 = n3231 & ~n5763 ;
  assign n9065 = n9064 ^ n3765 ^ n1969 ;
  assign n9066 = ( n555 & ~n1994 ) | ( n555 & n2408 ) | ( ~n1994 & n2408 ) ;
  assign n9067 = ( n2367 & n3428 ) | ( n2367 & ~n6379 ) | ( n3428 & ~n6379 ) ;
  assign n9068 = n9067 ^ n2498 ^ 1'b0 ;
  assign n9069 = n9066 | n9068 ;
  assign n9070 = ( n3999 & n4321 ) | ( n3999 & n9069 ) | ( n4321 & n9069 ) ;
  assign n9071 = n7236 ^ n3951 ^ 1'b0 ;
  assign n9072 = ( n3802 & ~n5589 ) | ( n3802 & n6077 ) | ( ~n5589 & n6077 ) ;
  assign n9073 = ( n755 & n836 ) | ( n755 & n5658 ) | ( n836 & n5658 ) ;
  assign n9074 = n5584 ^ n3569 ^ 1'b0 ;
  assign n9075 = ~n9073 & n9074 ;
  assign n9076 = ( n7725 & n9072 ) | ( n7725 & ~n9075 ) | ( n9072 & ~n9075 ) ;
  assign n9077 = n7655 ^ n1789 ^ 1'b0 ;
  assign n9078 = n4482 & n5020 ;
  assign n9079 = ~n4957 & n9078 ;
  assign n9080 = n4603 ^ n3546 ^ n2669 ;
  assign n9081 = ( n554 & n1947 ) | ( n554 & n9080 ) | ( n1947 & n9080 ) ;
  assign n9082 = ~n1437 & n5263 ;
  assign n9083 = n2368 ^ n1977 ^ n1356 ;
  assign n9084 = n9083 ^ n4748 ^ n3932 ;
  assign n9085 = n2261 & n4644 ;
  assign n9086 = n9084 & n9085 ;
  assign n9087 = ~n591 & n3832 ;
  assign n9088 = ( ~n9082 & n9086 ) | ( ~n9082 & n9087 ) | ( n9086 & n9087 ) ;
  assign n9089 = n2220 | n2913 ;
  assign n9090 = n6555 | n9089 ;
  assign n9091 = n9090 ^ n6784 ^ 1'b0 ;
  assign n9092 = n8939 ^ n3532 ^ 1'b0 ;
  assign n9093 = ~n1004 & n9092 ;
  assign n9094 = n9093 ^ n9033 ^ n7140 ;
  assign n9095 = ( n5046 & n5741 ) | ( n5046 & ~n9094 ) | ( n5741 & ~n9094 ) ;
  assign n9096 = ( n1552 & ~n1736 ) | ( n1552 & n7771 ) | ( ~n1736 & n7771 ) ;
  assign n9097 = ~n749 & n5679 ;
  assign n9098 = n3592 ^ n936 ^ 1'b0 ;
  assign n9099 = n2405 | n9098 ;
  assign n9100 = n9099 ^ n8487 ^ 1'b0 ;
  assign n9101 = n3278 | n3318 ;
  assign n9102 = ( ~n5677 & n6136 ) | ( ~n5677 & n9101 ) | ( n6136 & n9101 ) ;
  assign n9103 = n9100 & n9102 ;
  assign n9104 = x34 & ~n6523 ;
  assign n9105 = ~n9103 & n9104 ;
  assign n9106 = n886 & ~n3191 ;
  assign n9107 = ~n5359 & n7741 ;
  assign n9108 = ( n272 & ~n2279 ) | ( n272 & n9107 ) | ( ~n2279 & n9107 ) ;
  assign n9109 = n9108 ^ n7719 ^ 1'b0 ;
  assign n9110 = n9109 ^ n6306 ^ n3041 ;
  assign n9111 = n8860 ^ n5357 ^ n2027 ;
  assign n9112 = n9111 ^ n3761 ^ n900 ;
  assign n9113 = n5913 & ~n9112 ;
  assign n9114 = n9113 ^ n6270 ^ n1916 ;
  assign n9120 = ( n4626 & n4759 ) | ( n4626 & ~n4929 ) | ( n4759 & ~n4929 ) ;
  assign n9115 = n431 & ~n3933 ;
  assign n9116 = ~n2786 & n9115 ;
  assign n9117 = n6587 & ~n9116 ;
  assign n9118 = n9117 ^ x66 ^ 1'b0 ;
  assign n9119 = n9118 ^ n3556 ^ 1'b0 ;
  assign n9121 = n9120 ^ n9119 ^ 1'b0 ;
  assign n9122 = n973 & n9121 ;
  assign n9123 = n8509 ^ n6665 ^ 1'b0 ;
  assign n9124 = n1813 & n9123 ;
  assign n9125 = ~n2050 & n4801 ;
  assign n9126 = ( n9010 & n9124 ) | ( n9010 & n9125 ) | ( n9124 & n9125 ) ;
  assign n9129 = n7191 ^ n1338 ^ n1247 ;
  assign n9127 = ( n289 & n1504 ) | ( n289 & n2934 ) | ( n1504 & n2934 ) ;
  assign n9128 = x208 & ~n9127 ;
  assign n9130 = n9129 ^ n9128 ^ 1'b0 ;
  assign n9131 = n9130 ^ n7668 ^ n3738 ;
  assign n9132 = n9126 | n9131 ;
  assign n9133 = n389 & ~n2461 ;
  assign n9134 = n9133 ^ n1162 ^ 1'b0 ;
  assign n9135 = ~n461 & n3004 ;
  assign n9136 = ~n9134 & n9135 ;
  assign n9137 = n7210 & n9136 ;
  assign n9138 = n9137 ^ n6497 ^ 1'b0 ;
  assign n9139 = n6077 | n9138 ;
  assign n9140 = n9139 ^ n757 ^ 1'b0 ;
  assign n9141 = x26 & n9140 ;
  assign n9142 = n9132 | n9141 ;
  assign n9143 = n6470 & ~n8877 ;
  assign n9144 = n5520 ^ n5195 ^ 1'b0 ;
  assign n9145 = ~n4321 & n9144 ;
  assign n9146 = ~x82 & n9145 ;
  assign n9147 = ( n1691 & n4941 ) | ( n1691 & ~n5074 ) | ( n4941 & ~n5074 ) ;
  assign n9150 = n1458 & ~n5207 ;
  assign n9151 = n5135 & n9150 ;
  assign n9148 = n3410 ^ n2341 ^ 1'b0 ;
  assign n9149 = n1264 & n9148 ;
  assign n9152 = n9151 ^ n9149 ^ 1'b0 ;
  assign n9153 = ~n812 & n9152 ;
  assign n9154 = ( n2135 & ~n5435 ) | ( n2135 & n9153 ) | ( ~n5435 & n9153 ) ;
  assign n9155 = n1938 & ~n2389 ;
  assign n9156 = ~n3239 & n3951 ;
  assign n9157 = n5958 | n9156 ;
  assign n9158 = n9157 ^ n8827 ^ 1'b0 ;
  assign n9159 = n3862 ^ n561 ^ 1'b0 ;
  assign n9160 = n3418 ^ n587 ^ 1'b0 ;
  assign n9161 = ( ~n5954 & n9159 ) | ( ~n5954 & n9160 ) | ( n9159 & n9160 ) ;
  assign n9162 = n9161 ^ n7143 ^ 1'b0 ;
  assign n9163 = n7689 ^ n3245 ^ n1276 ;
  assign n9164 = x103 & n849 ;
  assign n9165 = n602 ^ n362 ^ 1'b0 ;
  assign n9166 = n9165 ^ n4750 ^ n2343 ;
  assign n9167 = n910 & n9166 ;
  assign n9168 = ~n5689 & n9167 ;
  assign n9169 = n4435 & ~n9168 ;
  assign n9170 = n7842 ^ n4873 ^ 1'b0 ;
  assign n9171 = x108 & n551 ;
  assign n9172 = n9171 ^ n8754 ^ 1'b0 ;
  assign n9173 = n6649 ^ n886 ^ 1'b0 ;
  assign n9174 = n3307 | n9173 ;
  assign n9175 = n9174 ^ n9156 ^ 1'b0 ;
  assign n9176 = n9172 | n9175 ;
  assign n9177 = n9176 ^ n642 ^ 1'b0 ;
  assign n9178 = ( n4051 & n9170 ) | ( n4051 & ~n9177 ) | ( n9170 & ~n9177 ) ;
  assign n9179 = n2077 & ~n2904 ;
  assign n9180 = n9179 ^ n2687 ^ 1'b0 ;
  assign n9181 = n9180 ^ n2611 ^ 1'b0 ;
  assign n9182 = ~n3154 & n9181 ;
  assign n9183 = n6196 & n9182 ;
  assign n9184 = n2771 & n9183 ;
  assign n9185 = n2230 & ~n2367 ;
  assign n9186 = n9185 ^ n1573 ^ 1'b0 ;
  assign n9187 = n9186 ^ n593 ^ 1'b0 ;
  assign n9188 = n2443 & ~n9187 ;
  assign n9189 = x201 & ~n4961 ;
  assign n9190 = n5205 ^ n360 ^ 1'b0 ;
  assign n9191 = x127 & ~n4585 ;
  assign n9192 = n9191 ^ n326 ^ 1'b0 ;
  assign n9193 = ~n9190 & n9192 ;
  assign n9194 = n6930 ^ n2785 ^ 1'b0 ;
  assign n9195 = x63 & n9194 ;
  assign n9196 = ( n9189 & ~n9193 ) | ( n9189 & n9195 ) | ( ~n9193 & n9195 ) ;
  assign n9197 = ( n807 & n916 ) | ( n807 & ~n1031 ) | ( n916 & ~n1031 ) ;
  assign n9198 = x141 & ~n9197 ;
  assign n9199 = n2730 & n9198 ;
  assign n9200 = n9199 ^ n2187 ^ n1591 ;
  assign n9201 = ( n1739 & n8608 ) | ( n1739 & n9200 ) | ( n8608 & n9200 ) ;
  assign n9207 = n4486 & ~n4866 ;
  assign n9208 = n9207 ^ n2872 ^ 1'b0 ;
  assign n9209 = n4799 & n9208 ;
  assign n9202 = ~n1726 & n2861 ;
  assign n9203 = n9202 ^ n3341 ^ 1'b0 ;
  assign n9204 = n9203 ^ n5575 ^ 1'b0 ;
  assign n9205 = ~n5767 & n9204 ;
  assign n9206 = n4182 & n9205 ;
  assign n9210 = n9209 ^ n9206 ^ 1'b0 ;
  assign n9211 = ( n660 & n4765 ) | ( n660 & n9052 ) | ( n4765 & n9052 ) ;
  assign n9212 = x110 & n4571 ;
  assign n9213 = ~n9211 & n9212 ;
  assign n9219 = n2107 ^ n1145 ^ n404 ;
  assign n9220 = n9219 ^ n5666 ^ 1'b0 ;
  assign n9215 = n552 & n3260 ;
  assign n9216 = ~n1749 & n9215 ;
  assign n9214 = ~n5231 & n7505 ;
  assign n9217 = n9216 ^ n9214 ^ 1'b0 ;
  assign n9218 = ( n616 & n2580 ) | ( n616 & ~n9217 ) | ( n2580 & ~n9217 ) ;
  assign n9221 = n9220 ^ n9218 ^ 1'b0 ;
  assign n9222 = n9213 | n9221 ;
  assign n9223 = ( n1299 & ~n3184 ) | ( n1299 & n6311 ) | ( ~n3184 & n6311 ) ;
  assign n9224 = n1214 & n9223 ;
  assign n9225 = n9224 ^ n4748 ^ 1'b0 ;
  assign n9226 = ( n2905 & n3072 ) | ( n2905 & n9225 ) | ( n3072 & n9225 ) ;
  assign n9227 = n5807 ^ n3960 ^ 1'b0 ;
  assign n9228 = n8995 ^ n1963 ^ n1592 ;
  assign n9229 = ( n9226 & ~n9227 ) | ( n9226 & n9228 ) | ( ~n9227 & n9228 ) ;
  assign n9230 = ( n5965 & n9149 ) | ( n5965 & n9229 ) | ( n9149 & n9229 ) ;
  assign n9231 = n7732 ^ n4064 ^ 1'b0 ;
  assign n9232 = x59 & n9231 ;
  assign n9233 = n9232 ^ n435 ^ 1'b0 ;
  assign n9234 = n5048 & n9233 ;
  assign n9235 = ~n3754 & n4924 ;
  assign n9236 = n789 & n9235 ;
  assign n9237 = n654 & n4550 ;
  assign n9238 = n9237 ^ n7274 ^ n7169 ;
  assign n9239 = ( n9234 & n9236 ) | ( n9234 & ~n9238 ) | ( n9236 & ~n9238 ) ;
  assign n9246 = ( ~n1415 & n4010 ) | ( ~n1415 & n6132 ) | ( n4010 & n6132 ) ;
  assign n9240 = n4879 ^ n1667 ^ 1'b0 ;
  assign n9241 = n4106 ^ n1043 ^ 1'b0 ;
  assign n9242 = n9240 & ~n9241 ;
  assign n9243 = n2208 | n2444 ;
  assign n9244 = n9243 ^ x178 ^ 1'b0 ;
  assign n9245 = n9242 & n9244 ;
  assign n9247 = n9246 ^ n9245 ^ 1'b0 ;
  assign n9248 = n9247 ^ n4872 ^ 1'b0 ;
  assign n9249 = ( n2444 & ~n2978 ) | ( n2444 & n5858 ) | ( ~n2978 & n5858 ) ;
  assign n9250 = ~n1674 & n6206 ;
  assign n9251 = ( n855 & n2317 ) | ( n855 & n9250 ) | ( n2317 & n9250 ) ;
  assign n9252 = n4544 ^ n867 ^ 1'b0 ;
  assign n9253 = n9252 ^ n2792 ^ 1'b0 ;
  assign n9254 = n2456 & ~n9253 ;
  assign n9255 = ( n3239 & n3424 ) | ( n3239 & ~n5363 ) | ( n3424 & ~n5363 ) ;
  assign n9256 = n9255 ^ n2119 ^ 1'b0 ;
  assign n9257 = n9256 ^ n8545 ^ n8453 ;
  assign n9258 = ( n5766 & n8502 ) | ( n5766 & n8644 ) | ( n8502 & n8644 ) ;
  assign n9259 = n9258 ^ n8986 ^ 1'b0 ;
  assign n9260 = n9259 ^ n7223 ^ n405 ;
  assign n9261 = n944 & ~n1239 ;
  assign n9262 = n9261 ^ n2189 ^ 1'b0 ;
  assign n9263 = n4629 & ~n6750 ;
  assign n9264 = n3330 & n9263 ;
  assign n9265 = ~n1042 & n1953 ;
  assign n9266 = n4238 ^ n1922 ^ 1'b0 ;
  assign n9267 = n9266 ^ n3508 ^ 1'b0 ;
  assign n9268 = ~n7464 & n9267 ;
  assign n9269 = n9265 & n9268 ;
  assign n9270 = ( n4933 & ~n9264 ) | ( n4933 & n9269 ) | ( ~n9264 & n9269 ) ;
  assign n9271 = n2145 & n2519 ;
  assign n9272 = n3288 | n6682 ;
  assign n9273 = n9271 | n9272 ;
  assign n9274 = n8828 | n9273 ;
  assign n9275 = n9274 ^ n8043 ^ n6560 ;
  assign n9276 = ( n1409 & n6683 ) | ( n1409 & ~n9275 ) | ( n6683 & ~n9275 ) ;
  assign n9277 = n8304 | n9276 ;
  assign n9278 = n9277 ^ n7634 ^ 1'b0 ;
  assign n9284 = n3366 | n7076 ;
  assign n9285 = n9284 ^ n5592 ^ 1'b0 ;
  assign n9282 = n8681 ^ n6213 ^ 1'b0 ;
  assign n9283 = ~n2780 & n9282 ;
  assign n9286 = n9285 ^ n9283 ^ 1'b0 ;
  assign n9287 = n9286 ^ n2933 ^ n2904 ;
  assign n9281 = x158 & ~n6290 ;
  assign n9288 = n9287 ^ n9281 ^ 1'b0 ;
  assign n9280 = n2688 | n4854 ;
  assign n9279 = ( n2585 & ~n4823 ) | ( n2585 & n5602 ) | ( ~n4823 & n5602 ) ;
  assign n9289 = n9288 ^ n9280 ^ n9279 ;
  assign n9290 = n6917 | n9289 ;
  assign n9291 = ( ~n4546 & n8802 ) | ( ~n4546 & n8913 ) | ( n8802 & n8913 ) ;
  assign n9292 = n1030 ^ n466 ^ 1'b0 ;
  assign n9299 = ( n2405 & ~n2478 ) | ( n2405 & n7626 ) | ( ~n2478 & n7626 ) ;
  assign n9300 = n9299 ^ n8103 ^ n6184 ;
  assign n9296 = n485 | n5813 ;
  assign n9297 = n3184 & ~n9296 ;
  assign n9293 = x156 & n3292 ;
  assign n9294 = n9293 ^ n4449 ^ n3856 ;
  assign n9295 = n9294 ^ n1986 ^ 1'b0 ;
  assign n9298 = n9297 ^ n9295 ^ 1'b0 ;
  assign n9301 = n9300 ^ n9298 ^ 1'b0 ;
  assign n9302 = n2757 | n3360 ;
  assign n9304 = ~n2009 & n3795 ;
  assign n9303 = x48 & ~n7461 ;
  assign n9305 = n9304 ^ n9303 ^ 1'b0 ;
  assign n9306 = ( ~n8392 & n9302 ) | ( ~n8392 & n9305 ) | ( n9302 & n9305 ) ;
  assign n9309 = n8200 ^ n650 ^ 1'b0 ;
  assign n9310 = n524 & n9309 ;
  assign n9311 = ~n3377 & n9310 ;
  assign n9308 = x123 & ~n468 ;
  assign n9312 = n9311 ^ n9308 ^ 1'b0 ;
  assign n9307 = n2201 & ~n8632 ;
  assign n9313 = n9312 ^ n9307 ^ 1'b0 ;
  assign n9314 = ( n6130 & ~n9306 ) | ( n6130 & n9313 ) | ( ~n9306 & n9313 ) ;
  assign n9315 = n3501 ^ n2050 ^ n2040 ;
  assign n9316 = ~n4905 & n9315 ;
  assign n9317 = ( ~n1187 & n2718 ) | ( ~n1187 & n9196 ) | ( n2718 & n9196 ) ;
  assign n9318 = n885 & ~n1652 ;
  assign n9319 = n9318 ^ n3824 ^ 1'b0 ;
  assign n9320 = ( n1867 & n4656 ) | ( n1867 & ~n9319 ) | ( n4656 & ~n9319 ) ;
  assign n9321 = n9320 ^ n5071 ^ n259 ;
  assign n9322 = ~n3278 & n9321 ;
  assign n9323 = n5336 ^ n750 ^ x88 ;
  assign n9324 = n1816 & n2574 ;
  assign n9325 = n9324 ^ n4369 ^ 1'b0 ;
  assign n9326 = ~n6501 & n9150 ;
  assign n9327 = n9326 ^ n8717 ^ 1'b0 ;
  assign n9330 = n946 & ~n7821 ;
  assign n9331 = ( ~n4932 & n8455 ) | ( ~n4932 & n9330 ) | ( n8455 & n9330 ) ;
  assign n9328 = n2629 ^ x10 ^ 1'b0 ;
  assign n9329 = n7373 & ~n9328 ;
  assign n9332 = n9331 ^ n9329 ^ 1'b0 ;
  assign n9333 = n7382 ^ n3325 ^ 1'b0 ;
  assign n9334 = n6919 & n9333 ;
  assign n9335 = x216 & ~n5089 ;
  assign n9336 = n4267 & n9335 ;
  assign n9337 = ( n3066 & ~n5565 ) | ( n3066 & n7698 ) | ( ~n5565 & n7698 ) ;
  assign n9338 = n6365 & ~n9337 ;
  assign n9339 = n9336 & n9338 ;
  assign n9340 = ( ~n2286 & n4873 ) | ( ~n2286 & n7939 ) | ( n4873 & n7939 ) ;
  assign n9341 = n6094 & ~n9340 ;
  assign n9342 = n1938 | n5842 ;
  assign n9346 = n2795 ^ x142 ^ 1'b0 ;
  assign n9347 = n1473 | n9346 ;
  assign n9348 = n9347 ^ n4119 ^ 1'b0 ;
  assign n9343 = n2258 ^ x116 ^ 1'b0 ;
  assign n9344 = x198 | n9343 ;
  assign n9345 = ~n3390 & n9344 ;
  assign n9349 = n9348 ^ n9345 ^ 1'b0 ;
  assign n9350 = n5940 & ~n9349 ;
  assign n9351 = n4337 ^ n2519 ^ n915 ;
  assign n9352 = n9351 ^ n4180 ^ x150 ;
  assign n9353 = n2757 | n6531 ;
  assign n9354 = n9352 & ~n9353 ;
  assign n9355 = n2802 | n3479 ;
  assign n9356 = n9354 & ~n9355 ;
  assign n9361 = n2786 ^ n502 ^ 1'b0 ;
  assign n9360 = n4494 ^ n2149 ^ 1'b0 ;
  assign n9357 = n3220 ^ n2972 ^ n2554 ;
  assign n9358 = ( n4182 & n6727 ) | ( n4182 & ~n9357 ) | ( n6727 & ~n9357 ) ;
  assign n9359 = ( n3113 & n7009 ) | ( n3113 & n9358 ) | ( n7009 & n9358 ) ;
  assign n9362 = n9361 ^ n9360 ^ n9359 ;
  assign n9365 = ( ~n940 & n1852 ) | ( ~n940 & n4908 ) | ( n1852 & n4908 ) ;
  assign n9363 = n2735 ^ n2559 ^ 1'b0 ;
  assign n9364 = ( ~n3401 & n3721 ) | ( ~n3401 & n9363 ) | ( n3721 & n9363 ) ;
  assign n9366 = n9365 ^ n9364 ^ 1'b0 ;
  assign n9367 = n9366 ^ n2994 ^ 1'b0 ;
  assign n9368 = ~n4513 & n9367 ;
  assign n9369 = n399 & n946 ;
  assign n9370 = n5741 | n9369 ;
  assign n9371 = n7797 ^ n1896 ^ 1'b0 ;
  assign n9372 = n320 & ~n9371 ;
  assign n9373 = n9372 ^ n3759 ^ 1'b0 ;
  assign n9374 = n9373 ^ n3898 ^ 1'b0 ;
  assign n9375 = n9374 ^ n7990 ^ 1'b0 ;
  assign n9376 = n6860 | n9375 ;
  assign n9377 = ~n4165 & n4970 ;
  assign n9378 = ( n2313 & n8430 ) | ( n2313 & n9377 ) | ( n8430 & n9377 ) ;
  assign n9379 = ( n1502 & n4409 ) | ( n1502 & ~n9378 ) | ( n4409 & ~n9378 ) ;
  assign n9380 = n9379 ^ n8777 ^ n536 ;
  assign n9381 = n700 | n3388 ;
  assign n9382 = n5929 & n8385 ;
  assign n9383 = ~n9381 & n9382 ;
  assign n9384 = n5840 ^ n4419 ^ 1'b0 ;
  assign n9385 = n9384 ^ n3650 ^ 1'b0 ;
  assign n9386 = ( n6745 & n7401 ) | ( n6745 & ~n7797 ) | ( n7401 & ~n7797 ) ;
  assign n9387 = ~n1372 & n6296 ;
  assign n9388 = n4006 ^ x98 ^ 1'b0 ;
  assign n9389 = n4893 | n9388 ;
  assign n9390 = n9309 & ~n9389 ;
  assign n9391 = n343 & ~n9390 ;
  assign n9392 = n9387 & n9391 ;
  assign n9393 = n9392 ^ n2904 ^ 1'b0 ;
  assign n9395 = n2175 & n3994 ;
  assign n9396 = n468 & n9395 ;
  assign n9394 = n6960 ^ n3109 ^ 1'b0 ;
  assign n9397 = n9396 ^ n9394 ^ n7182 ;
  assign n9398 = ~n5680 & n6402 ;
  assign n9399 = ~n1317 & n7820 ;
  assign n9400 = n7701 & n9399 ;
  assign n9401 = n8660 & n9400 ;
  assign n9402 = n9401 ^ n7285 ^ n3104 ;
  assign n9403 = ( n1243 & n1674 ) | ( n1243 & ~n1779 ) | ( n1674 & ~n1779 ) ;
  assign n9404 = n9403 ^ n4410 ^ 1'b0 ;
  assign n9405 = ~n2794 & n9404 ;
  assign n9406 = n9405 ^ n4575 ^ n2791 ;
  assign n9407 = n3917 & ~n4057 ;
  assign n9408 = n420 & n9407 ;
  assign n9409 = n4788 | n9408 ;
  assign n9410 = n915 | n9409 ;
  assign n9411 = n5316 | n9410 ;
  assign n9412 = n9406 & ~n9411 ;
  assign n9413 = n741 & ~n4517 ;
  assign n9414 = n4072 & ~n9413 ;
  assign n9415 = n1873 ^ x4 ^ 1'b0 ;
  assign n9416 = n1061 & ~n9415 ;
  assign n9417 = n9416 ^ n1576 ^ 1'b0 ;
  assign n9418 = ( n5126 & ~n6796 ) | ( n5126 & n9417 ) | ( ~n6796 & n9417 ) ;
  assign n9419 = ( n2972 & n9414 ) | ( n2972 & n9418 ) | ( n9414 & n9418 ) ;
  assign n9420 = n4856 ^ n1485 ^ n785 ;
  assign n9421 = n9420 ^ n4562 ^ 1'b0 ;
  assign n9422 = n9421 ^ n3689 ^ 1'b0 ;
  assign n9423 = ( x190 & n1181 ) | ( x190 & ~n1885 ) | ( n1181 & ~n1885 ) ;
  assign n9424 = n5451 & ~n9423 ;
  assign n9425 = n617 & ~n5902 ;
  assign n9426 = n9425 ^ n1644 ^ 1'b0 ;
  assign n9427 = n3973 & n9426 ;
  assign n9429 = n2230 ^ n1655 ^ 1'b0 ;
  assign n9428 = n864 & n7514 ;
  assign n9430 = n9429 ^ n9428 ^ 1'b0 ;
  assign n9431 = n4694 & n5138 ;
  assign n9432 = ( n8513 & ~n9430 ) | ( n8513 & n9431 ) | ( ~n9430 & n9431 ) ;
  assign n9433 = n396 | n652 ;
  assign n9434 = x66 & ~n9433 ;
  assign n9435 = n5374 & n9244 ;
  assign n9436 = n476 & n9435 ;
  assign n9437 = n2700 ^ n2519 ^ 1'b0 ;
  assign n9438 = ~n3341 & n9437 ;
  assign n9439 = x162 & n3962 ;
  assign n9440 = n9439 ^ n7552 ^ 1'b0 ;
  assign n9441 = n5968 ^ n4773 ^ 1'b0 ;
  assign n9442 = n9440 & n9441 ;
  assign n9443 = ~n5118 & n9442 ;
  assign n9444 = ~n9438 & n9443 ;
  assign n9445 = n431 ^ x238 ^ 1'b0 ;
  assign n9446 = x122 & ~n9445 ;
  assign n9447 = n4080 ^ n1610 ^ 1'b0 ;
  assign n9448 = ( ~x103 & n9446 ) | ( ~x103 & n9447 ) | ( n9446 & n9447 ) ;
  assign n9449 = n642 & ~n4838 ;
  assign n9450 = ( n1199 & ~n1420 ) | ( n1199 & n7160 ) | ( ~n1420 & n7160 ) ;
  assign n9456 = n3727 ^ n731 ^ 1'b0 ;
  assign n9451 = n3957 ^ n2529 ^ n485 ;
  assign n9452 = n435 & n9451 ;
  assign n9453 = n4851 & n4919 ;
  assign n9454 = n9452 & n9453 ;
  assign n9455 = n9454 ^ n8659 ^ n7075 ;
  assign n9457 = n9456 ^ n9455 ^ n1003 ;
  assign n9458 = n7185 ^ n455 ^ 1'b0 ;
  assign n9459 = n9403 ^ n1075 ^ 1'b0 ;
  assign n9460 = n8940 | n9459 ;
  assign n9461 = n8536 ^ n7463 ^ n1258 ;
  assign n9462 = ~n1991 & n2068 ;
  assign n9463 = n9462 ^ n1175 ^ 1'b0 ;
  assign n9464 = n3568 & ~n9463 ;
  assign n9465 = n9464 ^ n2663 ^ 1'b0 ;
  assign n9466 = ( ~n1776 & n2321 ) | ( ~n1776 & n9465 ) | ( n2321 & n9465 ) ;
  assign n9467 = ( n8190 & n8906 ) | ( n8190 & ~n9466 ) | ( n8906 & ~n9466 ) ;
  assign n9468 = ( ~n386 & n452 ) | ( ~n386 & n7195 ) | ( n452 & n7195 ) ;
  assign n9469 = n3633 & n6812 ;
  assign n9470 = ( n5489 & n5872 ) | ( n5489 & ~n9469 ) | ( n5872 & ~n9469 ) ;
  assign n9471 = ~n2846 & n5785 ;
  assign n9472 = ~n9470 & n9471 ;
  assign n9473 = n3334 & ~n6945 ;
  assign n9475 = ( n534 & n6323 ) | ( n534 & n7920 ) | ( n6323 & n7920 ) ;
  assign n9474 = ( n512 & ~n1109 ) | ( n512 & n4873 ) | ( ~n1109 & n4873 ) ;
  assign n9476 = n9475 ^ n9474 ^ n5634 ;
  assign n9477 = ( n4961 & ~n5003 ) | ( n4961 & n5313 ) | ( ~n5003 & n5313 ) ;
  assign n9478 = n9477 ^ n8734 ^ n1223 ;
  assign n9479 = n9478 ^ n2475 ^ n2205 ;
  assign n9480 = ( ~n4689 & n8153 ) | ( ~n4689 & n9479 ) | ( n8153 & n9479 ) ;
  assign n9481 = n962 ^ x48 ^ 1'b0 ;
  assign n9482 = x70 & ~n3118 ;
  assign n9483 = n3456 | n7911 ;
  assign n9484 = n9442 | n9483 ;
  assign n9486 = n2840 & ~n4274 ;
  assign n9487 = n3932 | n9486 ;
  assign n9488 = n2104 | n9487 ;
  assign n9485 = ~n3643 & n3750 ;
  assign n9489 = n9488 ^ n9485 ^ n6582 ;
  assign n9490 = n8122 & n9489 ;
  assign n9491 = ~n9484 & n9490 ;
  assign n9492 = ( n3509 & ~n4137 ) | ( n3509 & n9491 ) | ( ~n4137 & n9491 ) ;
  assign n9493 = n9482 & n9492 ;
  assign n9494 = n9493 ^ n5979 ^ 1'b0 ;
  assign n9495 = n1236 & ~n4382 ;
  assign n9496 = n9495 ^ n5364 ^ 1'b0 ;
  assign n9497 = ~n1875 & n7278 ;
  assign n9498 = n9242 ^ n6205 ^ n558 ;
  assign n9499 = n5032 ^ n5011 ^ n682 ;
  assign n9500 = ( n1046 & n8631 ) | ( n1046 & n9499 ) | ( n8631 & n9499 ) ;
  assign n9501 = n8658 ^ n459 ^ 1'b0 ;
  assign n9509 = x216 & n8604 ;
  assign n9510 = ~n1050 & n9509 ;
  assign n9503 = ( x48 & n3507 ) | ( x48 & n5132 ) | ( n3507 & n5132 ) ;
  assign n9504 = ~n6267 & n9503 ;
  assign n9505 = n9504 ^ n6415 ^ n2965 ;
  assign n9502 = ~n5620 & n7084 ;
  assign n9506 = n9505 ^ n9502 ^ 1'b0 ;
  assign n9507 = n4770 & ~n9506 ;
  assign n9508 = n9507 ^ n798 ^ 1'b0 ;
  assign n9511 = n9510 ^ n9508 ^ 1'b0 ;
  assign n9512 = n2699 & n9511 ;
  assign n9513 = n5532 ^ n1939 ^ 1'b0 ;
  assign n9514 = n9513 ^ n6859 ^ n5371 ;
  assign n9515 = n495 | n9514 ;
  assign n9516 = n6283 | n9515 ;
  assign n9517 = n5439 ^ n2230 ^ n2045 ;
  assign n9518 = n9517 ^ n6646 ^ 1'b0 ;
  assign n9519 = n9518 ^ n9405 ^ n6598 ;
  assign n9520 = n9519 ^ n6582 ^ 1'b0 ;
  assign n9521 = x243 & n3168 ;
  assign n9522 = ( n3894 & n6679 ) | ( n3894 & n9521 ) | ( n6679 & n9521 ) ;
  assign n9523 = n5014 ^ n3345 ^ 1'b0 ;
  assign n9524 = n6862 & ~n9523 ;
  assign n9525 = n2705 & n9524 ;
  assign n9526 = n4333 & n9525 ;
  assign n9527 = n6730 ^ n4083 ^ 1'b0 ;
  assign n9528 = n3303 | n8880 ;
  assign n9529 = n9527 & ~n9528 ;
  assign n9530 = ( ~n983 & n2687 ) | ( ~n983 & n9182 ) | ( n2687 & n9182 ) ;
  assign n9531 = ( n5407 & ~n7511 ) | ( n5407 & n9530 ) | ( ~n7511 & n9530 ) ;
  assign n9532 = n3323 ^ n1761 ^ 1'b0 ;
  assign n9533 = n9531 | n9532 ;
  assign n9534 = n9533 ^ n1208 ^ 1'b0 ;
  assign n9535 = n2032 & n3358 ;
  assign n9536 = n9535 ^ n8808 ^ n5551 ;
  assign n9542 = n8094 ^ n7802 ^ n3292 ;
  assign n9543 = n9542 ^ n2189 ^ 1'b0 ;
  assign n9538 = n7790 & n9119 ;
  assign n9539 = n9538 ^ n7070 ^ 1'b0 ;
  assign n9540 = n9539 ^ n9337 ^ n3757 ;
  assign n9537 = ~n3309 & n4808 ;
  assign n9541 = n9540 ^ n9537 ^ 1'b0 ;
  assign n9544 = n9543 ^ n9541 ^ n2286 ;
  assign n9545 = ~n1472 & n7599 ;
  assign n9546 = ( x173 & n4793 ) | ( x173 & n6822 ) | ( n4793 & n6822 ) ;
  assign n9547 = n9546 ^ n5347 ^ n2853 ;
  assign n9548 = n9547 ^ n9447 ^ 1'b0 ;
  assign n9549 = n6971 | n9548 ;
  assign n9550 = n2876 ^ n868 ^ 1'b0 ;
  assign n9551 = ~n6671 & n9550 ;
  assign n9552 = n9551 ^ x103 ^ 1'b0 ;
  assign n9553 = n7487 ^ n5352 ^ 1'b0 ;
  assign n9554 = n3526 | n4006 ;
  assign n9555 = n9554 ^ n6174 ^ n4611 ;
  assign n9556 = ( ~n3805 & n8731 ) | ( ~n3805 & n9555 ) | ( n8731 & n9555 ) ;
  assign n9557 = ( n9552 & ~n9553 ) | ( n9552 & n9556 ) | ( ~n9553 & n9556 ) ;
  assign n9558 = n5337 & n6395 ;
  assign n9559 = ~n1043 & n9558 ;
  assign n9560 = n1066 | n2267 ;
  assign n9561 = n9559 & ~n9560 ;
  assign n9562 = n9561 ^ n1353 ^ n1307 ;
  assign n9563 = n3917 & ~n9562 ;
  assign n9564 = ~n1287 & n7626 ;
  assign n9565 = n3805 ^ n3762 ^ 1'b0 ;
  assign n9566 = ~n9564 & n9565 ;
  assign n9567 = n9566 ^ x65 ^ 1'b0 ;
  assign n9568 = n481 & ~n1003 ;
  assign n9569 = n6330 | n9568 ;
  assign n9570 = n1158 ^ x213 ^ 1'b0 ;
  assign n9571 = n5750 | n9570 ;
  assign n9572 = x166 | n9571 ;
  assign n9573 = ~n9569 & n9572 ;
  assign n9574 = ~n9567 & n9573 ;
  assign n9575 = ( n8070 & ~n9563 ) | ( n8070 & n9574 ) | ( ~n9563 & n9574 ) ;
  assign n9576 = ~n5059 & n5111 ;
  assign n9577 = n3797 & ~n9576 ;
  assign n9578 = n3918 & n9577 ;
  assign n9588 = n9517 ^ n8097 ^ n1480 ;
  assign n9589 = ( n580 & ~n3748 ) | ( n580 & n5080 ) | ( ~n3748 & n5080 ) ;
  assign n9590 = ( n1385 & n4259 ) | ( n1385 & ~n9589 ) | ( n4259 & ~n9589 ) ;
  assign n9591 = ( n8675 & n9588 ) | ( n8675 & ~n9590 ) | ( n9588 & ~n9590 ) ;
  assign n9580 = ( n3536 & n4639 ) | ( n3536 & n4968 ) | ( n4639 & n4968 ) ;
  assign n9581 = n9580 ^ n3551 ^ n827 ;
  assign n9582 = n9581 ^ n1622 ^ 1'b0 ;
  assign n9583 = ~n1883 & n9582 ;
  assign n9584 = n3918 | n5342 ;
  assign n9585 = n9583 | n9584 ;
  assign n9579 = ( n2665 & n5285 ) | ( n2665 & ~n7588 ) | ( n5285 & ~n7588 ) ;
  assign n9586 = n9585 ^ n9579 ^ 1'b0 ;
  assign n9587 = n9586 ^ n5367 ^ n2745 ;
  assign n9592 = n9591 ^ n9587 ^ n5448 ;
  assign n9594 = ( x196 & ~n2710 ) | ( x196 & n3578 ) | ( ~n2710 & n3578 ) ;
  assign n9593 = n2333 & ~n6733 ;
  assign n9595 = n9594 ^ n9593 ^ n7795 ;
  assign n9596 = ~n7795 & n8737 ;
  assign n9597 = ( ~n1454 & n7172 ) | ( ~n1454 & n7208 ) | ( n7172 & n7208 ) ;
  assign n9598 = n3387 | n7145 ;
  assign n9599 = n8094 ^ n6470 ^ n5509 ;
  assign n9600 = ( n3305 & ~n9340 ) | ( n3305 & n9599 ) | ( ~n9340 & n9599 ) ;
  assign n9602 = n358 & n3511 ;
  assign n9603 = n9602 ^ n2252 ^ 1'b0 ;
  assign n9604 = n1543 & n9603 ;
  assign n9605 = n9604 ^ x128 ^ 1'b0 ;
  assign n9606 = n9605 ^ n4306 ^ 1'b0 ;
  assign n9601 = ( n1674 & n4051 ) | ( n1674 & n9524 ) | ( n4051 & n9524 ) ;
  assign n9607 = n9606 ^ n9601 ^ n2825 ;
  assign n9608 = n4064 ^ n1974 ^ 1'b0 ;
  assign n9609 = n1379 | n9608 ;
  assign n9610 = n9609 ^ n1192 ^ 1'b0 ;
  assign n9611 = n9610 ^ n3468 ^ n2524 ;
  assign n9612 = ~n4781 & n6323 ;
  assign n9613 = n2273 ^ x5 ^ 1'b0 ;
  assign n9614 = n4308 & ~n9613 ;
  assign n9615 = n9614 ^ n3311 ^ 1'b0 ;
  assign n9616 = ~n1883 & n4116 ;
  assign n9617 = ~n5528 & n7135 ;
  assign n9618 = ~n4081 & n9617 ;
  assign n9619 = n3465 & ~n5982 ;
  assign n9620 = ( n3319 & n9618 ) | ( n3319 & n9619 ) | ( n9618 & n9619 ) ;
  assign n9621 = ~n3286 & n6115 ;
  assign n9622 = ( x53 & ~n1529 ) | ( x53 & n5372 ) | ( ~n1529 & n5372 ) ;
  assign n9623 = ( n1278 & n6686 ) | ( n1278 & ~n7321 ) | ( n6686 & ~n7321 ) ;
  assign n9624 = ( n6483 & ~n6486 ) | ( n6483 & n9623 ) | ( ~n6486 & n9623 ) ;
  assign n9625 = x207 & ~n1331 ;
  assign n9626 = n9625 ^ n1876 ^ n903 ;
  assign n9627 = n5128 ^ n2793 ^ 1'b0 ;
  assign n9628 = n8097 | n9627 ;
  assign n9629 = n9628 ^ n5480 ^ 1'b0 ;
  assign n9630 = n7086 | n9629 ;
  assign n9631 = n9626 & ~n9630 ;
  assign n9632 = ( n1621 & ~n5030 ) | ( n1621 & n9108 ) | ( ~n5030 & n9108 ) ;
  assign n9633 = ( ~n1676 & n1935 ) | ( ~n1676 & n9632 ) | ( n1935 & n9632 ) ;
  assign n9634 = n3383 ^ n1810 ^ n429 ;
  assign n9635 = n8666 ^ n5667 ^ n5331 ;
  assign n9636 = n1973 & n8033 ;
  assign n9637 = ( n3046 & ~n9635 ) | ( n3046 & n9636 ) | ( ~n9635 & n9636 ) ;
  assign n9639 = n2774 & ~n4152 ;
  assign n9640 = n2607 & n9639 ;
  assign n9638 = n2369 & n4029 ;
  assign n9641 = n9640 ^ n9638 ^ 1'b0 ;
  assign n9642 = n3745 & n9641 ;
  assign n9643 = ~n1741 & n9642 ;
  assign n9644 = n6996 ^ n4147 ^ x247 ;
  assign n9645 = ~n2221 & n9644 ;
  assign n9646 = n9645 ^ n853 ^ 1'b0 ;
  assign n9647 = n2791 | n5452 ;
  assign n9648 = n2905 ^ x239 ^ 1'b0 ;
  assign n9649 = n9648 ^ n2731 ^ 1'b0 ;
  assign n9650 = n816 & ~n9649 ;
  assign n9651 = n6682 ^ n4993 ^ 1'b0 ;
  assign n9652 = n6269 & n9651 ;
  assign n9653 = n4518 ^ n4038 ^ n1385 ;
  assign n9654 = n4481 | n9653 ;
  assign n9657 = n1176 | n2880 ;
  assign n9658 = x179 | n9657 ;
  assign n9655 = n1134 ^ n1081 ^ n671 ;
  assign n9656 = n8551 & n9655 ;
  assign n9659 = n9658 ^ n9656 ^ 1'b0 ;
  assign n9660 = n9659 ^ n2730 ^ n2677 ;
  assign n9661 = n5961 ^ n3775 ^ n3721 ;
  assign n9662 = ~n9660 & n9661 ;
  assign n9663 = ( n5601 & n9654 ) | ( n5601 & n9662 ) | ( n9654 & n9662 ) ;
  assign n9664 = ( ~n763 & n4363 ) | ( ~n763 & n5656 ) | ( n4363 & n5656 ) ;
  assign n9665 = n7083 ^ n5797 ^ 1'b0 ;
  assign n9669 = ~n5473 & n5679 ;
  assign n9670 = n5034 & n9669 ;
  assign n9666 = n1592 ^ n1446 ^ 1'b0 ;
  assign n9667 = n9363 ^ n4452 ^ 1'b0 ;
  assign n9668 = ~n9666 & n9667 ;
  assign n9671 = n9670 ^ n9668 ^ 1'b0 ;
  assign n9672 = x31 & ~n9671 ;
  assign n9673 = n9672 ^ n3234 ^ 1'b0 ;
  assign n9674 = ~n7055 & n9673 ;
  assign n9675 = n3576 ^ n1881 ^ n1874 ;
  assign n9676 = n9675 ^ n560 ^ 1'b0 ;
  assign n9677 = n4036 | n9676 ;
  assign n9678 = ( n3627 & n5958 ) | ( n3627 & n8660 ) | ( n5958 & n8660 ) ;
  assign n9679 = n8372 ^ n414 ^ 1'b0 ;
  assign n9680 = n6580 | n9679 ;
  assign n9681 = n9535 ^ n6367 ^ 1'b0 ;
  assign n9682 = ~n2909 & n3846 ;
  assign n9683 = n9682 ^ n7098 ^ 1'b0 ;
  assign n9684 = n366 & ~n483 ;
  assign n9685 = n9684 ^ x138 ^ 1'b0 ;
  assign n9686 = n1191 & ~n9685 ;
  assign n9687 = n9686 ^ n1780 ^ 1'b0 ;
  assign n9688 = n9687 ^ n4738 ^ n4479 ;
  assign n9689 = ~n1868 & n7084 ;
  assign n9690 = n9689 ^ n8809 ^ 1'b0 ;
  assign n9691 = n9690 ^ n3459 ^ 1'b0 ;
  assign n9692 = ~n3650 & n8697 ;
  assign n9693 = n9692 ^ x108 ^ 1'b0 ;
  assign n9694 = ~n2502 & n5126 ;
  assign n9695 = ( ~n4438 & n7955 ) | ( ~n4438 & n9694 ) | ( n7955 & n9694 ) ;
  assign n9696 = ~n1097 & n9695 ;
  assign n9697 = n9693 & n9696 ;
  assign n9698 = n5494 ^ n2114 ^ 1'b0 ;
  assign n9699 = n533 & n9698 ;
  assign n9700 = n1533 ^ n1390 ^ 1'b0 ;
  assign n9701 = n9700 ^ n4842 ^ n827 ;
  assign n9702 = ( ~n3260 & n7943 ) | ( ~n3260 & n9701 ) | ( n7943 & n9701 ) ;
  assign n9703 = n3206 & n9702 ;
  assign n9710 = n6629 ^ n2928 ^ n575 ;
  assign n9704 = n3752 ^ n1802 ^ 1'b0 ;
  assign n9705 = ~n759 & n9704 ;
  assign n9706 = n4199 ^ n3402 ^ n2657 ;
  assign n9707 = n9705 & ~n9706 ;
  assign n9708 = n9707 ^ n7752 ^ 1'b0 ;
  assign n9709 = n9182 & n9708 ;
  assign n9711 = n9710 ^ n9709 ^ 1'b0 ;
  assign n9712 = ~n3456 & n5238 ;
  assign n9713 = ~n1325 & n4970 ;
  assign n9714 = n9713 ^ x4 ^ 1'b0 ;
  assign n9720 = x231 & n6640 ;
  assign n9721 = n3548 & n9720 ;
  assign n9719 = x15 & n3902 ;
  assign n9722 = n9721 ^ n9719 ^ 1'b0 ;
  assign n9723 = n9722 ^ n5765 ^ n396 ;
  assign n9715 = n2868 ^ n1836 ^ n841 ;
  assign n9716 = n4350 & n9150 ;
  assign n9717 = n9715 & n9716 ;
  assign n9718 = n9717 ^ n5242 ^ n2492 ;
  assign n9724 = n9723 ^ n9718 ^ n3276 ;
  assign n9725 = ( x94 & ~n2388 ) | ( x94 & n2687 ) | ( ~n2388 & n2687 ) ;
  assign n9726 = n9725 ^ n9594 ^ n1117 ;
  assign n9727 = n9726 ^ n8472 ^ n3858 ;
  assign n9729 = n634 & ~n2856 ;
  assign n9730 = ( n1996 & ~n4555 ) | ( n1996 & n9729 ) | ( ~n4555 & n9729 ) ;
  assign n9731 = n2936 | n7774 ;
  assign n9732 = n9730 | n9731 ;
  assign n9728 = n7846 | n9024 ;
  assign n9733 = n9732 ^ n9728 ^ 1'b0 ;
  assign n9734 = n1814 ^ n424 ^ 1'b0 ;
  assign n9735 = n6475 & n9734 ;
  assign n9736 = n9735 ^ n2744 ^ 1'b0 ;
  assign n9737 = ~n5316 & n9736 ;
  assign n9738 = ( n1031 & ~n7096 ) | ( n1031 & n9737 ) | ( ~n7096 & n9737 ) ;
  assign n9739 = ~n1340 & n4168 ;
  assign n9740 = n9738 & n9739 ;
  assign n9741 = x69 & x74 ;
  assign n9742 = n2610 & n9741 ;
  assign n9743 = n9742 ^ n5214 ^ n1484 ;
  assign n9745 = ( x208 & n1936 ) | ( x208 & ~n3125 ) | ( n1936 & ~n3125 ) ;
  assign n9744 = n2276 & ~n3478 ;
  assign n9746 = n9745 ^ n9744 ^ 1'b0 ;
  assign n9747 = n9746 ^ n6395 ^ 1'b0 ;
  assign n9748 = n3107 ^ n895 ^ 1'b0 ;
  assign n9749 = n9747 & ~n9748 ;
  assign n9750 = n4272 & n9749 ;
  assign n9751 = ~n9743 & n9750 ;
  assign n9752 = ( x34 & n3114 ) | ( x34 & n3305 ) | ( n3114 & n3305 ) ;
  assign n9753 = ~n774 & n9752 ;
  assign n9754 = n9753 ^ n4957 ^ 1'b0 ;
  assign n9755 = n9754 ^ n7622 ^ n2573 ;
  assign n9756 = ~x101 & n9755 ;
  assign n9757 = ~n3237 & n5138 ;
  assign n9758 = n5470 | n6192 ;
  assign n9759 = ( n5151 & n9757 ) | ( n5151 & ~n9758 ) | ( n9757 & ~n9758 ) ;
  assign n9760 = n8346 ^ n4682 ^ n4588 ;
  assign n9761 = n9760 ^ n4546 ^ 1'b0 ;
  assign n9769 = ( n381 & n1863 ) | ( n381 & ~n8935 ) | ( n1863 & ~n8935 ) ;
  assign n9762 = n3250 ^ n528 ^ 1'b0 ;
  assign n9763 = n3024 & n9762 ;
  assign n9764 = n9763 ^ n491 ^ 1'b0 ;
  assign n9765 = n2930 & ~n9764 ;
  assign n9766 = n9765 ^ n6138 ^ n2934 ;
  assign n9767 = ~n1268 & n9766 ;
  assign n9768 = ~n3953 & n9767 ;
  assign n9770 = n9769 ^ n9768 ^ 1'b0 ;
  assign n9771 = n2442 ^ n1806 ^ 1'b0 ;
  assign n9772 = n5188 & n9771 ;
  assign n9774 = n3478 ^ n2353 ^ 1'b0 ;
  assign n9775 = n1864 | n9774 ;
  assign n9773 = n2075 | n9576 ;
  assign n9776 = n9775 ^ n9773 ^ 1'b0 ;
  assign n9777 = ( n2470 & ~n9772 ) | ( n2470 & n9776 ) | ( ~n9772 & n9776 ) ;
  assign n9778 = ( n483 & n2059 ) | ( n483 & ~n5929 ) | ( n2059 & ~n5929 ) ;
  assign n9779 = ( n7264 & n8707 ) | ( n7264 & ~n9778 ) | ( n8707 & ~n9778 ) ;
  assign n9781 = n4306 ^ n3061 ^ n2957 ;
  assign n9782 = n4738 | n9781 ;
  assign n9780 = n2679 & ~n3790 ;
  assign n9783 = n9782 ^ n9780 ^ 1'b0 ;
  assign n9784 = ~n9779 & n9783 ;
  assign n9785 = ~n7464 & n7841 ;
  assign n9786 = n9785 ^ n7215 ^ 1'b0 ;
  assign n9789 = ( n306 & ~n881 ) | ( n306 & n3705 ) | ( ~n881 & n3705 ) ;
  assign n9787 = ~n3290 & n4100 ;
  assign n9788 = n1243 | n9787 ;
  assign n9790 = n9789 ^ n9788 ^ n9001 ;
  assign n9791 = ~n4045 & n9625 ;
  assign n9792 = n1477 & n9791 ;
  assign n9793 = n8941 | n9792 ;
  assign n9794 = ~x157 & n3647 ;
  assign n9795 = n9794 ^ n6878 ^ 1'b0 ;
  assign n9796 = n3366 ^ n3138 ^ 1'b0 ;
  assign n9797 = n9795 | n9796 ;
  assign n9803 = n1473 | n8203 ;
  assign n9801 = ~n5321 & n8212 ;
  assign n9798 = n6607 ^ n4854 ^ n847 ;
  assign n9799 = n9798 ^ n1576 ^ 1'b0 ;
  assign n9800 = n1405 & n9799 ;
  assign n9802 = n9801 ^ n9800 ^ 1'b0 ;
  assign n9804 = n9803 ^ n9802 ^ 1'b0 ;
  assign n9805 = ( n2293 & n7040 ) | ( n2293 & n8951 ) | ( n7040 & n8951 ) ;
  assign n9806 = n1801 & ~n4310 ;
  assign n9807 = n3632 & n9806 ;
  assign n9808 = ~n3325 & n4239 ;
  assign n9809 = n9808 ^ n3165 ^ 1'b0 ;
  assign n9810 = ( n2340 & ~n9807 ) | ( n2340 & n9809 ) | ( ~n9807 & n9809 ) ;
  assign n9811 = n1192 ^ n711 ^ 1'b0 ;
  assign n9812 = n8620 & ~n9811 ;
  assign n9813 = n9812 ^ n3545 ^ 1'b0 ;
  assign n9814 = n657 & n9813 ;
  assign n9815 = ~n795 & n7544 ;
  assign n9816 = n4935 & n9815 ;
  assign n9817 = n6320 & ~n8296 ;
  assign n9818 = n6022 ^ n2934 ^ n1804 ;
  assign n9819 = n1783 & ~n1961 ;
  assign n9820 = n9818 & n9819 ;
  assign n9821 = n9820 ^ n7766 ^ n2569 ;
  assign n9822 = n8512 ^ n7067 ^ 1'b0 ;
  assign n9823 = n1661 & n9822 ;
  assign n9824 = n4629 ^ n1838 ^ 1'b0 ;
  assign n9825 = ( n434 & n4854 ) | ( n434 & ~n6671 ) | ( n4854 & ~n6671 ) ;
  assign n9826 = n2705 & n9825 ;
  assign n9827 = n9826 ^ n1655 ^ 1'b0 ;
  assign n9828 = n9827 ^ n1559 ^ 1'b0 ;
  assign n9829 = ~n4708 & n9828 ;
  assign n9830 = ~n7744 & n9829 ;
  assign n9831 = n9824 & n9830 ;
  assign n9832 = n9831 ^ n6015 ^ 1'b0 ;
  assign n9833 = n7263 & ~n9832 ;
  assign n9834 = n430 | n5907 ;
  assign n9835 = n4793 & ~n9834 ;
  assign n9836 = ~n2417 & n4034 ;
  assign n9837 = n9836 ^ n855 ^ 1'b0 ;
  assign n9838 = n9835 | n9837 ;
  assign n9839 = n9838 ^ n441 ^ 1'b0 ;
  assign n9840 = ( ~n3781 & n5918 ) | ( ~n3781 & n9839 ) | ( n5918 & n9839 ) ;
  assign n9841 = n4173 ^ n2388 ^ n1095 ;
  assign n9842 = n9841 ^ n7306 ^ 1'b0 ;
  assign n9843 = ( x247 & n357 ) | ( x247 & ~n2479 ) | ( n357 & ~n2479 ) ;
  assign n9844 = n9843 ^ n2655 ^ 1'b0 ;
  assign n9845 = n2355 & ~n9844 ;
  assign n9846 = n4038 ^ n2721 ^ x45 ;
  assign n9847 = n9845 & n9846 ;
  assign n9848 = n9842 & n9847 ;
  assign n9849 = n9848 ^ n5299 ^ 1'b0 ;
  assign n9850 = n4175 & n4575 ;
  assign n9851 = n9850 ^ n3543 ^ 1'b0 ;
  assign n9853 = ( n1676 & ~n3225 ) | ( n1676 & n7464 ) | ( ~n3225 & n7464 ) ;
  assign n9854 = n678 & n4435 ;
  assign n9855 = ( n5353 & n7950 ) | ( n5353 & ~n8975 ) | ( n7950 & ~n8975 ) ;
  assign n9856 = ( n9853 & n9854 ) | ( n9853 & n9855 ) | ( n9854 & n9855 ) ;
  assign n9852 = n4335 ^ n3330 ^ n2563 ;
  assign n9857 = n9856 ^ n9852 ^ 1'b0 ;
  assign n9858 = n9851 | n9857 ;
  assign n9859 = ( n2255 & n6426 ) | ( n2255 & ~n9046 ) | ( n6426 & ~n9046 ) ;
  assign n9860 = ~n1652 & n9544 ;
  assign n9861 = n9860 ^ n7211 ^ 1'b0 ;
  assign n9864 = n3256 ^ n2225 ^ 1'b0 ;
  assign n9865 = n8120 & ~n9864 ;
  assign n9862 = n595 & ~n5435 ;
  assign n9863 = n9862 ^ n1254 ^ 1'b0 ;
  assign n9866 = n9865 ^ n9863 ^ n6608 ;
  assign n9867 = n9866 ^ n5583 ^ n2194 ;
  assign n9870 = n7724 ^ n5873 ^ 1'b0 ;
  assign n9868 = n2413 ^ n526 ^ n487 ;
  assign n9869 = n966 & n9868 ;
  assign n9871 = n9870 ^ n9869 ^ 1'b0 ;
  assign n9872 = n6582 ^ n374 ^ 1'b0 ;
  assign n9873 = n9872 ^ n6680 ^ 1'b0 ;
  assign n9874 = n3639 & n9873 ;
  assign n9875 = n2333 ^ n1845 ^ x22 ;
  assign n9876 = ~n820 & n9875 ;
  assign n9877 = ( n2444 & n2456 ) | ( n2444 & ~n9876 ) | ( n2456 & ~n9876 ) ;
  assign n9878 = ( n5323 & n5524 ) | ( n5323 & n9877 ) | ( n5524 & n9877 ) ;
  assign n9879 = n9878 ^ n8517 ^ 1'b0 ;
  assign n9881 = n5500 ^ n5479 ^ 1'b0 ;
  assign n9880 = n633 & ~n7846 ;
  assign n9882 = n9881 ^ n9880 ^ 1'b0 ;
  assign n9886 = n2357 ^ n1771 ^ n1637 ;
  assign n9887 = ( n847 & n4294 ) | ( n847 & ~n9886 ) | ( n4294 & ~n9886 ) ;
  assign n9883 = n631 & n6640 ;
  assign n9884 = n9883 ^ n4190 ^ 1'b0 ;
  assign n9885 = ~n1941 & n9884 ;
  assign n9888 = n9887 ^ n9885 ^ 1'b0 ;
  assign n9889 = n7540 ^ n6763 ^ n1240 ;
  assign n9890 = n1378 ^ n1292 ^ n1239 ;
  assign n9891 = n6753 ^ n1538 ^ 1'b0 ;
  assign n9892 = ~n1475 & n9891 ;
  assign n9893 = n9890 & n9892 ;
  assign n9894 = ~n6878 & n9893 ;
  assign n9895 = n8162 ^ n3716 ^ 1'b0 ;
  assign n9896 = n4868 | n6780 ;
  assign n9897 = ~n1097 & n5169 ;
  assign n9898 = ~n4531 & n5251 ;
  assign n9899 = n9898 ^ n2450 ^ 1'b0 ;
  assign n9903 = n3311 ^ n2616 ^ 1'b0 ;
  assign n9900 = ( ~n774 & n1714 ) | ( ~n774 & n2374 ) | ( n1714 & n2374 ) ;
  assign n9901 = n2850 | n9900 ;
  assign n9902 = ~n295 & n9901 ;
  assign n9904 = n9903 ^ n9902 ^ 1'b0 ;
  assign n9905 = ( n4318 & n6914 ) | ( n4318 & ~n9904 ) | ( n6914 & ~n9904 ) ;
  assign n9906 = n6947 ^ n1491 ^ 1'b0 ;
  assign n9907 = n7771 | n9906 ;
  assign n9908 = n9907 ^ n8318 ^ n5289 ;
  assign n9909 = ( n3049 & ~n9154 ) | ( n3049 & n9908 ) | ( ~n9154 & n9908 ) ;
  assign n9910 = n4738 | n7617 ;
  assign n9911 = n9910 ^ n9267 ^ n4726 ;
  assign n9912 = ~n3740 & n9911 ;
  assign n9913 = n5416 ^ n626 ^ 1'b0 ;
  assign n9914 = ~n9912 & n9913 ;
  assign n9915 = n9484 ^ n8848 ^ 1'b0 ;
  assign n9916 = x183 & ~n343 ;
  assign n9917 = ( n511 & n2782 ) | ( n511 & n6070 ) | ( n2782 & n6070 ) ;
  assign n9918 = n3551 & n9917 ;
  assign n9919 = n7698 | n9918 ;
  assign n9920 = ( n4010 & n4239 ) | ( n4010 & ~n9919 ) | ( n4239 & ~n9919 ) ;
  assign n9921 = n2182 ^ n1312 ^ n257 ;
  assign n9922 = n680 & ~n6943 ;
  assign n9923 = n2985 & ~n9587 ;
  assign n9924 = n9923 ^ n4713 ^ 1'b0 ;
  assign n9925 = n925 | n2735 ;
  assign n9926 = n8159 | n9925 ;
  assign n9927 = n9926 ^ n7814 ^ n716 ;
  assign n9928 = n9927 ^ n3732 ^ 1'b0 ;
  assign n9929 = n4384 & n9928 ;
  assign n9930 = n4439 ^ n3155 ^ 1'b0 ;
  assign n9931 = n9930 ^ n9607 ^ n6364 ;
  assign n9935 = n326 & n3002 ;
  assign n9936 = n9935 ^ n430 ^ 1'b0 ;
  assign n9937 = n9936 ^ n869 ^ 1'b0 ;
  assign n9938 = n5858 & ~n9937 ;
  assign n9932 = n9418 ^ n5537 ^ n3110 ;
  assign n9933 = n9932 ^ n2124 ^ x205 ;
  assign n9934 = ( n2415 & n9749 ) | ( n2415 & ~n9933 ) | ( n9749 & ~n9933 ) ;
  assign n9939 = n9938 ^ n9934 ^ 1'b0 ;
  assign n9940 = n820 | n9939 ;
  assign n9941 = n2548 ^ x227 ^ 1'b0 ;
  assign n9942 = n2619 | n3474 ;
  assign n9943 = n5936 | n9942 ;
  assign n9944 = n4432 ^ n1483 ^ n700 ;
  assign n9945 = ( n1099 & n1568 ) | ( n1099 & ~n1573 ) | ( n1568 & ~n1573 ) ;
  assign n9946 = n1692 & n3151 ;
  assign n9947 = n9946 ^ n1176 ^ 1'b0 ;
  assign n9948 = n6435 ^ n855 ^ 1'b0 ;
  assign n9949 = ~n6005 & n9948 ;
  assign n9950 = n9947 & n9949 ;
  assign n9951 = ~n9945 & n9950 ;
  assign n9952 = n1887 & ~n8211 ;
  assign n9953 = ~n1084 & n9952 ;
  assign n9954 = n2466 ^ n1721 ^ 1'b0 ;
  assign n9955 = n3243 & n9954 ;
  assign n9956 = n9953 & n9955 ;
  assign n9958 = x26 & n5442 ;
  assign n9959 = n937 & n9958 ;
  assign n9957 = n1778 & ~n6884 ;
  assign n9960 = n9959 ^ n9957 ^ 1'b0 ;
  assign n9961 = n2995 | n5950 ;
  assign n9964 = ( ~n485 & n943 ) | ( ~n485 & n3042 ) | ( n943 & n3042 ) ;
  assign n9965 = ( ~n2303 & n3776 ) | ( ~n2303 & n9964 ) | ( n3776 & n9964 ) ;
  assign n9962 = n1773 | n4095 ;
  assign n9963 = n9962 ^ n5016 ^ 1'b0 ;
  assign n9966 = n9965 ^ n9963 ^ x81 ;
  assign n9968 = x96 & ~n1374 ;
  assign n9969 = ~n973 & n9968 ;
  assign n9970 = n9969 ^ n1932 ^ n512 ;
  assign n9967 = n6870 & n8911 ;
  assign n9971 = n9970 ^ n9967 ^ 1'b0 ;
  assign n9972 = ( n2475 & ~n2478 ) | ( n2475 & n6795 ) | ( ~n2478 & n6795 ) ;
  assign n9973 = n9972 ^ n3075 ^ 1'b0 ;
  assign n9974 = ( n1913 & n4083 ) | ( n1913 & ~n4152 ) | ( n4083 & ~n4152 ) ;
  assign n9975 = ( n4695 & ~n9973 ) | ( n4695 & n9974 ) | ( ~n9973 & n9974 ) ;
  assign n9976 = n7396 ^ n4436 ^ n2775 ;
  assign n9977 = n7608 | n9897 ;
  assign n9978 = n9976 & ~n9977 ;
  assign n9979 = n4138 & n7818 ;
  assign n9980 = n1943 & n9979 ;
  assign n9981 = n9980 ^ n7756 ^ 1'b0 ;
  assign n9982 = n841 & n5214 ;
  assign n9983 = n9982 ^ n5604 ^ 1'b0 ;
  assign n9984 = n7239 & n9983 ;
  assign n9985 = n9984 ^ n3867 ^ 1'b0 ;
  assign n9986 = n2391 & n9985 ;
  assign n9994 = ( n1494 & n2960 ) | ( n1494 & n6868 ) | ( n2960 & n6868 ) ;
  assign n9987 = ~n3839 & n7373 ;
  assign n9988 = ~n579 & n5407 ;
  assign n9989 = n9988 ^ n3243 ^ n1556 ;
  assign n9990 = n5008 | n9989 ;
  assign n9991 = n9990 ^ n7808 ^ 1'b0 ;
  assign n9992 = n9991 ^ n773 ^ 1'b0 ;
  assign n9993 = ~n9987 & n9992 ;
  assign n9995 = n9994 ^ n9993 ^ 1'b0 ;
  assign n9996 = n9432 ^ n1046 ^ 1'b0 ;
  assign n9997 = n1643 & ~n6388 ;
  assign n10004 = n5984 ^ n4230 ^ n2052 ;
  assign n10005 = ( x170 & ~n695 ) | ( x170 & n2080 ) | ( ~n695 & n2080 ) ;
  assign n10006 = n10005 ^ n3247 ^ 1'b0 ;
  assign n10007 = n10004 & n10006 ;
  assign n10008 = x36 & n10007 ;
  assign n9998 = x3 & n8688 ;
  assign n9999 = ~n5398 & n9998 ;
  assign n10000 = ( n5207 & n8770 ) | ( n5207 & ~n9999 ) | ( n8770 & ~n9999 ) ;
  assign n10001 = n10000 ^ n791 ^ 1'b0 ;
  assign n10002 = n10001 ^ n8295 ^ x191 ;
  assign n10003 = n10002 ^ n3495 ^ n3397 ;
  assign n10009 = n10008 ^ n10003 ^ 1'b0 ;
  assign n10010 = n7592 ^ n3920 ^ n3752 ;
  assign n10011 = n9944 | n10010 ;
  assign n10012 = n7678 & ~n10011 ;
  assign n10013 = n8488 ^ n5363 ^ n4743 ;
  assign n10014 = n10013 ^ n6755 ^ n5462 ;
  assign n10016 = n1118 | n3362 ;
  assign n10017 = n10016 ^ n325 ^ 1'b0 ;
  assign n10018 = n5233 & n10017 ;
  assign n10015 = n7608 | n7843 ;
  assign n10019 = n10018 ^ n10015 ^ 1'b0 ;
  assign n10020 = n2286 ^ n2094 ^ 1'b0 ;
  assign n10021 = n4504 & ~n6607 ;
  assign n10022 = n10021 ^ n2356 ^ 1'b0 ;
  assign n10023 = ( n5958 & ~n6451 ) | ( n5958 & n8114 ) | ( ~n6451 & n8114 ) ;
  assign n10024 = ( ~n1188 & n1804 ) | ( ~n1188 & n9746 ) | ( n1804 & n9746 ) ;
  assign n10025 = ~n1791 & n2700 ;
  assign n10026 = n10025 ^ n4343 ^ 1'b0 ;
  assign n10027 = n4266 & ~n6476 ;
  assign n10028 = ( ~n329 & n4883 ) | ( ~n329 & n10027 ) | ( n4883 & n10027 ) ;
  assign n10029 = n9772 ^ n1409 ^ 1'b0 ;
  assign n10030 = ( ~n2948 & n10028 ) | ( ~n2948 & n10029 ) | ( n10028 & n10029 ) ;
  assign n10031 = n6551 ^ n5535 ^ n4242 ;
  assign n10032 = n10030 | n10031 ;
  assign n10033 = ( n9406 & n10026 ) | ( n9406 & ~n10032 ) | ( n10026 & ~n10032 ) ;
  assign n10034 = n3184 | n8585 ;
  assign n10035 = n3528 ^ n446 ^ 1'b0 ;
  assign n10036 = ~n6952 & n10035 ;
  assign n10037 = ~n6107 & n7787 ;
  assign n10038 = ( x196 & n7683 ) | ( x196 & ~n10037 ) | ( n7683 & ~n10037 ) ;
  assign n10039 = ( n5089 & n7282 ) | ( n5089 & n10038 ) | ( n7282 & n10038 ) ;
  assign n10040 = n3803 ^ n961 ^ 1'b0 ;
  assign n10041 = n5162 | n10040 ;
  assign n10042 = n1589 | n7121 ;
  assign n10043 = n10042 ^ n7410 ^ 1'b0 ;
  assign n10044 = ( n1412 & n3366 ) | ( n1412 & n10043 ) | ( n3366 & n10043 ) ;
  assign n10045 = ( n2950 & n4463 ) | ( n2950 & n9687 ) | ( n4463 & n9687 ) ;
  assign n10046 = n1152 | n5448 ;
  assign n10047 = n4123 & ~n10046 ;
  assign n10050 = n3162 ^ n2313 ^ 1'b0 ;
  assign n10048 = n1483 ^ n1111 ^ 1'b0 ;
  assign n10049 = ( n660 & ~n1873 ) | ( n660 & n10048 ) | ( ~n1873 & n10048 ) ;
  assign n10051 = n10050 ^ n10049 ^ 1'b0 ;
  assign n10052 = ~n8508 & n10051 ;
  assign n10053 = n7883 | n10052 ;
  assign n10054 = n5662 ^ n2540 ^ 1'b0 ;
  assign n10055 = ~n930 & n4097 ;
  assign n10056 = n10054 & n10055 ;
  assign n10057 = ( ~n865 & n941 ) | ( ~n865 & n10056 ) | ( n941 & n10056 ) ;
  assign n10058 = n7732 ^ n5521 ^ n3873 ;
  assign n10059 = n2985 ^ n1637 ^ 1'b0 ;
  assign n10060 = n431 & ~n10059 ;
  assign n10062 = n9320 ^ n6994 ^ n3844 ;
  assign n10063 = ( n310 & n874 ) | ( n310 & ~n1270 ) | ( n874 & ~n1270 ) ;
  assign n10064 = n10063 ^ n4923 ^ 1'b0 ;
  assign n10065 = n10062 | n10064 ;
  assign n10061 = ~n2255 & n3066 ;
  assign n10066 = n10065 ^ n10061 ^ 1'b0 ;
  assign n10067 = n9177 ^ n3054 ^ 1'b0 ;
  assign n10068 = ~n5740 & n9992 ;
  assign n10069 = n10068 ^ n8843 ^ 1'b0 ;
  assign n10070 = n1873 ^ n315 ^ 1'b0 ;
  assign n10071 = n1571 & ~n10070 ;
  assign n10072 = n3016 ^ n2778 ^ n2119 ;
  assign n10073 = ( ~n926 & n1464 ) | ( ~n926 & n8262 ) | ( n1464 & n8262 ) ;
  assign n10074 = ~n10072 & n10073 ;
  assign n10075 = n10071 & ~n10074 ;
  assign n10076 = ~x34 & n10075 ;
  assign n10078 = n5315 ^ n2943 ^ n556 ;
  assign n10077 = n5871 ^ n5766 ^ x185 ;
  assign n10079 = n10078 ^ n10077 ^ n262 ;
  assign n10080 = n5093 ^ n3125 ^ 1'b0 ;
  assign n10081 = ~n421 & n3711 ;
  assign n10082 = n10081 ^ n2815 ^ 1'b0 ;
  assign n10083 = ~n8400 & n10082 ;
  assign n10084 = ~n550 & n1287 ;
  assign n10085 = ~x149 & n10084 ;
  assign n10086 = ( n1537 & n1591 ) | ( n1537 & n10085 ) | ( n1591 & n10085 ) ;
  assign n10087 = n10086 ^ n4597 ^ 1'b0 ;
  assign n10088 = ~n748 & n7821 ;
  assign n10089 = n8294 ^ n4445 ^ 1'b0 ;
  assign n10090 = n8023 ^ n3299 ^ n1031 ;
  assign n10091 = n6247 ^ n3371 ^ n1051 ;
  assign n10092 = n5402 ^ n1511 ^ 1'b0 ;
  assign n10093 = n6155 | n10092 ;
  assign n10094 = n6949 ^ n4080 ^ 1'b0 ;
  assign n10095 = ( n5100 & n10093 ) | ( n5100 & n10094 ) | ( n10093 & n10094 ) ;
  assign n10096 = n10045 ^ n2646 ^ 1'b0 ;
  assign n10097 = n1562 ^ n1348 ^ x120 ;
  assign n10098 = n10097 ^ n5456 ^ n5149 ;
  assign n10106 = n365 & n2623 ;
  assign n10107 = n5800 & n10106 ;
  assign n10102 = ( n621 & ~n2355 ) | ( n621 & n2957 ) | ( ~n2355 & n2957 ) ;
  assign n10103 = ~n1729 & n3039 ;
  assign n10104 = n10102 & n10103 ;
  assign n10101 = n5633 | n7859 ;
  assign n10105 = n10104 ^ n10101 ^ 1'b0 ;
  assign n10099 = n5631 ^ n468 ^ 1'b0 ;
  assign n10100 = n10099 ^ n8885 ^ n1695 ;
  assign n10108 = n10107 ^ n10105 ^ n10100 ;
  assign n10109 = ~n10098 & n10108 ;
  assign n10110 = n3627 & n4296 ;
  assign n10111 = ~n7250 & n7331 ;
  assign n10112 = n10110 | n10111 ;
  assign n10113 = n5479 | n10112 ;
  assign n10114 = n8472 ^ n2306 ^ n644 ;
  assign n10118 = n4502 ^ x45 ^ 1'b0 ;
  assign n10119 = n5940 & ~n10118 ;
  assign n10120 = ( n6281 & ~n9969 ) | ( n6281 & n10119 ) | ( ~n9969 & n10119 ) ;
  assign n10115 = n4424 ^ n1323 ^ 1'b0 ;
  assign n10116 = n3783 & n10115 ;
  assign n10117 = n5317 & n10116 ;
  assign n10121 = n10120 ^ n10117 ^ 1'b0 ;
  assign n10122 = ( ~n7353 & n10114 ) | ( ~n7353 & n10121 ) | ( n10114 & n10121 ) ;
  assign n10123 = n7820 ^ n2160 ^ 1'b0 ;
  assign n10124 = n2849 & n10123 ;
  assign n10125 = ~n10122 & n10124 ;
  assign n10126 = n10125 ^ n8361 ^ n6884 ;
  assign n10127 = n6771 ^ n5347 ^ 1'b0 ;
  assign n10128 = ( n757 & ~n1014 ) | ( n757 & n3557 ) | ( ~n1014 & n3557 ) ;
  assign n10129 = n10128 ^ n3205 ^ n2948 ;
  assign n10130 = ( n1799 & n3491 ) | ( n1799 & n6705 ) | ( n3491 & n6705 ) ;
  assign n10131 = n1928 | n4419 ;
  assign n10132 = ~n10130 & n10131 ;
  assign n10133 = n10132 ^ n5397 ^ 1'b0 ;
  assign n10134 = ( n10127 & ~n10129 ) | ( n10127 & n10133 ) | ( ~n10129 & n10133 ) ;
  assign n10135 = ~n8382 & n10134 ;
  assign n10136 = ~n5862 & n10135 ;
  assign n10137 = n9110 ^ n8340 ^ n6759 ;
  assign n10138 = n9474 ^ n6048 ^ n5602 ;
  assign n10139 = ~n9038 & n9690 ;
  assign n10140 = n9112 ^ n449 ^ 1'b0 ;
  assign n10141 = n7142 | n10140 ;
  assign n10142 = n9551 ^ n4442 ^ 1'b0 ;
  assign n10143 = n10142 ^ n2858 ^ 1'b0 ;
  assign n10144 = n6375 | n10143 ;
  assign n10145 = n10144 ^ n7600 ^ 1'b0 ;
  assign n10146 = ( ~n2024 & n9273 ) | ( ~n2024 & n10145 ) | ( n9273 & n10145 ) ;
  assign n10147 = n10141 | n10146 ;
  assign n10148 = n10147 ^ n7410 ^ 1'b0 ;
  assign n10149 = n3015 ^ x123 ^ 1'b0 ;
  assign n10150 = n6551 & ~n7439 ;
  assign n10151 = ( n6621 & n10149 ) | ( n6621 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = n9285 ^ n3946 ^ n3100 ;
  assign n10153 = n10152 ^ n3684 ^ 1'b0 ;
  assign n10154 = n10151 & n10153 ;
  assign n10155 = n1050 & n1813 ;
  assign n10156 = n2443 & ~n4533 ;
  assign n10157 = n2108 | n10156 ;
  assign n10158 = n353 ^ x228 ^ 1'b0 ;
  assign n10159 = n10157 & n10158 ;
  assign n10160 = n10159 ^ n1708 ^ 1'b0 ;
  assign n10161 = n10160 ^ n1554 ^ 1'b0 ;
  assign n10165 = n303 & n3109 ;
  assign n10166 = ( n2694 & n5653 ) | ( n2694 & ~n10165 ) | ( n5653 & ~n10165 ) ;
  assign n10162 = n4051 ^ n930 ^ 1'b0 ;
  assign n10163 = n8437 & n10162 ;
  assign n10164 = n3684 & n10163 ;
  assign n10167 = n10166 ^ n10164 ^ 1'b0 ;
  assign n10168 = n9623 ^ n2808 ^ 1'b0 ;
  assign n10169 = n4593 | n10168 ;
  assign n10170 = n4756 & ~n10169 ;
  assign n10171 = ~n5846 & n10170 ;
  assign n10172 = n8104 ^ n2768 ^ 1'b0 ;
  assign n10173 = n5148 ^ n3508 ^ n3472 ;
  assign n10174 = n10173 ^ n9888 ^ n5238 ;
  assign n10176 = ( n1104 & n1680 ) | ( n1104 & ~n2868 ) | ( n1680 & ~n2868 ) ;
  assign n10175 = ~n1127 & n9691 ;
  assign n10177 = n10176 ^ n10175 ^ 1'b0 ;
  assign n10178 = n2501 | n4574 ;
  assign n10179 = n10178 ^ n7815 ^ n2805 ;
  assign n10180 = x114 & n3639 ;
  assign n10181 = ~n4897 & n10180 ;
  assign n10182 = x239 & n353 ;
  assign n10183 = n3852 & n10182 ;
  assign n10184 = n2704 & ~n10183 ;
  assign n10185 = ( n4834 & ~n10181 ) | ( n4834 & n10184 ) | ( ~n10181 & n10184 ) ;
  assign n10186 = ( n6457 & ~n7559 ) | ( n6457 & n10185 ) | ( ~n7559 & n10185 ) ;
  assign n10187 = n3114 & n10186 ;
  assign n10188 = n1086 | n3910 ;
  assign n10189 = n6132 ^ n1081 ^ 1'b0 ;
  assign n10190 = n3031 ^ n466 ^ 1'b0 ;
  assign n10191 = n1359 & n10190 ;
  assign n10192 = n5372 & ~n10191 ;
  assign n10193 = ( ~n7322 & n10189 ) | ( ~n7322 & n10192 ) | ( n10189 & n10192 ) ;
  assign n10197 = ( n1635 & ~n1752 ) | ( n1635 & n7165 ) | ( ~n1752 & n7165 ) ;
  assign n10198 = n5189 & n10197 ;
  assign n10199 = n10198 ^ n6286 ^ 1'b0 ;
  assign n10194 = ~n1564 & n3927 ;
  assign n10195 = n8267 ^ n6729 ^ n4310 ;
  assign n10196 = n10194 & n10195 ;
  assign n10200 = n10199 ^ n10196 ^ 1'b0 ;
  assign n10201 = ( ~n5097 & n5447 ) | ( ~n5097 & n7831 ) | ( n5447 & n7831 ) ;
  assign n10203 = n4499 | n9559 ;
  assign n10204 = n5209 & ~n10203 ;
  assign n10202 = ( ~n836 & n5130 ) | ( ~n836 & n7377 ) | ( n5130 & n7377 ) ;
  assign n10205 = n10204 ^ n10202 ^ 1'b0 ;
  assign n10206 = n1133 & ~n10205 ;
  assign n10207 = ~n5508 & n5645 ;
  assign n10211 = ( n1116 & n4265 ) | ( n1116 & ~n4538 ) | ( n4265 & ~n4538 ) ;
  assign n10208 = n1118 | n3261 ;
  assign n10209 = n10208 ^ n6188 ^ 1'b0 ;
  assign n10210 = n10209 ^ n8091 ^ n7625 ;
  assign n10212 = n10211 ^ n10210 ^ n8313 ;
  assign n10213 = n10212 ^ n2651 ^ 1'b0 ;
  assign n10214 = n8148 | n10213 ;
  assign n10215 = ( n5912 & n8498 ) | ( n5912 & ~n10214 ) | ( n8498 & ~n10214 ) ;
  assign n10216 = ( n2201 & n4538 ) | ( n2201 & ~n10215 ) | ( n4538 & ~n10215 ) ;
  assign n10217 = n10207 & ~n10216 ;
  assign n10218 = n10217 ^ n885 ^ 1'b0 ;
  assign n10219 = n1634 | n4185 ;
  assign n10220 = n4371 & ~n10219 ;
  assign n10221 = n4218 & ~n4871 ;
  assign n10222 = n4416 & n10221 ;
  assign n10223 = n3665 & ~n10222 ;
  assign n10224 = n8992 & n10223 ;
  assign n10225 = n5133 & n10224 ;
  assign n10226 = n9348 ^ n6155 ^ n3301 ;
  assign n10230 = n9530 ^ n421 ^ 1'b0 ;
  assign n10227 = n804 & n9901 ;
  assign n10228 = ( ~n1961 & n3232 ) | ( ~n1961 & n10227 ) | ( n3232 & n10227 ) ;
  assign n10229 = n10228 ^ n10072 ^ x102 ;
  assign n10231 = n10230 ^ n10229 ^ n1998 ;
  assign n10233 = n6632 ^ n3372 ^ n901 ;
  assign n10234 = ( ~n1385 & n9421 ) | ( ~n1385 & n10233 ) | ( n9421 & n10233 ) ;
  assign n10232 = n5745 & ~n6782 ;
  assign n10235 = n10234 ^ n10232 ^ 1'b0 ;
  assign n10236 = n2555 & n5416 ;
  assign n10239 = n9124 ^ n7467 ^ 1'b0 ;
  assign n10237 = n3360 ^ n2474 ^ 1'b0 ;
  assign n10238 = n7213 & n10237 ;
  assign n10240 = n10239 ^ n10238 ^ n5398 ;
  assign n10241 = n1153 & n2868 ;
  assign n10242 = n10241 ^ n2097 ^ 1'b0 ;
  assign n10243 = ( n4283 & ~n8379 ) | ( n4283 & n10242 ) | ( ~n8379 & n10242 ) ;
  assign n10244 = n3972 | n10243 ;
  assign n10245 = n10244 ^ n4206 ^ 1'b0 ;
  assign n10250 = ( n1449 & n1666 ) | ( n1449 & ~n5577 ) | ( n1666 & ~n5577 ) ;
  assign n10251 = n2074 | n10250 ;
  assign n10246 = n7402 & n9660 ;
  assign n10247 = n4393 & n10246 ;
  assign n10248 = n10247 ^ n4442 ^ n1229 ;
  assign n10249 = n10248 ^ n9096 ^ n3518 ;
  assign n10252 = n10251 ^ n10249 ^ 1'b0 ;
  assign n10253 = n6011 ^ n2808 ^ n1505 ;
  assign n10254 = n10253 ^ n4194 ^ n3240 ;
  assign n10255 = n1975 | n10254 ;
  assign n10256 = n1318 ^ n1078 ^ 1'b0 ;
  assign n10257 = ~n2956 & n10256 ;
  assign n10258 = n10257 ^ n1405 ^ 1'b0 ;
  assign n10259 = x48 | n10258 ;
  assign n10260 = n4054 ^ n1780 ^ 1'b0 ;
  assign n10261 = n10259 & ~n10260 ;
  assign n10267 = ~n9002 & n9746 ;
  assign n10268 = n10267 ^ n9642 ^ n3807 ;
  assign n10269 = n7425 & ~n10268 ;
  assign n10262 = n1916 ^ x8 ^ 1'b0 ;
  assign n10263 = ~n4574 & n10262 ;
  assign n10264 = n8986 ^ n6556 ^ n1299 ;
  assign n10265 = ( n340 & n10263 ) | ( n340 & ~n10264 ) | ( n10263 & ~n10264 ) ;
  assign n10266 = n7282 & ~n10265 ;
  assign n10270 = n10269 ^ n10266 ^ 1'b0 ;
  assign n10271 = n3643 ^ n3364 ^ 1'b0 ;
  assign n10272 = n3156 & n10271 ;
  assign n10273 = n10272 ^ n7355 ^ 1'b0 ;
  assign n10274 = n8347 ^ n6538 ^ n6206 ;
  assign n10275 = n10274 ^ n3798 ^ 1'b0 ;
  assign n10276 = n6406 & n10275 ;
  assign n10277 = n10276 ^ n8052 ^ 1'b0 ;
  assign n10278 = ~n4032 & n10277 ;
  assign n10279 = n5951 & n10278 ;
  assign n10280 = n10279 ^ n8821 ^ 1'b0 ;
  assign n10281 = n3786 | n10280 ;
  assign n10282 = n6816 ^ n4724 ^ n1418 ;
  assign n10283 = n10282 ^ n8739 ^ n769 ;
  assign n10284 = n4902 ^ n1384 ^ n1239 ;
  assign n10285 = ~n5318 & n10284 ;
  assign n10286 = n9746 & n10285 ;
  assign n10287 = n6705 | n7854 ;
  assign n10288 = ( n1064 & ~n3272 ) | ( n1064 & n5229 ) | ( ~n3272 & n5229 ) ;
  assign n10289 = ( n1567 & ~n6282 ) | ( n1567 & n10288 ) | ( ~n6282 & n10288 ) ;
  assign n10290 = n6694 ^ n822 ^ n776 ;
  assign n10291 = ~n10289 & n10290 ;
  assign n10292 = n10287 & n10291 ;
  assign n10293 = n1647 ^ n919 ^ 1'b0 ;
  assign n10294 = n2073 & ~n10293 ;
  assign n10295 = ~n8530 & n10294 ;
  assign n10296 = ~n3855 & n8004 ;
  assign n10297 = n10296 ^ n3583 ^ 1'b0 ;
  assign n10298 = n10297 ^ n2877 ^ 1'b0 ;
  assign n10299 = n7200 ^ n2846 ^ n2430 ;
  assign n10300 = n1838 ^ x17 ^ 1'b0 ;
  assign n10301 = n10300 ^ n3833 ^ n2362 ;
  assign n10302 = n5406 | n5880 ;
  assign n10303 = n10301 | n10302 ;
  assign n10304 = n10303 ^ n3846 ^ 1'b0 ;
  assign n10305 = n10299 & ~n10304 ;
  assign n10306 = n5794 ^ n2947 ^ n1843 ;
  assign n10307 = n10306 ^ n2995 ^ 1'b0 ;
  assign n10308 = n851 & n9149 ;
  assign n10309 = n6005 ^ n3844 ^ 1'b0 ;
  assign n10310 = n10309 ^ n8043 ^ 1'b0 ;
  assign n10311 = n1061 & n4973 ;
  assign n10312 = n10311 ^ n627 ^ 1'b0 ;
  assign n10313 = n331 & ~n10312 ;
  assign n10314 = n10313 ^ n6176 ^ 1'b0 ;
  assign n10315 = n3718 ^ n3297 ^ 1'b0 ;
  assign n10316 = n10315 ^ n10210 ^ n9987 ;
  assign n10317 = n8885 ^ n7076 ^ x133 ;
  assign n10318 = ( n1132 & ~n3805 ) | ( n1132 & n10317 ) | ( ~n3805 & n10317 ) ;
  assign n10319 = ~n6574 & n8513 ;
  assign n10320 = n5597 & n10319 ;
  assign n10321 = n10318 & ~n10320 ;
  assign n10322 = n10321 ^ n6279 ^ 1'b0 ;
  assign n10323 = n4027 & n10322 ;
  assign n10324 = ~n1621 & n10323 ;
  assign n10325 = n7087 ^ n3327 ^ x74 ;
  assign n10326 = n10325 ^ n8675 ^ 1'b0 ;
  assign n10327 = n7803 | n10326 ;
  assign n10328 = n10327 ^ n9116 ^ n2696 ;
  assign n10329 = ( ~n3471 & n4332 ) | ( ~n3471 & n6938 ) | ( n4332 & n6938 ) ;
  assign n10330 = n10329 ^ n4983 ^ n530 ;
  assign n10331 = ( n806 & n1011 ) | ( n806 & ~n3274 ) | ( n1011 & ~n3274 ) ;
  assign n10332 = n10331 ^ n6149 ^ 1'b0 ;
  assign n10333 = n10332 ^ n9792 ^ n3050 ;
  assign n10334 = n3229 ^ n2368 ^ 1'b0 ;
  assign n10335 = n10334 ^ n3536 ^ n2461 ;
  assign n10336 = n5388 & ~n7293 ;
  assign n10337 = n10336 ^ n3594 ^ 1'b0 ;
  assign n10338 = n4289 ^ n2338 ^ 1'b0 ;
  assign n10339 = n5439 & n10338 ;
  assign n10340 = ( ~n8848 & n10337 ) | ( ~n8848 & n10339 ) | ( n10337 & n10339 ) ;
  assign n10341 = n7281 & n10340 ;
  assign n10342 = ~n10335 & n10341 ;
  assign n10343 = x134 & n4965 ;
  assign n10344 = n305 & n10343 ;
  assign n10345 = n10344 ^ n3091 ^ 1'b0 ;
  assign n10346 = n10342 | n10345 ;
  assign n10347 = n10346 ^ n7164 ^ n1963 ;
  assign n10348 = ( n2024 & ~n7643 ) | ( n2024 & n9715 ) | ( ~n7643 & n9715 ) ;
  assign n10349 = n7293 ^ n6611 ^ 1'b0 ;
  assign n10350 = n3026 & ~n10349 ;
  assign n10351 = n10350 ^ n737 ^ 1'b0 ;
  assign n10352 = n6196 & n10351 ;
  assign n10353 = n10352 ^ n8008 ^ 1'b0 ;
  assign n10354 = n10353 ^ n6936 ^ n3830 ;
  assign n10356 = n2042 ^ n1863 ^ n1222 ;
  assign n10357 = n2059 & ~n10356 ;
  assign n10358 = n10357 ^ n6048 ^ 1'b0 ;
  assign n10355 = ( n1468 & n4896 ) | ( n1468 & ~n8574 ) | ( n4896 & ~n8574 ) ;
  assign n10359 = n10358 ^ n10355 ^ n7102 ;
  assign n10360 = n2865 ^ n445 ^ 1'b0 ;
  assign n10361 = ( n5027 & n7422 ) | ( n5027 & n8123 ) | ( n7422 & n8123 ) ;
  assign n10362 = n3633 ^ n3256 ^ 1'b0 ;
  assign n10363 = n5242 | n10362 ;
  assign n10364 = n9904 | n10363 ;
  assign n10365 = n5205 ^ n4883 ^ 1'b0 ;
  assign n10372 = n7814 ^ n7794 ^ n4725 ;
  assign n10366 = n4457 | n6274 ;
  assign n10367 = n604 | n10366 ;
  assign n10368 = n9580 ^ n4552 ^ 1'b0 ;
  assign n10369 = n10367 & ~n10368 ;
  assign n10370 = n10369 ^ n5940 ^ 1'b0 ;
  assign n10371 = ( n723 & n7482 ) | ( n723 & ~n10370 ) | ( n7482 & ~n10370 ) ;
  assign n10373 = n10372 ^ n10371 ^ n7187 ;
  assign n10376 = ( n2384 & n3066 ) | ( n2384 & ~n3203 ) | ( n3066 & ~n3203 ) ;
  assign n10375 = ~n3675 & n5116 ;
  assign n10377 = n10376 ^ n10375 ^ 1'b0 ;
  assign n10374 = ~n3734 & n8493 ;
  assign n10378 = n10377 ^ n10374 ^ 1'b0 ;
  assign n10379 = ( x95 & ~n388 ) | ( x95 & n5248 ) | ( ~n388 & n5248 ) ;
  assign n10380 = n10379 ^ n8551 ^ 1'b0 ;
  assign n10381 = n3330 | n4793 ;
  assign n10382 = n10381 ^ n3054 ^ 1'b0 ;
  assign n10383 = n10382 ^ n3802 ^ 1'b0 ;
  assign n10384 = n466 & ~n10383 ;
  assign n10385 = n10384 ^ n5252 ^ 1'b0 ;
  assign n10386 = n7596 & n10385 ;
  assign n10387 = n1053 | n2755 ;
  assign n10388 = ( n6164 & ~n6954 ) | ( n6164 & n10387 ) | ( ~n6954 & n10387 ) ;
  assign n10389 = n5679 ^ n5431 ^ n3180 ;
  assign n10390 = n5060 ^ n3278 ^ 1'b0 ;
  assign n10391 = n10389 & n10390 ;
  assign n10392 = n9789 & n10391 ;
  assign n10393 = ~n9153 & n10392 ;
  assign n10394 = ( n2510 & n6237 ) | ( n2510 & n10393 ) | ( n6237 & n10393 ) ;
  assign n10395 = ~n720 & n1377 ;
  assign n10396 = ~n2199 & n10395 ;
  assign n10397 = n6677 ^ n684 ^ 1'b0 ;
  assign n10398 = n10396 | n10397 ;
  assign n10399 = ( n2482 & n3180 ) | ( n2482 & ~n6264 ) | ( n3180 & ~n6264 ) ;
  assign n10400 = n10369 ^ n9901 ^ n7911 ;
  assign n10401 = ( n4338 & n10399 ) | ( n4338 & ~n10400 ) | ( n10399 & ~n10400 ) ;
  assign n10408 = n3127 ^ x15 ^ 1'b0 ;
  assign n10409 = ( ~n644 & n4010 ) | ( ~n644 & n10408 ) | ( n4010 & n10408 ) ;
  assign n10407 = n1197 & ~n1617 ;
  assign n10410 = n10409 ^ n10407 ^ 1'b0 ;
  assign n10402 = n2040 & n4331 ;
  assign n10403 = ~n2281 & n10402 ;
  assign n10404 = n10403 ^ n7701 ^ x132 ;
  assign n10405 = ( n5836 & n6844 ) | ( n5836 & n10404 ) | ( n6844 & n10404 ) ;
  assign n10406 = ~n1611 & n10405 ;
  assign n10411 = n10410 ^ n10406 ^ n1511 ;
  assign n10412 = n9232 ^ n5251 ^ 1'b0 ;
  assign n10413 = n10411 & ~n10412 ;
  assign n10414 = n2917 & ~n3099 ;
  assign n10415 = n10414 ^ n2221 ^ 1'b0 ;
  assign n10416 = n5112 ^ n4776 ^ n1217 ;
  assign n10417 = n10415 & ~n10416 ;
  assign n10418 = n10417 ^ n1433 ^ 1'b0 ;
  assign n10419 = n7573 ^ n3269 ^ n2808 ;
  assign n10420 = n2485 & ~n5416 ;
  assign n10421 = n10420 ^ n4211 ^ 1'b0 ;
  assign n10422 = ~n1814 & n10421 ;
  assign n10423 = ( ~x209 & n3479 ) | ( ~x209 & n8962 ) | ( n3479 & n8962 ) ;
  assign n10424 = n5567 & n10423 ;
  assign n10425 = ~n10422 & n10424 ;
  assign n10430 = ~n277 & n4908 ;
  assign n10431 = n10430 ^ n6423 ^ 1'b0 ;
  assign n10432 = ~n3880 & n10431 ;
  assign n10433 = n2477 | n10432 ;
  assign n10426 = n10007 ^ n4421 ^ 1'b0 ;
  assign n10427 = ( n3080 & ~n4436 ) | ( n3080 & n5440 ) | ( ~n4436 & n5440 ) ;
  assign n10428 = n10427 ^ n6395 ^ 1'b0 ;
  assign n10429 = n10426 | n10428 ;
  assign n10434 = n10433 ^ n10429 ^ 1'b0 ;
  assign n10435 = n3855 | n5522 ;
  assign n10436 = n1919 & ~n10435 ;
  assign n10437 = n1206 | n10436 ;
  assign n10438 = n8985 | n10437 ;
  assign n10439 = n10129 & n10438 ;
  assign n10440 = n1773 & n10439 ;
  assign n10441 = n3163 & ~n10440 ;
  assign n10442 = n10441 ^ n1349 ^ 1'b0 ;
  assign n10443 = ( n3648 & n6397 ) | ( n3648 & n7063 ) | ( n6397 & n7063 ) ;
  assign n10444 = ~n10442 & n10443 ;
  assign n10445 = ~n338 & n10444 ;
  assign n10446 = ~x183 & n1682 ;
  assign n10447 = n4787 & n4919 ;
  assign n10448 = n9854 & n10447 ;
  assign n10449 = n10448 ^ n879 ^ 1'b0 ;
  assign n10450 = n952 & ~n10449 ;
  assign n10451 = ( n2975 & n4349 ) | ( n2975 & n10450 ) | ( n4349 & n10450 ) ;
  assign n10452 = n8595 ^ n7934 ^ n3353 ;
  assign n10453 = n1236 | n3008 ;
  assign n10454 = n10453 ^ n374 ^ 1'b0 ;
  assign n10455 = n10454 ^ n2194 ^ 1'b0 ;
  assign n10456 = n8599 & n10455 ;
  assign n10457 = ( n6114 & ~n7184 ) | ( n6114 & n10456 ) | ( ~n7184 & n10456 ) ;
  assign n10458 = n3349 ^ n3068 ^ n951 ;
  assign n10459 = ~n5231 & n10458 ;
  assign n10460 = n10457 & n10459 ;
  assign n10461 = n4958 ^ n3435 ^ 1'b0 ;
  assign n10462 = ~n6462 & n10461 ;
  assign n10463 = n4527 & n10462 ;
  assign n10464 = n10463 ^ n4701 ^ n3839 ;
  assign n10467 = n2393 & n7217 ;
  assign n10468 = n10467 ^ n3994 ^ 1'b0 ;
  assign n10465 = n1279 & n1746 ;
  assign n10466 = n10465 ^ n2532 ^ 1'b0 ;
  assign n10469 = n10468 ^ n10466 ^ n7223 ;
  assign n10470 = ~n6528 & n8726 ;
  assign n10471 = ~n10469 & n10470 ;
  assign n10472 = n8458 | n9802 ;
  assign n10473 = ~n579 & n6186 ;
  assign n10474 = n10473 ^ n3498 ^ 1'b0 ;
  assign n10475 = ~n3992 & n5635 ;
  assign n10476 = n10475 ^ n4488 ^ 1'b0 ;
  assign n10478 = n8642 ^ n2123 ^ n1252 ;
  assign n10479 = ( n1897 & n9845 ) | ( n1897 & n10478 ) | ( n9845 & n10478 ) ;
  assign n10477 = ( n3422 & ~n3653 ) | ( n3422 & n4268 ) | ( ~n3653 & n4268 ) ;
  assign n10480 = n10479 ^ n10477 ^ n9413 ;
  assign n10481 = ( n5650 & n10476 ) | ( n5650 & ~n10480 ) | ( n10476 & ~n10480 ) ;
  assign n10482 = n3041 ^ n2299 ^ 1'b0 ;
  assign n10483 = ( n446 & n1174 ) | ( n446 & n3222 ) | ( n1174 & n3222 ) ;
  assign n10484 = n7722 ^ n5815 ^ 1'b0 ;
  assign n10485 = n10483 & n10484 ;
  assign n10486 = n10485 ^ n4166 ^ 1'b0 ;
  assign n10487 = n5276 | n10486 ;
  assign n10488 = ( n4329 & ~n5677 ) | ( n4329 & n10482 ) | ( ~n5677 & n10482 ) ;
  assign n10489 = n5000 ^ n2793 ^ 1'b0 ;
  assign n10495 = n5907 ^ n3289 ^ 1'b0 ;
  assign n10490 = n8620 ^ n518 ^ 1'b0 ;
  assign n10491 = n6043 ^ x191 ^ 1'b0 ;
  assign n10492 = n10490 | n10491 ;
  assign n10493 = n1984 & ~n10492 ;
  assign n10494 = ~n8079 & n10493 ;
  assign n10496 = n10495 ^ n10494 ^ n7540 ;
  assign n10497 = n2029 | n10496 ;
  assign n10498 = n10497 ^ n6415 ^ 1'b0 ;
  assign n10499 = ~n751 & n2258 ;
  assign n10500 = n10499 ^ n1254 ^ n502 ;
  assign n10501 = ( n8276 & n9033 ) | ( n8276 & n10500 ) | ( n9033 & n10500 ) ;
  assign n10503 = n8011 ^ n3732 ^ 1'b0 ;
  assign n10504 = n1706 & ~n10503 ;
  assign n10502 = ( n841 & ~n2029 ) | ( n841 & n3830 ) | ( ~n2029 & n3830 ) ;
  assign n10505 = n10504 ^ n10502 ^ 1'b0 ;
  assign n10506 = n9682 ^ n1409 ^ 1'b0 ;
  assign n10507 = n2523 & n5662 ;
  assign n10513 = ~n2566 & n8642 ;
  assign n10508 = n1287 ^ n429 ^ 1'b0 ;
  assign n10509 = n4763 & ~n10508 ;
  assign n10510 = n3947 ^ n1488 ^ 1'b0 ;
  assign n10511 = n10509 & n10510 ;
  assign n10512 = ~n3430 & n10511 ;
  assign n10514 = n10513 ^ n10512 ^ 1'b0 ;
  assign n10515 = n7518 ^ n6530 ^ 1'b0 ;
  assign n10516 = n1385 & n10515 ;
  assign n10518 = ( x112 & ~n299 ) | ( x112 & n3303 ) | ( ~n299 & n3303 ) ;
  assign n10519 = n10518 ^ n6818 ^ n1285 ;
  assign n10520 = n10519 ^ n3875 ^ n1090 ;
  assign n10521 = ( n4072 & ~n9603 ) | ( n4072 & n10520 ) | ( ~n9603 & n10520 ) ;
  assign n10522 = n9519 & ~n10521 ;
  assign n10523 = n6528 & n10522 ;
  assign n10517 = ( n2741 & ~n4506 ) | ( n2741 & n6871 ) | ( ~n4506 & n6871 ) ;
  assign n10524 = n10523 ^ n10517 ^ n5425 ;
  assign n10525 = n4635 & n8795 ;
  assign n10526 = n10525 ^ n8358 ^ 1'b0 ;
  assign n10527 = n3512 ^ n2683 ^ 1'b0 ;
  assign n10528 = ( n340 & n6015 ) | ( n340 & ~n10527 ) | ( n6015 & ~n10527 ) ;
  assign n10529 = n5476 ^ n4889 ^ n1961 ;
  assign n10530 = n10529 ^ n7592 ^ 1'b0 ;
  assign n10531 = ( ~n431 & n1906 ) | ( ~n431 & n2893 ) | ( n1906 & n2893 ) ;
  assign n10532 = n10531 ^ n2908 ^ n1580 ;
  assign n10534 = x132 | n2377 ;
  assign n10533 = n268 & n4728 ;
  assign n10535 = n10534 ^ n10533 ^ n2100 ;
  assign n10543 = ( n1903 & ~n2461 ) | ( n1903 & n3672 ) | ( ~n2461 & n3672 ) ;
  assign n10539 = n2743 | n5411 ;
  assign n10540 = n2438 | n10539 ;
  assign n10536 = ( ~n362 & n3512 ) | ( ~n362 & n6558 ) | ( n3512 & n6558 ) ;
  assign n10537 = ( n2119 & n2549 ) | ( n2119 & n10536 ) | ( n2549 & n10536 ) ;
  assign n10538 = ~n394 & n10537 ;
  assign n10541 = n10540 ^ n10538 ^ 1'b0 ;
  assign n10542 = n3075 | n10541 ;
  assign n10544 = n10543 ^ n10542 ^ 1'b0 ;
  assign n10545 = ( n9771 & n10535 ) | ( n9771 & ~n10544 ) | ( n10535 & ~n10544 ) ;
  assign n10546 = n1669 & ~n6176 ;
  assign n10547 = n3577 ^ n615 ^ 1'b0 ;
  assign n10548 = n6615 & n10547 ;
  assign n10549 = n9857 & n10548 ;
  assign n10550 = ( ~n1130 & n10546 ) | ( ~n1130 & n10549 ) | ( n10546 & n10549 ) ;
  assign n10551 = n3598 & ~n5235 ;
  assign n10554 = n4692 ^ n3482 ^ 1'b0 ;
  assign n10555 = n4684 & n10554 ;
  assign n10552 = ( n4036 & n5509 ) | ( n4036 & n5848 ) | ( n5509 & n5848 ) ;
  assign n10553 = ~n6705 & n10552 ;
  assign n10556 = n10555 ^ n10553 ^ n3508 ;
  assign n10557 = ( n1173 & ~n3106 ) | ( n1173 & n10556 ) | ( ~n3106 & n10556 ) ;
  assign n10558 = n1591 ^ n1331 ^ 1'b0 ;
  assign n10559 = x209 & ~n10558 ;
  assign n10560 = n7270 & n10559 ;
  assign n10561 = n10560 ^ n5688 ^ 1'b0 ;
  assign n10562 = n10561 ^ n7859 ^ n2351 ;
  assign n10563 = ( n10551 & n10557 ) | ( n10551 & ~n10562 ) | ( n10557 & ~n10562 ) ;
  assign n10564 = n4690 & ~n5289 ;
  assign n10565 = n10563 & ~n10564 ;
  assign n10566 = ( n5286 & ~n7897 ) | ( n5286 & n9336 ) | ( ~n7897 & n9336 ) ;
  assign n10567 = x31 & ~n10566 ;
  assign n10568 = n7190 & n10567 ;
  assign n10569 = ~n2349 & n10568 ;
  assign n10570 = n5082 ^ n2036 ^ n1537 ;
  assign n10571 = ~x133 & n10570 ;
  assign n10572 = n10571 ^ n4592 ^ n4413 ;
  assign n10573 = n3264 & ~n10572 ;
  assign n10574 = ~n9378 & n10559 ;
  assign n10575 = n10573 & n10574 ;
  assign n10587 = n8062 ^ x38 ^ 1'b0 ;
  assign n10588 = x106 & n10587 ;
  assign n10577 = n8638 ^ n6648 ^ x61 ;
  assign n10578 = n10577 ^ n2525 ^ 1'b0 ;
  assign n10579 = n2437 | n10578 ;
  assign n10580 = n10579 ^ n6321 ^ 1'b0 ;
  assign n10576 = n4677 & ~n5989 ;
  assign n10581 = n10580 ^ n10576 ^ 1'b0 ;
  assign n10584 = n5642 | n7750 ;
  assign n10582 = ~n1475 & n2056 ;
  assign n10583 = ~n2148 & n10582 ;
  assign n10585 = n10584 ^ n10583 ^ n1681 ;
  assign n10586 = n10581 & ~n10585 ;
  assign n10589 = n10588 ^ n10586 ^ 1'b0 ;
  assign n10590 = n6207 & ~n10589 ;
  assign n10591 = n10590 ^ n4363 ^ 1'b0 ;
  assign n10592 = n9473 ^ n3080 ^ n695 ;
  assign n10593 = ~n1294 & n4284 ;
  assign n10594 = n1317 | n3118 ;
  assign n10595 = n10593 & ~n10594 ;
  assign n10596 = ( n6866 & n10592 ) | ( n6866 & ~n10595 ) | ( n10592 & ~n10595 ) ;
  assign n10597 = n10596 ^ n9369 ^ n8475 ;
  assign n10598 = n1057 & ~n2904 ;
  assign n10599 = n6854 & n10598 ;
  assign n10600 = n10599 ^ n4060 ^ 1'b0 ;
  assign n10601 = ~n1202 & n10600 ;
  assign n10602 = n7867 & n10601 ;
  assign n10603 = n10602 ^ n1947 ^ 1'b0 ;
  assign n10604 = n4730 ^ x115 ^ 1'b0 ;
  assign n10605 = n5357 & ~n10604 ;
  assign n10606 = n2802 & n10605 ;
  assign n10607 = n871 | n10606 ;
  assign n10608 = n10607 ^ n1898 ^ 1'b0 ;
  assign n10609 = n7238 | n10608 ;
  assign n10610 = n8254 | n10609 ;
  assign n10611 = n6478 ^ n820 ^ 1'b0 ;
  assign n10612 = ~n3032 & n10611 ;
  assign n10613 = ( ~n3058 & n10610 ) | ( ~n3058 & n10612 ) | ( n10610 & n10612 ) ;
  assign n10614 = n1006 ^ x246 ^ 1'b0 ;
  assign n10615 = n1978 | n10614 ;
  assign n10616 = n8482 & ~n10615 ;
  assign n10617 = n1632 & n10616 ;
  assign n10619 = x186 & n545 ;
  assign n10620 = n10619 ^ n6395 ^ 1'b0 ;
  assign n10621 = n10620 ^ n8182 ^ 1'b0 ;
  assign n10618 = n3721 & n8644 ;
  assign n10622 = n10621 ^ n10618 ^ 1'b0 ;
  assign n10623 = n2276 & ~n8619 ;
  assign n10624 = n10623 ^ n6101 ^ n1555 ;
  assign n10625 = n8716 ^ n1601 ^ 1'b0 ;
  assign n10626 = n7409 & ~n10625 ;
  assign n10627 = n10626 ^ n6697 ^ n3313 ;
  assign n10628 = ( n5236 & ~n5669 ) | ( n5236 & n6729 ) | ( ~n5669 & n6729 ) ;
  assign n10629 = n1997 | n10628 ;
  assign n10630 = n10629 ^ n5403 ^ 1'b0 ;
  assign n10631 = n8620 ^ n5272 ^ n2890 ;
  assign n10633 = n1607 | n9246 ;
  assign n10632 = ~n468 & n1994 ;
  assign n10634 = n10633 ^ n10632 ^ 1'b0 ;
  assign n10635 = ~n8223 & n10634 ;
  assign n10636 = n10635 ^ n8685 ^ 1'b0 ;
  assign n10637 = ~n4765 & n7922 ;
  assign n10638 = n865 & n1921 ;
  assign n10639 = n3693 | n10416 ;
  assign n10640 = n10638 & n10639 ;
  assign n10641 = n10640 ^ n4091 ^ 1'b0 ;
  assign n10643 = n1175 & n2384 ;
  assign n10644 = n7823 & n10643 ;
  assign n10645 = n9146 & ~n10644 ;
  assign n10642 = n4744 & ~n8795 ;
  assign n10646 = n10645 ^ n10642 ^ 1'b0 ;
  assign n10647 = n9580 ^ n859 ^ 1'b0 ;
  assign n10648 = n10647 ^ n6433 ^ n3689 ;
  assign n10658 = n1906 ^ x3 ^ 1'b0 ;
  assign n10659 = n2382 & n10658 ;
  assign n10649 = n1458 & ~n5948 ;
  assign n10650 = n6809 & n10649 ;
  assign n10651 = n10650 ^ n9364 ^ 1'b0 ;
  assign n10652 = n7859 | n10651 ;
  assign n10655 = n673 ^ n609 ^ x63 ;
  assign n10653 = n2722 ^ n1186 ^ x158 ;
  assign n10654 = n10653 ^ n6563 ^ n2730 ;
  assign n10656 = n10655 ^ n10654 ^ 1'b0 ;
  assign n10657 = ( n6301 & n10652 ) | ( n6301 & n10656 ) | ( n10652 & n10656 ) ;
  assign n10660 = n10659 ^ n10657 ^ n4793 ;
  assign n10661 = ( n1451 & n10648 ) | ( n1451 & n10660 ) | ( n10648 & n10660 ) ;
  assign n10662 = n2036 & n8119 ;
  assign n10663 = n4582 & n10662 ;
  assign n10672 = ( n1858 & n2330 ) | ( n1858 & ~n8203 ) | ( n2330 & ~n8203 ) ;
  assign n10666 = x134 & ~n1446 ;
  assign n10667 = ~n2608 & n10666 ;
  assign n10668 = n2775 & n10667 ;
  assign n10669 = ( x214 & ~x231 ) | ( x214 & n10668 ) | ( ~x231 & n10668 ) ;
  assign n10670 = n10669 ^ n5370 ^ n1334 ;
  assign n10671 = n8999 & ~n10670 ;
  assign n10664 = n9996 & ~n10002 ;
  assign n10665 = n10664 ^ x148 ^ 1'b0 ;
  assign n10673 = n10672 ^ n10671 ^ n10665 ;
  assign n10674 = ( n951 & ~n4644 ) | ( n951 & n7783 ) | ( ~n4644 & n7783 ) ;
  assign n10675 = n8324 | n10674 ;
  assign n10676 = ( x210 & n4890 ) | ( x210 & ~n10675 ) | ( n4890 & ~n10675 ) ;
  assign n10677 = n10204 & n10676 ;
  assign n10678 = ( x151 & n7198 ) | ( x151 & n10677 ) | ( n7198 & n10677 ) ;
  assign n10679 = n4797 ^ n2244 ^ 1'b0 ;
  assign n10680 = n10679 ^ n7185 ^ 1'b0 ;
  assign n10681 = ( x10 & ~n462 ) | ( x10 & n1673 ) | ( ~n462 & n1673 ) ;
  assign n10682 = n2670 & n10681 ;
  assign n10683 = n1301 ^ n1051 ^ 1'b0 ;
  assign n10684 = n2680 | n10683 ;
  assign n10685 = n2512 & ~n10684 ;
  assign n10686 = ~n4728 & n10685 ;
  assign n10687 = n10686 ^ n8667 ^ 1'b0 ;
  assign n10688 = ~n10682 & n10687 ;
  assign n10689 = ( n4970 & n9073 ) | ( n4970 & ~n10688 ) | ( n9073 & ~n10688 ) ;
  assign n10690 = n9960 ^ n8953 ^ n2057 ;
  assign n10691 = n5002 ^ n1988 ^ n665 ;
  assign n10692 = n1283 | n10691 ;
  assign n10693 = ~n3420 & n5917 ;
  assign n10694 = n10693 ^ n280 ^ 1'b0 ;
  assign n10695 = n10694 ^ n5716 ^ n1470 ;
  assign n10696 = ( n2814 & n6244 ) | ( n2814 & ~n10695 ) | ( n6244 & ~n10695 ) ;
  assign n10697 = n4754 & n10696 ;
  assign n10698 = n10692 & n10697 ;
  assign n10699 = ( n4052 & n7537 ) | ( n4052 & n10698 ) | ( n7537 & n10698 ) ;
  assign n10700 = n4251 ^ n2894 ^ 1'b0 ;
  assign n10701 = ~n2646 & n10700 ;
  assign n10702 = n10701 ^ n6457 ^ n3336 ;
  assign n10703 = n5015 & n5846 ;
  assign n10705 = n4272 ^ n3989 ^ 1'b0 ;
  assign n10706 = n5683 & n10705 ;
  assign n10704 = ~n3830 & n9300 ;
  assign n10707 = n10706 ^ n10704 ^ 1'b0 ;
  assign n10708 = n6285 | n6297 ;
  assign n10709 = n10707 & ~n10708 ;
  assign n10710 = n8737 | n10709 ;
  assign n10711 = n1837 & ~n5078 ;
  assign n10712 = n1470 & n10711 ;
  assign n10713 = n6793 ^ n1986 ^ x7 ;
  assign n10714 = x82 & ~n3865 ;
  assign n10715 = n10714 ^ n9387 ^ n5121 ;
  assign n10719 = ( n2569 & ~n6891 ) | ( n2569 & n9306 ) | ( ~n6891 & n9306 ) ;
  assign n10720 = n5080 & ~n7442 ;
  assign n10721 = n10720 ^ n9447 ^ 1'b0 ;
  assign n10722 = ~n10719 & n10721 ;
  assign n10716 = n1560 | n10580 ;
  assign n10717 = n1655 & ~n10716 ;
  assign n10718 = n10483 & ~n10717 ;
  assign n10723 = n10722 ^ n10718 ^ 1'b0 ;
  assign n10724 = n8566 ^ n4201 ^ 1'b0 ;
  assign n10725 = n9126 ^ n8711 ^ 1'b0 ;
  assign n10726 = n10119 ^ n3569 ^ 1'b0 ;
  assign n10727 = n5175 & n10726 ;
  assign n10728 = n10727 ^ n3578 ^ 1'b0 ;
  assign n10729 = ( ~n6789 & n10725 ) | ( ~n6789 & n10728 ) | ( n10725 & n10728 ) ;
  assign n10730 = n10729 ^ n8169 ^ x102 ;
  assign n10731 = ~n3744 & n6846 ;
  assign n10732 = n2865 ^ n2779 ^ n1016 ;
  assign n10733 = ( ~n1511 & n6377 ) | ( ~n1511 & n10732 ) | ( n6377 & n10732 ) ;
  assign n10734 = n10733 ^ n3165 ^ 1'b0 ;
  assign n10735 = ~n2766 & n10734 ;
  assign n10736 = n6587 ^ n3490 ^ 1'b0 ;
  assign n10737 = n10736 ^ x248 ^ 1'b0 ;
  assign n10738 = ( n1362 & n4848 ) | ( n1362 & n6579 ) | ( n4848 & n6579 ) ;
  assign n10739 = ~n2795 & n4847 ;
  assign n10740 = n10738 | n10739 ;
  assign n10741 = n4946 | n8093 ;
  assign n10742 = n3604 & n4573 ;
  assign n10743 = n7892 ^ n2682 ^ 1'b0 ;
  assign n10744 = n818 | n10743 ;
  assign n10745 = n10744 ^ n2156 ^ 1'b0 ;
  assign n10746 = n3762 ^ n1603 ^ 1'b0 ;
  assign n10747 = ~n10745 & n10746 ;
  assign n10748 = n10747 ^ n2950 ^ 1'b0 ;
  assign n10749 = n6246 ^ n5500 ^ 1'b0 ;
  assign n10750 = n9344 & n10749 ;
  assign n10751 = ( n1838 & n2944 ) | ( n1838 & ~n5741 ) | ( n2944 & ~n5741 ) ;
  assign n10752 = n5484 ^ n1758 ^ 1'b0 ;
  assign n10753 = n1671 | n3732 ;
  assign n10754 = ( ~n1062 & n1445 ) | ( ~n1062 & n3219 ) | ( n1445 & n3219 ) ;
  assign n10755 = n10277 & ~n10754 ;
  assign n10756 = n5564 ^ n487 ^ 1'b0 ;
  assign n10757 = n4842 & ~n10756 ;
  assign n10758 = ~n6918 & n10278 ;
  assign n10759 = ~n8500 & n10758 ;
  assign n10766 = n3399 ^ n1926 ^ 1'b0 ;
  assign n10761 = n5529 ^ n4065 ^ 1'b0 ;
  assign n10760 = n2930 ^ n1047 ^ n285 ;
  assign n10762 = n10761 ^ n10760 ^ 1'b0 ;
  assign n10763 = n2136 & ~n10762 ;
  assign n10764 = n7716 ^ n5231 ^ 1'b0 ;
  assign n10765 = n10763 & ~n10764 ;
  assign n10767 = n10766 ^ n10765 ^ n5796 ;
  assign n10768 = n4721 & n8992 ;
  assign n10769 = n4340 & n10768 ;
  assign n10770 = n10769 ^ n4440 ^ 1'b0 ;
  assign n10773 = ~n4070 & n4622 ;
  assign n10771 = n8382 ^ n4850 ^ 1'b0 ;
  assign n10772 = n8282 & n10771 ;
  assign n10774 = n10773 ^ n10772 ^ 1'b0 ;
  assign n10775 = ( ~n2314 & n7017 ) | ( ~n2314 & n10774 ) | ( n7017 & n10774 ) ;
  assign n10777 = n8605 & ~n9608 ;
  assign n10776 = n5320 ^ n4223 ^ n3585 ;
  assign n10778 = n10777 ^ n10776 ^ 1'b0 ;
  assign n10779 = n9489 & ~n10778 ;
  assign n10780 = n6138 ^ n2362 ^ n2041 ;
  assign n10781 = ( n1828 & ~n3026 ) | ( n1828 & n10780 ) | ( ~n3026 & n10780 ) ;
  assign n10782 = n8769 | n10781 ;
  assign n10783 = n8186 | n10782 ;
  assign n10788 = ~n5673 & n7519 ;
  assign n10786 = n2445 ^ n434 ^ 1'b0 ;
  assign n10787 = ~n9378 & n10786 ;
  assign n10789 = n10788 ^ n10787 ^ 1'b0 ;
  assign n10784 = ~n2397 & n3875 ;
  assign n10785 = n3804 & n10784 ;
  assign n10790 = n10789 ^ n10785 ^ 1'b0 ;
  assign n10791 = n10783 & ~n10790 ;
  assign n10792 = ( ~n2282 & n4315 ) | ( ~n2282 & n4556 ) | ( n4315 & n4556 ) ;
  assign n10793 = n9988 ^ n7358 ^ n716 ;
  assign n10794 = ( ~n4212 & n10792 ) | ( ~n4212 & n10793 ) | ( n10792 & n10793 ) ;
  assign n10800 = ( n491 & n5284 ) | ( n491 & n6445 ) | ( n5284 & n6445 ) ;
  assign n10797 = n2068 & n2767 ;
  assign n10798 = n10797 ^ n4350 ^ n3471 ;
  assign n10795 = n1199 | n3141 ;
  assign n10796 = n10795 ^ n7431 ^ 1'b0 ;
  assign n10799 = n10798 ^ n10796 ^ n7433 ;
  assign n10801 = n10800 ^ n10799 ^ n4842 ;
  assign n10802 = n9552 ^ n9267 ^ 1'b0 ;
  assign n10803 = n1996 ^ x117 ^ 1'b0 ;
  assign n10804 = n10802 & n10803 ;
  assign n10805 = ~n2306 & n9246 ;
  assign n10806 = ~n5652 & n10805 ;
  assign n10807 = ~n4432 & n7446 ;
  assign n10808 = n10807 ^ n983 ^ 1'b0 ;
  assign n10809 = n4835 & ~n10808 ;
  assign n10810 = n10808 & n10809 ;
  assign n10811 = n9467 ^ n5551 ^ n3206 ;
  assign n10812 = ~n8335 & n9622 ;
  assign n10813 = n10812 ^ n4462 ^ 1'b0 ;
  assign n10814 = n926 | n2698 ;
  assign n10815 = n10814 ^ n2247 ^ 1'b0 ;
  assign n10816 = n10815 ^ n4723 ^ 1'b0 ;
  assign n10817 = n3462 & ~n10816 ;
  assign n10818 = n1223 & ~n10817 ;
  assign n10819 = n10671 & n10818 ;
  assign n10820 = n4956 ^ n4026 ^ 1'b0 ;
  assign n10821 = n10820 ^ n2437 ^ 1'b0 ;
  assign n10822 = ~n10819 & n10821 ;
  assign n10823 = n10569 ^ n3468 ^ n2344 ;
  assign n10824 = ( ~n841 & n1559 ) | ( ~n841 & n4346 ) | ( n1559 & n4346 ) ;
  assign n10825 = n6353 | n10656 ;
  assign n10826 = n10825 ^ n6194 ^ 1'b0 ;
  assign n10827 = n2476 ^ n2234 ^ n1945 ;
  assign n10828 = n3809 | n10827 ;
  assign n10829 = n7706 | n10828 ;
  assign n10830 = ~n4340 & n10829 ;
  assign n10831 = n10830 ^ n4704 ^ 1'b0 ;
  assign n10832 = x81 | n5926 ;
  assign n10833 = n10832 ^ n3814 ^ 1'b0 ;
  assign n10834 = n6873 ^ n1719 ^ 1'b0 ;
  assign n10835 = n10833 & n10834 ;
  assign n10836 = ~n6495 & n10835 ;
  assign n10837 = n5627 & ~n9530 ;
  assign n10838 = n6977 & n10837 ;
  assign n10839 = ( n6671 & n8084 ) | ( n6671 & ~n8383 ) | ( n8084 & ~n8383 ) ;
  assign n10840 = n8585 ^ n2956 ^ 1'b0 ;
  assign n10841 = n2413 & n7383 ;
  assign n10842 = n3289 & n10841 ;
  assign n10843 = ( n8315 & n10840 ) | ( n8315 & n10842 ) | ( n10840 & n10842 ) ;
  assign n10850 = n7762 ^ n5014 ^ n4185 ;
  assign n10844 = n4481 ^ n4217 ^ x106 ;
  assign n10845 = n10844 ^ n4271 ^ 1'b0 ;
  assign n10846 = ~n3309 & n10845 ;
  assign n10847 = n10846 ^ n6304 ^ 1'b0 ;
  assign n10848 = x81 & n10847 ;
  assign n10849 = ( n3690 & n8549 ) | ( n3690 & n10848 ) | ( n8549 & n10848 ) ;
  assign n10851 = n10850 ^ n10849 ^ n5656 ;
  assign n10852 = n10851 ^ n355 ^ 1'b0 ;
  assign n10853 = n2995 & ~n7444 ;
  assign n10854 = ~n7216 & n10853 ;
  assign n10855 = n3782 & n8624 ;
  assign n10856 = ~n937 & n10855 ;
  assign n10857 = ~n8285 & n10856 ;
  assign n10858 = n2889 & ~n8402 ;
  assign n10859 = n1430 & n6540 ;
  assign n10860 = ~n6630 & n10859 ;
  assign n10868 = ~n2791 & n6094 ;
  assign n10869 = n10868 ^ n615 ^ 1'b0 ;
  assign n10870 = ( ~n496 & n2140 ) | ( ~n496 & n10869 ) | ( n2140 & n10869 ) ;
  assign n10861 = n3840 ^ n1522 ^ 1'b0 ;
  assign n10862 = n6281 | n10861 ;
  assign n10863 = ( ~n4779 & n5962 ) | ( ~n4779 & n10862 ) | ( n5962 & n10862 ) ;
  assign n10864 = n5715 & n5988 ;
  assign n10865 = n1663 & n10864 ;
  assign n10866 = n10863 & ~n10865 ;
  assign n10867 = n10866 ^ n5286 ^ n1437 ;
  assign n10871 = n10870 ^ n10867 ^ 1'b0 ;
  assign n10872 = n3647 & n10871 ;
  assign n10873 = n5560 | n6481 ;
  assign n10874 = n2258 ^ n1906 ^ 1'b0 ;
  assign n10875 = n3923 & n10874 ;
  assign n10876 = n10875 ^ n285 ^ 1'b0 ;
  assign n10877 = n7006 | n10876 ;
  assign n10878 = n10877 ^ n984 ^ 1'b0 ;
  assign n10879 = ~n750 & n2994 ;
  assign n10880 = ~n3106 & n10879 ;
  assign n10881 = ( n409 & n5730 ) | ( n409 & ~n7080 ) | ( n5730 & ~n7080 ) ;
  assign n10882 = ~n3227 & n7410 ;
  assign n10883 = n3311 ^ n510 ^ 1'b0 ;
  assign n10884 = n9019 ^ n5149 ^ 1'b0 ;
  assign n10885 = n6308 ^ n879 ^ 1'b0 ;
  assign n10886 = n2456 & ~n3914 ;
  assign n10887 = ~n3062 & n10886 ;
  assign n10888 = n2730 & ~n10887 ;
  assign n10889 = n10264 ^ n6904 ^ 1'b0 ;
  assign n10890 = n10888 | n10889 ;
  assign n10891 = ( n1706 & n8779 ) | ( n1706 & ~n10890 ) | ( n8779 & ~n10890 ) ;
  assign n10892 = ~n4469 & n9661 ;
  assign n10893 = ~n8319 & n10892 ;
  assign n10900 = n7294 ^ n1592 ^ 1'b0 ;
  assign n10898 = ( n382 & ~n2856 ) | ( n382 & n8405 ) | ( ~n2856 & n8405 ) ;
  assign n10894 = n1844 | n1882 ;
  assign n10895 = n10894 ^ n3663 ^ 1'b0 ;
  assign n10896 = n2180 & n10895 ;
  assign n10897 = n5306 & n10896 ;
  assign n10899 = n10898 ^ n10897 ^ 1'b0 ;
  assign n10901 = n10900 ^ n10899 ^ n6254 ;
  assign n10902 = n10901 ^ n1488 ^ 1'b0 ;
  assign n10903 = ~n4591 & n6414 ;
  assign n10904 = n10903 ^ n2909 ^ n618 ;
  assign n10905 = ~n2628 & n2746 ;
  assign n10906 = n5411 & n10905 ;
  assign n10907 = ( n2391 & n10904 ) | ( n2391 & n10906 ) | ( n10904 & n10906 ) ;
  assign n10908 = ( n604 & ~n9065 ) | ( n604 & n10907 ) | ( ~n9065 & n10907 ) ;
  assign n10909 = n8586 ^ n6798 ^ n4105 ;
  assign n10910 = n1359 ^ n1192 ^ n1121 ;
  assign n10911 = n9315 ^ n2550 ^ 1'b0 ;
  assign n10912 = n7993 | n10911 ;
  assign n10913 = n4956 & ~n10912 ;
  assign n10914 = n2725 & n3436 ;
  assign n10915 = n1512 & n10914 ;
  assign n10916 = n10915 ^ n3352 ^ 1'b0 ;
  assign n10917 = n5514 & ~n10916 ;
  assign n10918 = n6283 ^ n5236 ^ 1'b0 ;
  assign n10919 = n10918 ^ n1400 ^ 1'b0 ;
  assign n10920 = n10917 | n10919 ;
  assign n10921 = ( n1735 & n2777 ) | ( n1735 & ~n3699 ) | ( n2777 & ~n3699 ) ;
  assign n10922 = n7444 | n10921 ;
  assign n10923 = n7781 & n10355 ;
  assign n10924 = n10923 ^ n7726 ^ 1'b0 ;
  assign n10925 = n10924 ^ n4409 ^ 1'b0 ;
  assign n10926 = n10000 ^ x162 ^ 1'b0 ;
  assign n10927 = n408 & ~n10926 ;
  assign n10928 = n8768 & n10927 ;
  assign n10929 = n5608 & n10928 ;
  assign n10937 = n1630 ^ n333 ^ 1'b0 ;
  assign n10938 = n2528 & ~n10937 ;
  assign n10939 = ( n4243 & n4471 ) | ( n4243 & n10938 ) | ( n4471 & n10938 ) ;
  assign n10933 = n464 | n693 ;
  assign n10934 = n1818 & ~n10933 ;
  assign n10935 = n10934 ^ n7458 ^ n2220 ;
  assign n10930 = ( x178 & n3341 ) | ( x178 & ~n5424 ) | ( n3341 & ~n5424 ) ;
  assign n10931 = n4329 | n10930 ;
  assign n10932 = n2498 & ~n10931 ;
  assign n10936 = n10935 ^ n10932 ^ n7170 ;
  assign n10940 = n10939 ^ n10936 ^ 1'b0 ;
  assign n10941 = n8864 & ~n10940 ;
  assign n10942 = ~n3459 & n9421 ;
  assign n10945 = ( ~n657 & n7924 ) | ( ~n657 & n9156 ) | ( n7924 & n9156 ) ;
  assign n10946 = n7698 ^ n6835 ^ n5565 ;
  assign n10947 = n10945 & ~n10946 ;
  assign n10948 = n7409 & ~n10947 ;
  assign n10943 = n10220 ^ x192 ^ 1'b0 ;
  assign n10944 = n6164 & ~n10943 ;
  assign n10949 = n10948 ^ n10944 ^ 1'b0 ;
  assign n10950 = n5687 ^ n4388 ^ 1'b0 ;
  assign n10951 = n2508 & n10950 ;
  assign n10952 = n8785 & ~n10951 ;
  assign n10953 = ( n4875 & ~n5008 ) | ( n4875 & n10918 ) | ( ~n5008 & n10918 ) ;
  assign n10954 = n9722 & ~n10953 ;
  assign n10955 = ~n3453 & n6377 ;
  assign n10956 = ( n2393 & n3032 ) | ( n2393 & ~n10955 ) | ( n3032 & ~n10955 ) ;
  assign n10957 = ( n544 & ~n10954 ) | ( n544 & n10956 ) | ( ~n10954 & n10956 ) ;
  assign n10958 = n10957 ^ n6472 ^ 1'b0 ;
  assign n10959 = n3136 | n9379 ;
  assign n10960 = n10959 ^ n8376 ^ 1'b0 ;
  assign n10966 = n6659 ^ n2529 ^ 1'b0 ;
  assign n10961 = n499 & n2968 ;
  assign n10963 = n4445 ^ n3873 ^ 1'b0 ;
  assign n10962 = x202 & n3401 ;
  assign n10964 = n10963 ^ n10962 ^ 1'b0 ;
  assign n10965 = n10961 & ~n10964 ;
  assign n10967 = n10966 ^ n10965 ^ 1'b0 ;
  assign n10968 = n2911 & ~n3385 ;
  assign n10969 = n7973 ^ n7814 ^ 1'b0 ;
  assign n10970 = n8953 & n10969 ;
  assign n10971 = ( ~n10440 & n10968 ) | ( ~n10440 & n10970 ) | ( n10968 & n10970 ) ;
  assign n10972 = ( n1027 & n1265 ) | ( n1027 & n3302 ) | ( n1265 & n3302 ) ;
  assign n10973 = ( n355 & n468 ) | ( n355 & ~n8520 ) | ( n468 & ~n8520 ) ;
  assign n10974 = n3030 & n6375 ;
  assign n10993 = n5823 | n7099 ;
  assign n10991 = n1776 & ~n6118 ;
  assign n10975 = ~n2735 & n6173 ;
  assign n10976 = ~n3381 & n10975 ;
  assign n10984 = ( n3089 & n5310 ) | ( n3089 & n5403 ) | ( n5310 & n5403 ) ;
  assign n10981 = ( n1779 & ~n2319 ) | ( n1779 & n4930 ) | ( ~n2319 & n4930 ) ;
  assign n10982 = ~n2003 & n10981 ;
  assign n10983 = n2163 & n10982 ;
  assign n10985 = n10984 ^ n10983 ^ n10013 ;
  assign n10978 = n2945 ^ n2408 ^ n2154 ;
  assign n10979 = n10978 ^ n5739 ^ n874 ;
  assign n10980 = n5288 & n10979 ;
  assign n10986 = n10985 ^ n10980 ^ 1'b0 ;
  assign n10987 = n10986 ^ n4350 ^ n1304 ;
  assign n10977 = ~n10110 & n10917 ;
  assign n10988 = n10987 ^ n10977 ^ 1'b0 ;
  assign n10989 = n3915 ^ n1574 ^ n929 ;
  assign n10990 = ( n10976 & ~n10988 ) | ( n10976 & n10989 ) | ( ~n10988 & n10989 ) ;
  assign n10992 = n10991 ^ n10990 ^ 1'b0 ;
  assign n10994 = n10993 ^ n10992 ^ n6193 ;
  assign n10995 = n6812 ^ n1926 ^ n894 ;
  assign n10996 = n10995 ^ n2771 ^ 1'b0 ;
  assign n10997 = n4310 ^ n3690 ^ n2135 ;
  assign n10998 = n10997 ^ n10456 ^ n6156 ;
  assign n10999 = ~n10996 & n10998 ;
  assign n11000 = ~n1372 & n10999 ;
  assign n11001 = ~n1608 & n2156 ;
  assign n11002 = n2972 & ~n3099 ;
  assign n11003 = n703 | n11002 ;
  assign n11004 = n10295 ^ n2554 ^ 1'b0 ;
  assign n11005 = n3271 & ~n11004 ;
  assign n11007 = n5449 ^ n394 ^ x168 ;
  assign n11006 = n480 & ~n2952 ;
  assign n11008 = n11007 ^ n11006 ^ n1452 ;
  assign n11009 = ( x248 & n8307 ) | ( x248 & n11008 ) | ( n8307 & n11008 ) ;
  assign n11016 = n2407 & ~n4552 ;
  assign n11015 = n1531 | n6683 ;
  assign n11017 = n11016 ^ n11015 ^ 1'b0 ;
  assign n11018 = ~n4574 & n11017 ;
  assign n11010 = n8872 ^ x97 ^ 1'b0 ;
  assign n11011 = x110 & n11010 ;
  assign n11012 = ~n3632 & n11011 ;
  assign n11013 = n2445 & n11012 ;
  assign n11014 = n10939 & ~n11013 ;
  assign n11019 = n11018 ^ n11014 ^ 1'b0 ;
  assign n11020 = n1468 ^ n584 ^ 1'b0 ;
  assign n11021 = n1440 | n11020 ;
  assign n11022 = ( n4265 & ~n7462 ) | ( n4265 & n11021 ) | ( ~n7462 & n11021 ) ;
  assign n11023 = n2823 & ~n11022 ;
  assign n11024 = n11023 ^ n459 ^ 1'b0 ;
  assign n11025 = n4876 | n11024 ;
  assign n11026 = n11019 | n11025 ;
  assign n11029 = x167 & ~n2738 ;
  assign n11030 = ( n1162 & n7195 ) | ( n1162 & n11029 ) | ( n7195 & n11029 ) ;
  assign n11027 = ( n2397 & ~n3696 ) | ( n2397 & n5737 ) | ( ~n3696 & n5737 ) ;
  assign n11028 = n8692 | n11027 ;
  assign n11031 = n11030 ^ n11028 ^ 1'b0 ;
  assign n11032 = n1813 & ~n7311 ;
  assign n11034 = ( n1258 & n4639 ) | ( n1258 & n8786 ) | ( n4639 & n8786 ) ;
  assign n11033 = n618 | n10850 ;
  assign n11035 = n11034 ^ n11033 ^ n1440 ;
  assign n11036 = n735 & ~n6362 ;
  assign n11037 = ~n1645 & n11036 ;
  assign n11038 = n7965 | n11037 ;
  assign n11039 = n11038 ^ n1260 ^ 1'b0 ;
  assign n11040 = n388 | n1926 ;
  assign n11041 = n11040 ^ n711 ^ 1'b0 ;
  assign n11042 = ( ~n1088 & n2164 ) | ( ~n1088 & n9320 ) | ( n2164 & n9320 ) ;
  assign n11043 = ( n2785 & ~n11041 ) | ( n2785 & n11042 ) | ( ~n11041 & n11042 ) ;
  assign n11044 = ( n4348 & n9172 ) | ( n4348 & n11043 ) | ( n9172 & n11043 ) ;
  assign n11045 = ( n3191 & n5573 ) | ( n3191 & n11044 ) | ( n5573 & n11044 ) ;
  assign n11046 = n2980 & n11045 ;
  assign n11047 = n11039 & n11046 ;
  assign n11048 = n3380 ^ n256 ^ 1'b0 ;
  assign n11049 = n11048 ^ n10317 ^ n2780 ;
  assign n11050 = ( n2016 & n3931 ) | ( n2016 & ~n11049 ) | ( n3931 & ~n11049 ) ;
  assign n11051 = n4977 ^ n4662 ^ n2994 ;
  assign n11055 = ( ~n295 & n1522 ) | ( ~n295 & n2670 ) | ( n1522 & n2670 ) ;
  assign n11056 = n6464 & n11055 ;
  assign n11057 = n11056 ^ n2844 ^ 1'b0 ;
  assign n11058 = n11057 ^ n9447 ^ 1'b0 ;
  assign n11052 = n5059 ^ n2050 ^ 1'b0 ;
  assign n11053 = n11052 ^ n5476 ^ n2946 ;
  assign n11054 = n10849 & n11053 ;
  assign n11059 = n11058 ^ n11054 ^ 1'b0 ;
  assign n11060 = n10723 ^ n4705 ^ 1'b0 ;
  assign n11061 = ~n6955 & n11060 ;
  assign n11062 = n2481 & n9438 ;
  assign n11063 = n1826 | n8735 ;
  assign n11064 = n6699 | n11063 ;
  assign n11065 = n2408 & n3429 ;
  assign n11066 = n11065 ^ n396 ^ 1'b0 ;
  assign n11067 = n11066 ^ n7544 ^ n3338 ;
  assign n11068 = n10626 | n11067 ;
  assign n11069 = n5724 ^ n4150 ^ n3254 ;
  assign n11070 = n7802 ^ n4194 ^ 1'b0 ;
  assign n11071 = n3844 | n10356 ;
  assign n11072 = n6707 & n11071 ;
  assign n11073 = x105 & n1338 ;
  assign n11074 = n11073 ^ n1134 ^ 1'b0 ;
  assign n11075 = n11074 ^ n7704 ^ n6169 ;
  assign n11076 = n8354 & n11075 ;
  assign n11077 = ~n10369 & n11076 ;
  assign n11078 = ( ~n3039 & n4882 ) | ( ~n3039 & n5454 ) | ( n4882 & n5454 ) ;
  assign n11079 = n11077 & n11078 ;
  assign n11080 = n11079 ^ n5755 ^ 1'b0 ;
  assign n11081 = n2538 & n11080 ;
  assign n11082 = n810 | n5216 ;
  assign n11083 = n11082 ^ n7599 ^ n5464 ;
  assign n11084 = ( x15 & ~n3000 ) | ( x15 & n5097 ) | ( ~n3000 & n5097 ) ;
  assign n11085 = n5136 & ~n11084 ;
  assign n11086 = n11085 ^ n1542 ^ 1'b0 ;
  assign n11087 = ( n1049 & ~n3946 ) | ( n1049 & n8374 ) | ( ~n3946 & n8374 ) ;
  assign n11088 = ( ~n1912 & n3475 ) | ( ~n1912 & n5295 ) | ( n3475 & n5295 ) ;
  assign n11089 = n11088 ^ n9629 ^ n5126 ;
  assign n11090 = n11089 ^ n7802 ^ 1'b0 ;
  assign n11091 = ( n2694 & n11087 ) | ( n2694 & ~n11090 ) | ( n11087 & ~n11090 ) ;
  assign n11092 = ( n11050 & n11086 ) | ( n11050 & n11091 ) | ( n11086 & n11091 ) ;
  assign n11094 = n7403 & n7892 ;
  assign n11095 = n1737 & n11094 ;
  assign n11093 = n284 & n5356 ;
  assign n11096 = n11095 ^ n11093 ^ n2161 ;
  assign n11097 = n5295 ^ n3655 ^ 1'b0 ;
  assign n11098 = n1269 & ~n11097 ;
  assign n11099 = n1796 & n11098 ;
  assign n11100 = ( n5310 & n10686 ) | ( n5310 & ~n11099 ) | ( n10686 & ~n11099 ) ;
  assign n11101 = n10200 ^ n303 ^ 1'b0 ;
  assign n11102 = n2761 | n11101 ;
  assign n11105 = n2970 ^ n2470 ^ 1'b0 ;
  assign n11106 = n2571 & ~n11105 ;
  assign n11107 = ( ~n2419 & n3033 ) | ( ~n2419 & n11106 ) | ( n3033 & n11106 ) ;
  assign n11103 = ( ~n1654 & n5753 ) | ( ~n1654 & n10855 ) | ( n5753 & n10855 ) ;
  assign n11104 = n11103 ^ n6063 ^ n3719 ;
  assign n11108 = n11107 ^ n11104 ^ n5062 ;
  assign n11109 = ( n1978 & n5065 ) | ( n1978 & ~n9148 ) | ( n5065 & ~n9148 ) ;
  assign n11110 = n3482 | n4480 ;
  assign n11111 = n11110 ^ n4129 ^ 1'b0 ;
  assign n11112 = n11111 ^ n11037 ^ n9465 ;
  assign n11113 = n1830 & n2719 ;
  assign n11114 = n11113 ^ n1757 ^ 1'b0 ;
  assign n11115 = n11112 & ~n11114 ;
  assign n11116 = ( ~x244 & n11109 ) | ( ~x244 & n11115 ) | ( n11109 & n11115 ) ;
  assign n11121 = n2571 ^ n303 ^ x239 ;
  assign n11120 = n5492 ^ n1522 ^ n506 ;
  assign n11122 = n11121 ^ n11120 ^ n10691 ;
  assign n11123 = n11122 ^ n6701 ^ 1'b0 ;
  assign n11124 = n6055 | n11123 ;
  assign n11117 = n4112 & n4322 ;
  assign n11118 = n11117 ^ n7094 ^ 1'b0 ;
  assign n11119 = n11118 ^ n6495 ^ n647 ;
  assign n11125 = n11124 ^ n11119 ^ 1'b0 ;
  assign n11126 = n3492 | n11125 ;
  assign n11134 = n10178 ^ n7154 ^ n3316 ;
  assign n11127 = n7102 ^ x98 ^ 1'b0 ;
  assign n11129 = n7897 ^ n3279 ^ 1'b0 ;
  assign n11128 = n4005 & n6886 ;
  assign n11130 = n11129 ^ n11128 ^ 1'b0 ;
  assign n11131 = ~n2718 & n11130 ;
  assign n11132 = ( n7782 & ~n7821 ) | ( n7782 & n11131 ) | ( ~n7821 & n11131 ) ;
  assign n11133 = n11127 | n11132 ;
  assign n11135 = n11134 ^ n11133 ^ 1'b0 ;
  assign n11136 = ( ~n4459 & n4556 ) | ( ~n4459 & n5449 ) | ( n4556 & n5449 ) ;
  assign n11137 = ~n448 & n11136 ;
  assign n11138 = n11137 ^ n8960 ^ 1'b0 ;
  assign n11139 = n5843 ^ n5122 ^ n2263 ;
  assign n11140 = n2967 ^ n1969 ^ 1'b0 ;
  assign n11141 = ( ~n5234 & n6500 ) | ( ~n5234 & n11140 ) | ( n6500 & n11140 ) ;
  assign n11142 = n10769 ^ n7642 ^ 1'b0 ;
  assign n11143 = ~n11141 & n11142 ;
  assign n11144 = n11143 ^ n2041 ^ 1'b0 ;
  assign n11148 = n3432 & ~n7449 ;
  assign n11145 = ~n2306 & n7972 ;
  assign n11146 = n1624 & n11145 ;
  assign n11147 = n11146 ^ n9208 ^ 1'b0 ;
  assign n11149 = n11148 ^ n11147 ^ n2081 ;
  assign n11150 = ~n1647 & n10284 ;
  assign n11151 = ( n7143 & n9147 ) | ( n7143 & n11150 ) | ( n9147 & n11150 ) ;
  assign n11154 = n1977 ^ n1595 ^ 1'b0 ;
  assign n11155 = ~n2788 & n11154 ;
  assign n11156 = ( n3556 & ~n10655 ) | ( n3556 & n11155 ) | ( ~n10655 & n11155 ) ;
  assign n11157 = n11156 ^ n1933 ^ n1911 ;
  assign n11152 = n4949 ^ n1680 ^ 1'b0 ;
  assign n11153 = n6285 | n11152 ;
  assign n11158 = n11157 ^ n11153 ^ 1'b0 ;
  assign n11159 = ( n1173 & n3585 ) | ( n1173 & n8548 ) | ( n3585 & n8548 ) ;
  assign n11160 = n1154 | n4341 ;
  assign n11161 = n11160 ^ n2527 ^ 1'b0 ;
  assign n11162 = n7922 & ~n11161 ;
  assign n11163 = n1682 & n4984 ;
  assign n11164 = ~n1866 & n11163 ;
  assign n11165 = n11164 ^ n9655 ^ 1'b0 ;
  assign n11166 = n11165 ^ n6511 ^ n999 ;
  assign n11167 = n5252 & n11166 ;
  assign n11168 = n3817 & n11167 ;
  assign n11169 = ~n5336 & n11168 ;
  assign n11170 = n7014 ^ n2035 ^ 1'b0 ;
  assign n11171 = n5560 & n11170 ;
  assign n11172 = n3928 ^ n3216 ^ 1'b0 ;
  assign n11173 = n11171 & ~n11172 ;
  assign n11174 = n11173 ^ n6246 ^ 1'b0 ;
  assign n11175 = n416 & n3645 ;
  assign n11176 = n5503 & n7518 ;
  assign n11177 = n11176 ^ n6021 ^ 1'b0 ;
  assign n11178 = n6064 & ~n11177 ;
  assign n11179 = ( n8851 & n11175 ) | ( n8851 & ~n11178 ) | ( n11175 & ~n11178 ) ;
  assign n11180 = n11179 ^ n3527 ^ 1'b0 ;
  assign n11181 = ~n5322 & n11180 ;
  assign n11182 = n1933 | n6307 ;
  assign n11183 = n11182 ^ n4077 ^ 1'b0 ;
  assign n11184 = n1173 & ~n2985 ;
  assign n11185 = n532 & n11184 ;
  assign n11186 = n11185 ^ n6921 ^ 1'b0 ;
  assign n11187 = ( n438 & n4025 ) | ( n438 & n11186 ) | ( n4025 & n11186 ) ;
  assign n11188 = n827 ^ x46 ^ 1'b0 ;
  assign n11189 = n6956 ^ n4244 ^ 1'b0 ;
  assign n11190 = ~n11188 & n11189 ;
  assign n11191 = n4646 ^ n2867 ^ 1'b0 ;
  assign n11192 = ( ~x230 & n2169 ) | ( ~x230 & n8370 ) | ( n2169 & n8370 ) ;
  assign n11193 = n11192 ^ n8188 ^ n3664 ;
  assign n11194 = ( n3821 & n11191 ) | ( n3821 & n11193 ) | ( n11191 & n11193 ) ;
  assign n11195 = n3100 | n4125 ;
  assign n11196 = n2388 & ~n11195 ;
  assign n11197 = ( n4845 & ~n8030 ) | ( n4845 & n11196 ) | ( ~n8030 & n11196 ) ;
  assign n11198 = ~n1717 & n8789 ;
  assign n11199 = n6897 & n11198 ;
  assign n11200 = n11199 ^ n10073 ^ 1'b0 ;
  assign n11201 = n4597 & ~n11200 ;
  assign n11202 = n11201 ^ n4040 ^ 1'b0 ;
  assign n11203 = n11197 & ~n11202 ;
  assign n11204 = n11194 & n11203 ;
  assign n11205 = n2217 ^ n2125 ^ n1074 ;
  assign n11206 = ( n6179 & n9313 ) | ( n6179 & ~n11205 ) | ( n9313 & ~n11205 ) ;
  assign n11207 = n2195 & n5507 ;
  assign n11208 = n950 & n2747 ;
  assign n11209 = ( n3601 & n5919 ) | ( n3601 & n11208 ) | ( n5919 & n11208 ) ;
  assign n11210 = n1324 & ~n4466 ;
  assign n11211 = ~n11209 & n11210 ;
  assign n11212 = n779 ^ x55 ^ 1'b0 ;
  assign n11213 = n11212 ^ n6382 ^ 1'b0 ;
  assign n11214 = n3337 & ~n5959 ;
  assign n11215 = ~n11213 & n11214 ;
  assign n11216 = n1016 & ~n11215 ;
  assign n11217 = ( n4479 & n5557 ) | ( n4479 & ~n7440 ) | ( n5557 & ~n7440 ) ;
  assign n11218 = n6640 ^ n2234 ^ 1'b0 ;
  assign n11219 = n3974 & n11218 ;
  assign n11220 = n3237 & ~n4471 ;
  assign n11221 = n11220 ^ n9450 ^ 1'b0 ;
  assign n11222 = n5492 ^ n5362 ^ n2029 ;
  assign n11223 = n11222 ^ n8880 ^ n3614 ;
  assign n11224 = ( n276 & n1214 ) | ( n276 & n1501 ) | ( n1214 & n1501 ) ;
  assign n11225 = n11224 ^ n3037 ^ n1580 ;
  assign n11226 = ( n7038 & n7698 ) | ( n7038 & ~n11225 ) | ( n7698 & ~n11225 ) ;
  assign n11227 = ~x225 & n2332 ;
  assign n11228 = n11227 ^ n1148 ^ 1'b0 ;
  assign n11229 = n2238 & n11228 ;
  assign n11230 = n11229 ^ n1405 ^ 1'b0 ;
  assign n11231 = n6279 ^ n4110 ^ n1798 ;
  assign n11232 = ~n6101 & n11231 ;
  assign n11233 = n11232 ^ n10056 ^ 1'b0 ;
  assign n11243 = n731 & n1963 ;
  assign n11244 = ~n1449 & n11243 ;
  assign n11241 = n9275 ^ n6275 ^ n2400 ;
  assign n11242 = ( ~n2270 & n4053 ) | ( ~n2270 & n11241 ) | ( n4053 & n11241 ) ;
  assign n11234 = n10468 ^ n8926 ^ 1'b0 ;
  assign n11235 = n3091 ^ n1277 ^ 1'b0 ;
  assign n11236 = ~n2014 & n11235 ;
  assign n11237 = n11236 ^ n5231 ^ 1'b0 ;
  assign n11238 = n11237 ^ n5038 ^ 1'b0 ;
  assign n11239 = ~n11234 & n11238 ;
  assign n11240 = ( n1705 & n4066 ) | ( n1705 & ~n11239 ) | ( n4066 & ~n11239 ) ;
  assign n11245 = n11244 ^ n11242 ^ n11240 ;
  assign n11246 = n2935 ^ n2530 ^ 1'b0 ;
  assign n11247 = n6146 ^ n4689 ^ 1'b0 ;
  assign n11248 = ( n2451 & n8618 ) | ( n2451 & n11247 ) | ( n8618 & n11247 ) ;
  assign n11249 = n11246 & ~n11248 ;
  assign n11250 = ( ~n3693 & n4636 ) | ( ~n3693 & n10007 ) | ( n4636 & n10007 ) ;
  assign n11253 = n841 & ~n8429 ;
  assign n11254 = n2227 & ~n11253 ;
  assign n11255 = n11254 ^ n11225 ^ 1'b0 ;
  assign n11256 = n4028 | n11255 ;
  assign n11257 = n11256 ^ n7770 ^ 1'b0 ;
  assign n11251 = x183 & ~n3715 ;
  assign n11252 = ( ~n3106 & n8128 ) | ( ~n3106 & n11251 ) | ( n8128 & n11251 ) ;
  assign n11258 = n11257 ^ n11252 ^ n9794 ;
  assign n11259 = n10754 ^ n3375 ^ 1'b0 ;
  assign n11260 = n7824 | n11259 ;
  assign n11261 = n8606 ^ n5880 ^ n3424 ;
  assign n11262 = n9009 ^ n5476 ^ n893 ;
  assign n11263 = n1877 & n11262 ;
  assign n11264 = n3100 & ~n8537 ;
  assign n11265 = n374 & n8478 ;
  assign n11266 = n11265 ^ n2634 ^ 1'b0 ;
  assign n11267 = ( ~n10029 & n11264 ) | ( ~n10029 & n11266 ) | ( n11264 & n11266 ) ;
  assign n11268 = n3991 ^ n2781 ^ 1'b0 ;
  assign n11269 = n4714 | n11268 ;
  assign n11270 = n6617 ^ n2931 ^ n1930 ;
  assign n11271 = n11270 ^ n2523 ^ 1'b0 ;
  assign n11272 = n1956 ^ n1342 ^ 1'b0 ;
  assign n11274 = x88 & n9581 ;
  assign n11275 = n11274 ^ n4049 ^ 1'b0 ;
  assign n11273 = ( n374 & ~n8992 ) | ( n374 & n9083 ) | ( ~n8992 & n9083 ) ;
  assign n11276 = n11275 ^ n11273 ^ n10986 ;
  assign n11277 = ~n8251 & n11276 ;
  assign n11278 = ( n2924 & ~n3543 ) | ( n2924 & n9030 ) | ( ~n3543 & n9030 ) ;
  assign n11279 = ( x229 & n1348 ) | ( x229 & ~n8911 ) | ( n1348 & ~n8911 ) ;
  assign n11280 = ~n11278 & n11279 ;
  assign n11281 = n9429 ^ n6764 ^ n1072 ;
  assign n11282 = n11281 ^ n5060 ^ 1'b0 ;
  assign n11283 = n2501 | n11282 ;
  assign n11284 = n8502 ^ x82 ^ 1'b0 ;
  assign n11285 = n5129 & ~n7415 ;
  assign n11286 = ( ~n3235 & n7022 ) | ( ~n3235 & n11285 ) | ( n7022 & n11285 ) ;
  assign n11287 = n376 & ~n11286 ;
  assign n11288 = ( x231 & n4951 ) | ( x231 & ~n9242 ) | ( n4951 & ~n9242 ) ;
  assign n11289 = ~n1039 & n5005 ;
  assign n11290 = n11289 ^ n2056 ^ 1'b0 ;
  assign n11291 = ( n297 & n572 ) | ( n297 & n1083 ) | ( n572 & n1083 ) ;
  assign n11292 = ~n3856 & n11291 ;
  assign n11293 = n10924 ^ n5468 ^ n4914 ;
  assign n11295 = ( n650 & n1658 ) | ( n650 & n2669 ) | ( n1658 & n2669 ) ;
  assign n11296 = n11295 ^ n7301 ^ n2564 ;
  assign n11297 = n3026 & ~n9721 ;
  assign n11298 = n11296 & n11297 ;
  assign n11294 = n11113 ^ n2868 ^ n1690 ;
  assign n11299 = n11298 ^ n11294 ^ n4240 ;
  assign n11306 = n1154 | n2682 ;
  assign n11307 = n11306 ^ n2595 ^ n2522 ;
  assign n11308 = n3805 & ~n11307 ;
  assign n11309 = n11308 ^ n2026 ^ 1'b0 ;
  assign n11300 = n898 ^ n428 ^ x65 ;
  assign n11301 = n11300 ^ n3272 ^ n336 ;
  assign n11302 = n1330 ^ n1283 ^ 1'b0 ;
  assign n11303 = ( ~n2415 & n11301 ) | ( ~n2415 & n11302 ) | ( n11301 & n11302 ) ;
  assign n11304 = x129 | n11303 ;
  assign n11305 = n11041 & n11304 ;
  assign n11310 = n11309 ^ n11305 ^ 1'b0 ;
  assign n11311 = n2767 | n3862 ;
  assign n11312 = n11311 ^ n3360 ^ 1'b0 ;
  assign n11313 = n5189 & ~n11247 ;
  assign n11314 = n1134 & ~n9717 ;
  assign n11315 = n11314 ^ n3966 ^ 1'b0 ;
  assign n11317 = n1753 | n2038 ;
  assign n11318 = n11317 ^ n5116 ^ 1'b0 ;
  assign n11316 = n3839 & ~n4010 ;
  assign n11319 = n11318 ^ n11316 ^ 1'b0 ;
  assign n11320 = ~n1473 & n1675 ;
  assign n11321 = n3197 & n11320 ;
  assign n11322 = n11321 ^ n5453 ^ 1'b0 ;
  assign n11323 = n11319 & n11322 ;
  assign n11324 = ( ~n1403 & n3619 ) | ( ~n1403 & n7947 ) | ( n3619 & n7947 ) ;
  assign n11325 = n709 & n11324 ;
  assign n11326 = n341 | n11325 ;
  assign n11327 = ~n4516 & n4644 ;
  assign n11328 = n9446 ^ n9341 ^ n2049 ;
  assign n11329 = n11327 & ~n11328 ;
  assign n11330 = ~n5666 & n11329 ;
  assign n11333 = n2391 ^ n637 ^ 1'b0 ;
  assign n11334 = n3021 | n11333 ;
  assign n11331 = ~n6296 & n7614 ;
  assign n11332 = n11331 ^ n5233 ^ 1'b0 ;
  assign n11335 = n11334 ^ n11332 ^ 1'b0 ;
  assign n11336 = n11335 ^ n1050 ^ 1'b0 ;
  assign n11337 = ( n2039 & n10057 ) | ( n2039 & n11336 ) | ( n10057 & n11336 ) ;
  assign n11338 = n11330 | n11337 ;
  assign n11339 = n1067 | n11338 ;
  assign n11340 = ( x161 & ~n699 ) | ( x161 & n1839 ) | ( ~n699 & n1839 ) ;
  assign n11341 = n10251 & ~n11340 ;
  assign n11342 = n3104 & ~n7377 ;
  assign n11343 = ~n10083 & n11342 ;
  assign n11344 = n9246 ^ n3943 ^ 1'b0 ;
  assign n11345 = ~n7870 & n11344 ;
  assign n11346 = n11345 ^ n9564 ^ 1'b0 ;
  assign n11347 = n7291 & ~n11346 ;
  assign n11348 = ( n334 & ~n2782 ) | ( n334 & n2836 ) | ( ~n2782 & n2836 ) ;
  assign n11358 = x102 & ~n3787 ;
  assign n11359 = n11358 ^ n2101 ^ 1'b0 ;
  assign n11354 = n7928 ^ n7070 ^ 1'b0 ;
  assign n11355 = n4081 & ~n11354 ;
  assign n11356 = n4173 & n11355 ;
  assign n11351 = n1683 & ~n4107 ;
  assign n11352 = n2082 & n11351 ;
  assign n11353 = ( ~n2273 & n4131 ) | ( ~n2273 & n11352 ) | ( n4131 & n11352 ) ;
  assign n11349 = ~n393 & n11222 ;
  assign n11350 = n11349 ^ n5664 ^ n1384 ;
  assign n11357 = n11356 ^ n11353 ^ n11350 ;
  assign n11360 = n11359 ^ n11357 ^ n1408 ;
  assign n11365 = n10456 ^ n7067 ^ n1158 ;
  assign n11362 = n3170 ^ n1816 ^ 1'b0 ;
  assign n11363 = n869 | n11362 ;
  assign n11361 = ~n259 & n6053 ;
  assign n11364 = n11363 ^ n11361 ^ 1'b0 ;
  assign n11366 = n11365 ^ n11364 ^ n2169 ;
  assign n11369 = ~n883 & n1255 ;
  assign n11370 = n11369 ^ n1776 ^ 1'b0 ;
  assign n11368 = n7070 ^ n6938 ^ n4242 ;
  assign n11367 = n9512 ^ n1429 ^ 1'b0 ;
  assign n11371 = n11370 ^ n11368 ^ n11367 ;
  assign n11378 = n314 | n6083 ;
  assign n11372 = n9695 ^ n963 ^ 1'b0 ;
  assign n11373 = n1028 | n11372 ;
  assign n11374 = ( ~n1513 & n6963 ) | ( ~n1513 & n11373 ) | ( n6963 & n11373 ) ;
  assign n11375 = n1683 & ~n6840 ;
  assign n11376 = n11375 ^ n2474 ^ 1'b0 ;
  assign n11377 = n11374 & n11376 ;
  assign n11379 = n11378 ^ n11377 ^ 1'b0 ;
  assign n11380 = n2845 & n7888 ;
  assign n11381 = n11380 ^ n4634 ^ 1'b0 ;
  assign n11382 = ( n4139 & n5547 ) | ( n4139 & ~n11381 ) | ( n5547 & ~n11381 ) ;
  assign n11383 = n8015 & n9632 ;
  assign n11384 = n2846 & n5945 ;
  assign n11385 = ( n6690 & n9721 ) | ( n6690 & n11384 ) | ( n9721 & n11384 ) ;
  assign n11386 = n9001 ^ n8385 ^ n1483 ;
  assign n11387 = n4112 ^ n3281 ^ 1'b0 ;
  assign n11388 = ~n2934 & n8429 ;
  assign n11389 = n11388 ^ n4591 ^ 1'b0 ;
  assign n11390 = ( ~n5310 & n11387 ) | ( ~n5310 & n11389 ) | ( n11387 & n11389 ) ;
  assign n11391 = n11390 ^ n10774 ^ 1'b0 ;
  assign n11392 = ( n3175 & n7492 ) | ( n3175 & ~n11391 ) | ( n7492 & ~n11391 ) ;
  assign n11393 = n10997 ^ n6625 ^ 1'b0 ;
  assign n11394 = n7201 & n11393 ;
  assign n11395 = n5523 & ~n7926 ;
  assign n11396 = ~n11364 & n11395 ;
  assign n11397 = n6989 ^ n5315 ^ 1'b0 ;
  assign n11398 = ~n11396 & n11397 ;
  assign n11399 = ~n3565 & n6497 ;
  assign n11400 = n11399 ^ n5162 ^ 1'b0 ;
  assign n11401 = n11400 ^ n8039 ^ 1'b0 ;
  assign n11402 = n773 ^ n574 ^ 1'b0 ;
  assign n11403 = n11266 | n11402 ;
  assign n11404 = n9524 & ~n11403 ;
  assign n11405 = n11404 ^ n5063 ^ 1'b0 ;
  assign n11406 = n8396 ^ n6196 ^ 1'b0 ;
  assign n11407 = n11405 | n11406 ;
  assign n11411 = ( n1289 & n2662 ) | ( n1289 & ~n5402 ) | ( n2662 & ~n5402 ) ;
  assign n11412 = n6531 ^ n1813 ^ 1'b0 ;
  assign n11413 = ( n2443 & ~n6070 ) | ( n2443 & n11412 ) | ( ~n6070 & n11412 ) ;
  assign n11414 = n11413 ^ n9174 ^ n3415 ;
  assign n11415 = n11414 ^ n9509 ^ 1'b0 ;
  assign n11416 = n11411 & n11415 ;
  assign n11408 = n8591 ^ n7538 ^ n6150 ;
  assign n11409 = n1372 | n9151 ;
  assign n11410 = n11408 & n11409 ;
  assign n11417 = n11416 ^ n11410 ^ 1'b0 ;
  assign n11418 = n4054 ^ n1229 ^ 1'b0 ;
  assign n11419 = n285 | n9098 ;
  assign n11420 = ( ~n2576 & n2802 ) | ( ~n2576 & n3839 ) | ( n2802 & n3839 ) ;
  assign n11421 = ~n3946 & n5153 ;
  assign n11422 = n4242 & n11421 ;
  assign n11423 = n11420 | n11422 ;
  assign n11424 = n11419 | n11423 ;
  assign n11425 = ~n5160 & n10673 ;
  assign n11426 = ~n995 & n11425 ;
  assign n11427 = n5962 ^ n4486 ^ x56 ;
  assign n11428 = n11427 ^ n3966 ^ n1284 ;
  assign n11429 = n8237 | n11428 ;
  assign n11430 = n581 | n11429 ;
  assign n11431 = n11430 ^ n8965 ^ 1'b0 ;
  assign n11432 = n9389 | n11431 ;
  assign n11433 = n1156 | n11432 ;
  assign n11434 = n11121 ^ n8374 ^ n1682 ;
  assign n11435 = n11434 ^ n7573 ^ 1'b0 ;
  assign n11436 = ~n10214 & n11080 ;
  assign n11437 = n11436 ^ n294 ^ 1'b0 ;
  assign n11438 = ~n1268 & n4465 ;
  assign n11439 = n11438 ^ n9107 ^ n785 ;
  assign n11440 = n9012 & n11439 ;
  assign n11441 = n9965 ^ n3943 ^ 1'b0 ;
  assign n11442 = n4141 ^ n2263 ^ 1'b0 ;
  assign n11443 = x97 & ~n11442 ;
  assign n11444 = ~n7744 & n11443 ;
  assign n11445 = ~n733 & n11444 ;
  assign n11446 = n3897 | n11445 ;
  assign n11447 = n1603 | n11446 ;
  assign n11448 = n11447 ^ n10736 ^ n6382 ;
  assign n11449 = n9405 ^ n7310 ^ 1'b0 ;
  assign n11456 = n6475 & ~n8573 ;
  assign n11457 = ~n7161 & n11456 ;
  assign n11450 = n3873 ^ x175 ^ 1'b0 ;
  assign n11451 = n652 & n11450 ;
  assign n11452 = n2518 | n3932 ;
  assign n11453 = n11451 | n11452 ;
  assign n11454 = n829 & ~n1269 ;
  assign n11455 = n11453 & ~n11454 ;
  assign n11458 = n11457 ^ n11455 ^ 1'b0 ;
  assign n11459 = ~n2903 & n4089 ;
  assign n11460 = n11459 ^ n1317 ^ n264 ;
  assign n11461 = n9852 | n11460 ;
  assign n11462 = ~n6269 & n8814 ;
  assign n11463 = n2699 & ~n7272 ;
  assign n11464 = n11463 ^ n2056 ^ 1'b0 ;
  assign n11465 = n9799 & n11464 ;
  assign n11466 = ~n2758 & n11465 ;
  assign n11467 = n475 | n9589 ;
  assign n11468 = ( ~n6895 & n7126 ) | ( ~n6895 & n11467 ) | ( n7126 & n11467 ) ;
  assign n11473 = n1712 & ~n2716 ;
  assign n11474 = n11473 ^ n11467 ^ 1'b0 ;
  assign n11469 = n10130 ^ n5584 ^ 1'b0 ;
  assign n11470 = n1196 | n5397 ;
  assign n11471 = ~n7490 & n11470 ;
  assign n11472 = ~n11469 & n11471 ;
  assign n11475 = n11474 ^ n11472 ^ n8953 ;
  assign n11476 = ( n1176 & n7741 ) | ( n1176 & ~n8810 ) | ( n7741 & ~n8810 ) ;
  assign n11477 = ~n1410 & n11476 ;
  assign n11478 = n11477 ^ n6660 ^ 1'b0 ;
  assign n11479 = n2600 & ~n11478 ;
  assign n11480 = ( n1581 & ~n1667 ) | ( n1581 & n4934 ) | ( ~n1667 & n4934 ) ;
  assign n11482 = n3335 | n3465 ;
  assign n11481 = n7671 ^ n5370 ^ n3101 ;
  assign n11483 = n11482 ^ n11481 ^ n2445 ;
  assign n11484 = ( n1066 & n11480 ) | ( n1066 & n11483 ) | ( n11480 & n11483 ) ;
  assign n11485 = n9380 ^ n4574 ^ 1'b0 ;
  assign n11486 = n4989 | n11485 ;
  assign n11487 = n7926 ^ n1521 ^ 1'b0 ;
  assign n11488 = n11487 ^ n1315 ^ n946 ;
  assign n11489 = n11488 ^ n8198 ^ 1'b0 ;
  assign n11490 = n3289 ^ n1566 ^ n1204 ;
  assign n11491 = n5352 ^ n4116 ^ 1'b0 ;
  assign n11492 = x208 & n11491 ;
  assign n11493 = ( ~n3903 & n4153 ) | ( ~n3903 & n11492 ) | ( n4153 & n11492 ) ;
  assign n11494 = ( n1252 & n11490 ) | ( n1252 & ~n11493 ) | ( n11490 & ~n11493 ) ;
  assign n11495 = n11494 ^ n9936 ^ n5357 ;
  assign n11496 = ~n9327 & n11495 ;
  assign n11497 = n5393 ^ n652 ^ 1'b0 ;
  assign n11498 = n1627 | n11497 ;
  assign n11499 = n6288 ^ n5043 ^ 1'b0 ;
  assign n11500 = n9432 | n11499 ;
  assign n11501 = ~n5424 & n8209 ;
  assign n11502 = n4977 | n11501 ;
  assign n11503 = n526 & ~n1444 ;
  assign n11504 = ( ~n4856 & n6196 ) | ( ~n4856 & n8122 ) | ( n6196 & n8122 ) ;
  assign n11505 = ( n2486 & ~n11503 ) | ( n2486 & n11504 ) | ( ~n11503 & n11504 ) ;
  assign n11506 = n10806 ^ n7318 ^ n1739 ;
  assign n11507 = n5416 ^ n3854 ^ 1'b0 ;
  assign n11508 = n11507 ^ n4929 ^ n1397 ;
  assign n11509 = n6589 ^ n4878 ^ 1'b0 ;
  assign n11510 = n11508 & n11509 ;
  assign n11511 = ~n607 & n4224 ;
  assign n11512 = n11511 ^ n3363 ^ 1'b0 ;
  assign n11513 = n11512 ^ n10228 ^ n3238 ;
  assign n11514 = n7632 & n11513 ;
  assign n11515 = n579 & n11514 ;
  assign n11516 = n7634 ^ n2042 ^ 1'b0 ;
  assign n11517 = ~n6323 & n11516 ;
  assign n11518 = n11517 ^ n7628 ^ n6534 ;
  assign n11519 = n5427 & ~n6887 ;
  assign n11521 = n1384 ^ n545 ^ 1'b0 ;
  assign n11522 = n9363 & ~n11521 ;
  assign n11523 = n11522 ^ n990 ^ 1'b0 ;
  assign n11520 = ~n5863 & n7377 ;
  assign n11524 = n11523 ^ n11520 ^ 1'b0 ;
  assign n11525 = ( n7048 & n11519 ) | ( n7048 & n11524 ) | ( n11519 & n11524 ) ;
  assign n11526 = n4727 & n9351 ;
  assign n11527 = n1033 & n11526 ;
  assign n11528 = n11527 ^ n7929 ^ 1'b0 ;
  assign n11531 = n2905 ^ n2488 ^ 1'b0 ;
  assign n11532 = n851 & ~n11531 ;
  assign n11529 = n6632 ^ n5059 ^ 1'b0 ;
  assign n11530 = n8835 & n11529 ;
  assign n11533 = n11532 ^ n11530 ^ n3561 ;
  assign n11536 = n4319 ^ n476 ^ 1'b0 ;
  assign n11534 = n7651 ^ n5228 ^ 1'b0 ;
  assign n11535 = ~n4008 & n11534 ;
  assign n11537 = n11536 ^ n11535 ^ 1'b0 ;
  assign n11538 = n8823 & n9026 ;
  assign n11539 = n7930 & n11538 ;
  assign n11540 = n1840 ^ n301 ^ 1'b0 ;
  assign n11541 = n11539 | n11540 ;
  assign n11543 = n6213 ^ n3830 ^ 1'b0 ;
  assign n11542 = n4986 | n7815 ;
  assign n11544 = n11543 ^ n11542 ^ n1874 ;
  assign n11545 = n9910 ^ n9219 ^ n496 ;
  assign n11546 = ( ~n747 & n2538 ) | ( ~n747 & n11545 ) | ( n2538 & n11545 ) ;
  assign n11547 = n10288 ^ n544 ^ 1'b0 ;
  assign n11548 = n11546 & ~n11547 ;
  assign n11549 = n8876 ^ n7757 ^ n6560 ;
  assign n11550 = n11549 ^ n4889 ^ x155 ;
  assign n11551 = n11550 ^ n2966 ^ 1'b0 ;
  assign n11552 = n8015 & n11551 ;
  assign n11553 = ~n8409 & n11552 ;
  assign n11554 = n8628 ^ n4072 ^ 1'b0 ;
  assign n11555 = n1054 & ~n8127 ;
  assign n11556 = n2333 & n11555 ;
  assign n11557 = n11556 ^ n2479 ^ n1031 ;
  assign n11558 = ~n3496 & n9268 ;
  assign n11559 = n11558 ^ n3430 ^ 1'b0 ;
  assign n11560 = ( ~n3763 & n7935 ) | ( ~n3763 & n11559 ) | ( n7935 & n11559 ) ;
  assign n11561 = n11560 ^ n6290 ^ 1'b0 ;
  assign n11564 = n3711 ^ n2143 ^ n1961 ;
  assign n11562 = n6023 | n7102 ;
  assign n11563 = n3954 & ~n11562 ;
  assign n11565 = n11564 ^ n11563 ^ n4862 ;
  assign n11566 = ( ~n677 & n1643 ) | ( ~n677 & n3868 ) | ( n1643 & n3868 ) ;
  assign n11567 = n11566 ^ n8518 ^ 1'b0 ;
  assign n11568 = n8413 | n11567 ;
  assign n11569 = n266 & n6441 ;
  assign n11570 = n11569 ^ n881 ^ 1'b0 ;
  assign n11571 = n11570 ^ n11190 ^ 1'b0 ;
  assign n11572 = n8893 ^ n3984 ^ 1'b0 ;
  assign n11573 = x181 & n2284 ;
  assign n11574 = n11573 ^ n4912 ^ 1'b0 ;
  assign n11575 = n11574 ^ n7774 ^ n4761 ;
  assign n11576 = n2745 & ~n3924 ;
  assign n11577 = ~n10808 & n11576 ;
  assign n11578 = ~n11575 & n11577 ;
  assign n11580 = n8577 ^ n2213 ^ 1'b0 ;
  assign n11579 = n4015 ^ n1698 ^ x246 ;
  assign n11581 = n11580 ^ n11579 ^ 1'b0 ;
  assign n11582 = n11581 ^ n10535 ^ 1'b0 ;
  assign n11583 = x212 & ~n11582 ;
  assign n11584 = n9433 ^ n3029 ^ 1'b0 ;
  assign n11585 = n11584 ^ n5307 ^ 1'b0 ;
  assign n11586 = n2750 & n5317 ;
  assign n11587 = n11586 ^ n4565 ^ 1'b0 ;
  assign n11588 = n11587 ^ n7300 ^ n2580 ;
  assign n11597 = ( n2576 & ~n4398 ) | ( n2576 & n8770 ) | ( ~n4398 & n8770 ) ;
  assign n11593 = ~n2252 & n3622 ;
  assign n11594 = n11593 ^ n3251 ^ 1'b0 ;
  assign n11589 = n763 | n6884 ;
  assign n11590 = n5992 ^ n2470 ^ n279 ;
  assign n11591 = ( n2714 & n11589 ) | ( n2714 & ~n11590 ) | ( n11589 & ~n11590 ) ;
  assign n11592 = ~n1162 & n11591 ;
  assign n11595 = n11594 ^ n11592 ^ n5599 ;
  assign n11596 = ~n8306 & n11595 ;
  assign n11598 = n11597 ^ n11596 ^ 1'b0 ;
  assign n11599 = n3360 & ~n6659 ;
  assign n11600 = n11599 ^ n5917 ^ n5682 ;
  assign n11601 = n7734 ^ n5029 ^ 1'b0 ;
  assign n11602 = n10167 & n11601 ;
  assign n11603 = ~n1854 & n11602 ;
  assign n11604 = ( n566 & n3391 ) | ( n566 & ~n11603 ) | ( n3391 & ~n11603 ) ;
  assign n11605 = ( n4536 & n10461 ) | ( n4536 & n11604 ) | ( n10461 & n11604 ) ;
  assign n11606 = n333 & ~n7698 ;
  assign n11607 = n11606 ^ n4612 ^ n4435 ;
  assign n11616 = n4154 & ~n10570 ;
  assign n11617 = n9589 & ~n11616 ;
  assign n11618 = n10569 & n11617 ;
  assign n11611 = n9197 ^ n3555 ^ 1'b0 ;
  assign n11612 = n2036 & n11611 ;
  assign n11613 = n11612 ^ n5685 ^ n3037 ;
  assign n11608 = n1663 | n2654 ;
  assign n11609 = n11608 ^ n1997 ^ 1'b0 ;
  assign n11610 = n6125 | n11609 ;
  assign n11614 = n11613 ^ n11610 ^ 1'b0 ;
  assign n11615 = n450 & ~n11614 ;
  assign n11619 = n11618 ^ n11615 ^ 1'b0 ;
  assign n11620 = n2338 ^ n1444 ^ n1054 ;
  assign n11621 = ~n11316 & n11620 ;
  assign n11622 = ( n2710 & ~n6324 ) | ( n2710 & n6904 ) | ( ~n6324 & n6904 ) ;
  assign n11623 = n11622 ^ n1380 ^ 1'b0 ;
  assign n11624 = n7895 ^ n5468 ^ 1'b0 ;
  assign n11625 = n4809 & ~n11624 ;
  assign n11626 = n8533 ^ n3200 ^ 1'b0 ;
  assign n11627 = n2455 & ~n11626 ;
  assign n11628 = ( ~n2841 & n11272 ) | ( ~n2841 & n11627 ) | ( n11272 & n11627 ) ;
  assign n11629 = n8977 ^ n8337 ^ 1'b0 ;
  assign n11630 = n3823 & ~n4600 ;
  assign n11631 = n1280 & n11630 ;
  assign n11632 = n3103 ^ n2369 ^ n406 ;
  assign n11633 = n11631 | n11632 ;
  assign n11634 = n3235 & ~n11633 ;
  assign n11635 = n7936 ^ n4238 ^ 1'b0 ;
  assign n11636 = n6685 ^ n2428 ^ 1'b0 ;
  assign n11637 = ~n11635 & n11636 ;
  assign n11638 = n10243 ^ n3335 ^ 1'b0 ;
  assign n11639 = ( n2800 & n11637 ) | ( n2800 & n11638 ) | ( n11637 & n11638 ) ;
  assign n11640 = x165 & n1117 ;
  assign n11641 = ~x216 & n11640 ;
  assign n11642 = n11641 ^ n11022 ^ n5092 ;
  assign n11643 = ( n11634 & n11639 ) | ( n11634 & ~n11642 ) | ( n11639 & ~n11642 ) ;
  assign n11644 = n3046 & ~n6227 ;
  assign n11645 = ( n1281 & n1690 ) | ( n1281 & ~n3402 ) | ( n1690 & ~n3402 ) ;
  assign n11646 = ( ~n2160 & n4041 ) | ( ~n2160 & n11645 ) | ( n4041 & n11645 ) ;
  assign n11647 = n1231 & n11646 ;
  assign n11648 = n9387 ^ x194 ^ 1'b0 ;
  assign n11649 = n11647 & n11648 ;
  assign n11650 = ( n2805 & ~n2972 ) | ( n2805 & n11649 ) | ( ~n2972 & n11649 ) ;
  assign n11651 = n11644 & ~n11650 ;
  assign n11652 = n4893 | n9259 ;
  assign n11653 = n6662 | n11652 ;
  assign n11654 = n5367 ^ n1390 ^ n905 ;
  assign n11655 = ~n1889 & n2383 ;
  assign n11656 = n11655 ^ n2542 ^ 1'b0 ;
  assign n11657 = n11656 ^ n1353 ^ 1'b0 ;
  assign n11658 = n2780 | n7841 ;
  assign n11659 = n11658 ^ n8605 ^ 1'b0 ;
  assign n11660 = ( n5910 & n11358 ) | ( n5910 & n11659 ) | ( n11358 & n11659 ) ;
  assign n11661 = ( n4162 & n8114 ) | ( n4162 & ~n11660 ) | ( n8114 & ~n11660 ) ;
  assign n11662 = ( ~n11654 & n11657 ) | ( ~n11654 & n11661 ) | ( n11657 & n11661 ) ;
  assign n11663 = n10530 ^ n9075 ^ 1'b0 ;
  assign n11664 = n8155 & ~n11663 ;
  assign n11665 = n2070 ^ n715 ^ 1'b0 ;
  assign n11666 = n1981 | n11665 ;
  assign n11667 = ( n3220 & n8757 ) | ( n3220 & ~n11666 ) | ( n8757 & ~n11666 ) ;
  assign n11668 = n11667 ^ n9396 ^ n7854 ;
  assign n11669 = n8090 & ~n11668 ;
  assign n11670 = ~n2339 & n7180 ;
  assign n11671 = ( n770 & n3776 ) | ( n770 & ~n6017 ) | ( n3776 & ~n6017 ) ;
  assign n11672 = ( ~n2923 & n4126 ) | ( ~n2923 & n11671 ) | ( n4126 & n11671 ) ;
  assign n11673 = n5979 ^ n3009 ^ 1'b0 ;
  assign n11674 = n10466 ^ n5520 ^ 1'b0 ;
  assign n11675 = ( n495 & ~n587 ) | ( n495 & n7770 ) | ( ~n587 & n7770 ) ;
  assign n11676 = n475 | n11675 ;
  assign n11677 = ( n7061 & n8913 ) | ( n7061 & n11676 ) | ( n8913 & n11676 ) ;
  assign n11678 = n2610 & ~n5726 ;
  assign n11679 = n11677 | n11678 ;
  assign n11680 = n1036 | n11159 ;
  assign n11681 = n6073 & n11115 ;
  assign n11682 = n8729 ^ n879 ^ 1'b0 ;
  assign n11683 = n3579 & ~n11682 ;
  assign n11684 = ~n11572 & n11683 ;
  assign n11685 = n9060 ^ n4721 ^ n4575 ;
  assign n11686 = n321 & ~n1247 ;
  assign n11687 = n11686 ^ n3206 ^ 1'b0 ;
  assign n11688 = n11685 & ~n11687 ;
  assign n11689 = n11688 ^ n1267 ^ 1'b0 ;
  assign n11690 = ~n4163 & n11689 ;
  assign n11692 = n4040 ^ n1891 ^ 1'b0 ;
  assign n11691 = n10240 ^ n9380 ^ n3761 ;
  assign n11693 = n11692 ^ n11691 ^ x213 ;
  assign n11694 = n3943 ^ n1278 ^ 1'b0 ;
  assign n11695 = n2778 & ~n10691 ;
  assign n11696 = n11695 ^ n3636 ^ 1'b0 ;
  assign n11697 = n11696 ^ n5204 ^ 1'b0 ;
  assign n11698 = n7052 & n11697 ;
  assign n11699 = x10 & n3449 ;
  assign n11700 = ( n1599 & n4789 ) | ( n1599 & ~n11699 ) | ( n4789 & ~n11699 ) ;
  assign n11701 = ~n3003 & n6684 ;
  assign n11702 = n6692 & ~n8540 ;
  assign n11703 = ( n11700 & ~n11701 ) | ( n11700 & n11702 ) | ( ~n11701 & n11702 ) ;
  assign n11709 = n2057 | n7531 ;
  assign n11710 = n11709 ^ n479 ^ 1'b0 ;
  assign n11704 = n6607 ^ n3306 ^ 1'b0 ;
  assign n11705 = x214 & n11704 ;
  assign n11706 = n8574 & n11705 ;
  assign n11707 = n11706 ^ n3472 ^ n2391 ;
  assign n11708 = n11707 ^ n7959 ^ 1'b0 ;
  assign n11711 = n11710 ^ n11708 ^ 1'b0 ;
  assign n11712 = n1375 | n11711 ;
  assign n11713 = ( n10717 & n11703 ) | ( n10717 & ~n11712 ) | ( n11703 & ~n11712 ) ;
  assign n11716 = n1091 & n1122 ;
  assign n11717 = n11716 ^ n9485 ^ 1'b0 ;
  assign n11718 = n627 & ~n11717 ;
  assign n11719 = ( ~n4839 & n6587 ) | ( ~n4839 & n11718 ) | ( n6587 & n11718 ) ;
  assign n11714 = n5320 ^ n508 ^ 1'b0 ;
  assign n11715 = n2286 & n11714 ;
  assign n11720 = n11719 ^ n11715 ^ 1'b0 ;
  assign n11721 = n399 | n1659 ;
  assign n11722 = n11721 ^ n3705 ^ 1'b0 ;
  assign n11723 = n11722 ^ n8951 ^ x45 ;
  assign n11724 = ~n9814 & n11723 ;
  assign n11725 = n2524 ^ n2249 ^ n1290 ;
  assign n11726 = n2477 ^ n1640 ^ 1'b0 ;
  assign n11727 = n3658 | n11726 ;
  assign n11728 = n11727 ^ n1434 ^ 1'b0 ;
  assign n11729 = n11725 | n11728 ;
  assign n11730 = n11729 ^ x128 ^ 1'b0 ;
  assign n11731 = n11730 ^ n7626 ^ 1'b0 ;
  assign n11732 = n4261 & ~n11731 ;
  assign n11733 = n3523 & n8390 ;
  assign n11734 = ~n6110 & n11733 ;
  assign n11735 = n1819 | n3682 ;
  assign n11736 = n327 & n6622 ;
  assign n11737 = ~n11735 & n11736 ;
  assign n11738 = n11737 ^ n5720 ^ 1'b0 ;
  assign n11739 = ~n8429 & n8763 ;
  assign n11740 = n4167 & ~n5969 ;
  assign n11741 = ( n6512 & n11739 ) | ( n6512 & ~n11740 ) | ( n11739 & ~n11740 ) ;
  assign n11742 = n8036 ^ n4302 ^ 1'b0 ;
  assign n11743 = ~n11741 & n11742 ;
  assign n11744 = ( ~n973 & n9344 ) | ( ~n973 & n11743 ) | ( n9344 & n11743 ) ;
  assign n11745 = ( ~n6109 & n7831 ) | ( ~n6109 & n9792 ) | ( n7831 & n9792 ) ;
  assign n11747 = ( n604 & n2283 ) | ( n604 & n3113 ) | ( n2283 & n3113 ) ;
  assign n11746 = ( n1539 & n2550 ) | ( n1539 & n7888 ) | ( n2550 & n7888 ) ;
  assign n11748 = n11747 ^ n11746 ^ 1'b0 ;
  assign n11749 = n7016 ^ n6238 ^ 1'b0 ;
  assign n11750 = n11748 & n11749 ;
  assign n11751 = n10409 ^ n1042 ^ 1'b0 ;
  assign n11752 = n4734 & n11751 ;
  assign n11753 = ~n4148 & n11752 ;
  assign n11754 = n11753 ^ n5202 ^ 1'b0 ;
  assign n11755 = n2091 | n11754 ;
  assign n11756 = n5320 & n11755 ;
  assign n11757 = n7542 ^ n4469 ^ 1'b0 ;
  assign n11760 = n4933 ^ n4025 ^ n2607 ;
  assign n11761 = ~n3315 & n11760 ;
  assign n11762 = n11761 ^ n597 ^ 1'b0 ;
  assign n11758 = n9130 ^ n2008 ^ 1'b0 ;
  assign n11759 = n11758 ^ n8019 ^ n3655 ;
  assign n11763 = n11762 ^ n11759 ^ 1'b0 ;
  assign n11764 = n11757 | n11763 ;
  assign n11765 = ~n822 & n4659 ;
  assign n11766 = n11765 ^ n2726 ^ n704 ;
  assign n11767 = x97 & n1068 ;
  assign n11768 = ( ~n3165 & n7526 ) | ( ~n3165 & n11767 ) | ( n7526 & n11767 ) ;
  assign n11769 = n11768 ^ n10004 ^ 1'b0 ;
  assign n11770 = n8599 ^ n7334 ^ n5496 ;
  assign n11771 = ( ~n11766 & n11769 ) | ( ~n11766 & n11770 ) | ( n11769 & n11770 ) ;
  assign n11772 = n11771 ^ x130 ^ 1'b0 ;
  assign n11773 = n3269 & n11772 ;
  assign n11774 = n5111 ^ n3851 ^ n987 ;
  assign n11775 = ~n2645 & n11774 ;
  assign n11776 = ( n496 & n4983 ) | ( n496 & n11775 ) | ( n4983 & n11775 ) ;
  assign n11777 = n4506 & ~n8534 ;
  assign n11778 = ( ~x132 & n3041 ) | ( ~x132 & n7713 ) | ( n3041 & n7713 ) ;
  assign n11779 = n11777 & ~n11778 ;
  assign n11780 = n11779 ^ n10514 ^ 1'b0 ;
  assign n11781 = n5124 ^ n4516 ^ n3278 ;
  assign n11782 = n5415 & n7748 ;
  assign n11783 = n4156 & ~n11782 ;
  assign n11784 = n11783 ^ n7856 ^ 1'b0 ;
  assign n11785 = n11212 | n11784 ;
  assign n11786 = n9098 ^ n7195 ^ 1'b0 ;
  assign n11787 = n3140 & n4378 ;
  assign n11788 = n2500 & ~n4989 ;
  assign n11789 = n11788 ^ n7206 ^ 1'b0 ;
  assign n11790 = n3509 | n11789 ;
  assign n11791 = ~n11155 & n11790 ;
  assign n11792 = n4378 ^ x154 ^ 1'b0 ;
  assign n11793 = n11289 | n11792 ;
  assign n11794 = ( n2205 & n3627 ) | ( n2205 & n6023 ) | ( n3627 & n6023 ) ;
  assign n11795 = ~n11793 & n11794 ;
  assign n11798 = n3205 & n3634 ;
  assign n11799 = ~n2410 & n11798 ;
  assign n11800 = n11799 ^ n946 ^ 1'b0 ;
  assign n11796 = n2705 | n4301 ;
  assign n11797 = ~n1977 & n11796 ;
  assign n11801 = n11800 ^ n11797 ^ 1'b0 ;
  assign n11802 = n11801 ^ n2201 ^ 1'b0 ;
  assign n11803 = ( n1709 & ~n11795 ) | ( n1709 & n11802 ) | ( ~n11795 & n11802 ) ;
  assign n11804 = ~n550 & n10995 ;
  assign n11805 = n749 & ~n11804 ;
  assign n11806 = n11805 ^ n584 ^ 1'b0 ;
  assign n11807 = n11806 ^ n968 ^ 1'b0 ;
  assign n11808 = n1222 ^ n533 ^ n449 ;
  assign n11809 = ( n4345 & n11807 ) | ( n4345 & n11808 ) | ( n11807 & n11808 ) ;
  assign n11810 = n8640 ^ n4322 ^ n459 ;
  assign n11813 = n10800 | n11130 ;
  assign n11811 = ( n2356 & ~n3604 ) | ( n2356 & n7254 ) | ( ~n3604 & n7254 ) ;
  assign n11812 = n2651 & ~n11811 ;
  assign n11814 = n11813 ^ n11812 ^ 1'b0 ;
  assign n11815 = n7949 ^ n1398 ^ 1'b0 ;
  assign n11816 = ~n5438 & n5728 ;
  assign n11817 = ~n11815 & n11816 ;
  assign n11818 = n9315 ^ n413 ^ 1'b0 ;
  assign n11819 = n10257 & ~n11818 ;
  assign n11820 = n11819 ^ n1654 ^ 1'b0 ;
  assign n11821 = ~n1206 & n11820 ;
  assign n11822 = n547 | n11231 ;
  assign n11823 = ~n11821 & n11822 ;
  assign n11824 = n614 & n6148 ;
  assign n11825 = n11824 ^ n2893 ^ 1'b0 ;
  assign n11826 = n4526 ^ n810 ^ 1'b0 ;
  assign n11827 = ( n1300 & n11825 ) | ( n1300 & ~n11826 ) | ( n11825 & ~n11826 ) ;
  assign n11828 = n6497 ^ n5503 ^ n4741 ;
  assign n11829 = n1878 | n3910 ;
  assign n11830 = n11829 ^ n2125 ^ 1'b0 ;
  assign n11831 = n7358 & n11830 ;
  assign n11832 = x22 & ~n5660 ;
  assign n11833 = n11832 ^ n3256 ^ 1'b0 ;
  assign n11834 = n11831 & ~n11833 ;
  assign n11835 = ~n5012 & n6364 ;
  assign n11836 = ~n11834 & n11835 ;
  assign n11837 = n11836 ^ n5507 ^ 1'b0 ;
  assign n11838 = ~n2345 & n8403 ;
  assign n11839 = n11837 | n11838 ;
  assign n11840 = n11839 ^ n4048 ^ 1'b0 ;
  assign n11841 = n3413 & ~n5992 ;
  assign n11842 = n3909 & ~n11841 ;
  assign n11843 = ~n1510 & n6021 ;
  assign n11844 = n11843 ^ n11505 ^ 1'b0 ;
  assign n11845 = x151 & n11844 ;
  assign n11846 = n1352 & ~n4214 ;
  assign n11847 = ~x58 & n11846 ;
  assign n11848 = n3476 ^ n511 ^ 1'b0 ;
  assign n11849 = n925 | n11848 ;
  assign n11850 = n11849 ^ n8538 ^ 1'b0 ;
  assign n11851 = ( ~n5217 & n11847 ) | ( ~n5217 & n11850 ) | ( n11847 & n11850 ) ;
  assign n11852 = n5956 & n7141 ;
  assign n11853 = n11852 ^ n1196 ^ 1'b0 ;
  assign n11854 = n11853 ^ n6587 ^ 1'b0 ;
  assign n11855 = n7357 & n11854 ;
  assign n11856 = n6331 & n11855 ;
  assign n11857 = ~n1385 & n11856 ;
  assign n11859 = n362 & n3813 ;
  assign n11860 = n3992 ^ n715 ^ 1'b0 ;
  assign n11861 = n11860 ^ n5489 ^ 1'b0 ;
  assign n11862 = n6353 & ~n11861 ;
  assign n11863 = ( n8482 & n11859 ) | ( n8482 & ~n11862 ) | ( n11859 & ~n11862 ) ;
  assign n11864 = n4404 & ~n11863 ;
  assign n11858 = n8339 ^ n6311 ^ 1'b0 ;
  assign n11865 = n11864 ^ n11858 ^ 1'b0 ;
  assign n11866 = n6812 ^ n5704 ^ 1'b0 ;
  assign n11867 = n11866 ^ n11769 ^ 1'b0 ;
  assign n11868 = n3031 & n11867 ;
  assign n11869 = n11868 ^ n9034 ^ x233 ;
  assign n11870 = n11673 & n11869 ;
  assign n11871 = n7950 & n11870 ;
  assign n11872 = n4423 ^ n3562 ^ n2774 ;
  assign n11873 = n11872 ^ n11043 ^ n3724 ;
  assign n11874 = ( n680 & n1067 ) | ( n680 & ~n1421 ) | ( n1067 & ~n1421 ) ;
  assign n11875 = n689 ^ n335 ^ 1'b0 ;
  assign n11876 = n11874 | n11875 ;
  assign n11877 = n11876 ^ n9088 ^ 1'b0 ;
  assign n11878 = ~n6626 & n11877 ;
  assign n11879 = n1225 ^ x14 ^ x5 ;
  assign n11880 = n9064 | n11879 ;
  assign n11881 = ( n570 & ~n3457 ) | ( n570 & n5521 ) | ( ~n3457 & n5521 ) ;
  assign n11882 = n2639 & ~n8762 ;
  assign n11883 = ~x109 & n11882 ;
  assign n11884 = ~n5195 & n5896 ;
  assign n11885 = n3728 & n11884 ;
  assign n11886 = n2724 | n11545 ;
  assign n11887 = ( ~n1524 & n4672 ) | ( ~n1524 & n11886 ) | ( n4672 & n11886 ) ;
  assign n11888 = n11887 ^ n5234 ^ n1589 ;
  assign n11889 = n6510 ^ n2527 ^ 1'b0 ;
  assign n11893 = n5507 ^ n2894 ^ 1'b0 ;
  assign n11894 = n11893 ^ n8614 ^ 1'b0 ;
  assign n11890 = n4332 ^ n3476 ^ 1'b0 ;
  assign n11891 = ~n5971 & n11890 ;
  assign n11892 = n10170 & ~n11891 ;
  assign n11895 = n11894 ^ n11892 ^ 1'b0 ;
  assign n11896 = n5223 | n11895 ;
  assign n11897 = ( n9113 & n9793 ) | ( n9113 & ~n11168 ) | ( n9793 & ~n11168 ) ;
  assign n11898 = n10648 ^ n6045 ^ 1'b0 ;
  assign n11899 = n9417 & ~n11898 ;
  assign n11900 = n4875 | n11899 ;
  assign n11901 = n11900 ^ n3803 ^ 1'b0 ;
  assign n11902 = n11901 ^ n11002 ^ n8683 ;
  assign n11903 = n2520 & n4941 ;
  assign n11904 = n11903 ^ n7907 ^ n5307 ;
  assign n11905 = ( ~n7243 & n10974 ) | ( ~n7243 & n11904 ) | ( n10974 & n11904 ) ;
  assign n11906 = n3711 & ~n5675 ;
  assign n11907 = n4549 & n11906 ;
  assign n11908 = n11907 ^ n855 ^ 1'b0 ;
  assign n11909 = x122 & ~n11908 ;
  assign n11910 = n3965 ^ n382 ^ 1'b0 ;
  assign n11911 = n11909 & n11910 ;
  assign n11912 = n11911 ^ n7921 ^ 1'b0 ;
  assign n11916 = n6023 & ~n10955 ;
  assign n11915 = ( n1569 & n6646 ) | ( n1569 & n11405 ) | ( n6646 & n11405 ) ;
  assign n11913 = n4229 | n5937 ;
  assign n11914 = n5210 & ~n11913 ;
  assign n11917 = n11916 ^ n11915 ^ n11914 ;
  assign n11920 = ~n297 & n3114 ;
  assign n11921 = ~n1214 & n11920 ;
  assign n11922 = n2781 & ~n11921 ;
  assign n11923 = n11922 ^ n2676 ^ 1'b0 ;
  assign n11924 = n10130 | n11923 ;
  assign n11919 = n7522 & n10763 ;
  assign n11925 = n11924 ^ n11919 ^ n5671 ;
  assign n11926 = n3761 & n11925 ;
  assign n11927 = ~n1939 & n11926 ;
  assign n11928 = n11927 ^ n6689 ^ 1'b0 ;
  assign n11929 = n468 & n11928 ;
  assign n11918 = ~n1978 & n10791 ;
  assign n11930 = n11929 ^ n11918 ^ 1'b0 ;
  assign n11931 = n11656 ^ n8447 ^ 1'b0 ;
  assign n11932 = ~n11930 & n11931 ;
  assign n11933 = n9169 | n9779 ;
  assign n11934 = n8327 & ~n11933 ;
  assign n11935 = ~n2226 & n4677 ;
  assign n11936 = n2082 & n11935 ;
  assign n11937 = n5401 ^ n2575 ^ 1'b0 ;
  assign n11938 = n4137 ^ n2409 ^ 1'b0 ;
  assign n11939 = n11938 ^ n4150 ^ 1'b0 ;
  assign n11940 = n11937 | n11939 ;
  assign n11941 = n11940 ^ n10072 ^ n3781 ;
  assign n11942 = n6995 & n11941 ;
  assign n11943 = ( n3526 & ~n4708 ) | ( n3526 & n11942 ) | ( ~n4708 & n11942 ) ;
  assign n11946 = n3251 ^ n1953 ^ n1464 ;
  assign n11945 = n10961 ^ n5466 ^ 1'b0 ;
  assign n11947 = n11946 ^ n11945 ^ n6651 ;
  assign n11948 = n7731 & ~n11947 ;
  assign n11944 = ~n5144 & n8279 ;
  assign n11949 = n11948 ^ n11944 ^ 1'b0 ;
  assign n11950 = n4889 & ~n8011 ;
  assign n11951 = n11950 ^ n4607 ^ 1'b0 ;
  assign n11952 = n4114 ^ n1372 ^ 1'b0 ;
  assign n11953 = ~n6797 & n11952 ;
  assign n11954 = n3578 ^ n3142 ^ 1'b0 ;
  assign n11955 = n11954 ^ n2789 ^ n2127 ;
  assign n11956 = ( ~n4453 & n11953 ) | ( ~n4453 & n11955 ) | ( n11953 & n11955 ) ;
  assign n11957 = n11956 ^ n11750 ^ n5299 ;
  assign n11958 = ( x203 & n3009 ) | ( x203 & ~n5373 ) | ( n3009 & ~n5373 ) ;
  assign n11959 = n8705 ^ n2655 ^ n1478 ;
  assign n11960 = n11959 ^ n577 ^ 1'b0 ;
  assign n11961 = n11958 | n11960 ;
  assign n11962 = ~n11700 & n11961 ;
  assign n11963 = n2528 | n11962 ;
  assign n11964 = n8011 ^ n4919 ^ n3286 ;
  assign n11965 = n10880 ^ n7559 ^ 1'b0 ;
  assign n11966 = n5987 & n7613 ;
  assign n11967 = n3813 & n11966 ;
  assign n11968 = n11967 ^ x239 ^ 1'b0 ;
  assign n11969 = ( n6796 & ~n7104 ) | ( n6796 & n7223 ) | ( ~n7104 & n7223 ) ;
  assign n11976 = ~n8175 & n8372 ;
  assign n11977 = ( ~n4718 & n6979 ) | ( ~n4718 & n11976 ) | ( n6979 & n11976 ) ;
  assign n11971 = n1140 & n3247 ;
  assign n11970 = n1850 | n7709 ;
  assign n11972 = n11971 ^ n11970 ^ 1'b0 ;
  assign n11973 = n3881 | n7965 ;
  assign n11974 = n11973 ^ n9256 ^ 1'b0 ;
  assign n11975 = ~n11972 & n11974 ;
  assign n11978 = n11977 ^ n11975 ^ 1'b0 ;
  assign n11979 = n11635 ^ n8083 ^ n2317 ;
  assign n11980 = n11979 ^ n4806 ^ n640 ;
  assign n11981 = n8700 ^ n1475 ^ 1'b0 ;
  assign n11982 = ~n1401 & n11981 ;
  assign n11983 = n3831 & ~n7992 ;
  assign n11984 = ~n11982 & n11983 ;
  assign n11985 = n3322 ^ n2600 ^ 1'b0 ;
  assign n11986 = n3907 & ~n11985 ;
  assign n11987 = n554 | n3096 ;
  assign n11988 = n11987 ^ n10498 ^ n7810 ;
  assign n11989 = n9153 ^ n2576 ^ 1'b0 ;
  assign n11990 = ( ~n1901 & n6058 ) | ( ~n1901 & n7352 ) | ( n6058 & n7352 ) ;
  assign n11991 = x15 & n11990 ;
  assign n11992 = n1655 & n11991 ;
  assign n11993 = n11284 ^ n9489 ^ n7026 ;
  assign n11994 = n2689 ^ n514 ^ 1'b0 ;
  assign n11995 = n1381 & n11994 ;
  assign n11996 = n5991 & ~n11995 ;
  assign n11998 = ( n771 & n810 ) | ( n771 & n6507 ) | ( n810 & n6507 ) ;
  assign n11999 = ( n3323 & n8408 ) | ( n3323 & n11998 ) | ( n8408 & n11998 ) ;
  assign n12000 = n11999 ^ n5089 ^ 1'b0 ;
  assign n11997 = n9605 ^ n4417 ^ n2904 ;
  assign n12001 = n12000 ^ n11997 ^ n8603 ;
  assign n12002 = ~n2657 & n6815 ;
  assign n12003 = ~n2803 & n12002 ;
  assign n12004 = n3951 ^ n857 ^ 1'b0 ;
  assign n12005 = n12003 | n12004 ;
  assign n12006 = n12005 ^ n5468 ^ 1'b0 ;
  assign n12007 = n8245 & ~n12006 ;
  assign n12008 = n12007 ^ n6253 ^ 1'b0 ;
  assign n12009 = n2686 & n11534 ;
  assign n12010 = n6697 ^ n3876 ^ 1'b0 ;
  assign n12011 = n4141 ^ n2021 ^ 1'b0 ;
  assign n12012 = n7698 & ~n8027 ;
  assign n12013 = n11146 ^ n1108 ^ 1'b0 ;
  assign n12014 = ( ~n2819 & n12012 ) | ( ~n2819 & n12013 ) | ( n12012 & n12013 ) ;
  assign n12015 = ( n6806 & ~n12011 ) | ( n6806 & n12014 ) | ( ~n12011 & n12014 ) ;
  assign n12016 = ( n1367 & ~n2059 ) | ( n1367 & n12015 ) | ( ~n2059 & n12015 ) ;
  assign n12017 = n5652 & ~n8768 ;
  assign n12018 = n12017 ^ n8012 ^ 1'b0 ;
  assign n12019 = ( ~n6064 & n10405 ) | ( ~n6064 & n11074 ) | ( n10405 & n11074 ) ;
  assign n12020 = n7000 ^ n4619 ^ 1'b0 ;
  assign n12021 = n12020 ^ n8448 ^ n4726 ;
  assign n12022 = n1171 & ~n4825 ;
  assign n12023 = n12022 ^ n8508 ^ 1'b0 ;
  assign n12024 = ~n11680 & n12023 ;
  assign n12027 = ( ~x92 & n1828 ) | ( ~x92 & n2030 ) | ( n1828 & n2030 ) ;
  assign n12028 = n12027 ^ n3325 ^ n1949 ;
  assign n12025 = n4509 ^ n1664 ^ 1'b0 ;
  assign n12026 = n10670 | n12025 ;
  assign n12029 = n12028 ^ n12026 ^ n8394 ;
  assign n12030 = n12029 ^ n2415 ^ 1'b0 ;
  assign n12031 = n2299 ^ n1570 ^ n816 ;
  assign n12032 = x251 & n12031 ;
  assign n12033 = x233 | n10466 ;
  assign n12034 = n2106 & ~n11851 ;
  assign n12035 = n12033 & n12034 ;
  assign n12036 = n7364 ^ n3553 ^ 1'b0 ;
  assign n12037 = n3462 | n12036 ;
  assign n12038 = n4167 & ~n9715 ;
  assign n12039 = n7327 ^ n1438 ^ 1'b0 ;
  assign n12040 = n12038 | n12039 ;
  assign n12041 = n3875 ^ n2498 ^ 1'b0 ;
  assign n12042 = n12041 ^ n7865 ^ 1'b0 ;
  assign n12043 = ~n6564 & n10277 ;
  assign n12044 = ~n409 & n2369 ;
  assign n12045 = n12044 ^ n2694 ^ 1'b0 ;
  assign n12046 = n12045 ^ n3325 ^ 1'b0 ;
  assign n12047 = n12046 ^ n2525 ^ n2286 ;
  assign n12051 = n8949 ^ n8740 ^ 1'b0 ;
  assign n12048 = n2870 & n9841 ;
  assign n12049 = n9878 | n12048 ;
  assign n12050 = n12049 ^ n6955 ^ 1'b0 ;
  assign n12052 = n12051 ^ n12050 ^ 1'b0 ;
  assign n12053 = ( ~n585 & n4366 ) | ( ~n585 & n7055 ) | ( n4366 & n7055 ) ;
  assign n12054 = n2345 & n12053 ;
  assign n12055 = ~n2903 & n3438 ;
  assign n12056 = n6955 & n12055 ;
  assign n12057 = n2071 | n12056 ;
  assign n12058 = n12054 | n12057 ;
  assign n12059 = ( ~n470 & n1562 ) | ( ~n470 & n3043 ) | ( n1562 & n3043 ) ;
  assign n12060 = n12059 ^ n5820 ^ 1'b0 ;
  assign n12061 = n12060 ^ n7421 ^ 1'b0 ;
  assign n12062 = n4177 & n8646 ;
  assign n12063 = n7308 & n10504 ;
  assign n12064 = n12063 ^ n3110 ^ 1'b0 ;
  assign n12065 = ~n2854 & n8911 ;
  assign n12066 = n12064 & n12065 ;
  assign n12067 = ( n6602 & n12062 ) | ( n6602 & n12066 ) | ( n12062 & n12066 ) ;
  assign n12068 = n7243 & n8250 ;
  assign n12069 = n12068 ^ n2469 ^ 1'b0 ;
  assign n12070 = n625 & n12069 ;
  assign n12071 = n12070 ^ n6531 ^ n4333 ;
  assign n12072 = n12071 ^ n5620 ^ n5451 ;
  assign n12073 = ( n5649 & ~n7098 ) | ( n5649 & n8950 ) | ( ~n7098 & n8950 ) ;
  assign n12074 = n898 & n1084 ;
  assign n12075 = n2492 & n12074 ;
  assign n12076 = n12075 ^ n8527 ^ 1'b0 ;
  assign n12077 = ( ~n1887 & n8313 ) | ( ~n1887 & n9377 ) | ( n8313 & n9377 ) ;
  assign n12078 = n2551 | n5637 ;
  assign n12079 = n5132 | n6355 ;
  assign n12080 = n12079 ^ n9377 ^ 1'b0 ;
  assign n12081 = ( x96 & n5038 ) | ( x96 & n12080 ) | ( n5038 & n12080 ) ;
  assign n12082 = ~n9620 & n12081 ;
  assign n12083 = n12082 ^ n5589 ^ 1'b0 ;
  assign n12084 = n9752 ^ n2146 ^ 1'b0 ;
  assign n12085 = n12084 ^ n6399 ^ 1'b0 ;
  assign n12086 = n4935 ^ n2726 ^ x243 ;
  assign n12087 = n12086 ^ n838 ^ 1'b0 ;
  assign n12088 = ( n3034 & n3717 ) | ( n3034 & ~n6969 ) | ( n3717 & ~n6969 ) ;
  assign n12089 = ~n733 & n12088 ;
  assign n12090 = n12087 & n12089 ;
  assign n12091 = n4334 | n6958 ;
  assign n12092 = n12091 ^ n2666 ^ 1'b0 ;
  assign n12093 = ( n2444 & n4671 ) | ( n2444 & ~n6367 ) | ( n4671 & ~n6367 ) ;
  assign n12094 = n12093 ^ n2169 ^ 1'b0 ;
  assign n12095 = n8888 & n12094 ;
  assign n12096 = n12092 & n12095 ;
  assign n12097 = n6111 | n7039 ;
  assign n12098 = n12096 & ~n12097 ;
  assign n12099 = ~n2027 & n5422 ;
  assign n12100 = n12098 & n12099 ;
  assign n12101 = n4214 ^ n2434 ^ x128 ;
  assign n12102 = ~n9370 & n12101 ;
  assign n12103 = n12100 & n12102 ;
  assign n12104 = n5779 | n9831 ;
  assign n12105 = n5416 & ~n11278 ;
  assign n12106 = n4346 ^ n3972 ^ n3813 ;
  assign n12107 = n10495 ^ n600 ^ 1'b0 ;
  assign n12108 = n615 & ~n12107 ;
  assign n12109 = n2306 & n12108 ;
  assign n12110 = ( n1353 & ~n1989 ) | ( n1353 & n2723 ) | ( ~n1989 & n2723 ) ;
  assign n12111 = n12110 ^ n2824 ^ n2092 ;
  assign n12112 = n5541 ^ n1497 ^ 1'b0 ;
  assign n12113 = n12111 & ~n12112 ;
  assign n12114 = n12113 ^ n5199 ^ n5085 ;
  assign n12115 = ~n9197 & n12114 ;
  assign n12116 = ~n6159 & n12115 ;
  assign n12117 = ( n12106 & ~n12109 ) | ( n12106 & n12116 ) | ( ~n12109 & n12116 ) ;
  assign n12118 = n258 & ~n12117 ;
  assign n12119 = n4688 | n7922 ;
  assign n12120 = n12119 ^ n11487 ^ 1'b0 ;
  assign n12121 = n303 & ~n6994 ;
  assign n12122 = n12121 ^ x8 ^ 1'b0 ;
  assign n12123 = n7470 | n12003 ;
  assign n12124 = n373 | n12123 ;
  assign n12125 = n9771 ^ n1287 ^ 1'b0 ;
  assign n12126 = n12125 ^ n8103 ^ n993 ;
  assign n12127 = n10670 ^ n6510 ^ x3 ;
  assign n12128 = ~n7824 & n8868 ;
  assign n12129 = n9710 & n12128 ;
  assign n12130 = ( n2709 & n5804 ) | ( n2709 & ~n12129 ) | ( n5804 & ~n12129 ) ;
  assign n12131 = ~n7732 & n12130 ;
  assign n12132 = ( n957 & n5471 ) | ( n957 & ~n8284 ) | ( n5471 & ~n8284 ) ;
  assign n12133 = n6328 & ~n12132 ;
  assign n12134 = n5359 ^ n3844 ^ 1'b0 ;
  assign n12135 = n1148 | n12134 ;
  assign n12136 = n8534 ^ n259 ^ 1'b0 ;
  assign n12137 = ~n2043 & n12136 ;
  assign n12138 = ~n12135 & n12137 ;
  assign n12139 = ~n9033 & n12138 ;
  assign n12140 = ( n8110 & ~n12133 ) | ( n8110 & n12139 ) | ( ~n12133 & n12139 ) ;
  assign n12145 = n1567 | n7103 ;
  assign n12146 = n12145 ^ n3518 ^ 1'b0 ;
  assign n12147 = ( n5310 & n7571 ) | ( n5310 & ~n12146 ) | ( n7571 & ~n12146 ) ;
  assign n12141 = n1759 | n7877 ;
  assign n12142 = n12141 ^ n2714 ^ 1'b0 ;
  assign n12143 = n12142 ^ n4359 ^ n2086 ;
  assign n12144 = ~n10902 & n12143 ;
  assign n12148 = n12147 ^ n12144 ^ 1'b0 ;
  assign n12149 = n4930 ^ n1140 ^ 1'b0 ;
  assign n12150 = n1491 | n12149 ;
  assign n12151 = n5868 | n12150 ;
  assign n12152 = n1312 & ~n12151 ;
  assign n12153 = n12152 ^ n4323 ^ 1'b0 ;
  assign n12154 = x71 & ~n12153 ;
  assign n12155 = n1743 ^ n1353 ^ 1'b0 ;
  assign n12156 = n11656 ^ n9463 ^ 1'b0 ;
  assign n12157 = n8370 & ~n12156 ;
  assign n12158 = n3459 | n4760 ;
  assign n12159 = n12157 | n12158 ;
  assign n12160 = ( ~n6906 & n10728 ) | ( ~n6906 & n12159 ) | ( n10728 & n12159 ) ;
  assign n12161 = ( n1529 & ~n2680 ) | ( n1529 & n5521 ) | ( ~n2680 & n5521 ) ;
  assign n12162 = n6543 & n12161 ;
  assign n12164 = n4589 ^ n4285 ^ n2070 ;
  assign n12165 = n1061 & ~n12164 ;
  assign n12166 = n6212 & n12165 ;
  assign n12163 = n10780 ^ n5006 ^ 1'b0 ;
  assign n12167 = n12166 ^ n12163 ^ 1'b0 ;
  assign n12168 = ( n2448 & ~n2467 ) | ( n2448 & n8019 ) | ( ~n2467 & n8019 ) ;
  assign n12169 = x126 & n7454 ;
  assign n12170 = ~n12168 & n12169 ;
  assign n12171 = n12170 ^ n10804 ^ 1'b0 ;
  assign n12172 = n961 & n5087 ;
  assign n12173 = ~n11476 & n12172 ;
  assign n12175 = n5136 & n5431 ;
  assign n12174 = ( n3135 & n4673 ) | ( n3135 & n6727 ) | ( n4673 & n6727 ) ;
  assign n12176 = n12175 ^ n12174 ^ n7123 ;
  assign n12177 = n2557 ^ n1050 ^ 1'b0 ;
  assign n12178 = n5126 | n6546 ;
  assign n12179 = n908 | n12178 ;
  assign n12180 = ~n12177 & n12179 ;
  assign n12181 = n11146 | n12180 ;
  assign n12182 = n9268 ^ n8638 ^ n1053 ;
  assign n12183 = n10976 | n12182 ;
  assign n12184 = n2442 ^ n1267 ^ 1'b0 ;
  assign n12185 = n12184 ^ n3690 ^ 1'b0 ;
  assign n12186 = n7146 | n12185 ;
  assign n12187 = n9842 | n12186 ;
  assign n12188 = n12187 ^ n3159 ^ 1'b0 ;
  assign n12189 = ~n943 & n6572 ;
  assign n12190 = n12189 ^ n2276 ^ 1'b0 ;
  assign n12191 = n1705 & n3546 ;
  assign n12192 = n7952 & n12191 ;
  assign n12193 = ( n3989 & ~n4912 ) | ( n3989 & n5364 ) | ( ~n4912 & n5364 ) ;
  assign n12194 = ( n8472 & n11359 ) | ( n8472 & n12193 ) | ( n11359 & n12193 ) ;
  assign n12195 = n12194 ^ n5378 ^ x186 ;
  assign n12196 = n12195 ^ n8422 ^ n1347 ;
  assign n12197 = ( n12190 & n12192 ) | ( n12190 & ~n12196 ) | ( n12192 & ~n12196 ) ;
  assign n12198 = ~n4381 & n7726 ;
  assign n12199 = n8290 & n12198 ;
  assign n12200 = n12199 ^ n5458 ^ 1'b0 ;
  assign n12201 = n12200 ^ n8324 ^ 1'b0 ;
  assign n12202 = n4247 & ~n5265 ;
  assign n12203 = n881 & n12202 ;
  assign n12204 = ( ~n939 & n5076 ) | ( ~n939 & n12203 ) | ( n5076 & n12203 ) ;
  assign n12205 = ( n1588 & n2438 ) | ( n1588 & n7237 ) | ( n2438 & n7237 ) ;
  assign n12210 = n5838 ^ n1241 ^ x12 ;
  assign n12206 = n3872 ^ n2014 ^ 1'b0 ;
  assign n12207 = n1822 & n12206 ;
  assign n12208 = ~n2553 & n6468 ;
  assign n12209 = ~n12207 & n12208 ;
  assign n12211 = n12210 ^ n12209 ^ 1'b0 ;
  assign n12212 = n12205 & ~n12211 ;
  assign n12213 = ( ~n3358 & n7650 ) | ( ~n3358 & n11614 ) | ( n7650 & n11614 ) ;
  assign n12214 = n1919 | n2896 ;
  assign n12215 = n12214 ^ n2592 ^ 1'b0 ;
  assign n12216 = n12215 ^ n8940 ^ n5303 ;
  assign n12218 = n1470 | n10655 ;
  assign n12219 = n903 | n12218 ;
  assign n12220 = n12219 ^ n4966 ^ 1'b0 ;
  assign n12217 = n869 | n4505 ;
  assign n12221 = n12220 ^ n12217 ^ 1'b0 ;
  assign n12222 = ( n5470 & n9316 ) | ( n5470 & ~n10004 ) | ( n9316 & ~n10004 ) ;
  assign n12223 = n12222 ^ n7953 ^ n6618 ;
  assign n12224 = n3740 & n10373 ;
  assign n12225 = n8894 & n12224 ;
  assign n12226 = n3452 ^ x19 ^ 1'b0 ;
  assign n12227 = n6279 ^ n4449 ^ n1557 ;
  assign n12228 = n12226 & n12227 ;
  assign n12229 = n12228 ^ n4460 ^ 1'b0 ;
  assign n12230 = ~n5125 & n8408 ;
  assign n12231 = n3080 | n4986 ;
  assign n12232 = n12231 ^ n2287 ^ 1'b0 ;
  assign n12233 = n4073 & ~n12232 ;
  assign n12234 = n12233 ^ n9655 ^ 1'b0 ;
  assign n12235 = n3709 | n6228 ;
  assign n12236 = n4503 & ~n12235 ;
  assign n12237 = n12236 ^ n4066 ^ n1663 ;
  assign n12238 = n12234 & n12237 ;
  assign n12239 = ~n12230 & n12238 ;
  assign n12240 = ~n1822 & n4260 ;
  assign n12241 = n5584 & n5685 ;
  assign n12242 = n12240 & n12241 ;
  assign n12243 = n2085 & ~n4478 ;
  assign n12244 = ~n6347 & n12243 ;
  assign n12245 = ( n1268 & n2759 ) | ( n1268 & ~n12244 ) | ( n2759 & ~n12244 ) ;
  assign n12246 = n12242 | n12245 ;
  assign n12250 = n2125 & ~n6534 ;
  assign n12251 = ( n1221 & n1920 ) | ( n1221 & ~n11843 ) | ( n1920 & ~n11843 ) ;
  assign n12252 = n12251 ^ n3696 ^ n2528 ;
  assign n12253 = ~n3802 & n12252 ;
  assign n12254 = n12250 & n12253 ;
  assign n12255 = ~n9066 & n12254 ;
  assign n12247 = n496 & n8210 ;
  assign n12248 = n12247 ^ n11684 ^ 1'b0 ;
  assign n12249 = n1953 & ~n12248 ;
  assign n12256 = n12255 ^ n12249 ^ 1'b0 ;
  assign n12257 = n307 & ~n2280 ;
  assign n12258 = n8637 & n12257 ;
  assign n12259 = n1684 & n6937 ;
  assign n12260 = ~n4119 & n12259 ;
  assign n12261 = n1732 & n12260 ;
  assign n12262 = ( n3110 & n5199 ) | ( n3110 & n6804 ) | ( n5199 & n6804 ) ;
  assign n12263 = ~n618 & n12262 ;
  assign n12264 = n5456 & ~n12263 ;
  assign n12265 = n12019 & n12264 ;
  assign n12266 = ( n4434 & ~n4445 ) | ( n4434 & n6175 ) | ( ~n4445 & n6175 ) ;
  assign n12267 = n12266 ^ n12233 ^ n1709 ;
  assign n12268 = n3744 ^ n3706 ^ 1'b0 ;
  assign n12269 = n1532 & n12268 ;
  assign n12272 = n9420 ^ n1470 ^ 1'b0 ;
  assign n12270 = ( n492 & ~n9410 ) | ( n492 & n12219 ) | ( ~n9410 & n12219 ) ;
  assign n12271 = n9200 & n12270 ;
  assign n12273 = n12272 ^ n12271 ^ 1'b0 ;
  assign n12274 = ( n7388 & ~n12269 ) | ( n7388 & n12273 ) | ( ~n12269 & n12273 ) ;
  assign n12278 = ( n3247 & n3693 ) | ( n3247 & n11937 ) | ( n3693 & n11937 ) ;
  assign n12279 = n12278 ^ n3638 ^ 1'b0 ;
  assign n12280 = ~n1408 & n12279 ;
  assign n12281 = n12280 ^ n3204 ^ 1'b0 ;
  assign n12275 = n6291 & n8297 ;
  assign n12276 = ~n2538 & n12275 ;
  assign n12277 = n12276 ^ n6272 ^ 1'b0 ;
  assign n12282 = n12281 ^ n12277 ^ n6458 ;
  assign n12283 = n12282 ^ n9165 ^ n5914 ;
  assign n12284 = n3782 ^ n1080 ^ 1'b0 ;
  assign n12285 = n9708 & ~n12284 ;
  assign n12286 = x73 & n4139 ;
  assign n12287 = n12286 ^ n5849 ^ 1'b0 ;
  assign n12288 = n10002 & ~n12287 ;
  assign n12296 = n7762 ^ n7216 ^ n703 ;
  assign n12297 = n12296 ^ n1169 ^ 1'b0 ;
  assign n12298 = n468 & ~n12297 ;
  assign n12294 = n10763 ^ n5365 ^ 1'b0 ;
  assign n12295 = n2845 & n12294 ;
  assign n12289 = n2700 ^ n1504 ^ 1'b0 ;
  assign n12290 = n3803 & n12289 ;
  assign n12291 = n12290 ^ n4978 ^ 1'b0 ;
  assign n12292 = n3627 ^ n3371 ^ 1'b0 ;
  assign n12293 = n12291 & n12292 ;
  assign n12299 = n12298 ^ n12295 ^ n12293 ;
  assign n12300 = ( ~n2547 & n3250 ) | ( ~n2547 & n12299 ) | ( n3250 & n12299 ) ;
  assign n12301 = n9766 ^ n7686 ^ 1'b0 ;
  assign n12302 = n12301 ^ n10215 ^ n9189 ;
  assign n12303 = ~n3032 & n5456 ;
  assign n12304 = n12303 ^ n966 ^ 1'b0 ;
  assign n12305 = n798 | n6562 ;
  assign n12306 = n3204 | n12305 ;
  assign n12307 = ~n12304 & n12306 ;
  assign n12308 = n12307 ^ n6658 ^ 1'b0 ;
  assign n12309 = n2861 & n12308 ;
  assign n12312 = ( n2793 & ~n3166 ) | ( n2793 & n6793 ) | ( ~n3166 & n6793 ) ;
  assign n12313 = n12312 ^ n5666 ^ 1'b0 ;
  assign n12314 = ( n1233 & n6162 ) | ( n1233 & ~n12313 ) | ( n6162 & ~n12313 ) ;
  assign n12310 = n7366 ^ n1202 ^ n1027 ;
  assign n12311 = n12310 ^ n4604 ^ n1211 ;
  assign n12315 = n12314 ^ n12311 ^ n1855 ;
  assign n12316 = n1816 & n2655 ;
  assign n12317 = n5800 & n12316 ;
  assign n12319 = n1938 & ~n11235 ;
  assign n12318 = n8649 & n12045 ;
  assign n12320 = n12319 ^ n12318 ^ 1'b0 ;
  assign n12321 = n12317 | n12320 ;
  assign n12322 = n444 | n12321 ;
  assign n12323 = ( ~n405 & n7713 ) | ( ~n405 & n9070 ) | ( n7713 & n9070 ) ;
  assign n12324 = n11777 & ~n12323 ;
  assign n12325 = n12324 ^ n3089 ^ 1'b0 ;
  assign n12326 = n4043 & n7154 ;
  assign n12335 = n1749 & ~n6856 ;
  assign n12327 = ( ~n1365 & n2478 ) | ( ~n1365 & n5796 ) | ( n2478 & n5796 ) ;
  assign n12328 = ~n370 & n3738 ;
  assign n12329 = n12327 & n12328 ;
  assign n12330 = n6188 ^ n3409 ^ 1'b0 ;
  assign n12331 = n1276 | n12330 ;
  assign n12332 = n988 | n12331 ;
  assign n12333 = n561 | n12332 ;
  assign n12334 = n12329 & n12333 ;
  assign n12336 = n12335 ^ n12334 ^ 1'b0 ;
  assign n12337 = n2201 & ~n3305 ;
  assign n12338 = ( ~n574 & n10133 ) | ( ~n574 & n12337 ) | ( n10133 & n12337 ) ;
  assign n12339 = n9678 ^ n3026 ^ 1'b0 ;
  assign n12340 = ~n1348 & n1512 ;
  assign n12341 = n2461 & n12340 ;
  assign n12342 = n12341 ^ n9668 ^ 1'b0 ;
  assign n12343 = n598 & ~n4073 ;
  assign n12344 = n5660 | n12343 ;
  assign n12345 = n12342 & ~n12344 ;
  assign n12346 = n10672 ^ n2977 ^ 1'b0 ;
  assign n12347 = x69 & ~n12346 ;
  assign n12348 = ( ~n4248 & n4351 ) | ( ~n4248 & n5111 ) | ( n4351 & n5111 ) ;
  assign n12349 = n12347 & ~n12348 ;
  assign n12350 = ~n1228 & n12349 ;
  assign n12351 = n2634 & n6295 ;
  assign n12352 = n4473 | n6211 ;
  assign n12353 = n2234 | n12352 ;
  assign n12354 = n12353 ^ n4606 ^ 1'b0 ;
  assign n12355 = n12351 & ~n12354 ;
  assign n12356 = n6331 ^ n561 ^ 1'b0 ;
  assign n12357 = ( ~n799 & n4434 ) | ( ~n799 & n7460 ) | ( n4434 & n7460 ) ;
  assign n12359 = n6374 ^ n4821 ^ 1'b0 ;
  assign n12358 = n4644 & n5137 ;
  assign n12360 = n12359 ^ n12358 ^ 1'b0 ;
  assign n12361 = n12357 & ~n12360 ;
  assign n12362 = ~n12356 & n12361 ;
  assign n12363 = ( n6160 & n9568 ) | ( n6160 & n12362 ) | ( n9568 & n12362 ) ;
  assign n12364 = ( n4214 & n10206 ) | ( n4214 & ~n12363 ) | ( n10206 & ~n12363 ) ;
  assign n12366 = n9518 ^ n1906 ^ 1'b0 ;
  assign n12365 = n6231 ^ n1477 ^ 1'b0 ;
  assign n12367 = n12366 ^ n12365 ^ 1'b0 ;
  assign n12368 = n8958 & n12367 ;
  assign n12369 = n10694 ^ n3584 ^ 1'b0 ;
  assign n12370 = n12369 ^ n10018 ^ 1'b0 ;
  assign n12371 = n4072 & ~n12370 ;
  assign n12372 = ( ~n3079 & n4032 ) | ( ~n3079 & n6101 ) | ( n4032 & n6101 ) ;
  assign n12373 = n12372 ^ n11199 ^ n9482 ;
  assign n12374 = n10411 & n12373 ;
  assign n12388 = n6534 ^ n2712 ^ 1'b0 ;
  assign n12384 = n3499 | n5100 ;
  assign n12385 = ( n1247 & n4794 ) | ( n1247 & ~n12384 ) | ( n4794 & ~n12384 ) ;
  assign n12380 = n3816 ^ x42 ^ 1'b0 ;
  assign n12379 = n4928 & n9521 ;
  assign n12381 = n12380 ^ n12379 ^ 1'b0 ;
  assign n12378 = n6597 ^ n6432 ^ n1784 ;
  assign n12382 = n12381 ^ n12378 ^ 1'b0 ;
  assign n12383 = n2822 & n12382 ;
  assign n12386 = n12385 ^ n12383 ^ n1604 ;
  assign n12375 = x25 & ~n2019 ;
  assign n12376 = n3088 & n12375 ;
  assign n12377 = n8330 & ~n12376 ;
  assign n12387 = n12386 ^ n12377 ^ 1'b0 ;
  assign n12389 = n12388 ^ n12387 ^ 1'b0 ;
  assign n12390 = ( n652 & ~n4809 ) | ( n652 & n7710 ) | ( ~n4809 & n7710 ) ;
  assign n12391 = n12390 ^ n10361 ^ 1'b0 ;
  assign n12392 = n3565 | n7963 ;
  assign n12393 = n7927 | n12392 ;
  assign n12395 = n3738 & ~n6312 ;
  assign n12396 = n12395 ^ n899 ^ 1'b0 ;
  assign n12394 = n5660 ^ n2750 ^ n1857 ;
  assign n12397 = n12396 ^ n12394 ^ n3457 ;
  assign n12400 = ( ~n2683 & n5685 ) | ( ~n2683 & n6629 ) | ( n5685 & n6629 ) ;
  assign n12398 = n4557 & ~n5969 ;
  assign n12399 = n12398 ^ n1658 ^ 1'b0 ;
  assign n12401 = n12400 ^ n12399 ^ n1935 ;
  assign n12402 = ~n2223 & n10655 ;
  assign n12403 = n12401 & n12402 ;
  assign n12404 = n4003 ^ n832 ^ 1'b0 ;
  assign n12405 = n10986 ^ n305 ^ 1'b0 ;
  assign n12406 = ~n4593 & n12405 ;
  assign n12407 = ( ~n7024 & n8122 ) | ( ~n7024 & n12406 ) | ( n8122 & n12406 ) ;
  assign n12408 = n12407 ^ n989 ^ 1'b0 ;
  assign n12409 = ~n9481 & n12408 ;
  assign n12410 = n3608 ^ n996 ^ 1'b0 ;
  assign n12411 = ( n6152 & n9794 ) | ( n6152 & ~n12410 ) | ( n9794 & ~n12410 ) ;
  assign n12412 = n9482 ^ n3228 ^ 1'b0 ;
  assign n12413 = n12411 | n12412 ;
  assign n12420 = n12142 ^ n8110 ^ 1'b0 ;
  assign n12414 = ( n1705 & n3029 ) | ( n1705 & n3641 ) | ( n3029 & n3641 ) ;
  assign n12415 = n6286 ^ n5753 ^ n4839 ;
  assign n12416 = n12414 | n12415 ;
  assign n12417 = n12416 ^ n10674 ^ 1'b0 ;
  assign n12418 = n12417 ^ n7300 ^ n4725 ;
  assign n12419 = n4356 & ~n12418 ;
  assign n12421 = n12420 ^ n12419 ^ n1630 ;
  assign n12422 = n10259 ^ n8698 ^ n5111 ;
  assign n12423 = n11196 ^ n7157 ^ n6886 ;
  assign n12424 = n12423 ^ n9635 ^ 1'b0 ;
  assign n12425 = n2746 ^ n1029 ^ 1'b0 ;
  assign n12426 = ( ~n8870 & n12424 ) | ( ~n8870 & n12425 ) | ( n12424 & n12425 ) ;
  assign n12428 = n8901 ^ n7819 ^ n5327 ;
  assign n12429 = ~n9124 & n12428 ;
  assign n12427 = ~n1176 & n6216 ;
  assign n12430 = n12429 ^ n12427 ^ 1'b0 ;
  assign n12431 = ~n8705 & n12430 ;
  assign n12432 = ~n12426 & n12431 ;
  assign n12433 = ( n1278 & ~n3543 ) | ( n1278 & n6962 ) | ( ~n3543 & n6962 ) ;
  assign n12434 = ( n5100 & n7643 ) | ( n5100 & ~n9068 ) | ( n7643 & ~n9068 ) ;
  assign n12435 = n12433 | n12434 ;
  assign n12436 = n12435 ^ n1819 ^ 1'b0 ;
  assign n12437 = n11860 ^ n9615 ^ n3141 ;
  assign n12438 = n11052 & n12437 ;
  assign n12439 = n11246 ^ n4374 ^ 1'b0 ;
  assign n12440 = n9588 ^ n3103 ^ 1'b0 ;
  assign n12441 = n9524 & ~n12440 ;
  assign n12442 = n7104 ^ n5869 ^ n4331 ;
  assign n12443 = ( n5038 & n10746 ) | ( n5038 & n12442 ) | ( n10746 & n12442 ) ;
  assign n12444 = n8120 | n9086 ;
  assign n12445 = n6113 | n10049 ;
  assign n12446 = n4512 & ~n12445 ;
  assign n12447 = ( ~n2448 & n4417 ) | ( ~n2448 & n6831 ) | ( n4417 & n6831 ) ;
  assign n12448 = n1321 & ~n1776 ;
  assign n12449 = ~n1828 & n12448 ;
  assign n12450 = n9590 ^ n8699 ^ n6575 ;
  assign n12451 = ~n4904 & n12450 ;
  assign n12452 = n12451 ^ n3131 ^ 1'b0 ;
  assign n12453 = n548 | n3133 ;
  assign n12454 = n12453 ^ n4025 ^ 1'b0 ;
  assign n12455 = n12454 ^ n12089 ^ 1'b0 ;
  assign n12456 = ( n841 & n2325 ) | ( n841 & n3216 ) | ( n2325 & n3216 ) ;
  assign n12457 = n12456 ^ n10363 ^ 1'b0 ;
  assign n12458 = n3019 | n12457 ;
  assign n12459 = n12458 ^ n5089 ^ 1'b0 ;
  assign n12460 = n3915 ^ n3819 ^ 1'b0 ;
  assign n12461 = ~n2871 & n8414 ;
  assign n12462 = n12461 ^ n10030 ^ 1'b0 ;
  assign n12463 = n12462 ^ n2401 ^ 1'b0 ;
  assign n12464 = n9722 & n12463 ;
  assign n12465 = ( n5730 & n12460 ) | ( n5730 & n12464 ) | ( n12460 & n12464 ) ;
  assign n12466 = n6229 | n12465 ;
  assign n12467 = n9155 ^ n2808 ^ 1'b0 ;
  assign n12469 = ( n857 & n3543 ) | ( n857 & ~n6146 ) | ( n3543 & ~n6146 ) ;
  assign n12468 = n396 | n10085 ;
  assign n12470 = n12469 ^ n12468 ^ 1'b0 ;
  assign n12471 = n12470 ^ n5574 ^ 1'b0 ;
  assign n12472 = n12467 & n12471 ;
  assign n12473 = n12472 ^ n1340 ^ 1'b0 ;
  assign n12474 = n6640 & ~n12473 ;
  assign n12475 = n8176 & n8939 ;
  assign n12476 = n5097 & n12475 ;
  assign n12481 = n1547 ^ n983 ^ 1'b0 ;
  assign n12482 = ~n4090 & n12481 ;
  assign n12483 = n12482 ^ n2255 ^ 1'b0 ;
  assign n12480 = ( x62 & n372 ) | ( x62 & ~n2085 ) | ( n372 & ~n2085 ) ;
  assign n12477 = n7595 ^ n3245 ^ n636 ;
  assign n12478 = n12477 ^ n6362 ^ n4163 ;
  assign n12479 = ~n576 & n12478 ;
  assign n12484 = n12483 ^ n12480 ^ n12479 ;
  assign n12485 = n9900 ^ n2238 ^ n608 ;
  assign n12486 = n5916 ^ n5885 ^ 1'b0 ;
  assign n12487 = n12485 & ~n12486 ;
  assign n12488 = n6349 & ~n12487 ;
  assign n12489 = ( n9803 & n12129 ) | ( n9803 & ~n12488 ) | ( n12129 & ~n12488 ) ;
  assign n12497 = n2383 & ~n3998 ;
  assign n12498 = ~n1255 & n12497 ;
  assign n12499 = n745 & ~n3788 ;
  assign n12500 = ~n1605 & n12499 ;
  assign n12501 = n12498 | n12500 ;
  assign n12502 = n12501 ^ n3180 ^ 1'b0 ;
  assign n12503 = ( n5342 & n7476 ) | ( n5342 & ~n12502 ) | ( n7476 & ~n12502 ) ;
  assign n12504 = n2995 | n12503 ;
  assign n12490 = n8859 ^ n2807 ^ 1'b0 ;
  assign n12491 = n7769 & ~n12490 ;
  assign n12492 = n12491 ^ n8124 ^ n5034 ;
  assign n12493 = n12492 ^ n5995 ^ 1'b0 ;
  assign n12494 = n4773 ^ n4763 ^ 1'b0 ;
  assign n12495 = n12493 & n12494 ;
  assign n12496 = ~n1876 & n12495 ;
  assign n12505 = n12504 ^ n12496 ^ 1'b0 ;
  assign n12506 = n9799 & n12505 ;
  assign n12507 = n7382 ^ n5513 ^ 1'b0 ;
  assign n12508 = n1435 & n9856 ;
  assign n12509 = n5766 ^ n3163 ^ 1'b0 ;
  assign n12510 = ( n7270 & ~n10229 ) | ( n7270 & n12509 ) | ( ~n10229 & n12509 ) ;
  assign n12511 = n8465 | n9994 ;
  assign n12512 = n12510 | n12511 ;
  assign n12514 = n853 & n3572 ;
  assign n12515 = n8304 & n12514 ;
  assign n12513 = x58 & n629 ;
  assign n12516 = n12515 ^ n12513 ^ 1'b0 ;
  assign n12517 = ( x216 & n8487 ) | ( x216 & ~n10073 ) | ( n8487 & ~n10073 ) ;
  assign n12518 = n12517 ^ n9557 ^ 1'b0 ;
  assign n12519 = ~n11371 & n12518 ;
  assign n12520 = n4308 & ~n5293 ;
  assign n12521 = n12520 ^ n2109 ^ 1'b0 ;
  assign n12522 = n4906 ^ n1256 ^ n625 ;
  assign n12523 = n2563 & n12522 ;
  assign n12524 = n1353 & n12523 ;
  assign n12532 = ( n761 & n1545 ) | ( n761 & n1857 ) | ( n1545 & n1857 ) ;
  assign n12533 = ( n1475 & ~n4335 ) | ( n1475 & n12532 ) | ( ~n4335 & n12532 ) ;
  assign n12534 = x230 & n12533 ;
  assign n12535 = n12534 ^ n4886 ^ 1'b0 ;
  assign n12525 = ( ~n2148 & n7838 ) | ( ~n2148 & n8392 ) | ( n7838 & n8392 ) ;
  assign n12526 = ( x102 & ~n585 ) | ( x102 & n809 ) | ( ~n585 & n809 ) ;
  assign n12527 = n8528 | n11995 ;
  assign n12528 = ( ~n4793 & n5994 ) | ( ~n4793 & n12527 ) | ( n5994 & n12527 ) ;
  assign n12529 = n12528 ^ x213 ^ 1'b0 ;
  assign n12530 = n12526 & n12529 ;
  assign n12531 = ~n12525 & n12530 ;
  assign n12536 = n12535 ^ n12531 ^ 1'b0 ;
  assign n12537 = n4223 & ~n12536 ;
  assign n12539 = n7036 ^ n481 ^ x194 ;
  assign n12538 = n11376 ^ n7561 ^ n3996 ;
  assign n12540 = n12539 ^ n12538 ^ n4818 ;
  assign n12546 = n8919 ^ n6228 ^ n4041 ;
  assign n12547 = n12546 ^ n3311 ^ 1'b0 ;
  assign n12541 = n11937 ^ n6641 ^ n1020 ;
  assign n12542 = n12541 ^ n3984 ^ 1'b0 ;
  assign n12543 = ~n642 & n12542 ;
  assign n12544 = n12543 ^ n6321 ^ 1'b0 ;
  assign n12545 = n11620 & ~n12544 ;
  assign n12548 = n12547 ^ n12545 ^ 1'b0 ;
  assign n12549 = n11291 ^ n4231 ^ x34 ;
  assign n12550 = ~n6219 & n12549 ;
  assign n12551 = n12550 ^ n9498 ^ 1'b0 ;
  assign n12552 = n393 & n12551 ;
  assign n12553 = n9947 & n12552 ;
  assign n12554 = n12548 & n12553 ;
  assign n12555 = n704 & ~n7464 ;
  assign n12556 = n12555 ^ n2170 ^ 1'b0 ;
  assign n12557 = n12556 ^ n573 ^ 1'b0 ;
  assign n12558 = ~n2968 & n12557 ;
  assign n12559 = n12554 | n12558 ;
  assign n12560 = n6162 | n12559 ;
  assign n12561 = n12122 ^ n10524 ^ n2040 ;
  assign n12562 = ( n575 & ~n1537 ) | ( n575 & n1690 ) | ( ~n1537 & n1690 ) ;
  assign n12563 = ( n3238 & ~n3465 ) | ( n3238 & n12562 ) | ( ~n3465 & n12562 ) ;
  assign n12564 = n9474 ^ n4603 ^ n3732 ;
  assign n12565 = n12563 & ~n12564 ;
  assign n12568 = n2705 & n9244 ;
  assign n12569 = ~n2032 & n12568 ;
  assign n12567 = n1475 | n7886 ;
  assign n12570 = n12569 ^ n12567 ^ 1'b0 ;
  assign n12566 = n8425 ^ n5899 ^ 1'b0 ;
  assign n12571 = n12570 ^ n12566 ^ n12541 ;
  assign n12572 = n6319 ^ n779 ^ 1'b0 ;
  assign n12573 = ~n3363 & n4048 ;
  assign n12574 = ~n5082 & n12573 ;
  assign n12575 = n2623 | n12574 ;
  assign n12576 = n642 ^ x90 ^ x49 ;
  assign n12577 = n12576 ^ n3069 ^ n2500 ;
  assign n12578 = ( n989 & n5233 ) | ( n989 & ~n5850 ) | ( n5233 & ~n5850 ) ;
  assign n12579 = ( n9024 & ~n12577 ) | ( n9024 & n12578 ) | ( ~n12577 & n12578 ) ;
  assign n12580 = n2004 | n12579 ;
  assign n12581 = ( n2175 & n12295 ) | ( n2175 & ~n12580 ) | ( n12295 & ~n12580 ) ;
  assign n12582 = n7637 & ~n12581 ;
  assign n12583 = ~n6560 & n6733 ;
  assign n12584 = n12583 ^ n7478 ^ 1'b0 ;
  assign n12585 = n6346 | n12584 ;
  assign n12586 = n9994 ^ n4391 ^ x198 ;
  assign n12594 = ( ~x233 & n3888 ) | ( ~x233 & n4849 ) | ( n3888 & n4849 ) ;
  assign n12595 = ( n952 & ~n2676 ) | ( n952 & n5749 ) | ( ~n2676 & n5749 ) ;
  assign n12596 = n12594 & n12595 ;
  assign n12592 = ~n943 & n3692 ;
  assign n12593 = n12592 ^ n1908 ^ 1'b0 ;
  assign n12589 = n2560 ^ n1601 ^ 1'b0 ;
  assign n12590 = n438 & ~n12589 ;
  assign n12587 = n2388 | n8041 ;
  assign n12588 = n2971 | n12587 ;
  assign n12591 = n12590 ^ n12588 ^ n4677 ;
  assign n12597 = n12596 ^ n12593 ^ n12591 ;
  assign n12598 = n11808 ^ n11443 ^ 1'b0 ;
  assign n12599 = ( n2333 & n10010 ) | ( n2333 & ~n12598 ) | ( n10010 & ~n12598 ) ;
  assign n12600 = ~n868 & n4720 ;
  assign n12601 = n1121 & n12600 ;
  assign n12602 = n12601 ^ x48 ^ 1'b0 ;
  assign n12603 = n6514 | n7785 ;
  assign n12604 = n12602 | n12603 ;
  assign n12607 = n12210 ^ n5285 ^ x44 ;
  assign n12605 = n6173 ^ n4198 ^ 1'b0 ;
  assign n12606 = n12605 ^ n5998 ^ n4803 ;
  assign n12608 = n12607 ^ n12606 ^ 1'b0 ;
  assign n12609 = ~n11927 & n12608 ;
  assign n12610 = n11291 ^ n10849 ^ n3644 ;
  assign n12611 = ( n12300 & n12483 ) | ( n12300 & n12610 ) | ( n12483 & n12610 ) ;
  assign n12612 = ( n1671 & n3460 ) | ( n1671 & ~n4806 ) | ( n3460 & ~n4806 ) ;
  assign n12613 = ( n1014 & n3702 ) | ( n1014 & n12612 ) | ( n3702 & n12612 ) ;
  assign n12614 = n4137 ^ n1305 ^ n962 ;
  assign n12615 = n12614 ^ n2949 ^ 1'b0 ;
  assign n12616 = n12615 ^ n12287 ^ n1121 ;
  assign n12617 = n2153 | n2502 ;
  assign n12618 = ( n2939 & n4978 ) | ( n2939 & n12617 ) | ( n4978 & n12617 ) ;
  assign n12619 = n10620 ^ n2892 ^ 1'b0 ;
  assign n12620 = ( ~n7874 & n8903 ) | ( ~n7874 & n10745 ) | ( n8903 & n10745 ) ;
  assign n12621 = n1250 & ~n4963 ;
  assign n12622 = ( n2057 & n12620 ) | ( n2057 & n12621 ) | ( n12620 & n12621 ) ;
  assign n12623 = n7541 & ~n8130 ;
  assign n12624 = ~n7903 & n12623 ;
  assign n12625 = n2073 & ~n12624 ;
  assign n12626 = n12625 ^ n11977 ^ 1'b0 ;
  assign n12627 = n5402 ^ n4498 ^ 1'b0 ;
  assign n12628 = n12627 ^ n4068 ^ 1'b0 ;
  assign n12629 = ~n4978 & n10954 ;
  assign n12630 = n12629 ^ n11298 ^ 1'b0 ;
  assign n12633 = n1848 | n6375 ;
  assign n12634 = n12633 ^ n9875 ^ 1'b0 ;
  assign n12635 = n12634 ^ n11580 ^ n1632 ;
  assign n12631 = n6475 ^ n1155 ^ 1'b0 ;
  assign n12632 = n481 & n12631 ;
  assign n12636 = n12635 ^ n12632 ^ 1'b0 ;
  assign n12637 = n10722 ^ n1861 ^ 1'b0 ;
  assign n12638 = ~n905 & n12637 ;
  assign n12639 = ( ~n6420 & n12062 ) | ( ~n6420 & n12638 ) | ( n12062 & n12638 ) ;
  assign n12640 = n9695 ^ n4167 ^ n660 ;
  assign n12641 = n7174 ^ n4906 ^ 1'b0 ;
  assign n12642 = ~n12640 & n12641 ;
  assign n12643 = n2790 | n6911 ;
  assign n12644 = n12642 | n12643 ;
  assign n12645 = n8124 | n8940 ;
  assign n12646 = n7843 | n11090 ;
  assign n12647 = ~n9572 & n12646 ;
  assign n12648 = x227 & ~n1168 ;
  assign n12649 = n5658 ^ n4215 ^ n716 ;
  assign n12650 = n560 | n12649 ;
  assign n12651 = n7477 | n12650 ;
  assign n12652 = n8652 ^ n6853 ^ 1'b0 ;
  assign n12653 = ~n8538 & n12652 ;
  assign n12654 = n12653 ^ n7752 ^ 1'b0 ;
  assign n12655 = ( ~n10334 & n12651 ) | ( ~n10334 & n12654 ) | ( n12651 & n12654 ) ;
  assign n12656 = n12648 & ~n12655 ;
  assign n12657 = n6648 ^ n4620 ^ 1'b0 ;
  assign n12658 = n11650 ^ n3063 ^ n680 ;
  assign n12659 = n10004 ^ n9635 ^ n9512 ;
  assign n12660 = n12659 ^ n8850 ^ n808 ;
  assign n12661 = n9089 | n12660 ;
  assign n12662 = ~n706 & n8210 ;
  assign n12663 = n12662 ^ n597 ^ 1'b0 ;
  assign n12664 = n10382 ^ n9486 ^ 1'b0 ;
  assign n12665 = n1830 & ~n12664 ;
  assign n12667 = ~n4875 & n6421 ;
  assign n12668 = ~x162 & n12667 ;
  assign n12669 = ( n2363 & ~n2559 ) | ( n2363 & n3913 ) | ( ~n2559 & n3913 ) ;
  assign n12670 = n4973 & n12669 ;
  assign n12671 = n8705 | n12670 ;
  assign n12672 = n12668 & ~n12671 ;
  assign n12673 = n12672 ^ n1205 ^ x202 ;
  assign n12666 = n8296 & n11034 ;
  assign n12674 = n12673 ^ n12666 ^ n9463 ;
  assign n12675 = n7125 ^ n4737 ^ n1403 ;
  assign n12676 = n7972 & n12675 ;
  assign n12677 = ~n716 & n12676 ;
  assign n12678 = n8764 | n12677 ;
  assign n12679 = n4821 | n12678 ;
  assign n12681 = n11029 ^ n964 ^ 1'b0 ;
  assign n12682 = n683 | n12681 ;
  assign n12683 = ( n1581 & n3475 ) | ( n1581 & n12682 ) | ( n3475 & n12682 ) ;
  assign n12684 = ( ~n2388 & n4051 ) | ( ~n2388 & n12683 ) | ( n4051 & n12683 ) ;
  assign n12685 = n587 & n12684 ;
  assign n12680 = n1659 | n12465 ;
  assign n12686 = n12685 ^ n12680 ^ 1'b0 ;
  assign n12687 = ( n2022 & n4621 ) | ( n2022 & n4727 ) | ( n4621 & n4727 ) ;
  assign n12688 = n12687 ^ n12086 ^ n6000 ;
  assign n12689 = ~n8573 & n12688 ;
  assign n12690 = n1604 & n12689 ;
  assign n12691 = x44 & ~n8053 ;
  assign n12692 = n12690 & n12691 ;
  assign n12696 = ( ~n8383 & n8758 ) | ( ~n8383 & n10494 ) | ( n8758 & n10494 ) ;
  assign n12693 = n8068 | n12454 ;
  assign n12694 = n12693 ^ n8297 ^ 1'b0 ;
  assign n12695 = ~n11859 & n12694 ;
  assign n12697 = n12696 ^ n12695 ^ 1'b0 ;
  assign n12698 = ~n2033 & n12697 ;
  assign n12699 = n12698 ^ n6434 ^ 1'b0 ;
  assign n12700 = ( ~n3079 & n5716 ) | ( ~n3079 & n10468 ) | ( n5716 & n10468 ) ;
  assign n12702 = n11725 ^ n4741 ^ n1097 ;
  assign n12701 = n8811 ^ n7797 ^ 1'b0 ;
  assign n12703 = n12702 ^ n12701 ^ n4444 ;
  assign n12704 = ~n1080 & n3104 ;
  assign n12705 = n12704 ^ n2434 ^ 1'b0 ;
  assign n12706 = ( n12700 & n12703 ) | ( n12700 & n12705 ) | ( n12703 & n12705 ) ;
  assign n12707 = n6123 & ~n7055 ;
  assign n12708 = n6818 & n7992 ;
  assign n12709 = n12708 ^ n9738 ^ 1'b0 ;
  assign n12710 = n11460 & ~n12709 ;
  assign n12711 = n7561 & n12710 ;
  assign n12712 = ~n2805 & n7135 ;
  assign n12713 = n12712 ^ n5921 ^ 1'b0 ;
  assign n12714 = n12713 ^ n3257 ^ n2254 ;
  assign n12715 = n6502 ^ n6497 ^ n2283 ;
  assign n12716 = ( n7411 & ~n8399 ) | ( n7411 & n12715 ) | ( ~n8399 & n12715 ) ;
  assign n12717 = n12716 ^ n12709 ^ n10951 ;
  assign n12718 = n619 | n8907 ;
  assign n12719 = n12718 ^ n12052 ^ n2594 ;
  assign n12720 = n4142 & ~n7143 ;
  assign n12721 = n1064 & n12720 ;
  assign n12722 = n6013 ^ n1808 ^ 1'b0 ;
  assign n12723 = n6534 & ~n12722 ;
  assign n12724 = n12723 ^ n5295 ^ 1'b0 ;
  assign n12725 = n1855 & ~n12724 ;
  assign n12726 = ~n3415 & n5820 ;
  assign n12727 = n338 & ~n4799 ;
  assign n12728 = n12727 ^ x125 ^ 1'b0 ;
  assign n12729 = ( n3559 & n7189 ) | ( n3559 & n12728 ) | ( n7189 & n12728 ) ;
  assign n12730 = ( n11052 & n12726 ) | ( n11052 & ~n12729 ) | ( n12726 & ~n12729 ) ;
  assign n12732 = n5685 ^ x24 ^ 1'b0 ;
  assign n12733 = ~n2794 & n12732 ;
  assign n12731 = ~n3804 & n9218 ;
  assign n12734 = n12733 ^ n12731 ^ 1'b0 ;
  assign n12735 = n9803 & ~n12734 ;
  assign n12736 = n5228 ^ n4346 ^ n1111 ;
  assign n12737 = n12736 ^ n4898 ^ 1'b0 ;
  assign n12738 = n5461 ^ n1307 ^ 1'b0 ;
  assign n12739 = n12738 ^ n4143 ^ 1'b0 ;
  assign n12740 = ( n2740 & n3076 ) | ( n2740 & ~n12045 ) | ( n3076 & ~n12045 ) ;
  assign n12741 = n9129 ^ n8394 ^ n1752 ;
  assign n12742 = n9378 & ~n12741 ;
  assign n12743 = n12740 & ~n12742 ;
  assign n12744 = n751 & n12743 ;
  assign n12745 = n3425 ^ n905 ^ n332 ;
  assign n12746 = ( n11790 & n11821 ) | ( n11790 & n12745 ) | ( n11821 & n12745 ) ;
  assign n12747 = ( n1810 & n2840 ) | ( n1810 & ~n8887 ) | ( n2840 & ~n8887 ) ;
  assign n12748 = ~n3833 & n5035 ;
  assign n12749 = n1795 & n11576 ;
  assign n12750 = n12749 ^ n4686 ^ 1'b0 ;
  assign n12751 = ( n5680 & n10638 ) | ( n5680 & ~n12750 ) | ( n10638 & ~n12750 ) ;
  assign n12752 = n10800 & n12751 ;
  assign n12753 = ( ~n4845 & n12748 ) | ( ~n4845 & n12752 ) | ( n12748 & n12752 ) ;
  assign n12754 = n9620 ^ x87 ^ 1'b0 ;
  assign n12755 = n2430 & ~n10756 ;
  assign n12761 = n8593 ^ n1844 ^ n1582 ;
  assign n12756 = n1048 ^ n446 ^ 1'b0 ;
  assign n12757 = n12756 ^ n8015 ^ n7833 ;
  assign n12758 = ~n8894 & n12757 ;
  assign n12759 = ~n8295 & n12758 ;
  assign n12760 = n10887 | n12759 ;
  assign n12762 = n12761 ^ n12760 ^ 1'b0 ;
  assign n12763 = n6337 ^ n4440 ^ n3327 ;
  assign n12764 = n7752 ^ n2825 ^ n576 ;
  assign n12765 = n838 | n1759 ;
  assign n12766 = n12764 & ~n12765 ;
  assign n12767 = n12766 ^ n1169 ^ n748 ;
  assign n12768 = n1197 & ~n9419 ;
  assign n12769 = ~n7403 & n12768 ;
  assign n12770 = n3795 | n11757 ;
  assign n12771 = n4763 | n12770 ;
  assign n12780 = n2764 ^ n940 ^ 1'b0 ;
  assign n12772 = n416 | n1953 ;
  assign n12773 = n12772 ^ n1051 ^ 1'b0 ;
  assign n12774 = n5529 ^ n1983 ^ 1'b0 ;
  assign n12775 = n12773 & ~n12774 ;
  assign n12776 = ( n5451 & ~n12121 ) | ( n5451 & n12775 ) | ( ~n12121 & n12775 ) ;
  assign n12777 = n12776 ^ n11916 ^ n11088 ;
  assign n12778 = n12777 ^ n1832 ^ 1'b0 ;
  assign n12779 = n4416 | n12778 ;
  assign n12781 = n12780 ^ n12779 ^ 1'b0 ;
  assign n12782 = n6152 ^ n4474 ^ 1'b0 ;
  assign n12783 = n2788 & ~n12782 ;
  assign n12784 = ~n4014 & n9130 ;
  assign n12785 = n5989 | n10634 ;
  assign n12792 = n4757 ^ n3985 ^ 1'b0 ;
  assign n12787 = n1357 | n2457 ;
  assign n12788 = n316 & ~n12787 ;
  assign n12789 = n3746 | n12788 ;
  assign n12786 = ( ~n847 & n3880 ) | ( ~n847 & n11303 ) | ( n3880 & n11303 ) ;
  assign n12790 = n12789 ^ n12786 ^ n6837 ;
  assign n12791 = n1494 | n12790 ;
  assign n12793 = n12792 ^ n12791 ^ 1'b0 ;
  assign n12794 = n5216 & n7929 ;
  assign n12795 = n12794 ^ n5741 ^ 1'b0 ;
  assign n12796 = ( ~n5356 & n5825 ) | ( ~n5356 & n12795 ) | ( n5825 & n12795 ) ;
  assign n12797 = n12796 ^ n5202 ^ 1'b0 ;
  assign n12798 = n2401 ^ n936 ^ 1'b0 ;
  assign n12799 = n373 & n12798 ;
  assign n12800 = n12799 ^ n1852 ^ 1'b0 ;
  assign n12801 = n12800 ^ n9599 ^ n550 ;
  assign n12805 = n3004 ^ n1661 ^ 1'b0 ;
  assign n12802 = n575 | n3455 ;
  assign n12803 = n12802 ^ n6030 ^ 1'b0 ;
  assign n12804 = n6628 & n12803 ;
  assign n12806 = n12805 ^ n12804 ^ 1'b0 ;
  assign n12807 = ~n8896 & n12806 ;
  assign n12808 = n5439 ^ n1090 ^ 1'b0 ;
  assign n12809 = x3 & ~n12808 ;
  assign n12810 = ~n3583 & n12809 ;
  assign n12811 = ~n5049 & n12810 ;
  assign n12812 = n12811 ^ n7509 ^ 1'b0 ;
  assign n12818 = n4017 ^ n1581 ^ 1'b0 ;
  assign n12819 = x142 & n12818 ;
  assign n12820 = ( n3457 & ~n5003 ) | ( n3457 & n12819 ) | ( ~n5003 & n12819 ) ;
  assign n12813 = ( n2823 & ~n5714 ) | ( n2823 & n8433 ) | ( ~n5714 & n8433 ) ;
  assign n12814 = n12813 ^ n5418 ^ 1'b0 ;
  assign n12815 = ( x208 & n4754 ) | ( x208 & n12814 ) | ( n4754 & n12814 ) ;
  assign n12816 = n5289 ^ n1512 ^ 1'b0 ;
  assign n12817 = n12815 & ~n12816 ;
  assign n12821 = n12820 ^ n12817 ^ 1'b0 ;
  assign n12822 = n12821 ^ n10183 ^ 1'b0 ;
  assign n12823 = n11459 ^ n6311 ^ n503 ;
  assign n12824 = n8465 & ~n12823 ;
  assign n12825 = n5445 & n7841 ;
  assign n12826 = ~n12605 & n12825 ;
  assign n12827 = n11767 ^ n6647 ^ 1'b0 ;
  assign n12828 = n12826 | n12827 ;
  assign n12829 = n12824 | n12828 ;
  assign n12830 = n6630 & n12829 ;
  assign n12831 = n7289 ^ n1964 ^ 1'b0 ;
  assign n12832 = n12831 ^ n7817 ^ n7558 ;
  assign n12833 = ~n2374 & n4635 ;
  assign n12834 = n12833 ^ n586 ^ 1'b0 ;
  assign n12835 = n2730 & n4107 ;
  assign n12836 = n4620 & n8910 ;
  assign n12837 = ~n12835 & n12836 ;
  assign n12842 = n11306 ^ n1488 ^ 1'b0 ;
  assign n12843 = n3159 | n12842 ;
  assign n12840 = ( ~n1346 & n7018 ) | ( ~n1346 & n12372 ) | ( n7018 & n12372 ) ;
  assign n12838 = n783 & ~n3187 ;
  assign n12839 = n5136 & n12838 ;
  assign n12841 = n12840 ^ n12839 ^ 1'b0 ;
  assign n12844 = n12843 ^ n12841 ^ 1'b0 ;
  assign n12845 = n12837 | n12844 ;
  assign n12846 = ~n3688 & n9309 ;
  assign n12847 = n12846 ^ n332 ^ 1'b0 ;
  assign n12848 = n355 & ~n12847 ;
  assign n12849 = ~n11171 & n12848 ;
  assign n12850 = n8651 & ~n12849 ;
  assign n12851 = n12393 ^ n11666 ^ 1'b0 ;
  assign n12852 = n9005 ^ n6349 ^ n2205 ;
  assign n12853 = n12852 ^ n10008 ^ n7048 ;
  assign n12854 = n3947 | n10866 ;
  assign n12855 = n12854 ^ n11303 ^ 1'b0 ;
  assign n12856 = n12535 ^ x187 ^ 1'b0 ;
  assign n12857 = n7708 & n12856 ;
  assign n12858 = n2041 & n7655 ;
  assign n12859 = n12858 ^ n4015 ^ 1'b0 ;
  assign n12860 = ( n6809 & n11356 ) | ( n6809 & n12859 ) | ( n11356 & n12859 ) ;
  assign n12861 = n7207 ^ n5357 ^ 1'b0 ;
  assign n12862 = n12861 ^ n764 ^ 1'b0 ;
  assign n12863 = n12862 ^ n11727 ^ 1'b0 ;
  assign n12864 = n10324 | n12863 ;
  assign n12865 = n5848 & ~n7096 ;
  assign n12866 = ~n12864 & n12865 ;
  assign n12867 = ( n5221 & ~n9147 ) | ( n5221 & n11816 ) | ( ~n9147 & n11816 ) ;
  assign n12868 = ( n2830 & n6395 ) | ( n2830 & n12450 ) | ( n6395 & n12450 ) ;
  assign n12869 = n5371 & ~n7216 ;
  assign n12870 = n5877 | n12869 ;
  assign n12871 = n12870 ^ n11817 ^ 1'b0 ;
  assign n12872 = x23 & ~n5949 ;
  assign n12873 = n10183 & n12872 ;
  assign n12874 = ( n1305 & n6468 ) | ( n1305 & n12873 ) | ( n6468 & n12873 ) ;
  assign n12875 = n11972 ^ n2847 ^ 1'b0 ;
  assign n12878 = n1448 & n6390 ;
  assign n12879 = n1673 & n12878 ;
  assign n12876 = n6358 ^ n4156 ^ n2994 ;
  assign n12877 = ~n3587 & n12876 ;
  assign n12880 = n12879 ^ n12877 ^ 1'b0 ;
  assign n12881 = n10176 ^ n5753 ^ n4848 ;
  assign n12882 = ~n1475 & n12881 ;
  assign n12883 = n12882 ^ n289 ^ 1'b0 ;
  assign n12884 = n12883 ^ n1370 ^ 1'b0 ;
  assign n12885 = n408 & ~n7302 ;
  assign n12886 = n2566 & n12885 ;
  assign n12887 = n7983 ^ n7638 ^ n266 ;
  assign n12888 = n12887 ^ n7195 ^ 1'b0 ;
  assign n12895 = n491 & ~n1821 ;
  assign n12896 = n2211 & n12895 ;
  assign n12897 = n4085 & n12896 ;
  assign n12898 = n3509 & ~n12897 ;
  assign n12899 = n12898 ^ n5480 ^ 1'b0 ;
  assign n12900 = n12899 ^ n4251 ^ 1'b0 ;
  assign n12901 = n1010 & n12900 ;
  assign n12902 = n12901 ^ n8931 ^ n8769 ;
  assign n12889 = n9625 ^ n5102 ^ n358 ;
  assign n12890 = n3562 ^ n3448 ^ 1'b0 ;
  assign n12891 = n2514 | n12890 ;
  assign n12892 = n1351 | n12891 ;
  assign n12893 = n1854 | n12892 ;
  assign n12894 = ( ~n1822 & n12889 ) | ( ~n1822 & n12893 ) | ( n12889 & n12893 ) ;
  assign n12903 = n12902 ^ n12894 ^ n10519 ;
  assign n12904 = ( n331 & n5587 ) | ( n331 & n7068 ) | ( n5587 & n7068 ) ;
  assign n12905 = n12247 & n12904 ;
  assign n12908 = n1932 & n9331 ;
  assign n12906 = n5795 ^ n3928 ^ n634 ;
  assign n12907 = n12906 ^ n10017 ^ n8369 ;
  assign n12909 = n12908 ^ n12907 ^ 1'b0 ;
  assign n12910 = n2764 | n8845 ;
  assign n12911 = n12910 ^ n11607 ^ 1'b0 ;
  assign n12912 = n3503 & n12911 ;
  assign n12913 = n1281 ^ n541 ^ 1'b0 ;
  assign n12914 = n12053 ^ n6173 ^ n702 ;
  assign n12915 = n12914 ^ n4107 ^ n649 ;
  assign n12916 = n3973 & n12915 ;
  assign n12917 = n10387 & n12916 ;
  assign n12918 = n5082 & ~n5633 ;
  assign n12919 = ~n8437 & n12918 ;
  assign n12920 = n4323 | n9304 ;
  assign n12921 = n2972 & ~n12920 ;
  assign n12922 = ( n2538 & n4835 ) | ( n2538 & n12921 ) | ( n4835 & n12921 ) ;
  assign n12923 = ~n12919 & n12922 ;
  assign n12924 = n11691 & n12923 ;
  assign n12927 = n2287 & ~n9555 ;
  assign n12925 = ~n1297 & n8165 ;
  assign n12926 = n10464 & n12925 ;
  assign n12928 = n12927 ^ n12926 ^ 1'b0 ;
  assign n12932 = n2569 ^ x82 ^ 1'b0 ;
  assign n12933 = n9344 & ~n12932 ;
  assign n12931 = n11800 ^ n736 ^ n483 ;
  assign n12929 = n9113 ^ n6659 ^ n1289 ;
  assign n12930 = n795 | n12929 ;
  assign n12934 = n12933 ^ n12931 ^ n12930 ;
  assign n12935 = n9789 ^ n3054 ^ 1'b0 ;
  assign n12936 = ( n7926 & ~n11039 ) | ( n7926 & n12935 ) | ( ~n11039 & n12935 ) ;
  assign n12937 = ( n521 & ~n1948 ) | ( n521 & n4457 ) | ( ~n1948 & n4457 ) ;
  assign n12938 = n12937 ^ n11461 ^ 1'b0 ;
  assign n12939 = n1861 & ~n11251 ;
  assign n12940 = ( n1098 & ~n8362 ) | ( n1098 & n8740 ) | ( ~n8362 & n8740 ) ;
  assign n12941 = ( ~n4753 & n6225 ) | ( ~n4753 & n8366 ) | ( n6225 & n8366 ) ;
  assign n12942 = n12941 ^ n4571 ^ 1'b0 ;
  assign n12943 = n12940 | n12942 ;
  assign n12945 = n10169 | n10239 ;
  assign n12946 = n12945 ^ n5669 ^ 1'b0 ;
  assign n12944 = ~n1978 & n9556 ;
  assign n12947 = n12946 ^ n12944 ^ 1'b0 ;
  assign n12948 = ( x225 & ~n9855 ) | ( x225 & n9984 ) | ( ~n9855 & n9984 ) ;
  assign n12951 = ~n2768 & n9043 ;
  assign n12952 = ~n9015 & n12951 ;
  assign n12949 = n7149 & n8688 ;
  assign n12950 = n12949 ^ n9247 ^ 1'b0 ;
  assign n12953 = n12952 ^ n12950 ^ n5873 ;
  assign n12954 = ( ~n1589 & n1830 ) | ( ~n1589 & n1938 ) | ( n1830 & n1938 ) ;
  assign n12957 = x88 | n1771 ;
  assign n12956 = ~n1064 & n5085 ;
  assign n12958 = n12957 ^ n12956 ^ 1'b0 ;
  assign n12955 = ( n5029 & ~n6620 ) | ( n5029 & n11564 ) | ( ~n6620 & n11564 ) ;
  assign n12959 = n12958 ^ n12955 ^ 1'b0 ;
  assign n12960 = ( n3285 & n4436 ) | ( n3285 & n8108 ) | ( n4436 & n8108 ) ;
  assign n12961 = n8659 ^ n7511 ^ 1'b0 ;
  assign n12962 = n12960 | n12961 ;
  assign n12963 = n9802 ^ n6986 ^ 1'b0 ;
  assign n12964 = n4724 & ~n9086 ;
  assign n12965 = ~n12963 & n12964 ;
  assign n12966 = n777 | n3281 ;
  assign n12967 = n12966 ^ n11146 ^ 1'b0 ;
  assign n12968 = n12967 ^ n2364 ^ 1'b0 ;
  assign n12969 = ~n10606 & n12968 ;
  assign n12970 = n6938 ^ n3100 ^ 1'b0 ;
  assign n12971 = n9473 ^ n3507 ^ x43 ;
  assign n12972 = n12971 ^ n1448 ^ 1'b0 ;
  assign n12973 = n11166 ^ n6883 ^ 1'b0 ;
  assign n12974 = ( n2945 & ~n3542 ) | ( n2945 & n6369 ) | ( ~n3542 & n6369 ) ;
  assign n12975 = n12974 ^ n5235 ^ 1'b0 ;
  assign n12976 = n12973 & n12975 ;
  assign n12977 = n692 | n8483 ;
  assign n12978 = ( n2840 & n6269 ) | ( n2840 & ~n12977 ) | ( n6269 & ~n12977 ) ;
  assign n12979 = n9663 ^ n4066 ^ 1'b0 ;
  assign n12980 = ~n12978 & n12979 ;
  assign n12981 = n12976 & n12980 ;
  assign n12983 = n5763 | n6019 ;
  assign n12984 = n12983 ^ n10802 ^ 1'b0 ;
  assign n12982 = n6557 & ~n11387 ;
  assign n12985 = n12984 ^ n12982 ^ 1'b0 ;
  assign n12986 = ~n3616 & n5070 ;
  assign n12987 = n3191 & n5445 ;
  assign n12988 = n12986 & n12987 ;
  assign n12989 = ( ~n4442 & n10499 ) | ( ~n4442 & n12502 ) | ( n10499 & n12502 ) ;
  assign n12990 = n12989 ^ n6716 ^ n6121 ;
  assign n12991 = ( x232 & n2697 ) | ( x232 & n2709 ) | ( n2697 & n2709 ) ;
  assign n12992 = n7260 ^ n5585 ^ n2277 ;
  assign n12993 = ( n1046 & ~n9661 ) | ( n1046 & n12992 ) | ( ~n9661 & n12992 ) ;
  assign n12994 = ~n12991 & n12993 ;
  assign n12995 = n12994 ^ n11348 ^ 1'b0 ;
  assign n12996 = n12121 ^ n12113 ^ n8667 ;
  assign n12997 = ( ~n6073 & n8422 ) | ( ~n6073 & n12996 ) | ( n8422 & n12996 ) ;
  assign n12998 = ( n12990 & n12995 ) | ( n12990 & ~n12997 ) | ( n12995 & ~n12997 ) ;
  assign n12999 = n1714 & n12628 ;
  assign n13000 = n7415 ^ n5695 ^ n1337 ;
  assign n13001 = n6486 ^ n1907 ^ x32 ;
  assign n13002 = ( n4859 & ~n12991 ) | ( n4859 & n13001 ) | ( ~n12991 & n13001 ) ;
  assign n13003 = n13000 | n13002 ;
  assign n13004 = n2651 & ~n7061 ;
  assign n13005 = n6955 & n13004 ;
  assign n13006 = n13005 ^ n2100 ^ 1'b0 ;
  assign n13007 = n5408 & n13006 ;
  assign n13008 = n10130 ^ n8292 ^ 1'b0 ;
  assign n13009 = n6977 | n13008 ;
  assign n13010 = ( ~n4153 & n4421 ) | ( ~n4153 & n13009 ) | ( n4421 & n13009 ) ;
  assign n13011 = n11521 ^ n9959 ^ n7375 ;
  assign n13012 = ( ~x210 & n4251 ) | ( ~x210 & n8408 ) | ( n4251 & n8408 ) ;
  assign n13013 = n11089 ^ n9701 ^ 1'b0 ;
  assign n13014 = n13012 | n13013 ;
  assign n13015 = ~n10062 & n13014 ;
  assign n13016 = n8740 ^ n8088 ^ 1'b0 ;
  assign n13017 = n10121 ^ n6718 ^ 1'b0 ;
  assign n13018 = n13017 ^ n10197 ^ 1'b0 ;
  assign n13029 = n9947 ^ n1136 ^ 1'b0 ;
  assign n13030 = n7928 & n13029 ;
  assign n13027 = n12069 ^ n2878 ^ 1'b0 ;
  assign n13028 = n13027 ^ n10770 ^ 1'b0 ;
  assign n13031 = n13030 ^ n13028 ^ 1'b0 ;
  assign n13032 = n1088 & n13031 ;
  assign n13019 = ( n732 & ~n4219 ) | ( n732 & n9232 ) | ( ~n4219 & n9232 ) ;
  assign n13020 = ( n4933 & n6369 ) | ( n4933 & n13019 ) | ( n6369 & n13019 ) ;
  assign n13021 = n10386 | n13020 ;
  assign n13022 = n4268 ^ n1616 ^ n578 ;
  assign n13023 = n13022 ^ n7555 ^ 1'b0 ;
  assign n13024 = n12869 ^ n11811 ^ n5238 ;
  assign n13025 = ( ~n10226 & n13023 ) | ( ~n10226 & n13024 ) | ( n13023 & n13024 ) ;
  assign n13026 = ~n13021 & n13025 ;
  assign n13033 = n13032 ^ n13026 ^ 1'b0 ;
  assign n13034 = n7612 ^ n7523 ^ 1'b0 ;
  assign n13035 = n9767 & n9789 ;
  assign n13036 = n13035 ^ n5049 ^ 1'b0 ;
  assign n13037 = n13034 & n13036 ;
  assign n13038 = n13037 ^ n8853 ^ 1'b0 ;
  assign n13039 = ( ~x133 & x238 ) | ( ~x133 & n3643 ) | ( x238 & n3643 ) ;
  assign n13040 = ~n1475 & n13039 ;
  assign n13041 = n13040 ^ n731 ^ 1'b0 ;
  assign n13042 = ( ~n1487 & n3874 ) | ( ~n1487 & n6608 ) | ( n3874 & n6608 ) ;
  assign n13043 = ( n9312 & ~n10042 ) | ( n9312 & n13042 ) | ( ~n10042 & n13042 ) ;
  assign n13044 = n13043 ^ n2548 ^ 1'b0 ;
  assign n13045 = n13044 ^ n12260 ^ 1'b0 ;
  assign n13046 = ( n1449 & n1557 ) | ( n1449 & n3131 ) | ( n1557 & n3131 ) ;
  assign n13047 = x163 & n2998 ;
  assign n13048 = n8289 & n13047 ;
  assign n13049 = n3504 | n13048 ;
  assign n13050 = n692 | n13049 ;
  assign n13051 = n13050 ^ n2051 ^ 1'b0 ;
  assign n13052 = ( n9982 & n13046 ) | ( n9982 & ~n13051 ) | ( n13046 & ~n13051 ) ;
  assign n13053 = n7537 ^ n3485 ^ 1'b0 ;
  assign n13054 = ~n5352 & n13053 ;
  assign n13055 = n13054 ^ n8337 ^ 1'b0 ;
  assign n13056 = ( n7166 & n11117 ) | ( n7166 & n12819 ) | ( n11117 & n12819 ) ;
  assign n13057 = ( n652 & ~n4870 ) | ( n652 & n13056 ) | ( ~n4870 & n13056 ) ;
  assign n13058 = x48 & n13057 ;
  assign n13059 = n13055 & n13058 ;
  assign n13060 = n4928 & ~n13059 ;
  assign n13061 = ~n9295 & n13060 ;
  assign n13062 = n13052 & ~n13061 ;
  assign n13063 = ~n9620 & n12955 ;
  assign n13064 = ~n4532 & n13063 ;
  assign n13065 = ( n1024 & n2725 ) | ( n1024 & n11103 ) | ( n2725 & n11103 ) ;
  assign n13066 = ( n431 & n1985 ) | ( n431 & ~n13065 ) | ( n1985 & ~n13065 ) ;
  assign n13067 = n1421 & n1458 ;
  assign n13068 = ~n5664 & n13067 ;
  assign n13069 = n13068 ^ n3309 ^ 1'b0 ;
  assign n13070 = ~n13066 & n13069 ;
  assign n13071 = n12021 & ~n13070 ;
  assign n13075 = n3671 ^ n3033 ^ 1'b0 ;
  assign n13076 = n13075 ^ n7447 ^ 1'b0 ;
  assign n13072 = n1449 & ~n7731 ;
  assign n13073 = n13072 ^ n8743 ^ 1'b0 ;
  assign n13074 = ( n2234 & n7379 ) | ( n2234 & ~n13073 ) | ( n7379 & ~n13073 ) ;
  assign n13077 = n13076 ^ n13074 ^ n12306 ;
  assign n13078 = n10714 ^ n9526 ^ 1'b0 ;
  assign n13079 = n13077 | n13078 ;
  assign n13080 = ( n3449 & ~n6653 ) | ( n3449 & n7651 ) | ( ~n6653 & n7651 ) ;
  assign n13081 = ~n771 & n13080 ;
  assign n13082 = n13081 ^ n3123 ^ 1'b0 ;
  assign n13083 = ~n1066 & n7671 ;
  assign n13084 = n13082 & n13083 ;
  assign n13085 = n13011 ^ n12347 ^ 1'b0 ;
  assign n13086 = n12562 ^ n9129 ^ 1'b0 ;
  assign n13087 = n4414 ^ n976 ^ 1'b0 ;
  assign n13088 = n13086 & ~n13087 ;
  assign n13089 = ( n360 & n12921 ) | ( n360 & ~n13042 ) | ( n12921 & ~n13042 ) ;
  assign n13090 = n5622 & ~n6698 ;
  assign n13091 = n13090 ^ n11129 ^ 1'b0 ;
  assign n13100 = n5675 ^ n4066 ^ 1'b0 ;
  assign n13101 = n4821 & n13100 ;
  assign n13099 = n656 & ~n8528 ;
  assign n13102 = n13101 ^ n13099 ^ 1'b0 ;
  assign n13093 = n6006 ^ x216 ^ 1'b0 ;
  assign n13094 = n7949 & n13093 ;
  assign n13092 = n5613 ^ n4175 ^ n3173 ;
  assign n13095 = n13094 ^ n13092 ^ 1'b0 ;
  assign n13096 = n1391 & ~n13095 ;
  assign n13097 = n2719 ^ n2134 ^ 1'b0 ;
  assign n13098 = n13096 & n13097 ;
  assign n13103 = n13102 ^ n13098 ^ 1'b0 ;
  assign n13104 = n291 & n10187 ;
  assign n13105 = ( x105 & n3016 ) | ( x105 & ~n3563 ) | ( n3016 & ~n3563 ) ;
  assign n13106 = n13105 ^ n1921 ^ 1'b0 ;
  assign n13107 = n629 & n13106 ;
  assign n13108 = n11953 ^ n8325 ^ n1480 ;
  assign n13109 = ( n5448 & n13107 ) | ( n5448 & n13108 ) | ( n13107 & n13108 ) ;
  assign n13110 = n11309 ^ n7541 ^ n5438 ;
  assign n13111 = n1301 & n10181 ;
  assign n13112 = n7905 ^ n6718 ^ n3026 ;
  assign n13113 = n13112 ^ n12616 ^ 1'b0 ;
  assign n13114 = ( n1378 & ~n2218 ) | ( n1378 & n7566 ) | ( ~n2218 & n7566 ) ;
  assign n13115 = ~n3147 & n5794 ;
  assign n13116 = n13115 ^ n8399 ^ n2457 ;
  assign n13117 = x131 & n13116 ;
  assign n13118 = n13117 ^ n4747 ^ 1'b0 ;
  assign n13122 = n4770 ^ n2234 ^ n1961 ;
  assign n13119 = ~n3456 & n11041 ;
  assign n13120 = n384 & n13119 ;
  assign n13121 = ~n10427 & n13120 ;
  assign n13123 = n13122 ^ n13121 ^ n3397 ;
  assign n13124 = ~n8405 & n12990 ;
  assign n13125 = n13124 ^ n9881 ^ 1'b0 ;
  assign n13127 = n1261 & ~n10655 ;
  assign n13126 = ~n2226 & n7136 ;
  assign n13128 = n13127 ^ n13126 ^ 1'b0 ;
  assign n13129 = n5070 | n13128 ;
  assign n13130 = n680 | n10824 ;
  assign n13131 = n3502 | n5291 ;
  assign n13132 = n9798 ^ n5387 ^ 1'b0 ;
  assign n13133 = n4570 & n13132 ;
  assign n13134 = n13054 ^ x191 ^ 1'b0 ;
  assign n13135 = n5916 & n13134 ;
  assign n13136 = n13133 & n13135 ;
  assign n13137 = ~x140 & n13136 ;
  assign n13138 = n4934 ^ n841 ^ 1'b0 ;
  assign n13139 = n8517 ^ n4248 ^ 1'b0 ;
  assign n13140 = ~n3245 & n7658 ;
  assign n13141 = n13140 ^ n2876 ^ 1'b0 ;
  assign n13142 = n10076 ^ n3556 ^ 1'b0 ;
  assign n13143 = n13141 & n13142 ;
  assign n13145 = ( n1793 & n4257 ) | ( n1793 & n7949 ) | ( n4257 & n7949 ) ;
  assign n13144 = n12899 ^ n4873 ^ 1'b0 ;
  assign n13146 = n13145 ^ n13144 ^ n755 ;
  assign n13147 = ( n481 & n964 ) | ( n481 & n966 ) | ( n964 & n966 ) ;
  assign n13148 = n13147 ^ n10165 ^ n1205 ;
  assign n13149 = ( n4529 & ~n7700 ) | ( n4529 & n13148 ) | ( ~n7700 & n13148 ) ;
  assign n13150 = ~n3985 & n13149 ;
  assign n13151 = n12864 ^ n12716 ^ n1124 ;
  assign n13152 = n13151 ^ n8192 ^ 1'b0 ;
  assign n13153 = n1771 | n3008 ;
  assign n13154 = n4968 & ~n13153 ;
  assign n13155 = n13154 ^ n2884 ^ 1'b0 ;
  assign n13156 = n13155 ^ n1130 ^ 1'b0 ;
  assign n13157 = n9724 ^ n8110 ^ n5470 ;
  assign n13159 = n853 & ~n3546 ;
  assign n13160 = ~n2504 & n13159 ;
  assign n13158 = n6384 ^ n391 ^ 1'b0 ;
  assign n13161 = n13160 ^ n13158 ^ 1'b0 ;
  assign n13162 = ~n2934 & n7670 ;
  assign n13163 = n11776 ^ n9432 ^ n3491 ;
  assign n13164 = n9396 & ~n11269 ;
  assign n13165 = ( ~n1545 & n4970 ) | ( ~n1545 & n12815 ) | ( n4970 & n12815 ) ;
  assign n13166 = ~n1130 & n9576 ;
  assign n13167 = n13166 ^ n2203 ^ x40 ;
  assign n13168 = n10968 ^ n4119 ^ n3166 ;
  assign n13169 = n13168 ^ n10074 ^ n3340 ;
  assign n13170 = n13167 & n13169 ;
  assign n13172 = n1433 ^ n1149 ^ 1'b0 ;
  assign n13173 = x7 & n13172 ;
  assign n13174 = ~n9111 & n13173 ;
  assign n13175 = n13174 ^ n3653 ^ 1'b0 ;
  assign n13171 = n4601 & n5748 ;
  assign n13176 = n13175 ^ n13171 ^ 1'b0 ;
  assign n13177 = n2226 | n8880 ;
  assign n13178 = n3214 ^ n995 ^ 1'b0 ;
  assign n13179 = n13177 & ~n13178 ;
  assign n13180 = n13179 ^ n9180 ^ n967 ;
  assign n13181 = n8405 ^ n4053 ^ n2643 ;
  assign n13182 = n12380 ^ n725 ^ 1'b0 ;
  assign n13183 = n4167 | n13182 ;
  assign n13184 = n10384 & ~n13183 ;
  assign n13185 = n2244 & n13184 ;
  assign n13186 = ( ~n5537 & n13181 ) | ( ~n5537 & n13185 ) | ( n13181 & n13185 ) ;
  assign n13187 = n2119 | n2794 ;
  assign n13188 = n13187 ^ n7413 ^ n6061 ;
  assign n13189 = ~n1246 & n1968 ;
  assign n13190 = n13189 ^ n2168 ^ 1'b0 ;
  assign n13191 = n12700 ^ n4409 ^ n2596 ;
  assign n13192 = ( ~n12384 & n13190 ) | ( ~n12384 & n13191 ) | ( n13190 & n13191 ) ;
  assign n13193 = n3018 & n6786 ;
  assign n13194 = n13193 ^ n12530 ^ 1'b0 ;
  assign n13195 = n13194 ^ n7168 ^ 1'b0 ;
  assign n13196 = n10339 ^ n9394 ^ 1'b0 ;
  assign n13197 = ( n941 & n1745 ) | ( n941 & ~n11841 ) | ( n1745 & ~n11841 ) ;
  assign n13198 = n13197 ^ n5639 ^ 1'b0 ;
  assign n13199 = n10939 & ~n13198 ;
  assign n13200 = ( ~n1045 & n7343 ) | ( ~n1045 & n9678 ) | ( n7343 & n9678 ) ;
  assign n13201 = n13200 ^ n673 ^ 1'b0 ;
  assign n13202 = n5132 ^ n780 ^ 1'b0 ;
  assign n13203 = ~n2126 & n13202 ;
  assign n13204 = n12177 ^ n9003 ^ n5343 ;
  assign n13205 = n11469 & ~n13204 ;
  assign n13206 = n2903 | n13205 ;
  assign n13207 = n6220 | n12773 ;
  assign n13208 = n1440 | n9855 ;
  assign n13209 = n13208 ^ n12280 ^ n1090 ;
  assign n13210 = x179 & n2752 ;
  assign n13211 = n2376 & n13210 ;
  assign n13212 = ( ~n7717 & n12472 ) | ( ~n7717 & n13211 ) | ( n12472 & n13211 ) ;
  assign n13213 = ~n4108 & n8574 ;
  assign n13214 = n281 & n13213 ;
  assign n13215 = n4187 & ~n9069 ;
  assign n13216 = n13215 ^ n11453 ^ 1'b0 ;
  assign n13217 = ( n10095 & ~n10152 ) | ( n10095 & n11977 ) | ( ~n10152 & n11977 ) ;
  assign n13218 = ( n6718 & n13216 ) | ( n6718 & ~n13217 ) | ( n13216 & ~n13217 ) ;
  assign n13219 = ( n2688 & n9191 ) | ( n2688 & ~n10896 ) | ( n9191 & ~n10896 ) ;
  assign n13220 = n12480 ^ n4484 ^ n1683 ;
  assign n13221 = n13220 ^ n6628 ^ 1'b0 ;
  assign n13222 = n4322 & n13221 ;
  assign n13223 = ~n5097 & n5953 ;
  assign n13224 = n6341 & ~n10745 ;
  assign n13225 = ~n13223 & n13224 ;
  assign n13226 = n5733 ^ n3919 ^ x114 ;
  assign n13227 = ( ~n1475 & n2947 ) | ( ~n1475 & n3958 ) | ( n2947 & n3958 ) ;
  assign n13228 = n13227 ^ n3228 ^ n971 ;
  assign n13229 = ( n1199 & ~n3450 ) | ( n1199 & n13228 ) | ( ~n3450 & n13228 ) ;
  assign n13230 = ~n13226 & n13229 ;
  assign n13231 = n12254 & n13230 ;
  assign n13232 = n7194 ^ n4106 ^ x166 ;
  assign n13233 = n13232 ^ n12556 ^ n750 ;
  assign n13234 = n13233 ^ n6129 ^ n5500 ;
  assign n13235 = n2750 ^ n2301 ^ 1'b0 ;
  assign n13236 = n4239 & n13235 ;
  assign n13237 = n13236 ^ n6047 ^ 1'b0 ;
  assign n13238 = n5234 ^ n5118 ^ 1'b0 ;
  assign n13239 = n13238 ^ n3169 ^ 1'b0 ;
  assign n13240 = n13237 | n13239 ;
  assign n13241 = n7306 ^ n4401 ^ 1'b0 ;
  assign n13242 = ( n2376 & ~n6937 ) | ( n2376 & n13241 ) | ( ~n6937 & n13241 ) ;
  assign n13243 = n7102 | n9514 ;
  assign n13244 = n1236 & ~n13243 ;
  assign n13245 = ( ~x46 & n3094 ) | ( ~x46 & n13244 ) | ( n3094 & n13244 ) ;
  assign n13246 = ( n2977 & n13242 ) | ( n2977 & n13245 ) | ( n13242 & n13245 ) ;
  assign n13255 = n6138 ^ n3713 ^ 1'b0 ;
  assign n13256 = ( n5486 & n12627 ) | ( n5486 & ~n13255 ) | ( n12627 & ~n13255 ) ;
  assign n13257 = n13256 ^ n3118 ^ n2263 ;
  assign n13247 = n7492 ^ n4332 ^ 1'b0 ;
  assign n13248 = ~n4796 & n13247 ;
  assign n13249 = ( n313 & n1221 ) | ( n313 & ~n1959 ) | ( n1221 & ~n1959 ) ;
  assign n13250 = ( ~n2949 & n5744 ) | ( ~n2949 & n13249 ) | ( n5744 & n13249 ) ;
  assign n13251 = ( x82 & ~n10906 ) | ( x82 & n13250 ) | ( ~n10906 & n13250 ) ;
  assign n13252 = ( ~x63 & n13248 ) | ( ~x63 & n13251 ) | ( n13248 & n13251 ) ;
  assign n13253 = n4777 & ~n13252 ;
  assign n13254 = n13253 ^ n2301 ^ 1'b0 ;
  assign n13258 = n13257 ^ n13254 ^ n13155 ;
  assign n13259 = ~x182 & n1145 ;
  assign n13262 = ( n1140 & n2132 ) | ( n1140 & ~n5850 ) | ( n2132 & ~n5850 ) ;
  assign n13263 = n13262 ^ n7679 ^ 1'b0 ;
  assign n13260 = n4691 ^ n2357 ^ x56 ;
  assign n13261 = n1883 | n13260 ;
  assign n13264 = n13263 ^ n13261 ^ 1'b0 ;
  assign n13265 = n13264 ^ n4730 ^ 1'b0 ;
  assign n13266 = ~n715 & n13265 ;
  assign n13267 = n11484 ^ n6003 ^ 1'b0 ;
  assign n13268 = ~n8573 & n13267 ;
  assign n13272 = x180 & ~n3937 ;
  assign n13269 = n4684 & ~n9005 ;
  assign n13270 = n1717 & n13269 ;
  assign n13271 = ~n1923 & n13270 ;
  assign n13273 = n13272 ^ n13271 ^ n10841 ;
  assign n13274 = ( n2403 & n2858 ) | ( n2403 & ~n6133 ) | ( n2858 & ~n6133 ) ;
  assign n13275 = n12900 & ~n13274 ;
  assign n13276 = ~x109 & n13275 ;
  assign n13277 = n13276 ^ n10527 ^ n1900 ;
  assign n13278 = n2859 | n6360 ;
  assign n13279 = ( ~n4278 & n4301 ) | ( ~n4278 & n12210 ) | ( n4301 & n12210 ) ;
  assign n13280 = n13279 ^ n8763 ^ 1'b0 ;
  assign n13281 = n12549 | n13280 ;
  assign n13282 = n7429 ^ n6433 ^ n2401 ;
  assign n13283 = n13282 ^ n1978 ^ 1'b0 ;
  assign n13284 = n8355 | n13283 ;
  assign n13285 = n1122 & ~n13284 ;
  assign n13286 = ( n13278 & n13281 ) | ( n13278 & ~n13285 ) | ( n13281 & ~n13285 ) ;
  assign n13287 = n13286 ^ n4618 ^ 1'b0 ;
  assign n13288 = ~n631 & n4359 ;
  assign n13289 = ( n1290 & n6771 ) | ( n1290 & ~n13288 ) | ( n6771 & ~n13288 ) ;
  assign n13290 = n13289 ^ n8697 ^ n7840 ;
  assign n13292 = n766 & ~n11536 ;
  assign n13293 = n13292 ^ n2394 ^ 1'b0 ;
  assign n13291 = ( ~n2774 & n4787 ) | ( ~n2774 & n7411 ) | ( n4787 & n7411 ) ;
  assign n13294 = n13293 ^ n13291 ^ n8240 ;
  assign n13295 = n3186 & n11121 ;
  assign n13296 = x56 & ~n13295 ;
  assign n13297 = n13296 ^ n7828 ^ n3586 ;
  assign n13298 = n10546 ^ n3520 ^ 1'b0 ;
  assign n13299 = n6697 & n13298 ;
  assign n13300 = n10918 ^ n3744 ^ 1'b0 ;
  assign n13301 = n2950 & n13300 ;
  assign n13302 = x120 & n2182 ;
  assign n13303 = n13302 ^ n2437 ^ 1'b0 ;
  assign n13304 = n9691 ^ n3061 ^ 1'b0 ;
  assign n13305 = n13303 & n13304 ;
  assign n13308 = ( ~n4323 & n8880 ) | ( ~n4323 & n9024 ) | ( n8880 & n9024 ) ;
  assign n13307 = ( ~n1879 & n5202 ) | ( ~n1879 & n9219 ) | ( n5202 & n9219 ) ;
  assign n13309 = n13308 ^ n13307 ^ n1352 ;
  assign n13306 = n4671 | n4935 ;
  assign n13310 = n13309 ^ n13306 ^ n1411 ;
  assign n13311 = n11560 & ~n13310 ;
  assign n13312 = ~n13305 & n13311 ;
  assign n13313 = n13301 & n13312 ;
  assign n13314 = n9223 ^ n2308 ^ 1'b0 ;
  assign n13315 = n7696 ^ n5112 ^ n5073 ;
  assign n13316 = ( ~n10093 & n13314 ) | ( ~n10093 & n13315 ) | ( n13314 & n13315 ) ;
  assign n13317 = ( ~n3954 & n6334 ) | ( ~n3954 & n6681 ) | ( n6334 & n6681 ) ;
  assign n13318 = ~n8460 & n13317 ;
  assign n13319 = n13318 ^ n7984 ^ 1'b0 ;
  assign n13320 = n13319 ^ n10028 ^ 1'b0 ;
  assign n13321 = n13316 | n13320 ;
  assign n13322 = ~n11563 & n13321 ;
  assign n13323 = n12937 ^ n11734 ^ n2697 ;
  assign n13324 = n388 | n8340 ;
  assign n13325 = n6520 ^ n2686 ^ 1'b0 ;
  assign n13326 = n12348 & ~n13325 ;
  assign n13327 = ( n4875 & ~n10052 ) | ( n4875 & n13326 ) | ( ~n10052 & n13326 ) ;
  assign n13328 = n1983 ^ x212 ^ 1'b0 ;
  assign n13329 = x105 & ~n13252 ;
  assign n13330 = n13329 ^ n12900 ^ 1'b0 ;
  assign n13331 = n13330 ^ n5945 ^ 1'b0 ;
  assign n13332 = n13331 ^ n9616 ^ 1'b0 ;
  assign n13337 = n3393 | n12075 ;
  assign n13334 = n8369 ^ n4821 ^ n3206 ;
  assign n13333 = ~n899 & n9143 ;
  assign n13335 = n13334 ^ n13333 ^ 1'b0 ;
  assign n13336 = n13335 ^ n11144 ^ n1116 ;
  assign n13338 = n13337 ^ n13336 ^ n3178 ;
  assign n13339 = n5392 ^ n2943 ^ 1'b0 ;
  assign n13340 = n13339 ^ n11631 ^ n430 ;
  assign n13341 = n3792 | n6906 ;
  assign n13342 = ( ~n855 & n3063 ) | ( ~n855 & n13341 ) | ( n3063 & n13341 ) ;
  assign n13343 = ~n6125 & n13342 ;
  assign n13344 = n5042 & n13343 ;
  assign n13345 = ( n276 & n2450 ) | ( n276 & n5497 ) | ( n2450 & n5497 ) ;
  assign n13346 = n2828 & ~n13345 ;
  assign n13347 = n12593 & n13346 ;
  assign n13348 = n2509 | n13347 ;
  assign n13349 = n2884 & ~n13348 ;
  assign n13351 = n1267 | n5022 ;
  assign n13350 = n2234 & ~n9354 ;
  assign n13352 = n13351 ^ n13350 ^ 1'b0 ;
  assign n13358 = n2825 & n8555 ;
  assign n13353 = n3718 ^ n3663 ^ 1'b0 ;
  assign n13354 = ~n3817 & n13353 ;
  assign n13355 = ~n841 & n1398 ;
  assign n13356 = ~n13354 & n13355 ;
  assign n13357 = n5275 & ~n13356 ;
  assign n13359 = n13358 ^ n13357 ^ 1'b0 ;
  assign n13362 = n683 | n9220 ;
  assign n13363 = n626 | n13362 ;
  assign n13360 = n5767 ^ n3966 ^ 1'b0 ;
  assign n13361 = n10036 & n13360 ;
  assign n13364 = n13363 ^ n13361 ^ n12651 ;
  assign n13365 = n1024 | n8070 ;
  assign n13368 = ( n1124 & n5459 ) | ( n1124 & ~n11696 ) | ( n5459 & ~n11696 ) ;
  assign n13366 = n1346 | n11825 ;
  assign n13367 = n13366 ^ n698 ^ 1'b0 ;
  assign n13369 = n13368 ^ n13367 ^ n11831 ;
  assign n13370 = n8294 ^ n1624 ^ 1'b0 ;
  assign n13371 = n12524 | n13370 ;
  assign n13372 = n2365 & n4910 ;
  assign n13373 = n13372 ^ n2947 ^ 1'b0 ;
  assign n13375 = n4921 & n8477 ;
  assign n13374 = n2845 & ~n7395 ;
  assign n13376 = n13375 ^ n13374 ^ 1'b0 ;
  assign n13377 = ( n1039 & n4308 ) | ( n1039 & ~n13376 ) | ( n4308 & ~n13376 ) ;
  assign n13378 = n6174 ^ n5710 ^ 1'b0 ;
  assign n13379 = ~n5981 & n13378 ;
  assign n13380 = n1095 | n13379 ;
  assign n13381 = n9986 & n13380 ;
  assign n13382 = n13381 ^ n11560 ^ 1'b0 ;
  assign n13386 = n632 & ~n3280 ;
  assign n13384 = n5302 ^ n1476 ^ 1'b0 ;
  assign n13385 = n561 & ~n13384 ;
  assign n13383 = n2574 & ~n6273 ;
  assign n13387 = n13386 ^ n13385 ^ n13383 ;
  assign n13388 = n8529 ^ n7411 ^ n1109 ;
  assign n13389 = n6258 & n13388 ;
  assign n13390 = ~n8247 & n13389 ;
  assign n13391 = n4819 | n13390 ;
  assign n13392 = n1588 | n9151 ;
  assign n13393 = n3957 | n13392 ;
  assign n13394 = n4270 ^ n1130 ^ 1'b0 ;
  assign n13395 = n5136 & ~n7484 ;
  assign n13396 = n13395 ^ n3065 ^ 1'b0 ;
  assign n13397 = ~n2213 & n13396 ;
  assign n13398 = n13397 ^ n12861 ^ 1'b0 ;
  assign n13399 = ~n812 & n13398 ;
  assign n13400 = ~n13394 & n13399 ;
  assign n13401 = n2227 & ~n13400 ;
  assign n13402 = n6629 ^ n3779 ^ 1'b0 ;
  assign n13403 = n793 | n2357 ;
  assign n13404 = n13403 ^ n8620 ^ 1'b0 ;
  assign n13405 = n1244 & ~n9049 ;
  assign n13406 = n13405 ^ n553 ^ n353 ;
  assign n13407 = n12849 ^ n3598 ^ 1'b0 ;
  assign n13408 = ~n8637 & n13407 ;
  assign n13409 = n13408 ^ n910 ^ 1'b0 ;
  assign n13410 = ~n4153 & n13409 ;
  assign n13411 = n13406 & n13410 ;
  assign n13412 = n13411 ^ n8705 ^ 1'b0 ;
  assign n13413 = n9339 | n9449 ;
  assign n13414 = n13412 | n13413 ;
  assign n13415 = ( n2021 & n2626 ) | ( n2021 & n7842 ) | ( n2626 & n7842 ) ;
  assign n13416 = n13415 ^ n8495 ^ n7984 ;
  assign n13417 = ~n6570 & n13416 ;
  assign n13418 = ( n1042 & n2788 ) | ( n1042 & ~n7243 ) | ( n2788 & ~n7243 ) ;
  assign n13419 = n7146 ^ n3026 ^ x114 ;
  assign n13420 = n13419 ^ n6340 ^ n5316 ;
  assign n13421 = n13418 | n13420 ;
  assign n13422 = n12665 | n13421 ;
  assign n13423 = ~n1768 & n2628 ;
  assign n13424 = n3004 ^ n2571 ^ 1'b0 ;
  assign n13425 = ( ~n6551 & n13423 ) | ( ~n6551 & n13424 ) | ( n13423 & n13424 ) ;
  assign n13426 = n13127 ^ n4671 ^ 1'b0 ;
  assign n13427 = ~n7921 & n13426 ;
  assign n13431 = n6960 ^ n4129 ^ n3094 ;
  assign n13428 = ~n7107 & n11507 ;
  assign n13429 = n13428 ^ n5679 ^ 1'b0 ;
  assign n13430 = n11373 | n13429 ;
  assign n13432 = n13431 ^ n13430 ^ n6152 ;
  assign n13433 = ( n4932 & n5357 ) | ( n4932 & n9631 ) | ( n5357 & n9631 ) ;
  assign n13434 = n13433 ^ n13207 ^ 1'b0 ;
  assign n13435 = n1098 | n5853 ;
  assign n13436 = n13435 ^ n10445 ^ n3787 ;
  assign n13437 = x160 & ~n3165 ;
  assign n13438 = n10267 & n13437 ;
  assign n13439 = n5874 & n7834 ;
  assign n13440 = n5549 & n13439 ;
  assign n13441 = n13438 & n13440 ;
  assign n13442 = n9632 & ~n10245 ;
  assign n13443 = n13442 ^ n277 ^ 1'b0 ;
  assign n13444 = n13441 & ~n13443 ;
  assign n13445 = n5697 & n10050 ;
  assign n13446 = n11646 ^ n5567 ^ n3219 ;
  assign n13447 = ( n5271 & n6358 ) | ( n5271 & ~n13446 ) | ( n6358 & ~n13446 ) ;
  assign n13448 = n5910 & ~n13447 ;
  assign n13449 = n11650 ^ n7241 ^ 1'b0 ;
  assign n13450 = ( ~n4841 & n5452 ) | ( ~n4841 & n8730 ) | ( n5452 & n8730 ) ;
  assign n13451 = ~n962 & n13450 ;
  assign n13452 = n13451 ^ n5011 ^ 1'b0 ;
  assign n13453 = x60 & ~n13452 ;
  assign n13454 = n617 & n13453 ;
  assign n13462 = n7104 ^ n3075 ^ x97 ;
  assign n13458 = n4001 & ~n5816 ;
  assign n13459 = n13458 ^ n4064 ^ 1'b0 ;
  assign n13456 = n4390 ^ n3125 ^ n2305 ;
  assign n13457 = n13456 ^ n8175 ^ n5320 ;
  assign n13460 = n13459 ^ n13457 ^ x199 ;
  assign n13455 = n997 | n1738 ;
  assign n13461 = n13460 ^ n13455 ^ 1'b0 ;
  assign n13463 = n13462 ^ n13461 ^ n12590 ;
  assign n13464 = n3787 & ~n8453 ;
  assign n13466 = n7086 ^ n5699 ^ n4844 ;
  assign n13465 = x158 & n4349 ;
  assign n13467 = n13466 ^ n13465 ^ 1'b0 ;
  assign n13468 = ( n1036 & n7554 ) | ( n1036 & n13467 ) | ( n7554 & n13467 ) ;
  assign n13469 = n3658 ^ n845 ^ 1'b0 ;
  assign n13470 = n10932 ^ n3785 ^ 1'b0 ;
  assign n13471 = n13469 & ~n13470 ;
  assign n13472 = n13427 & n13471 ;
  assign n13473 = n13472 ^ n12489 ^ 1'b0 ;
  assign n13474 = x237 & ~n10653 ;
  assign n13475 = ~n1776 & n8620 ;
  assign n13476 = n13475 ^ n11185 ^ 1'b0 ;
  assign n13477 = n9881 ^ n1149 ^ 1'b0 ;
  assign n13478 = n4560 ^ x89 ^ 1'b0 ;
  assign n13479 = ( n5816 & ~n13477 ) | ( n5816 & n13478 ) | ( ~n13477 & n13478 ) ;
  assign n13480 = n4796 & ~n4996 ;
  assign n13481 = n7748 ^ n6531 ^ 1'b0 ;
  assign n13482 = ~n13480 & n13481 ;
  assign n13484 = ( n2390 & n2544 ) | ( n2390 & ~n3791 ) | ( n2544 & ~n3791 ) ;
  assign n13485 = n13484 ^ n4284 ^ 1'b0 ;
  assign n13486 = ~n5112 & n13485 ;
  assign n13483 = n3026 & n3147 ;
  assign n13487 = n13486 ^ n13483 ^ 1'b0 ;
  assign n13488 = n9596 ^ n5176 ^ 1'b0 ;
  assign n13489 = ~n2178 & n3493 ;
  assign n13490 = n13489 ^ n1501 ^ 1'b0 ;
  assign n13491 = n13490 ^ n4509 ^ 1'b0 ;
  assign n13492 = n2851 | n13491 ;
  assign n13493 = ~n2667 & n8470 ;
  assign n13494 = ~n13492 & n13493 ;
  assign n13495 = n13494 ^ n11644 ^ n11032 ;
  assign n13496 = n5276 ^ n4662 ^ x45 ;
  assign n13497 = n3279 ^ n1012 ^ n447 ;
  assign n13498 = n995 & ~n13497 ;
  assign n13499 = n13498 ^ n8772 ^ 1'b0 ;
  assign n13500 = n8348 | n13499 ;
  assign n13501 = n12871 ^ n4041 ^ n3076 ;
  assign n13502 = ~n9018 & n13027 ;
  assign n13503 = n13502 ^ n3016 ^ 1'b0 ;
  assign n13504 = n4046 & n13503 ;
  assign n13505 = n6441 & n13504 ;
  assign n13506 = ( n1743 & ~n4318 ) | ( n1743 & n5169 ) | ( ~n4318 & n5169 ) ;
  assign n13507 = ~n10492 & n13506 ;
  assign n13508 = ( ~n3214 & n5020 ) | ( ~n3214 & n11019 ) | ( n5020 & n11019 ) ;
  assign n13509 = ( n1864 & ~n5811 ) | ( n1864 & n9964 ) | ( ~n5811 & n9964 ) ;
  assign n13510 = ( x132 & ~n938 ) | ( x132 & n13509 ) | ( ~n938 & n13509 ) ;
  assign n13511 = n10057 | n13510 ;
  assign n13512 = n12280 | n13511 ;
  assign n13513 = n6294 ^ n3941 ^ 1'b0 ;
  assign n13514 = n490 & ~n3818 ;
  assign n13515 = n2026 | n13514 ;
  assign n13516 = n739 | n13515 ;
  assign n13517 = n7260 & n13516 ;
  assign n13518 = ~n9043 & n13517 ;
  assign n13519 = n13518 ^ n2971 ^ 1'b0 ;
  assign n13520 = n11064 & ~n13519 ;
  assign n13522 = n738 & ~n3648 ;
  assign n13523 = ( n3888 & n13250 ) | ( n3888 & ~n13522 ) | ( n13250 & ~n13522 ) ;
  assign n13524 = n13523 ^ n9541 ^ n1554 ;
  assign n13521 = ( n4230 & n7044 ) | ( n4230 & n7353 ) | ( n7044 & n7353 ) ;
  assign n13525 = n13524 ^ n13521 ^ n7410 ;
  assign n13533 = n4579 ^ n1680 ^ 1'b0 ;
  assign n13534 = ~n4917 & n13533 ;
  assign n13535 = n9964 | n12289 ;
  assign n13536 = n13535 ^ n7401 ^ 1'b0 ;
  assign n13537 = n13536 ^ n1873 ^ 1'b0 ;
  assign n13538 = n13534 & n13537 ;
  assign n13539 = n13538 ^ n4807 ^ n2704 ;
  assign n13526 = n1719 | n7334 ;
  assign n13527 = ( ~x143 & n2032 ) | ( ~x143 & n4150 ) | ( n2032 & n4150 ) ;
  assign n13528 = ( n5246 & n5707 ) | ( n5246 & n13527 ) | ( n5707 & n13527 ) ;
  assign n13529 = ( ~n2107 & n5735 ) | ( ~n2107 & n13528 ) | ( n5735 & n13528 ) ;
  assign n13530 = n5720 & ~n13529 ;
  assign n13531 = n13530 ^ n3372 ^ 1'b0 ;
  assign n13532 = n13526 | n13531 ;
  assign n13540 = n13539 ^ n13532 ^ 1'b0 ;
  assign n13543 = n9129 ^ n842 ^ 1'b0 ;
  assign n13544 = n365 & n13543 ;
  assign n13545 = n13544 ^ n6148 ^ n5395 ;
  assign n13541 = ( x103 & n1186 ) | ( x103 & n1859 ) | ( n1186 & n1859 ) ;
  assign n13542 = n4350 & n13541 ;
  assign n13546 = n13545 ^ n13542 ^ 1'b0 ;
  assign n13547 = n2121 ^ n1408 ^ 1'b0 ;
  assign n13548 = x81 | n13547 ;
  assign n13549 = ( ~n1033 & n10645 ) | ( ~n1033 & n13548 ) | ( n10645 & n13548 ) ;
  assign n13550 = n13549 ^ n5521 ^ 1'b0 ;
  assign n13551 = n5571 & ~n13550 ;
  assign n13552 = n11560 ^ n1921 ^ n272 ;
  assign n13553 = ~n6175 & n10679 ;
  assign n13554 = ( n293 & ~n1175 ) | ( n293 & n6047 ) | ( ~n1175 & n6047 ) ;
  assign n13555 = n4505 ^ n3664 ^ 1'b0 ;
  assign n13556 = ~n13554 & n13555 ;
  assign n13557 = n12150 ^ n3903 ^ n3286 ;
  assign n13558 = n13556 & ~n13557 ;
  assign n13559 = n13558 ^ n7689 ^ 1'b0 ;
  assign n13563 = n3056 ^ n1966 ^ n483 ;
  assign n13560 = n8262 & ~n11079 ;
  assign n13561 = n13560 ^ n506 ^ 1'b0 ;
  assign n13562 = n11791 | n13561 ;
  assign n13564 = n13563 ^ n13562 ^ 1'b0 ;
  assign n13565 = n10869 ^ n5559 ^ 1'b0 ;
  assign n13566 = ~n8719 & n13565 ;
  assign n13567 = ( ~n1974 & n8538 ) | ( ~n1974 & n13566 ) | ( n8538 & n13566 ) ;
  assign n13568 = n4937 ^ n3914 ^ n475 ;
  assign n13569 = ( n2247 & ~n12895 ) | ( n2247 & n13568 ) | ( ~n12895 & n13568 ) ;
  assign n13570 = ~n10542 & n13569 ;
  assign n13571 = ( n3012 & ~n3444 ) | ( n3012 & n6682 ) | ( ~n3444 & n6682 ) ;
  assign n13572 = n13571 ^ n9034 ^ 1'b0 ;
  assign n13573 = ( ~n988 & n9111 ) | ( ~n988 & n13522 ) | ( n9111 & n13522 ) ;
  assign n13574 = n13573 ^ n9334 ^ n1431 ;
  assign n13575 = n13574 ^ n7822 ^ 1'b0 ;
  assign n13576 = n13575 ^ n6887 ^ 1'b0 ;
  assign n13577 = n5210 | n13576 ;
  assign n13578 = n6648 & n7315 ;
  assign n13579 = n13578 ^ n5573 ^ 1'b0 ;
  assign n13580 = ~n12157 & n13579 ;
  assign n13581 = n2059 ^ x57 ^ x4 ;
  assign n13582 = n6690 & n13581 ;
  assign n13584 = n4346 ^ x42 ^ 1'b0 ;
  assign n13585 = n6224 & ~n13584 ;
  assign n13586 = n13585 ^ n5723 ^ 1'b0 ;
  assign n13587 = n5514 | n13586 ;
  assign n13588 = ( n11659 & n12705 ) | ( n11659 & n13587 ) | ( n12705 & n13587 ) ;
  assign n13583 = n11845 ^ n566 ^ 1'b0 ;
  assign n13589 = n13588 ^ n13583 ^ n4025 ;
  assign n13590 = ( n8929 & n13582 ) | ( n8929 & ~n13589 ) | ( n13582 & ~n13589 ) ;
  assign n13591 = ( n2637 & n2930 ) | ( n2637 & n4656 ) | ( n2930 & n4656 ) ;
  assign n13592 = n9300 & ~n13591 ;
  assign n13593 = n3177 & n13592 ;
  assign n13594 = ~n330 & n10371 ;
  assign n13595 = ~n13593 & n13594 ;
  assign n13596 = n6567 & n13595 ;
  assign n13597 = n13129 ^ n12300 ^ n2180 ;
  assign n13598 = n5248 ^ n2566 ^ n1075 ;
  assign n13599 = ( n5118 & n11289 ) | ( n5118 & n13598 ) | ( n11289 & n13598 ) ;
  assign n13600 = n13599 ^ n4841 ^ 1'b0 ;
  assign n13601 = ( n2821 & n3031 ) | ( n2821 & n4645 ) | ( n3031 & n4645 ) ;
  assign n13602 = n4749 & n13601 ;
  assign n13603 = n13602 ^ n1601 ^ 1'b0 ;
  assign n13604 = ( n1383 & ~n12544 ) | ( n1383 & n13448 ) | ( ~n12544 & n13448 ) ;
  assign n13605 = ( n3717 & n9769 ) | ( n3717 & ~n12617 ) | ( n9769 & ~n12617 ) ;
  assign n13606 = x34 & n5386 ;
  assign n13607 = ~n13605 & n13606 ;
  assign n13608 = n13015 | n13607 ;
  assign n13609 = n13608 ^ x209 ^ 1'b0 ;
  assign n13610 = n5510 | n10916 ;
  assign n13611 = n5217 | n13610 ;
  assign n13612 = n10327 & ~n13611 ;
  assign n13613 = ( x251 & ~n6557 ) | ( x251 & n8323 ) | ( ~n6557 & n8323 ) ;
  assign n13614 = n13613 ^ n4741 ^ n2722 ;
  assign n13615 = n11075 & n11467 ;
  assign n13616 = n3872 & n13615 ;
  assign n13617 = ( n7225 & n13614 ) | ( n7225 & ~n13616 ) | ( n13614 & ~n13616 ) ;
  assign n13622 = n802 | n4232 ;
  assign n13623 = x142 & n13622 ;
  assign n13624 = n13623 ^ n11453 ^ n4546 ;
  assign n13618 = n5813 | n10065 ;
  assign n13619 = n13618 ^ n9159 ^ 1'b0 ;
  assign n13620 = n1145 & ~n13619 ;
  assign n13621 = n13620 ^ n13305 ^ 1'b0 ;
  assign n13625 = n13624 ^ n13621 ^ n976 ;
  assign n13626 = n5489 & ~n6215 ;
  assign n13627 = n13626 ^ n7853 ^ 1'b0 ;
  assign n13628 = ~n8559 & n13627 ;
  assign n13629 = n5136 & ~n13628 ;
  assign n13630 = n10275 ^ n9861 ^ 1'b0 ;
  assign n13631 = n10234 | n13630 ;
  assign n13632 = n1926 | n4562 ;
  assign n13633 = n13632 ^ n8842 ^ 1'b0 ;
  assign n13634 = n9745 ^ n479 ^ 1'b0 ;
  assign n13635 = ~n2847 & n13634 ;
  assign n13636 = n13635 ^ n6617 ^ n6060 ;
  assign n13637 = n5903 | n11289 ;
  assign n13638 = n6869 & ~n13637 ;
  assign n13639 = n8379 ^ n5201 ^ n1665 ;
  assign n13640 = n13639 ^ n10286 ^ 1'b0 ;
  assign n13641 = n13638 | n13640 ;
  assign n13642 = n5334 ^ n901 ^ 1'b0 ;
  assign n13643 = n13642 ^ n3472 ^ 1'b0 ;
  assign n13644 = n600 & ~n3509 ;
  assign n13645 = ~n5436 & n13644 ;
  assign n13646 = n2765 ^ n2651 ^ 1'b0 ;
  assign n13647 = n13646 ^ n1125 ^ 1'b0 ;
  assign n13648 = n4310 & n13647 ;
  assign n13649 = n5265 & n13648 ;
  assign n13650 = n13649 ^ n4059 ^ 1'b0 ;
  assign n13651 = ( ~n4379 & n13497 ) | ( ~n4379 & n13650 ) | ( n13497 & n13650 ) ;
  assign n13652 = n2647 & n11880 ;
  assign n13653 = ~n348 & n13652 ;
  assign n13654 = n1284 ^ n1156 ^ 1'b0 ;
  assign n13655 = n1054 & n13654 ;
  assign n13656 = n8878 & n13655 ;
  assign n13657 = n13656 ^ n2449 ^ 1'b0 ;
  assign n13658 = ~n7427 & n13657 ;
  assign n13659 = n8790 & n13658 ;
  assign n13660 = n7943 ^ n3617 ^ n1521 ;
  assign n13661 = n8194 & n13660 ;
  assign n13662 = n12795 ^ n2520 ^ x11 ;
  assign n13666 = n4474 ^ n3661 ^ 1'b0 ;
  assign n13667 = ( n3759 & n6022 ) | ( n3759 & n7716 ) | ( n6022 & n7716 ) ;
  assign n13668 = ( ~n3075 & n13666 ) | ( ~n3075 & n13667 ) | ( n13666 & n13667 ) ;
  assign n13664 = n890 & n1045 ;
  assign n13663 = n1964 & ~n8023 ;
  assign n13665 = n13664 ^ n13663 ^ 1'b0 ;
  assign n13669 = n13668 ^ n13665 ^ n9757 ;
  assign n13671 = n3737 & ~n12433 ;
  assign n13672 = n13671 ^ n2270 ^ 1'b0 ;
  assign n13670 = n2273 & n4491 ;
  assign n13673 = n13672 ^ n13670 ^ 1'b0 ;
  assign n13674 = n13673 ^ n9549 ^ n7544 ;
  assign n13675 = n13118 ^ n6594 ^ x175 ;
  assign n13676 = n3296 & ~n3870 ;
  assign n13677 = n6355 ^ n3495 ^ 1'b0 ;
  assign n13678 = n12741 & n13677 ;
  assign n13679 = ~n11358 & n13678 ;
  assign n13680 = n13679 ^ n3301 ^ 1'b0 ;
  assign n13681 = n13676 | n13680 ;
  assign n13686 = n9108 & ~n13368 ;
  assign n13682 = ~n2206 & n8389 ;
  assign n13683 = n13682 ^ n316 ^ 1'b0 ;
  assign n13684 = ~n8558 & n13683 ;
  assign n13685 = n9417 & ~n13684 ;
  assign n13687 = n13686 ^ n13685 ^ n483 ;
  assign n13688 = n7447 ^ n3195 ^ 1'b0 ;
  assign n13689 = n13687 & ~n13688 ;
  assign n13690 = n2712 | n6030 ;
  assign n13691 = n13690 ^ n8757 ^ 1'b0 ;
  assign n13692 = ( n799 & ~n6645 ) | ( n799 & n10763 ) | ( ~n6645 & n10763 ) ;
  assign n13693 = n13692 ^ n3542 ^ 1'b0 ;
  assign n13694 = n13693 ^ n6797 ^ n1938 ;
  assign n13695 = n2970 | n13694 ;
  assign n13696 = n1016 | n13309 ;
  assign n13697 = n13696 ^ n7209 ^ 1'b0 ;
  assign n13698 = n13697 ^ n12974 ^ n1769 ;
  assign n13699 = n13698 ^ n5444 ^ 1'b0 ;
  assign n13700 = n13699 ^ n10177 ^ 1'b0 ;
  assign n13701 = n1243 & n13700 ;
  assign n13702 = n4036 | n4180 ;
  assign n13703 = ~n10780 & n13702 ;
  assign n13704 = n9662 | n11281 ;
  assign n13705 = n2191 ^ n1328 ^ 1'b0 ;
  assign n13706 = ~n6215 & n13705 ;
  assign n13707 = n3699 | n5025 ;
  assign n13708 = n13707 ^ n4727 ^ 1'b0 ;
  assign n13709 = n13706 & n13708 ;
  assign n13710 = n13709 ^ n2998 ^ 1'b0 ;
  assign n13711 = ~n4739 & n13710 ;
  assign n13712 = n1037 | n13711 ;
  assign n13713 = n7515 & ~n13571 ;
  assign n13714 = ( n5701 & n11826 ) | ( n5701 & n13713 ) | ( n11826 & n13713 ) ;
  assign n13721 = n4557 & ~n10120 ;
  assign n13715 = n5239 ^ n2599 ^ 1'b0 ;
  assign n13716 = n6974 | n13715 ;
  assign n13717 = n9304 ^ n688 ^ n410 ;
  assign n13718 = n13717 ^ n1245 ^ 1'b0 ;
  assign n13719 = ( n1995 & n3406 ) | ( n1995 & n13718 ) | ( n3406 & n13718 ) ;
  assign n13720 = ( ~n4119 & n13716 ) | ( ~n4119 & n13719 ) | ( n13716 & n13719 ) ;
  assign n13722 = n13721 ^ n13720 ^ n8250 ;
  assign n13723 = n4783 & ~n13722 ;
  assign n13724 = n9396 ^ n6699 ^ n3839 ;
  assign n13725 = n13724 ^ n2783 ^ n1294 ;
  assign n13726 = ~n4819 & n10216 ;
  assign n13727 = n9136 ^ n3962 ^ 1'b0 ;
  assign n13728 = n11058 | n13727 ;
  assign n13729 = n5332 | n12784 ;
  assign n13732 = n4556 ^ n1333 ^ 1'b0 ;
  assign n13733 = ~n5362 & n13732 ;
  assign n13734 = ( ~n650 & n4874 ) | ( ~n650 & n13733 ) | ( n4874 & n13733 ) ;
  assign n13730 = n5671 | n9175 ;
  assign n13731 = n13730 ^ n4179 ^ 1'b0 ;
  assign n13735 = n13734 ^ n13731 ^ n5947 ;
  assign n13736 = n7724 ^ n3437 ^ 1'b0 ;
  assign n13737 = n13735 & ~n13736 ;
  assign n13738 = n7734 ^ n6657 ^ n521 ;
  assign n13739 = n5828 ^ n555 ^ 1'b0 ;
  assign n13740 = n13738 & n13739 ;
  assign n13741 = ( ~n1016 & n10074 ) | ( ~n1016 & n13740 ) | ( n10074 & n13740 ) ;
  assign n13742 = n13741 ^ n10506 ^ n5229 ;
  assign n13743 = n2359 & ~n3202 ;
  assign n13744 = n13742 & ~n13743 ;
  assign n13745 = ( x140 & n13737 ) | ( x140 & n13744 ) | ( n13737 & n13744 ) ;
  assign n13750 = ( n3091 & n6876 ) | ( n3091 & ~n12881 ) | ( n6876 & ~n12881 ) ;
  assign n13747 = n9229 ^ n3960 ^ 1'b0 ;
  assign n13748 = n1092 | n13747 ;
  assign n13746 = n725 & n3372 ;
  assign n13749 = n13748 ^ n13746 ^ 1'b0 ;
  assign n13751 = n13750 ^ n13749 ^ n7172 ;
  assign n13754 = n7787 ^ n2913 ^ 1'b0 ;
  assign n13755 = n2629 | n13754 ;
  assign n13756 = n13755 ^ n10648 ^ 1'b0 ;
  assign n13757 = n2563 & ~n13756 ;
  assign n13752 = n4464 & n8188 ;
  assign n13753 = ( n3226 & n7215 ) | ( n3226 & n13752 ) | ( n7215 & n13752 ) ;
  assign n13758 = n13757 ^ n13753 ^ n1786 ;
  assign n13759 = n13758 ^ n8800 ^ n4526 ;
  assign n13760 = n4088 & ~n6624 ;
  assign n13761 = ( n2036 & n3312 ) | ( n2036 & n7128 ) | ( n3312 & n7128 ) ;
  assign n13762 = n13760 & n13761 ;
  assign n13763 = n10172 & n13762 ;
  assign n13764 = ( n4287 & n7427 ) | ( n4287 & n7533 ) | ( n7427 & n7533 ) ;
  assign n13765 = n2907 & n4677 ;
  assign n13766 = n13764 & n13765 ;
  assign n13767 = n13766 ^ n6092 ^ 1'b0 ;
  assign n13768 = n5589 | n13767 ;
  assign n13769 = n9624 & ~n13768 ;
  assign n13770 = n7971 & n13769 ;
  assign n13771 = n4605 ^ n1046 ^ 1'b0 ;
  assign n13772 = n13771 ^ n13434 ^ n4360 ;
  assign n13773 = n13772 ^ n5850 ^ 1'b0 ;
  assign n13774 = n13770 | n13773 ;
  assign n13779 = ~n834 & n7371 ;
  assign n13780 = n6560 & n13779 ;
  assign n13778 = n6629 ^ n2400 ^ 1'b0 ;
  assign n13775 = n1957 & n2184 ;
  assign n13776 = ~n1212 & n13775 ;
  assign n13777 = n13776 ^ n7217 ^ n4789 ;
  assign n13781 = n13780 ^ n13778 ^ n13777 ;
  assign n13782 = n11193 ^ n7701 ^ 1'b0 ;
  assign n13783 = ~n6228 & n13782 ;
  assign n13784 = n2365 ^ n1044 ^ 1'b0 ;
  assign n13785 = ~n8051 & n13784 ;
  assign n13786 = n13785 ^ n8066 ^ 1'b0 ;
  assign n13787 = n11476 ^ n639 ^ 1'b0 ;
  assign n13788 = n1749 & n5995 ;
  assign n13789 = ~n8282 & n13788 ;
  assign n13790 = n13789 ^ n13166 ^ 1'b0 ;
  assign n13791 = ~n13787 & n13790 ;
  assign n13792 = n3774 & n6994 ;
  assign n13793 = n13792 ^ n7860 ^ 1'b0 ;
  assign n13794 = n3313 & n13793 ;
  assign n13795 = ~n6218 & n13794 ;
  assign n13796 = n13795 ^ n1547 ^ 1'b0 ;
  assign n13797 = n13549 & ~n13796 ;
  assign n13798 = n8735 | n13797 ;
  assign n13799 = n2070 ^ n1409 ^ 1'b0 ;
  assign n13800 = n13799 ^ n2000 ^ n307 ;
  assign n13801 = ( n1333 & n5222 ) | ( n1333 & n13800 ) | ( n5222 & n13800 ) ;
  assign n13802 = n1340 | n1444 ;
  assign n13803 = n6995 & ~n13802 ;
  assign n13804 = ( n980 & n2518 ) | ( n980 & n13467 ) | ( n2518 & n13467 ) ;
  assign n13805 = ~n4538 & n4726 ;
  assign n13806 = n13804 & n13805 ;
  assign n13807 = n13806 ^ n9093 ^ n782 ;
  assign n13809 = n4008 | n5349 ;
  assign n13810 = n13809 ^ n1952 ^ 1'b0 ;
  assign n13808 = n4917 | n11998 ;
  assign n13811 = n13810 ^ n13808 ^ 1'b0 ;
  assign n13812 = n938 & n1839 ;
  assign n13813 = n13812 ^ n9491 ^ n6789 ;
  assign n13814 = n13535 ^ n12515 ^ n10446 ;
  assign n13815 = n13814 ^ n6209 ^ n2928 ;
  assign n13816 = ~n258 & n2004 ;
  assign n13817 = n13816 ^ n7600 ^ 1'b0 ;
  assign n13818 = ( ~n1284 & n4724 ) | ( ~n1284 & n13817 ) | ( n4724 & n13817 ) ;
  assign n13819 = ( n5785 & n13719 ) | ( n5785 & n13818 ) | ( n13719 & n13818 ) ;
  assign n13820 = n8423 | n13819 ;
  assign n13831 = n1759 & ~n8818 ;
  assign n13827 = n958 & ~n6917 ;
  assign n13828 = n13827 ^ n5500 ^ 1'b0 ;
  assign n13829 = n1405 & n13828 ;
  assign n13830 = n5046 & n13829 ;
  assign n13832 = n13831 ^ n13830 ^ n7990 ;
  assign n13826 = ~n357 & n9069 ;
  assign n13833 = n13832 ^ n13826 ^ 1'b0 ;
  assign n13834 = n10054 | n13833 ;
  assign n13821 = n13147 ^ n477 ^ 1'b0 ;
  assign n13822 = ~n2464 & n13821 ;
  assign n13823 = ~n4235 & n13822 ;
  assign n13824 = n13823 ^ n9973 ^ 1'b0 ;
  assign n13825 = n4364 | n13824 ;
  assign n13835 = n13834 ^ n13825 ^ 1'b0 ;
  assign n13836 = n1301 | n10141 ;
  assign n13837 = n1655 ^ n1121 ^ 1'b0 ;
  assign n13838 = n13837 ^ n3313 ^ 1'b0 ;
  assign n13839 = n2221 ^ n541 ^ 1'b0 ;
  assign n13840 = n11564 | n13839 ;
  assign n13841 = n4030 & n4637 ;
  assign n13842 = n13841 ^ n12968 ^ n7308 ;
  assign n13843 = n1934 & ~n3924 ;
  assign n13844 = n9294 ^ n6562 ^ n2443 ;
  assign n13845 = n9919 & ~n13844 ;
  assign n13846 = ~n13843 & n13845 ;
  assign n13847 = n2287 & ~n3366 ;
  assign n13848 = ~n12958 & n13847 ;
  assign n13849 = n11312 ^ n5915 ^ x232 ;
  assign n13850 = ~n3857 & n8744 ;
  assign n13851 = n13850 ^ n11572 ^ n9491 ;
  assign n13852 = ~n783 & n5585 ;
  assign n13853 = n13731 ^ n2336 ^ 1'b0 ;
  assign n13854 = n4730 ^ n4546 ^ 1'b0 ;
  assign n13855 = n13207 ^ n1881 ^ 1'b0 ;
  assign n13866 = n5125 ^ n416 ^ 1'b0 ;
  assign n13867 = n1359 & n13866 ;
  assign n13868 = n13867 ^ n7513 ^ 1'b0 ;
  assign n13863 = n2328 | n3807 ;
  assign n13864 = n12780 | n13863 ;
  assign n13865 = n6642 & n13864 ;
  assign n13869 = n13868 ^ n13865 ^ 1'b0 ;
  assign n13856 = ~n4600 & n7149 ;
  assign n13857 = ( n2167 & n3892 ) | ( n2167 & n11291 ) | ( n3892 & n11291 ) ;
  assign n13858 = n3771 | n13857 ;
  assign n13859 = n13858 ^ n4066 ^ 1'b0 ;
  assign n13860 = n3010 & ~n13092 ;
  assign n13861 = ~n13859 & n13860 ;
  assign n13862 = n13856 & ~n13861 ;
  assign n13870 = n13869 ^ n13862 ^ 1'b0 ;
  assign n13872 = n10572 ^ n5020 ^ 1'b0 ;
  assign n13873 = n4494 | n13872 ;
  assign n13871 = n8385 & n11109 ;
  assign n13874 = n13873 ^ n13871 ^ n11407 ;
  assign n13875 = ~n611 & n8282 ;
  assign n13876 = n10636 & n13875 ;
  assign n13877 = n13876 ^ n764 ^ 1'b0 ;
  assign n13878 = ( n5435 & n8128 ) | ( n5435 & ~n8740 ) | ( n8128 & ~n8740 ) ;
  assign n13879 = ( n547 & ~n4751 ) | ( n547 & n6807 ) | ( ~n4751 & n6807 ) ;
  assign n13880 = n9956 | n13879 ;
  assign n13881 = n3268 | n13880 ;
  assign n13882 = ( n2225 & n7969 ) | ( n2225 & n9961 ) | ( n7969 & n9961 ) ;
  assign n13883 = n999 & ~n12401 ;
  assign n13884 = ~n13882 & n13883 ;
  assign n13885 = n1906 & n12070 ;
  assign n13886 = n5950 & n13885 ;
  assign n13887 = ~n5637 & n13886 ;
  assign n13888 = n10477 ^ n1981 ^ 1'b0 ;
  assign n13889 = n13888 ^ n2143 ^ 1'b0 ;
  assign n13890 = n4815 & ~n13889 ;
  assign n13893 = n5373 & n11258 ;
  assign n13894 = n13893 ^ n361 ^ 1'b0 ;
  assign n13891 = ( n384 & n9141 ) | ( n384 & ~n13657 ) | ( n9141 & ~n13657 ) ;
  assign n13892 = n8422 | n13891 ;
  assign n13895 = n13894 ^ n13892 ^ n2362 ;
  assign n13896 = n1011 & ~n5294 ;
  assign n13897 = ~n12485 & n13896 ;
  assign n13898 = ( n4993 & n7017 ) | ( n4993 & ~n13897 ) | ( n7017 & ~n13897 ) ;
  assign n13899 = ( n561 & ~n9070 ) | ( n561 & n13898 ) | ( ~n9070 & n13898 ) ;
  assign n13900 = n7579 & ~n12411 ;
  assign n13901 = n6797 & n13900 ;
  assign n13905 = ( x22 & n2119 ) | ( x22 & n2413 ) | ( n2119 & n2413 ) ;
  assign n13902 = x30 & ~n5349 ;
  assign n13903 = n13902 ^ n2709 ^ 1'b0 ;
  assign n13904 = n13903 ^ n2210 ^ 1'b0 ;
  assign n13906 = n13905 ^ n13904 ^ n13811 ;
  assign n13907 = n1881 | n7615 ;
  assign n13908 = n13907 ^ n6962 ^ 1'b0 ;
  assign n13909 = n4863 & n13908 ;
  assign n13910 = n10519 ^ n8887 ^ n4007 ;
  assign n13911 = n13910 ^ n12446 ^ n1776 ;
  assign n13912 = n13909 & ~n13911 ;
  assign n13913 = n13912 ^ n12576 ^ 1'b0 ;
  assign n13914 = ( n4398 & ~n11847 ) | ( n4398 & n11897 ) | ( ~n11847 & n11897 ) ;
  assign n13915 = n7750 ^ n6935 ^ n841 ;
  assign n13916 = x146 & ~n1187 ;
  assign n13919 = x184 & n866 ;
  assign n13920 = n1945 & n13919 ;
  assign n13921 = n13920 ^ n2532 ^ n992 ;
  assign n13917 = n5331 ^ n755 ^ 1'b0 ;
  assign n13918 = n10404 & n13917 ;
  assign n13922 = n13921 ^ n13918 ^ 1'b0 ;
  assign n13923 = n13916 & n13922 ;
  assign n13924 = n9654 & n13923 ;
  assign n13925 = n13915 & n13924 ;
  assign n13933 = n1155 & n3429 ;
  assign n13934 = n13933 ^ n2952 ^ 1'b0 ;
  assign n13935 = ( ~n9881 & n10660 ) | ( ~n9881 & n13934 ) | ( n10660 & n13934 ) ;
  assign n13926 = n4612 & ~n5081 ;
  assign n13927 = n13926 ^ n11956 ^ 1'b0 ;
  assign n13928 = ~n1844 & n2785 ;
  assign n13929 = n1059 & n13928 ;
  assign n13930 = x109 & ~n13929 ;
  assign n13931 = n13930 ^ n8463 ^ 1'b0 ;
  assign n13932 = ( n7600 & n13927 ) | ( n7600 & n13931 ) | ( n13927 & n13931 ) ;
  assign n13936 = n13935 ^ n13932 ^ 1'b0 ;
  assign n13938 = n1666 & ~n2362 ;
  assign n13937 = n7686 & ~n9097 ;
  assign n13939 = n13938 ^ n13937 ^ 1'b0 ;
  assign n13940 = n4027 ^ n3116 ^ n2280 ;
  assign n13941 = ~n4316 & n13940 ;
  assign n13942 = n5605 ^ n4410 ^ n2754 ;
  assign n13943 = n13942 ^ n9084 ^ 1'b0 ;
  assign n13944 = n5682 & ~n8716 ;
  assign n13945 = ~n3395 & n13944 ;
  assign n13946 = n13945 ^ n7375 ^ 1'b0 ;
  assign n13947 = ( n8523 & ~n13943 ) | ( n8523 & n13946 ) | ( ~n13943 & n13946 ) ;
  assign n13948 = n3131 ^ x63 ^ 1'b0 ;
  assign n13949 = n686 | n5401 ;
  assign n13950 = n2093 & ~n13949 ;
  assign n13951 = ( x0 & n1844 ) | ( x0 & n6441 ) | ( n1844 & n6441 ) ;
  assign n13952 = ~n13950 & n13951 ;
  assign n13953 = n13952 ^ n649 ^ 1'b0 ;
  assign n13954 = n11544 ^ n3735 ^ 1'b0 ;
  assign n13955 = n3690 | n12754 ;
  assign n13956 = n4568 & ~n13955 ;
  assign n13957 = n1134 | n8093 ;
  assign n13958 = n13957 ^ n2486 ^ 1'b0 ;
  assign n13959 = n5725 & ~n11592 ;
  assign n13960 = ~n3289 & n13959 ;
  assign n13961 = x222 & n11528 ;
  assign n13962 = n9625 ^ n3883 ^ 1'b0 ;
  assign n13963 = n12447 ^ n7296 ^ n5020 ;
  assign n13964 = ( n838 & n3634 ) | ( n838 & n13341 ) | ( n3634 & n13341 ) ;
  assign n13965 = n11266 | n13964 ;
  assign n13966 = n13965 ^ n2299 ^ 1'b0 ;
  assign n13967 = n4047 | n13692 ;
  assign n13968 = n7083 | n13967 ;
  assign n13969 = n11359 ^ n7489 ^ n818 ;
  assign n13970 = ( n4168 & n6282 ) | ( n4168 & ~n13183 ) | ( n6282 & ~n13183 ) ;
  assign n13971 = n8834 & n13970 ;
  assign n13972 = n13969 & n13971 ;
  assign n13974 = n7713 & ~n8558 ;
  assign n13975 = n7462 & n13974 ;
  assign n13973 = n7167 & ~n12222 ;
  assign n13976 = n13975 ^ n13973 ^ 1'b0 ;
  assign n13977 = n13976 ^ x3 ^ 1'b0 ;
  assign n13978 = n3621 | n12677 ;
  assign n13979 = n1427 & ~n1656 ;
  assign n13980 = ~n510 & n13979 ;
  assign n13981 = n13980 ^ n1579 ^ 1'b0 ;
  assign n13982 = n4368 & ~n13981 ;
  assign n13983 = n13982 ^ n10753 ^ n4127 ;
  assign n13984 = n5709 & n10706 ;
  assign n13985 = n7903 ^ n7095 ^ n4208 ;
  assign n13986 = n1742 & ~n3427 ;
  assign n13987 = ( n9309 & n13985 ) | ( n9309 & ~n13986 ) | ( n13985 & ~n13986 ) ;
  assign n13988 = n13104 & n13987 ;
  assign n13989 = n13988 ^ n12507 ^ 1'b0 ;
  assign n13994 = ~n3338 & n5449 ;
  assign n13995 = ( n6117 & ~n6553 ) | ( n6117 & n13994 ) | ( ~n6553 & n13994 ) ;
  assign n13993 = ( n3503 & n5953 ) | ( n3503 & n6626 ) | ( n5953 & n6626 ) ;
  assign n13996 = n13995 ^ n13993 ^ n977 ;
  assign n13990 = n8513 ^ n5539 ^ n4065 ;
  assign n13991 = n3339 | n13990 ;
  assign n13992 = n13991 ^ n10468 ^ 1'b0 ;
  assign n13997 = n13996 ^ n13992 ^ 1'b0 ;
  assign n13998 = ~n11102 & n12959 ;
  assign n13999 = ~n10331 & n13998 ;
  assign n14001 = x55 | n9343 ;
  assign n14002 = n14001 ^ n3856 ^ 1'b0 ;
  assign n14003 = n3155 & ~n14002 ;
  assign n14000 = n3010 & n6299 ;
  assign n14004 = n14003 ^ n14000 ^ 1'b0 ;
  assign n14005 = n10150 | n12028 ;
  assign n14006 = n10504 | n14005 ;
  assign n14011 = n10420 ^ n1873 ^ 1'b0 ;
  assign n14012 = ~n4552 & n14011 ;
  assign n14007 = n13837 ^ n7324 ^ n1994 ;
  assign n14008 = ( n413 & n10026 ) | ( n413 & ~n14007 ) | ( n10026 & ~n14007 ) ;
  assign n14009 = n14008 ^ n8162 ^ 1'b0 ;
  assign n14010 = n13276 | n14009 ;
  assign n14013 = n14012 ^ n14010 ^ n10826 ;
  assign n14014 = n5456 ^ n5274 ^ n576 ;
  assign n14015 = x41 & n3834 ;
  assign n14016 = n14015 ^ n3226 ^ 1'b0 ;
  assign n14017 = n6919 & n14016 ;
  assign n14018 = n10016 & n14017 ;
  assign n14019 = ( n3465 & n6788 ) | ( n3465 & n14018 ) | ( n6788 & n14018 ) ;
  assign n14020 = ( n4040 & n6677 ) | ( n4040 & ~n13734 ) | ( n6677 & ~n13734 ) ;
  assign n14025 = n4478 ^ n2819 ^ 1'b0 ;
  assign n14026 = ~n5770 & n14025 ;
  assign n14027 = n9853 & n14026 ;
  assign n14021 = n1292 | n4435 ;
  assign n14022 = ~n7766 & n14021 ;
  assign n14023 = ~n1480 & n14022 ;
  assign n14024 = n14023 ^ n3906 ^ 1'b0 ;
  assign n14028 = n14027 ^ n14024 ^ 1'b0 ;
  assign n14029 = n9416 ^ n2238 ^ n416 ;
  assign n14030 = n14029 ^ n11387 ^ n8294 ;
  assign n14031 = ( ~x158 & n7966 ) | ( ~x158 & n14030 ) | ( n7966 & n14030 ) ;
  assign n14032 = n14031 ^ n10116 ^ 1'b0 ;
  assign n14033 = n6380 ^ n2685 ^ 1'b0 ;
  assign n14034 = n4759 & n14033 ;
  assign n14035 = ~n4214 & n13372 ;
  assign n14036 = ~n14034 & n14035 ;
  assign n14037 = n8110 & ~n13704 ;
  assign n14038 = n5212 & n14037 ;
  assign n14039 = n284 | n8617 ;
  assign n14040 = n14039 ^ n6387 ^ 1'b0 ;
  assign n14041 = n12757 ^ n6923 ^ n3289 ;
  assign n14042 = n378 & n8947 ;
  assign n14043 = n14042 ^ n9517 ^ 1'b0 ;
  assign n14044 = n3268 & n14043 ;
  assign n14045 = ( n14040 & n14041 ) | ( n14040 & ~n14044 ) | ( n14041 & ~n14044 ) ;
  assign n14053 = n7566 | n7881 ;
  assign n14051 = ( n9475 & n10288 ) | ( n9475 & ~n13938 ) | ( n10288 & ~n13938 ) ;
  assign n14052 = n14051 ^ n7571 ^ n1683 ;
  assign n14046 = n485 | n1499 ;
  assign n14047 = n14046 ^ n2909 ^ 1'b0 ;
  assign n14048 = n3891 | n14047 ;
  assign n14049 = n7735 & ~n14048 ;
  assign n14050 = ( n11284 & n12922 ) | ( n11284 & ~n14049 ) | ( n12922 & ~n14049 ) ;
  assign n14054 = n14053 ^ n14052 ^ n14050 ;
  assign n14055 = n8273 ^ n5933 ^ 1'b0 ;
  assign n14056 = ( ~n1866 & n3015 ) | ( ~n1866 & n14055 ) | ( n3015 & n14055 ) ;
  assign n14057 = n3453 | n12313 ;
  assign n14058 = n4935 & ~n14057 ;
  assign n14059 = n14058 ^ n12738 ^ n4959 ;
  assign n14060 = n8405 & n12893 ;
  assign n14061 = n6019 ^ n335 ^ 1'b0 ;
  assign n14062 = x206 & ~n2904 ;
  assign n14063 = n14062 ^ x5 ^ 1'b0 ;
  assign n14064 = ~n13272 & n14063 ;
  assign n14065 = n14061 & ~n14064 ;
  assign n14066 = n13748 ^ n7127 ^ 1'b0 ;
  assign n14067 = n3314 & n14066 ;
  assign n14068 = n10446 ^ n7884 ^ n2113 ;
  assign n14069 = ~n8367 & n11625 ;
  assign n14070 = n14068 & n14069 ;
  assign n14071 = n10934 ^ n2657 ^ 1'b0 ;
  assign n14072 = n2149 & n14071 ;
  assign n14073 = n2637 & ~n11121 ;
  assign n14074 = n14072 & n14073 ;
  assign n14075 = ~n11185 & n14074 ;
  assign n14076 = ~n1685 & n4544 ;
  assign n14077 = n5436 ^ n2355 ^ n2333 ;
  assign n14078 = ~n577 & n10290 ;
  assign n14079 = n14078 ^ n1616 ^ 1'b0 ;
  assign n14080 = ( ~n14076 & n14077 ) | ( ~n14076 & n14079 ) | ( n14077 & n14079 ) ;
  assign n14081 = ~n13629 & n14080 ;
  assign n14082 = n7245 & n12728 ;
  assign n14083 = ( n3326 & ~n5633 ) | ( n3326 & n6297 ) | ( ~n5633 & n6297 ) ;
  assign n14084 = n7067 & n14083 ;
  assign n14085 = n11339 & n14084 ;
  assign n14086 = n3809 | n8292 ;
  assign n14087 = ( n939 & n5592 ) | ( n939 & ~n14086 ) | ( n5592 & ~n14086 ) ;
  assign n14089 = ~n362 & n552 ;
  assign n14090 = ~n9900 & n14089 ;
  assign n14088 = ~n1132 & n2620 ;
  assign n14091 = n14090 ^ n14088 ^ 1'b0 ;
  assign n14092 = n14091 ^ n3485 ^ 1'b0 ;
  assign n14093 = ~n14087 & n14092 ;
  assign n14094 = ( n4925 & n9484 ) | ( n4925 & n9715 ) | ( n9484 & n9715 ) ;
  assign n14099 = n3892 ^ n2913 ^ 1'b0 ;
  assign n14098 = ( n295 & ~n2340 ) | ( n295 & n4641 ) | ( ~n2340 & n4641 ) ;
  assign n14100 = n14099 ^ n14098 ^ n12252 ;
  assign n14095 = n6213 ^ x215 ^ 1'b0 ;
  assign n14096 = n1598 & ~n14095 ;
  assign n14097 = n14096 ^ n8400 ^ 1'b0 ;
  assign n14101 = n14100 ^ n14097 ^ n6252 ;
  assign n14102 = n12558 ^ n4670 ^ n3251 ;
  assign n14103 = n14101 | n14102 ;
  assign n14104 = n14094 | n14103 ;
  assign n14105 = ( ~n405 & n5827 ) | ( ~n405 & n8188 ) | ( n5827 & n8188 ) ;
  assign n14106 = ( n4907 & n6081 ) | ( n4907 & ~n14105 ) | ( n6081 & ~n14105 ) ;
  assign n14107 = n4887 ^ n2698 ^ 1'b0 ;
  assign n14108 = n8402 & n14107 ;
  assign n14109 = ( n3345 & n4771 ) | ( n3345 & ~n10885 ) | ( n4771 & ~n10885 ) ;
  assign n14110 = n4782 & n11566 ;
  assign n14111 = n14110 ^ n9377 ^ 1'b0 ;
  assign n14112 = n10214 ^ n6761 ^ 1'b0 ;
  assign n14113 = ~n6461 & n14112 ;
  assign n14114 = n2793 | n13135 ;
  assign n14115 = n3583 & ~n3724 ;
  assign n14116 = n10107 ^ n6991 ^ 1'b0 ;
  assign n14117 = n11735 & ~n14116 ;
  assign n14118 = n1395 | n3933 ;
  assign n14119 = n14118 ^ n6233 ^ 1'b0 ;
  assign n14120 = ~n1311 & n14119 ;
  assign n14121 = n13882 ^ n13819 ^ 1'b0 ;
  assign n14122 = n7621 & n12780 ;
  assign n14123 = n1268 & n3931 ;
  assign n14124 = n14123 ^ n8139 ^ 1'b0 ;
  assign n14125 = ( n4462 & n9287 ) | ( n4462 & n14124 ) | ( n9287 & n14124 ) ;
  assign n14126 = n13749 ^ n1102 ^ n357 ;
  assign n14127 = ( ~n734 & n4427 ) | ( ~n734 & n7702 ) | ( n4427 & n7702 ) ;
  assign n14128 = n405 & n496 ;
  assign n14129 = n12682 ^ n291 ^ 1'b0 ;
  assign n14130 = n9814 ^ n5355 ^ 1'b0 ;
  assign n14131 = ( ~n11427 & n11988 ) | ( ~n11427 & n14130 ) | ( n11988 & n14130 ) ;
  assign n14132 = ( ~n5424 & n5545 ) | ( ~n5424 & n7980 ) | ( n5545 & n7980 ) ;
  assign n14133 = n2983 ^ x180 ^ 1'b0 ;
  assign n14134 = n14133 ^ n11069 ^ n684 ;
  assign n14135 = ( n1186 & n14132 ) | ( n1186 & n14134 ) | ( n14132 & n14134 ) ;
  assign n14136 = n5912 & n8571 ;
  assign n14137 = n12023 & n14136 ;
  assign n14138 = n14137 ^ n12955 ^ 1'b0 ;
  assign n14140 = ~n5459 & n6202 ;
  assign n14141 = ( ~n7810 & n14016 ) | ( ~n7810 & n14140 ) | ( n14016 & n14140 ) ;
  assign n14139 = ( n2963 & n5219 ) | ( n2963 & ~n7185 ) | ( n5219 & ~n7185 ) ;
  assign n14142 = n14141 ^ n14139 ^ n548 ;
  assign n14143 = n487 | n1638 ;
  assign n14144 = n9147 & ~n11959 ;
  assign n14145 = n14144 ^ n3141 ^ 1'b0 ;
  assign n14146 = n14143 & n14145 ;
  assign n14148 = n2571 ^ n1828 ^ n1458 ;
  assign n14147 = n12478 ^ n11157 ^ 1'b0 ;
  assign n14149 = n14148 ^ n14147 ^ 1'b0 ;
  assign n14150 = ~n8800 & n14149 ;
  assign n14155 = ~n1574 & n3294 ;
  assign n14156 = n11041 | n14155 ;
  assign n14151 = n13733 ^ n1705 ^ 1'b0 ;
  assign n14152 = ~n11684 & n14151 ;
  assign n14153 = n14152 ^ n3015 ^ 1'b0 ;
  assign n14154 = n14153 ^ n11420 ^ n9878 ;
  assign n14157 = n14156 ^ n14154 ^ n703 ;
  assign n14159 = n4923 ^ n3089 ^ n1427 ;
  assign n14160 = n14159 ^ n11576 ^ 1'b0 ;
  assign n14158 = n1135 & n13367 ;
  assign n14161 = n14160 ^ n14158 ^ 1'b0 ;
  assign n14163 = n2145 ^ n1372 ^ n940 ;
  assign n14162 = n5184 | n7941 ;
  assign n14164 = n14163 ^ n14162 ^ 1'b0 ;
  assign n14165 = n1576 & n12525 ;
  assign n14166 = n14165 ^ n13345 ^ 1'b0 ;
  assign n14167 = n14164 & n14166 ;
  assign n14168 = n693 & ~n10130 ;
  assign n14175 = ( n1882 & ~n1935 ) | ( n1882 & n5110 ) | ( ~n1935 & n5110 ) ;
  assign n14169 = n5229 ^ n3242 ^ 1'b0 ;
  assign n14170 = n5064 & ~n14169 ;
  assign n14171 = n8798 & n14170 ;
  assign n14172 = ~n3362 & n14171 ;
  assign n14173 = n14172 ^ n1363 ^ 1'b0 ;
  assign n14174 = n14173 ^ n7225 ^ 1'b0 ;
  assign n14176 = n14175 ^ n14174 ^ 1'b0 ;
  assign n14177 = n8024 & ~n14176 ;
  assign n14178 = ( n1647 & n14168 ) | ( n1647 & n14177 ) | ( n14168 & n14177 ) ;
  assign n14179 = n7088 ^ n2442 ^ 1'b0 ;
  assign n14180 = n14179 ^ n1689 ^ n1454 ;
  assign n14181 = n7329 ^ n6120 ^ 1'b0 ;
  assign n14182 = n13282 & n14181 ;
  assign n14183 = ( n477 & n1562 ) | ( n477 & ~n4619 ) | ( n1562 & ~n4619 ) ;
  assign n14184 = n14183 ^ n12871 ^ n12203 ;
  assign n14191 = n1405 & ~n7452 ;
  assign n14192 = n715 & n14191 ;
  assign n14193 = n10963 & ~n14192 ;
  assign n14188 = ( n4104 & ~n6707 ) | ( n4104 & n7094 ) | ( ~n6707 & n7094 ) ;
  assign n14189 = ( n2062 & n8905 ) | ( n2062 & ~n14188 ) | ( n8905 & ~n14188 ) ;
  assign n14185 = n3857 & ~n7803 ;
  assign n14186 = ~n2164 & n14185 ;
  assign n14187 = n6316 | n14186 ;
  assign n14190 = n14189 ^ n14187 ^ 1'b0 ;
  assign n14194 = n14193 ^ n14190 ^ n5567 ;
  assign n14195 = ( ~n1403 & n8398 ) | ( ~n1403 & n9358 ) | ( n8398 & n9358 ) ;
  assign n14196 = n14195 ^ n11862 ^ 1'b0 ;
  assign n14199 = n3384 ^ n1374 ^ 1'b0 ;
  assign n14197 = n4497 ^ n2864 ^ n619 ;
  assign n14198 = n5827 & ~n14197 ;
  assign n14200 = n14199 ^ n14198 ^ 1'b0 ;
  assign n14201 = n1796 | n10269 ;
  assign n14202 = n964 | n12702 ;
  assign n14203 = n2692 & ~n14202 ;
  assign n14204 = n14203 ^ n10906 ^ n3792 ;
  assign n14205 = n12788 ^ n8324 ^ n7529 ;
  assign n14206 = n8995 ^ n8273 ^ n4243 ;
  assign n14207 = ( n13229 & n14205 ) | ( n13229 & n14206 ) | ( n14205 & n14206 ) ;
  assign n14214 = n9331 ^ n4916 ^ n583 ;
  assign n14208 = n12605 ^ n6110 ^ n979 ;
  assign n14209 = n2119 & ~n7748 ;
  assign n14210 = n1199 & n14209 ;
  assign n14211 = n14208 | n14210 ;
  assign n14212 = n14211 ^ n8519 ^ 1'b0 ;
  assign n14213 = ~n2596 & n14212 ;
  assign n14215 = n14214 ^ n14213 ^ 1'b0 ;
  assign n14216 = n10181 | n12265 ;
  assign n14217 = n434 | n14216 ;
  assign n14218 = n9904 ^ n3075 ^ n1738 ;
  assign n14220 = n1163 | n5807 ;
  assign n14219 = n9228 & ~n11212 ;
  assign n14221 = n14220 ^ n14219 ^ 1'b0 ;
  assign n14222 = n9054 | n14221 ;
  assign n14223 = n14222 ^ n3182 ^ 1'b0 ;
  assign n14224 = n9821 ^ n4952 ^ n4378 ;
  assign n14225 = n9562 ^ n4763 ^ 1'b0 ;
  assign n14226 = ~n5933 & n14225 ;
  assign n14227 = n5092 & n14226 ;
  assign n14228 = ~n12462 & n14227 ;
  assign n14229 = n4345 | n14228 ;
  assign n14230 = n14224 & ~n14229 ;
  assign n14231 = n10906 | n11270 ;
  assign n14232 = n14231 ^ n7494 ^ 1'b0 ;
  assign n14233 = n14232 ^ n8090 ^ 1'b0 ;
  assign n14235 = n7485 ^ x113 ^ 1'b0 ;
  assign n14236 = n14235 ^ n550 ^ 1'b0 ;
  assign n14237 = n870 & n14236 ;
  assign n14238 = n14237 ^ n12562 ^ 1'b0 ;
  assign n14239 = ~n4993 & n14238 ;
  assign n14234 = n771 | n10668 ;
  assign n14240 = n14239 ^ n14234 ^ 1'b0 ;
  assign n14241 = n14240 ^ n8739 ^ n1843 ;
  assign n14242 = n8199 | n10436 ;
  assign n14243 = n3765 & ~n14242 ;
  assign n14247 = x177 & ~n8438 ;
  assign n14248 = n3868 & ~n11849 ;
  assign n14249 = ~n2907 & n14248 ;
  assign n14250 = n14247 & ~n14249 ;
  assign n14251 = n14250 ^ n6294 ^ 1'b0 ;
  assign n14252 = n8649 ^ n5683 ^ 1'b0 ;
  assign n14253 = n14251 & n14252 ;
  assign n14244 = ( x187 & n2142 ) | ( x187 & n4945 ) | ( n2142 & n4945 ) ;
  assign n14245 = n3144 & ~n14244 ;
  assign n14246 = ~n8945 & n14245 ;
  assign n14254 = n14253 ^ n14246 ^ 1'b0 ;
  assign n14255 = n14254 ^ n8410 ^ 1'b0 ;
  assign n14256 = n14226 ^ n3402 ^ n2119 ;
  assign n14257 = ~n6123 & n14256 ;
  assign n14258 = n14257 ^ n4573 ^ 1'b0 ;
  assign n14259 = n14258 ^ n8561 ^ 1'b0 ;
  assign n14260 = n6087 & ~n14259 ;
  assign n14261 = n11644 & n14260 ;
  assign n14267 = x79 & n1004 ;
  assign n14264 = n5315 | n12823 ;
  assign n14265 = n11849 & ~n14264 ;
  assign n14266 = ( x90 & ~n1594 ) | ( x90 & n14265 ) | ( ~n1594 & n14265 ) ;
  assign n14262 = n5183 ^ n1113 ^ n768 ;
  assign n14263 = n14262 ^ n5231 ^ n3753 ;
  assign n14268 = n14267 ^ n14266 ^ n14263 ;
  assign n14272 = n2263 & ~n6732 ;
  assign n14273 = n14272 ^ n3831 ^ 1'b0 ;
  assign n14274 = ( n3323 & n11760 ) | ( n3323 & n14273 ) | ( n11760 & n14273 ) ;
  assign n14271 = n649 & ~n2610 ;
  assign n14275 = n14274 ^ n14271 ^ 1'b0 ;
  assign n14270 = n3162 | n4146 ;
  assign n14269 = n2731 & ~n7398 ;
  assign n14276 = n14275 ^ n14270 ^ n14269 ;
  assign n14277 = n4533 & ~n5473 ;
  assign n14278 = n14277 ^ n2849 ^ 1'b0 ;
  assign n14279 = n6220 ^ n3325 ^ 1'b0 ;
  assign n14280 = ~n3555 & n5074 ;
  assign n14281 = n14132 & n14280 ;
  assign n14282 = n14281 ^ n8550 ^ 1'b0 ;
  assign n14283 = ( n1444 & n14279 ) | ( n1444 & ~n14282 ) | ( n14279 & ~n14282 ) ;
  assign n14284 = n8930 ^ n8151 ^ 1'b0 ;
  assign n14285 = n14284 ^ n10310 ^ 1'b0 ;
  assign n14286 = n5438 | n6560 ;
  assign n14287 = n14286 ^ n11316 ^ 1'b0 ;
  assign n14295 = n12111 ^ n1451 ^ 1'b0 ;
  assign n14296 = x188 & n14295 ;
  assign n14292 = n1476 & n8599 ;
  assign n14288 = ( n699 & ~n3933 ) | ( n699 & n7682 ) | ( ~n3933 & n7682 ) ;
  assign n14289 = n11631 ^ n6600 ^ 1'b0 ;
  assign n14290 = n14288 & n14289 ;
  assign n14291 = ~n5380 & n14290 ;
  assign n14293 = n14292 ^ n14291 ^ 1'b0 ;
  assign n14294 = n3677 & n14293 ;
  assign n14297 = n14296 ^ n14294 ^ 1'b0 ;
  assign n14298 = n6233 ^ n5150 ^ 1'b0 ;
  assign n14299 = n10889 | n14298 ;
  assign n14300 = n14299 ^ n11896 ^ 1'b0 ;
  assign n14301 = n6149 & n7474 ;
  assign n14302 = n2509 & n14301 ;
  assign n14303 = n9208 ^ n6150 ^ 1'b0 ;
  assign n14304 = n1676 & ~n14303 ;
  assign n14305 = ~n14302 & n14304 ;
  assign n14306 = n14305 ^ n8827 ^ 1'b0 ;
  assign n14307 = n6969 & n7738 ;
  assign n14308 = ( n9876 & n14306 ) | ( n9876 & ~n14307 ) | ( n14306 & ~n14307 ) ;
  assign n14309 = ( n10363 & ~n14083 ) | ( n10363 & n14308 ) | ( ~n14083 & n14308 ) ;
  assign n14311 = ( n2822 & n5784 ) | ( n2822 & ~n11701 ) | ( n5784 & ~n11701 ) ;
  assign n14312 = n14311 ^ n2876 ^ x69 ;
  assign n14310 = n3528 & ~n6074 ;
  assign n14313 = n14312 ^ n14310 ^ n3748 ;
  assign n14314 = n6299 ^ n733 ^ 1'b0 ;
  assign n14315 = n14314 ^ n14206 ^ n8024 ;
  assign n14316 = ( n1385 & n6565 ) | ( n1385 & ~n11645 ) | ( n6565 & ~n11645 ) ;
  assign n14317 = n7391 ^ n4002 ^ 1'b0 ;
  assign n14318 = n3178 & ~n14317 ;
  assign n14319 = n14318 ^ n8198 ^ 1'b0 ;
  assign n14320 = n14319 ^ n7889 ^ n1226 ;
  assign n14321 = ( n2148 & ~n14316 ) | ( n2148 & n14320 ) | ( ~n14316 & n14320 ) ;
  assign n14322 = ~n14315 & n14321 ;
  assign n14323 = n5899 & n14322 ;
  assign n14324 = ( n4077 & n4331 ) | ( n4077 & n6911 ) | ( n4331 & n6911 ) ;
  assign n14325 = n438 & ~n4812 ;
  assign n14326 = n6889 & ~n7401 ;
  assign n14327 = n9060 & n14326 ;
  assign n14328 = ( ~n399 & n14325 ) | ( ~n399 & n14327 ) | ( n14325 & n14327 ) ;
  assign n14329 = n7408 ^ n1903 ^ 1'b0 ;
  assign n14330 = ~n318 & n14329 ;
  assign n14331 = n14330 ^ n4034 ^ 1'b0 ;
  assign n14332 = ( n1102 & n1773 ) | ( n1102 & ~n14331 ) | ( n1773 & ~n14331 ) ;
  assign n14333 = n4311 & ~n7462 ;
  assign n14334 = n7558 ^ n7366 ^ n3330 ;
  assign n14335 = n6848 ^ n2793 ^ 1'b0 ;
  assign n14336 = ~n3309 & n14335 ;
  assign n14337 = n14336 ^ n1487 ^ 1'b0 ;
  assign n14338 = ~n5146 & n14337 ;
  assign n14339 = n14338 ^ n3816 ^ 1'b0 ;
  assign n14340 = ~n2803 & n10885 ;
  assign n14341 = n12823 ^ n6169 ^ 1'b0 ;
  assign n14342 = n14341 ^ n3859 ^ 1'b0 ;
  assign n14343 = n3113 ^ n1506 ^ 1'b0 ;
  assign n14344 = n2639 & ~n14343 ;
  assign n14345 = n14344 ^ n4869 ^ n2359 ;
  assign n14346 = ( n5183 & ~n11262 ) | ( n5183 & n14345 ) | ( ~n11262 & n14345 ) ;
  assign n14347 = n13406 ^ n12122 ^ n4109 ;
  assign n14349 = n2171 & ~n3949 ;
  assign n14348 = n5945 & ~n11806 ;
  assign n14350 = n14349 ^ n14348 ^ 1'b0 ;
  assign n14351 = n14350 ^ n9724 ^ n3043 ;
  assign n14352 = n11190 & ~n14351 ;
  assign n14353 = n6373 ^ n4364 ^ 1'b0 ;
  assign n14354 = ( n6009 & ~n9982 ) | ( n6009 & n14353 ) | ( ~n9982 & n14353 ) ;
  assign n14355 = n14354 ^ n5304 ^ 1'b0 ;
  assign n14356 = n9332 | n14355 ;
  assign n14357 = n3330 & ~n4974 ;
  assign n14358 = n14357 ^ n1294 ^ 1'b0 ;
  assign n14359 = n11804 ^ n9431 ^ 1'b0 ;
  assign n14360 = n5574 & n14359 ;
  assign n14361 = n14360 ^ n3380 ^ 1'b0 ;
  assign n14362 = ( n1101 & ~n14358 ) | ( n1101 & n14361 ) | ( ~n14358 & n14361 ) ;
  assign n14365 = n8327 ^ n3992 ^ n1165 ;
  assign n14366 = n14365 ^ n1800 ^ 1'b0 ;
  assign n14363 = n9973 ^ n3575 ^ 1'b0 ;
  assign n14364 = ~n5473 & n14363 ;
  assign n14367 = n14366 ^ n14364 ^ 1'b0 ;
  assign n14368 = ~n5724 & n14367 ;
  assign n14369 = ( n391 & n9499 ) | ( n391 & n9530 ) | ( n9499 & n9530 ) ;
  assign n14370 = ( ~n2683 & n14368 ) | ( ~n2683 & n14369 ) | ( n14368 & n14369 ) ;
  assign n14371 = n533 & ~n14370 ;
  assign n14373 = n11121 ^ n4609 ^ n4090 ;
  assign n14374 = n14373 ^ n2952 ^ n1165 ;
  assign n14372 = n2276 & n3088 ;
  assign n14375 = n14374 ^ n14372 ^ n8695 ;
  assign n14376 = ~n6665 & n11213 ;
  assign n14377 = n14376 ^ n894 ^ 1'b0 ;
  assign n14378 = n4797 & n14377 ;
  assign n14379 = n14378 ^ n3111 ^ 1'b0 ;
  assign n14380 = n12974 | n14379 ;
  assign n14382 = n7852 ^ n4008 ^ n2074 ;
  assign n14381 = n4376 ^ n4173 ^ n554 ;
  assign n14383 = n14382 ^ n14381 ^ n678 ;
  assign n14384 = n8607 ^ n8111 ^ 1'b0 ;
  assign n14385 = n6690 & n14384 ;
  assign n14389 = n7285 ^ n5779 ^ n1180 ;
  assign n14390 = ( ~n687 & n11472 ) | ( ~n687 & n14389 ) | ( n11472 & n14389 ) ;
  assign n14386 = n6463 & ~n7914 ;
  assign n14387 = n14386 ^ n10513 ^ 1'b0 ;
  assign n14388 = n12959 & ~n14387 ;
  assign n14391 = n14390 ^ n14388 ^ n10483 ;
  assign n14392 = ~n1423 & n9798 ;
  assign n14393 = ~n5068 & n14392 ;
  assign n14397 = n345 & n12891 ;
  assign n14394 = x112 & n2868 ;
  assign n14395 = ~n5567 & n14394 ;
  assign n14396 = ( n1004 & n2008 ) | ( n1004 & ~n14395 ) | ( n2008 & ~n14395 ) ;
  assign n14398 = n14397 ^ n14396 ^ 1'b0 ;
  assign n14399 = n14393 | n14398 ;
  assign n14400 = n10078 ^ n9465 ^ 1'b0 ;
  assign n14401 = n4004 & ~n14400 ;
  assign n14402 = n6486 ^ n5196 ^ n3585 ;
  assign n14403 = n14401 | n14402 ;
  assign n14404 = n14403 ^ n7315 ^ 1'b0 ;
  assign n14405 = n4284 ^ n1974 ^ 1'b0 ;
  assign n14406 = n1664 & n14405 ;
  assign n14407 = n8083 ^ n7769 ^ n587 ;
  assign n14408 = n9612 ^ n2743 ^ 1'b0 ;
  assign n14409 = ~n8890 & n14408 ;
  assign n14410 = n7158 ^ n4530 ^ 1'b0 ;
  assign n14411 = ( n14407 & n14409 ) | ( n14407 & n14410 ) | ( n14409 & n14410 ) ;
  assign n14412 = n14406 & n14411 ;
  assign n14413 = ~n11381 & n14412 ;
  assign n14414 = ~n2567 & n3844 ;
  assign n14415 = ~x14 & n14414 ;
  assign n14416 = n8465 ^ n3483 ^ 1'b0 ;
  assign n14417 = n3791 & ~n14416 ;
  assign n14418 = ( ~x21 & n946 ) | ( ~x21 & n6176 ) | ( n946 & n6176 ) ;
  assign n14419 = n14418 ^ n9131 ^ n2206 ;
  assign n14420 = n1517 | n10794 ;
  assign n14421 = n6442 | n14420 ;
  assign n14422 = ( n3321 & ~n14269 ) | ( n3321 & n14421 ) | ( ~n14269 & n14421 ) ;
  assign n14423 = ~n5982 & n6174 ;
  assign n14424 = ~n10167 & n14423 ;
  assign n14425 = n8383 ^ n6271 ^ 1'b0 ;
  assign n14426 = n14425 ^ n5006 ^ 1'b0 ;
  assign n14427 = n8394 ^ n6910 ^ n4759 ;
  assign n14428 = ~n10738 & n14427 ;
  assign n14429 = n13753 ^ n3093 ^ 1'b0 ;
  assign n14430 = n14429 ^ n11645 ^ 1'b0 ;
  assign n14431 = ~n12092 & n14430 ;
  assign n14432 = n14431 ^ n1422 ^ 1'b0 ;
  assign n14434 = ~n3184 & n3479 ;
  assign n14435 = ~n2685 & n14434 ;
  assign n14433 = n9174 ^ n7657 ^ 1'b0 ;
  assign n14436 = n14435 ^ n14433 ^ 1'b0 ;
  assign n14437 = n14034 & ~n14436 ;
  assign n14438 = ~n14432 & n14437 ;
  assign n14439 = n14087 ^ n12569 ^ n597 ;
  assign n14440 = n10413 & ~n14439 ;
  assign n14441 = n14440 ^ n4214 ^ 1'b0 ;
  assign n14442 = n4863 & n14441 ;
  assign n14443 = n3609 & n14442 ;
  assign n14444 = ( n6353 & ~n11205 ) | ( n6353 & n11313 ) | ( ~n11205 & n11313 ) ;
  assign n14448 = n1558 | n2856 ;
  assign n14449 = n14448 ^ n1503 ^ 1'b0 ;
  assign n14445 = n8981 ^ n7342 ^ n3765 ;
  assign n14446 = ( n2927 & n3361 ) | ( n2927 & n14445 ) | ( n3361 & n14445 ) ;
  assign n14447 = ~n8080 & n14446 ;
  assign n14450 = n14449 ^ n14447 ^ 1'b0 ;
  assign n14451 = n6478 ^ n864 ^ 1'b0 ;
  assign n14452 = n5332 & ~n14451 ;
  assign n14453 = n8973 & n14452 ;
  assign n14454 = n14450 & n14453 ;
  assign n14455 = n516 & n4065 ;
  assign n14456 = n4137 | n9184 ;
  assign n14457 = n3157 | n14456 ;
  assign n14458 = ( n3555 & n7523 ) | ( n3555 & n14457 ) | ( n7523 & n14457 ) ;
  assign n14459 = n14458 ^ n7399 ^ 1'b0 ;
  assign n14460 = n3488 ^ n3205 ^ n693 ;
  assign n14461 = n8214 ^ n1334 ^ 1'b0 ;
  assign n14462 = n13228 ^ n10129 ^ 1'b0 ;
  assign n14463 = ( n6996 & n7821 ) | ( n6996 & ~n14462 ) | ( n7821 & ~n14462 ) ;
  assign n14464 = ( n10063 & n10961 ) | ( n10063 & ~n14463 ) | ( n10961 & ~n14463 ) ;
  assign n14465 = n14464 ^ n4766 ^ 1'b0 ;
  assign n14466 = ~n5105 & n13856 ;
  assign n14467 = n1592 & n14466 ;
  assign n14468 = n14201 | n14467 ;
  assign n14469 = n3411 | n14468 ;
  assign n14470 = ( n2182 & ~n2560 ) | ( n2182 & n3830 ) | ( ~n2560 & n3830 ) ;
  assign n14471 = n14470 ^ n4673 ^ n822 ;
  assign n14472 = ( n1278 & ~n3559 ) | ( n1278 & n8810 ) | ( ~n3559 & n8810 ) ;
  assign n14473 = n6737 & ~n11570 ;
  assign n14474 = ( ~n4924 & n12378 ) | ( ~n4924 & n13780 ) | ( n12378 & n13780 ) ;
  assign n14475 = n5682 & ~n14474 ;
  assign n14476 = n14473 & n14475 ;
  assign n14477 = ( ~x67 & n6464 ) | ( ~x67 & n14476 ) | ( n6464 & n14476 ) ;
  assign n14478 = n6626 ^ n2192 ^ n1297 ;
  assign n14479 = ~n10306 & n14478 ;
  assign n14480 = n2933 & n13295 ;
  assign n14481 = n14480 ^ n767 ^ 1'b0 ;
  assign n14482 = n4765 & ~n8186 ;
  assign n14483 = ~n13690 & n14482 ;
  assign n14484 = ~n4215 & n13544 ;
  assign n14485 = n14484 ^ n9120 ^ 1'b0 ;
  assign n14486 = n6996 | n14485 ;
  assign n14487 = ~x188 & n450 ;
  assign n14488 = n3779 ^ n2677 ^ 1'b0 ;
  assign n14489 = n14487 & n14488 ;
  assign n14493 = n2978 & ~n7217 ;
  assign n14494 = n12163 & n14493 ;
  assign n14490 = n4141 | n7670 ;
  assign n14491 = n14490 ^ n2097 ^ 1'b0 ;
  assign n14492 = n14491 ^ n10719 ^ 1'b0 ;
  assign n14495 = n14494 ^ n14492 ^ 1'b0 ;
  assign n14496 = n14489 & ~n14495 ;
  assign n14499 = n6574 ^ n4104 ^ n4100 ;
  assign n14497 = n5545 ^ n1646 ^ 1'b0 ;
  assign n14498 = n5129 | n14497 ;
  assign n14500 = n14499 ^ n14498 ^ 1'b0 ;
  assign n14501 = n14496 & n14500 ;
  assign n14505 = n12400 ^ n4875 ^ 1'b0 ;
  assign n14506 = n4510 & n14505 ;
  assign n14507 = n14506 ^ n9799 ^ n6451 ;
  assign n14502 = ( n284 & n4407 ) | ( n284 & n5446 ) | ( n4407 & n5446 ) ;
  assign n14503 = n3100 | n14502 ;
  assign n14504 = n5166 & ~n14503 ;
  assign n14508 = n14507 ^ n14504 ^ n9197 ;
  assign n14509 = n10263 ^ n5942 ^ n2464 ;
  assign n14510 = n10917 ^ n7764 ^ 1'b0 ;
  assign n14511 = n14509 & n14510 ;
  assign n14512 = n632 & ~n1352 ;
  assign n14513 = n3903 & n14512 ;
  assign n14514 = n12580 & ~n14513 ;
  assign n14515 = n14514 ^ n2553 ^ 1'b0 ;
  assign n14516 = n14515 ^ n7083 ^ n1600 ;
  assign n14517 = n14516 ^ n13248 ^ n9758 ;
  assign n14518 = n5366 & n8870 ;
  assign n14519 = n355 & ~n1009 ;
  assign n14520 = n9003 & n14519 ;
  assign n14521 = n1968 & ~n3849 ;
  assign n14522 = n14520 & n14521 ;
  assign n14523 = ( ~n3563 & n14518 ) | ( ~n3563 & n14522 ) | ( n14518 & n14522 ) ;
  assign n14524 = n4624 & ~n6482 ;
  assign n14525 = n7903 & n14524 ;
  assign n14526 = n4391 & ~n13452 ;
  assign n14527 = n14526 ^ n4809 ^ 1'b0 ;
  assign n14528 = n11751 & n14527 ;
  assign n14529 = n9114 ^ n5130 ^ 1'b0 ;
  assign n14530 = ( n3392 & ~n12881 ) | ( n3392 & n14449 ) | ( ~n12881 & n14449 ) ;
  assign n14531 = n905 & n7831 ;
  assign n14533 = n8604 ^ n4864 ^ x66 ;
  assign n14532 = x47 & n11328 ;
  assign n14534 = n14533 ^ n14532 ^ n3431 ;
  assign n14535 = n14531 & ~n14534 ;
  assign n14538 = n1367 ^ n1108 ^ 1'b0 ;
  assign n14539 = n3796 & ~n14538 ;
  assign n14536 = n1814 | n5567 ;
  assign n14537 = ~n14342 & n14536 ;
  assign n14540 = n14539 ^ n14537 ^ 1'b0 ;
  assign n14541 = ~n8304 & n14540 ;
  assign n14542 = n7742 ^ n3360 ^ n695 ;
  assign n14543 = ( n4124 & n13708 ) | ( n4124 & ~n14542 ) | ( n13708 & ~n14542 ) ;
  assign n14544 = n14543 ^ n11196 ^ n9868 ;
  assign n14545 = n6696 ^ n4185 ^ 1'b0 ;
  assign n14546 = n14544 & ~n14545 ;
  assign n14547 = x28 & n14546 ;
  assign n14548 = ( n1123 & ~n4533 ) | ( n1123 & n5992 ) | ( ~n4533 & n5992 ) ;
  assign n14549 = n6509 & ~n14548 ;
  assign n14550 = n14549 ^ n4926 ^ 1'b0 ;
  assign n14551 = n1957 & n14550 ;
  assign n14552 = n10000 ^ n5236 ^ 1'b0 ;
  assign n14553 = n3133 | n10844 ;
  assign n14554 = n4567 | n14553 ;
  assign n14555 = n13306 & n14554 ;
  assign n14556 = ~n3480 & n8905 ;
  assign n14557 = n14556 ^ n5236 ^ 1'b0 ;
  assign n14558 = n14557 ^ n11358 ^ n5344 ;
  assign n14559 = n5262 | n9374 ;
  assign n14560 = n5532 | n14467 ;
  assign n14561 = n14559 | n14560 ;
  assign n14562 = ~n3048 & n8793 ;
  assign n14563 = n13102 & n14562 ;
  assign n14564 = n13706 ^ n3968 ^ 1'b0 ;
  assign n14565 = n14563 & ~n14564 ;
  assign n14566 = n7665 & ~n12289 ;
  assign n14567 = n816 & n2749 ;
  assign n14568 = n14567 ^ n9947 ^ 1'b0 ;
  assign n14569 = ( n11843 & ~n12147 ) | ( n11843 & n14568 ) | ( ~n12147 & n14568 ) ;
  assign n14570 = n5813 ^ n2132 ^ 1'b0 ;
  assign n14571 = n1566 & n14570 ;
  assign n14578 = ( n5844 & ~n9498 ) | ( n5844 & n11127 ) | ( ~n9498 & n11127 ) ;
  assign n14579 = n14578 ^ n6023 ^ n1380 ;
  assign n14573 = n10848 ^ n10458 ^ n3818 ;
  assign n14574 = n12748 & ~n14573 ;
  assign n14575 = n14574 ^ n7526 ^ 1'b0 ;
  assign n14576 = ( n2286 & n5286 ) | ( n2286 & ~n14575 ) | ( n5286 & ~n14575 ) ;
  assign n14572 = n4095 | n4690 ;
  assign n14577 = n14576 ^ n14572 ^ 1'b0 ;
  assign n14580 = n14579 ^ n14577 ^ 1'b0 ;
  assign n14581 = ~n11260 & n14580 ;
  assign n14582 = n1506 & n14581 ;
  assign n14583 = n11019 ^ x82 ^ 1'b0 ;
  assign n14584 = n483 & n7203 ;
  assign n14585 = n14584 ^ n675 ^ 1'b0 ;
  assign n14587 = n3425 ^ n1144 ^ 1'b0 ;
  assign n14586 = n2152 & ~n5228 ;
  assign n14588 = n14587 ^ n14586 ^ n860 ;
  assign n14589 = n8483 ^ n4673 ^ 1'b0 ;
  assign n14590 = x66 & n14589 ;
  assign n14591 = n7831 & n14590 ;
  assign n14592 = ~n13022 & n14591 ;
  assign n14593 = n7264 & ~n14592 ;
  assign n14594 = n14593 ^ n831 ^ 1'b0 ;
  assign n14595 = n3512 | n3713 ;
  assign n14596 = n11381 ^ n7485 ^ 1'b0 ;
  assign n14597 = n14596 ^ n1054 ^ 1'b0 ;
  assign n14598 = n14595 & ~n14597 ;
  assign n14602 = n731 | n6376 ;
  assign n14603 = n14602 ^ n5707 ^ n679 ;
  assign n14599 = n3225 | n7039 ;
  assign n14600 = n7101 & ~n14599 ;
  assign n14601 = x109 & n14600 ;
  assign n14604 = n14603 ^ n14601 ^ n477 ;
  assign n14605 = n13956 ^ n12071 ^ 1'b0 ;
  assign n14606 = ~n11605 & n14605 ;
  assign n14607 = n5007 ^ n4261 ^ 1'b0 ;
  assign n14608 = n11707 | n11962 ;
  assign n14609 = n14607 & ~n14608 ;
  assign n14610 = n1249 ^ n357 ^ 1'b0 ;
  assign n14611 = n3977 & n14610 ;
  assign n14612 = n14462 & n14611 ;
  assign n14613 = n14612 ^ n12096 ^ 1'b0 ;
  assign n14614 = n14613 ^ n11227 ^ n5973 ;
  assign n14615 = n1939 | n9642 ;
  assign n14616 = n10547 ^ n481 ^ 1'b0 ;
  assign n14617 = ~n346 & n14616 ;
  assign n14618 = n14617 ^ n12624 ^ n6246 ;
  assign n14619 = n3702 & ~n4549 ;
  assign n14620 = n4101 & n14619 ;
  assign n14621 = ~n4587 & n6511 ;
  assign n14622 = n14620 | n14621 ;
  assign n14623 = n14618 & ~n14622 ;
  assign n14624 = n4604 ^ n299 ^ 1'b0 ;
  assign n14625 = ( n2238 & n5294 ) | ( n2238 & n7366 ) | ( n5294 & n7366 ) ;
  assign n14626 = n14624 | n14625 ;
  assign n14627 = n1795 | n14626 ;
  assign n14628 = ( n8571 & ~n8801 ) | ( n8571 & n14627 ) | ( ~n8801 & n14627 ) ;
  assign n14629 = n7818 & n13718 ;
  assign n14630 = n14628 & n14629 ;
  assign n14631 = n9403 | n13940 ;
  assign n14632 = n14631 ^ n11684 ^ 1'b0 ;
  assign n14633 = n11907 ^ n9510 ^ n7926 ;
  assign n14634 = n14633 ^ n9321 ^ n1109 ;
  assign n14635 = ~n8953 & n9093 ;
  assign n14636 = ( n7129 & n10637 ) | ( n7129 & ~n14635 ) | ( n10637 & ~n14635 ) ;
  assign n14637 = n736 & ~n6799 ;
  assign n14638 = n14637 ^ n13388 ^ 1'b0 ;
  assign n14639 = n11041 ^ n2476 ^ n1102 ;
  assign n14640 = ~n8770 & n9853 ;
  assign n14641 = ~n2139 & n2770 ;
  assign n14642 = ( n12322 & ~n14640 ) | ( n12322 & n14641 ) | ( ~n14640 & n14641 ) ;
  assign n14643 = n4030 ^ n3991 ^ 1'b0 ;
  assign n14644 = ~n10887 & n14643 ;
  assign n14647 = ~n1749 & n6857 ;
  assign n14648 = ( n5981 & n6066 ) | ( n5981 & n14647 ) | ( n6066 & n14647 ) ;
  assign n14645 = n4446 | n5964 ;
  assign n14646 = n14645 ^ x4 ^ 1'b0 ;
  assign n14649 = n14648 ^ n14646 ^ n2725 ;
  assign n14650 = n14644 & n14649 ;
  assign n14651 = n14650 ^ n10001 ^ 1'b0 ;
  assign n14652 = n8055 ^ n2020 ^ 1'b0 ;
  assign n14653 = n14652 ^ n8861 ^ n4042 ;
  assign n14654 = ( n1283 & n6623 ) | ( n1283 & ~n8361 ) | ( n6623 & ~n8361 ) ;
  assign n14655 = n14654 ^ n13918 ^ 1'b0 ;
  assign n14656 = ( n10209 & n10398 ) | ( n10209 & n11571 ) | ( n10398 & n11571 ) ;
  assign n14657 = n8396 ^ n4536 ^ n3465 ;
  assign n14658 = ( n2575 & ~n7769 ) | ( n2575 & n7980 ) | ( ~n7769 & n7980 ) ;
  assign n14659 = ~n4947 & n14658 ;
  assign n14660 = ~n14657 & n14659 ;
  assign n14661 = ( ~n5148 & n14354 ) | ( ~n5148 & n14660 ) | ( n14354 & n14660 ) ;
  assign n14662 = n6831 & n9170 ;
  assign n14663 = ~n5739 & n14662 ;
  assign n14664 = n10156 ^ n7953 ^ n7424 ;
  assign n14665 = n14664 ^ n4574 ^ n3932 ;
  assign n14666 = n8103 ^ n3220 ^ n2297 ;
  assign n14667 = n6387 & ~n12719 ;
  assign n14668 = n13275 & ~n14667 ;
  assign n14669 = ~x43 & n14668 ;
  assign n14670 = ~n1140 & n3104 ;
  assign n14671 = n14670 ^ n8433 ^ 1'b0 ;
  assign n14672 = ( n1975 & n2550 ) | ( n1975 & ~n14671 ) | ( n2550 & ~n14671 ) ;
  assign n14673 = n8729 & ~n8927 ;
  assign n14674 = n14673 ^ n4226 ^ 1'b0 ;
  assign n14675 = n11534 & n14674 ;
  assign n14676 = n14672 | n14675 ;
  assign n14677 = n2555 & ~n6527 ;
  assign n14678 = n14245 ^ n11013 ^ 1'b0 ;
  assign n14679 = ( n4929 & n9562 ) | ( n4929 & n10170 ) | ( n9562 & n10170 ) ;
  assign n14680 = ~n8413 & n12606 ;
  assign n14681 = n14680 ^ n2116 ^ 1'b0 ;
  assign n14682 = n14679 & n14681 ;
  assign n14683 = n13144 ^ n4169 ^ 1'b0 ;
  assign n14684 = n9752 | n14683 ;
  assign n14685 = n2691 & n9129 ;
  assign n14686 = n14685 ^ n1510 ^ 1'b0 ;
  assign n14687 = ~n1616 & n14686 ;
  assign n14688 = ( ~n2631 & n4723 ) | ( ~n2631 & n12921 ) | ( n4723 & n12921 ) ;
  assign n14689 = n14688 ^ n5087 ^ 1'b0 ;
  assign n14690 = n9742 ^ n6556 ^ 1'b0 ;
  assign n14691 = ( n10054 & ~n14325 ) | ( n10054 & n14690 ) | ( ~n14325 & n14690 ) ;
  assign n14692 = ( n5909 & n14689 ) | ( n5909 & ~n14691 ) | ( n14689 & ~n14691 ) ;
  assign n14695 = n10050 | n12110 ;
  assign n14693 = n13144 ^ n3930 ^ 1'b0 ;
  assign n14694 = n11915 | n14693 ;
  assign n14696 = n14695 ^ n14694 ^ n5978 ;
  assign n14697 = n4091 | n9704 ;
  assign n14698 = ( n3318 & n5767 ) | ( n3318 & n14697 ) | ( n5767 & n14697 ) ;
  assign n14699 = n12086 ^ n7544 ^ 1'b0 ;
  assign n14700 = n2907 & n14699 ;
  assign n14701 = ( n7304 & n14698 ) | ( n7304 & ~n14700 ) | ( n14698 & ~n14700 ) ;
  assign n14702 = ( n13237 & n13886 ) | ( n13237 & ~n14701 ) | ( n13886 & ~n14701 ) ;
  assign n14704 = n13307 ^ n8996 ^ n6682 ;
  assign n14705 = n14704 ^ n13502 ^ 1'b0 ;
  assign n14703 = n6666 ^ n4040 ^ 1'b0 ;
  assign n14706 = n14705 ^ n14703 ^ n690 ;
  assign n14708 = n8698 & ~n12092 ;
  assign n14709 = n14708 ^ n11765 ^ 1'b0 ;
  assign n14710 = n9914 & n14709 ;
  assign n14707 = n10543 ^ n10428 ^ n2206 ;
  assign n14711 = n14710 ^ n14707 ^ 1'b0 ;
  assign n14712 = x46 & ~n14711 ;
  assign n14716 = n3931 ^ n1370 ^ 1'b0 ;
  assign n14717 = ~n420 & n14716 ;
  assign n14715 = n13148 ^ n2241 ^ 1'b0 ;
  assign n14713 = n10185 ^ n687 ^ 1'b0 ;
  assign n14714 = x231 & n14713 ;
  assign n14718 = n14717 ^ n14715 ^ n14714 ;
  assign n14719 = n2068 & ~n3339 ;
  assign n14720 = n4053 & n14719 ;
  assign n14721 = ( n4054 & n4315 ) | ( n4054 & n8754 ) | ( n4315 & n8754 ) ;
  assign n14722 = n14721 ^ n10546 ^ n3860 ;
  assign n14723 = n14722 ^ n9730 ^ n2276 ;
  assign n14724 = ~n2673 & n7379 ;
  assign n14725 = ~n783 & n14724 ;
  assign n14726 = n8373 ^ n5344 ^ 1'b0 ;
  assign n14727 = n14725 & ~n14726 ;
  assign n14728 = n14727 ^ n8618 ^ n3551 ;
  assign n14729 = n4821 ^ n3251 ^ n2027 ;
  assign n14730 = n13994 ^ n7658 ^ 1'b0 ;
  assign n14731 = n6164 & n14730 ;
  assign n14732 = n6417 & n14731 ;
  assign n14736 = n4749 & n12798 ;
  assign n14737 = ~x248 & n14736 ;
  assign n14738 = n5585 | n5938 ;
  assign n14739 = n14737 & ~n14738 ;
  assign n14735 = n12683 ^ n8729 ^ n1529 ;
  assign n14740 = n14739 ^ n14735 ^ 1'b0 ;
  assign n14733 = n9174 ^ n4079 ^ n1063 ;
  assign n14734 = n13904 & n14733 ;
  assign n14741 = n14740 ^ n14734 ^ 1'b0 ;
  assign n14742 = ( n2905 & n7341 ) | ( n2905 & n14741 ) | ( n7341 & n14741 ) ;
  assign n14743 = n2925 & ~n14742 ;
  assign n14744 = n14732 & n14743 ;
  assign n14749 = ( ~n903 & n3792 ) | ( ~n903 & n7518 ) | ( n3792 & n7518 ) ;
  assign n14745 = n1897 ^ n516 ^ 1'b0 ;
  assign n14746 = n13439 ^ n10230 ^ 1'b0 ;
  assign n14747 = n14745 & ~n14746 ;
  assign n14748 = ~n10695 & n14747 ;
  assign n14750 = n14749 ^ n14748 ^ 1'b0 ;
  assign n14751 = n14750 ^ n4959 ^ 1'b0 ;
  assign n14752 = n3407 & ~n14751 ;
  assign n14753 = ( n4842 & n13626 ) | ( n4842 & ~n14752 ) | ( n13626 & ~n14752 ) ;
  assign n14754 = n2116 | n2779 ;
  assign n14755 = n14753 & ~n14754 ;
  assign n14763 = ( ~n1981 & n7317 ) | ( ~n1981 & n11414 ) | ( n7317 & n11414 ) ;
  assign n14757 = n5508 | n14267 ;
  assign n14758 = n14757 ^ n6150 ^ 1'b0 ;
  assign n14759 = n2333 | n14758 ;
  assign n14760 = n11117 ^ n5116 ^ n3814 ;
  assign n14761 = n6336 & n14760 ;
  assign n14762 = ~n14759 & n14761 ;
  assign n14764 = n14763 ^ n14762 ^ n13075 ;
  assign n14756 = n581 | n5522 ;
  assign n14765 = n14764 ^ n14756 ^ 1'b0 ;
  assign n14766 = ( n294 & n1749 ) | ( n294 & n2985 ) | ( n1749 & n2985 ) ;
  assign n14767 = n14766 ^ x101 ^ 1'b0 ;
  assign n14768 = ~n1176 & n14767 ;
  assign n14769 = ~n9120 & n14768 ;
  assign n14777 = ~n4398 & n8926 ;
  assign n14778 = n14777 ^ n12991 ^ 1'b0 ;
  assign n14773 = n4251 ^ n1236 ^ 1'b0 ;
  assign n14774 = n5953 & ~n14773 ;
  assign n14771 = n12805 ^ n2832 ^ n1597 ;
  assign n14772 = n7260 & n14771 ;
  assign n14775 = n14774 ^ n14772 ^ 1'b0 ;
  assign n14770 = n259 | n7558 ;
  assign n14776 = n14775 ^ n14770 ^ 1'b0 ;
  assign n14779 = n14778 ^ n14776 ^ x234 ;
  assign n14780 = n13864 ^ n5135 ^ n2697 ;
  assign n14781 = n4719 & ~n14780 ;
  assign n14782 = n14781 ^ x219 ^ 1'b0 ;
  assign n14783 = n14782 ^ n10721 ^ 1'b0 ;
  assign n14784 = n2082 | n4183 ;
  assign n14785 = n2184 | n14784 ;
  assign n14786 = n9016 ^ n4856 ^ 1'b0 ;
  assign n14790 = n3266 ^ n2785 ^ n1454 ;
  assign n14791 = ( n3974 & n7800 ) | ( n3974 & n14790 ) | ( n7800 & n14790 ) ;
  assign n14792 = ( ~n3250 & n3771 ) | ( ~n3250 & n14791 ) | ( n3771 & n14791 ) ;
  assign n14787 = n1403 ^ n1250 ^ n865 ;
  assign n14788 = n5439 & n14787 ;
  assign n14789 = n14788 ^ n481 ^ 1'b0 ;
  assign n14793 = n14792 ^ n14789 ^ n9610 ;
  assign n14794 = n11629 | n14793 ;
  assign n14795 = n7190 | n14794 ;
  assign n14796 = n14786 | n14795 ;
  assign n14797 = n2540 | n14796 ;
  assign n14798 = ( n4137 & n6669 ) | ( n4137 & ~n14362 ) | ( n6669 & ~n14362 ) ;
  assign n14799 = n5065 & n6174 ;
  assign n14800 = n14799 ^ n12467 ^ n2639 ;
  assign n14801 = x226 & n5817 ;
  assign n14802 = ~n367 & n14801 ;
  assign n14803 = n14802 ^ n4224 ^ 1'b0 ;
  assign n14804 = n6955 | n14803 ;
  assign n14805 = n14804 ^ n6941 ^ n2955 ;
  assign n14806 = n13232 ^ n9177 ^ n8230 ;
  assign n14807 = n4987 ^ n3358 ^ x97 ;
  assign n14808 = n14807 ^ n3260 ^ n1645 ;
  assign n14809 = n12240 ^ n1244 ^ 1'b0 ;
  assign n14810 = n14808 | n14809 ;
  assign n14811 = n3535 & ~n14810 ;
  assign n14812 = n10408 | n14811 ;
  assign n14813 = ( n13903 & n14806 ) | ( n13903 & ~n14812 ) | ( n14806 & ~n14812 ) ;
  assign n14821 = n2524 ^ n1559 ^ 1'b0 ;
  assign n14818 = n3392 & n9271 ;
  assign n14819 = ~n4634 & n14818 ;
  assign n14820 = n14819 ^ n10031 ^ 1'b0 ;
  assign n14814 = ~n6222 & n8766 ;
  assign n14815 = n2169 & n14814 ;
  assign n14816 = n14815 ^ n3209 ^ 1'b0 ;
  assign n14817 = n14816 ^ n14254 ^ n8099 ;
  assign n14822 = n14821 ^ n14820 ^ n14817 ;
  assign n14823 = ~n1325 & n12020 ;
  assign n14824 = n12075 & n14823 ;
  assign n14825 = n10739 & ~n14824 ;
  assign n14826 = n14825 ^ n14682 ^ 1'b0 ;
  assign n14827 = n3791 | n9647 ;
  assign n14828 = n12736 ^ n5357 ^ 1'b0 ;
  assign n14829 = n12046 ^ n8917 ^ n1913 ;
  assign n14830 = ~n1742 & n14829 ;
  assign n14831 = n12627 & n14830 ;
  assign n14832 = n4805 & n14831 ;
  assign n14833 = n11556 ^ n11251 ^ n10128 ;
  assign n14834 = n4858 ^ n832 ^ 1'b0 ;
  assign n14835 = ( n14832 & n14833 ) | ( n14832 & ~n14834 ) | ( n14833 & ~n14834 ) ;
  assign n14837 = n10761 ^ n2714 ^ 1'b0 ;
  assign n14838 = n5560 & ~n14837 ;
  assign n14836 = ( x142 & n4658 ) | ( x142 & n6636 ) | ( n4658 & n6636 ) ;
  assign n14839 = n14838 ^ n14836 ^ n12766 ;
  assign n14840 = n14839 ^ n9188 ^ 1'b0 ;
  assign n14841 = n3824 | n14840 ;
  assign n14842 = n14841 ^ n6430 ^ n879 ;
  assign n14843 = n6173 ^ n1964 ^ n1106 ;
  assign n14844 = n8527 ^ n4204 ^ 1'b0 ;
  assign n14845 = n665 & ~n14844 ;
  assign n14846 = n14843 & n14845 ;
  assign n14847 = n5193 & ~n11194 ;
  assign n14848 = ( n2899 & ~n3171 ) | ( n2899 & n4088 ) | ( ~n3171 & n4088 ) ;
  assign n14849 = n12485 ^ n1051 ^ 1'b0 ;
  assign n14850 = n14848 & ~n14849 ;
  assign n14851 = n14850 ^ n1438 ^ 1'b0 ;
  assign n14852 = ( n3739 & ~n6124 ) | ( n3739 & n6204 ) | ( ~n6124 & n6204 ) ;
  assign n14853 = n14852 ^ n11327 ^ n6983 ;
  assign n14854 = n14853 ^ n6818 ^ n950 ;
  assign n14855 = n3499 & ~n14854 ;
  assign n14856 = n7990 & n14855 ;
  assign n14858 = n7999 ^ n6823 ^ n6374 ;
  assign n14857 = n8059 | n8256 ;
  assign n14859 = n14858 ^ n14857 ^ n6901 ;
  assign n14860 = n11339 ^ n4067 ^ 1'b0 ;
  assign n14861 = n12371 & n14860 ;
  assign n14862 = n8427 & n11979 ;
  assign n14863 = n14695 ^ n10502 ^ 1'b0 ;
  assign n14864 = n14863 ^ n12995 ^ 1'b0 ;
  assign n14865 = n13394 & ~n14864 ;
  assign n14866 = n1352 & ~n11847 ;
  assign n14867 = n14866 ^ n6697 ^ n4670 ;
  assign n14868 = x203 & n5973 ;
  assign n14869 = n3844 | n14868 ;
  assign n14870 = n636 ^ n461 ^ 1'b0 ;
  assign n14871 = ~n4117 & n14870 ;
  assign n14872 = ~n6369 & n14871 ;
  assign n14873 = ( n6740 & ~n12726 ) | ( n6740 & n14872 ) | ( ~n12726 & n14872 ) ;
  assign n14874 = n14873 ^ n12050 ^ n4363 ;
  assign n14875 = n3722 & n14874 ;
  assign n14876 = n11737 ^ n7916 ^ 1'b0 ;
  assign n14877 = x71 & ~n3607 ;
  assign n14878 = n10278 ^ n770 ^ 1'b0 ;
  assign n14879 = n4349 ^ n2607 ^ 1'b0 ;
  assign n14880 = n2445 | n14879 ;
  assign n14881 = ( n3372 & ~n13905 ) | ( n3372 & n14633 ) | ( ~n13905 & n14633 ) ;
  assign n14882 = n2527 & ~n14881 ;
  assign n14883 = n14882 ^ n14461 ^ 1'b0 ;
  assign n14884 = n14883 ^ n6774 ^ 1'b0 ;
  assign n14885 = n3501 & n14884 ;
  assign n14886 = n4433 | n8888 ;
  assign n14887 = n14886 ^ n4832 ^ n1941 ;
  assign n14906 = ( n1020 & ~n4352 ) | ( n1020 & n4747 ) | ( ~n4352 & n4747 ) ;
  assign n14907 = ( n2233 & ~n7743 ) | ( n2233 & n14906 ) | ( ~n7743 & n14906 ) ;
  assign n14903 = n10926 ^ n5544 ^ 1'b0 ;
  assign n14904 = n9876 | n14903 ;
  assign n14905 = n14904 ^ n11185 ^ n2688 ;
  assign n14897 = n3015 ^ n1586 ^ 1'b0 ;
  assign n14895 = n2004 ^ n1964 ^ 1'b0 ;
  assign n14896 = ~n3374 & n14895 ;
  assign n14898 = n14897 ^ n14896 ^ 1'b0 ;
  assign n14899 = ( ~n1567 & n4066 ) | ( ~n1567 & n14898 ) | ( n4066 & n14898 ) ;
  assign n14900 = n8397 & ~n14899 ;
  assign n14894 = n4117 ^ n3992 ^ n2195 ;
  assign n14901 = n14900 ^ n14894 ^ n2588 ;
  assign n14890 = n14001 ^ n5730 ^ n3734 ;
  assign n14891 = n14890 ^ n9275 ^ 1'b0 ;
  assign n14888 = n14829 ^ n7352 ^ 1'b0 ;
  assign n14889 = n9954 & ~n14888 ;
  assign n14892 = n14891 ^ n14889 ^ 1'b0 ;
  assign n14893 = n2559 | n14892 ;
  assign n14902 = n14901 ^ n14893 ^ 1'b0 ;
  assign n14908 = n14907 ^ n14905 ^ n14902 ;
  assign n14909 = n5923 & n9915 ;
  assign n14910 = n13879 & ~n14909 ;
  assign n14911 = n14910 ^ n11508 ^ 1'b0 ;
  assign n14912 = n14478 & n14911 ;
  assign n14913 = ( n3701 & ~n4156 ) | ( n3701 & n9825 ) | ( ~n4156 & n9825 ) ;
  assign n14914 = n14913 ^ n4556 ^ n1773 ;
  assign n14915 = n1409 & ~n6500 ;
  assign n14916 = n6595 ^ n5680 ^ n1947 ;
  assign n14917 = n8169 ^ n3195 ^ 1'b0 ;
  assign n14918 = n14916 | n14917 ;
  assign n14919 = n14915 | n14918 ;
  assign n14920 = n14914 & n14919 ;
  assign n14921 = ~n2946 & n7860 ;
  assign n14922 = n3080 & n14921 ;
  assign n14923 = n287 | n861 ;
  assign n14924 = n14923 ^ n5093 ^ 1'b0 ;
  assign n14925 = ~n487 & n14924 ;
  assign n14926 = n14925 ^ n4470 ^ 1'b0 ;
  assign n14927 = n14926 ^ n4271 ^ 1'b0 ;
  assign n14928 = n6136 ^ n521 ^ 1'b0 ;
  assign n14929 = n7146 | n14928 ;
  assign n14930 = n8974 | n14929 ;
  assign n14931 = n5210 ^ n2573 ^ 1'b0 ;
  assign n14932 = ( n1265 & ~n3839 ) | ( n1265 & n5804 ) | ( ~n3839 & n5804 ) ;
  assign n14935 = ( n2654 & n4642 ) | ( n2654 & n5014 ) | ( n4642 & n5014 ) ;
  assign n14933 = n6097 & n9945 ;
  assign n14934 = n4121 & n14933 ;
  assign n14936 = n14935 ^ n14934 ^ 1'b0 ;
  assign n14937 = ( ~n10194 & n14932 ) | ( ~n10194 & n14936 ) | ( n14932 & n14936 ) ;
  assign n14938 = n4882 & n8362 ;
  assign n14939 = ~n10675 & n14938 ;
  assign n14940 = n3872 & n14939 ;
  assign n14941 = n5446 | n10688 ;
  assign n14942 = n13996 | n14941 ;
  assign n14943 = n7201 ^ n1140 ^ 1'b0 ;
  assign n14944 = x6 & ~n14943 ;
  assign n14945 = n6201 & n11534 ;
  assign n14946 = ~n14944 & n14945 ;
  assign n14947 = n10474 ^ n7318 ^ n1866 ;
  assign n14948 = ~n2782 & n7467 ;
  assign n14949 = n2500 & ~n14948 ;
  assign n14950 = n4502 & n14949 ;
  assign n14951 = ~n7458 & n14373 ;
  assign n14952 = n14951 ^ n13826 ^ 1'b0 ;
  assign n14953 = ( n13306 & ~n14950 ) | ( n13306 & n14952 ) | ( ~n14950 & n14952 ) ;
  assign n14954 = n14953 ^ n6438 ^ 1'b0 ;
  assign n14955 = n9405 ^ n6076 ^ n5992 ;
  assign n14956 = ~n5896 & n9134 ;
  assign n14957 = n14956 ^ n5388 ^ 1'b0 ;
  assign n14958 = ( n4144 & n6701 ) | ( n4144 & n12150 ) | ( n6701 & n12150 ) ;
  assign n14959 = n14958 ^ x24 ^ 1'b0 ;
  assign n14960 = n14959 ^ n12869 ^ 1'b0 ;
  assign n14961 = n13713 ^ n8802 ^ 1'b0 ;
  assign n14962 = n10207 & ~n14961 ;
  assign n14963 = n9739 ^ n5389 ^ 1'b0 ;
  assign n14964 = n14963 ^ n3720 ^ 1'b0 ;
  assign n14965 = n14962 & n14964 ;
  assign n14966 = n2620 & n2629 ;
  assign n14967 = n4409 ^ n3360 ^ 1'b0 ;
  assign n14968 = ~n1246 & n14967 ;
  assign n14969 = n7436 ^ n1863 ^ n337 ;
  assign n14970 = n2112 & n12838 ;
  assign n14971 = n2956 | n3240 ;
  assign n14972 = n12648 | n14971 ;
  assign n14973 = ~n6231 & n14972 ;
  assign n14974 = n926 & n14086 ;
  assign n14975 = n12026 ^ n10572 ^ x109 ;
  assign n14976 = n12656 & ~n14975 ;
  assign n14977 = n14976 ^ n10201 ^ 1'b0 ;
  assign n14978 = n11323 ^ n8099 ^ n4876 ;
  assign n14980 = n8551 ^ n2793 ^ 1'b0 ;
  assign n14981 = n5276 | n14980 ;
  assign n14979 = n11492 ^ n8045 ^ 1'b0 ;
  assign n14982 = n14981 ^ n14979 ^ 1'b0 ;
  assign n14987 = n5188 ^ n4163 ^ 1'b0 ;
  assign n14988 = ~n10252 & n14987 ;
  assign n14983 = n1786 & ~n2508 ;
  assign n14984 = n14983 ^ n4506 ^ 1'b0 ;
  assign n14985 = ( n6991 & n9430 ) | ( n6991 & ~n14984 ) | ( n9430 & ~n14984 ) ;
  assign n14986 = ~n10105 & n14985 ;
  assign n14989 = n14988 ^ n14986 ^ 1'b0 ;
  assign n14990 = ( n3736 & n10018 ) | ( n3736 & n11041 ) | ( n10018 & n11041 ) ;
  assign n14995 = ( n783 & n8397 ) | ( n783 & ~n9429 ) | ( n8397 & ~n9429 ) ;
  assign n14991 = n10769 ^ n4148 ^ n488 ;
  assign n14992 = n14991 ^ n11757 ^ 1'b0 ;
  assign n14993 = n14992 ^ n8421 ^ 1'b0 ;
  assign n14994 = x10 | n14993 ;
  assign n14996 = n14995 ^ n14994 ^ 1'b0 ;
  assign n14997 = n11169 ^ n9399 ^ 1'b0 ;
  assign n14998 = n9295 & n14997 ;
  assign n15000 = n9613 ^ n995 ^ 1'b0 ;
  assign n15001 = n6621 & ~n15000 ;
  assign n14999 = n5855 | n9379 ;
  assign n15002 = n15001 ^ n14999 ^ 1'b0 ;
  assign n15003 = ~x21 & n15002 ;
  assign n15004 = n15003 ^ n13703 ^ 1'b0 ;
  assign n15005 = n7129 & ~n8520 ;
  assign n15006 = ~n1086 & n8315 ;
  assign n15007 = ~n1678 & n15006 ;
  assign n15008 = n15007 ^ n1493 ^ x220 ;
  assign n15009 = ~n488 & n3364 ;
  assign n15010 = ~n2759 & n5017 ;
  assign n15011 = n9203 & n15010 ;
  assign n15012 = ( n15008 & n15009 ) | ( n15008 & n15011 ) | ( n15009 & n15011 ) ;
  assign n15013 = x21 & n15012 ;
  assign n15014 = n15005 & n15013 ;
  assign n15015 = n11901 ^ n5160 ^ 1'b0 ;
  assign n15016 = n10978 ^ n1576 ^ n1474 ;
  assign n15017 = n15016 ^ n10389 ^ 1'b0 ;
  assign n15018 = ~n1974 & n10127 ;
  assign n15019 = n3456 & n15018 ;
  assign n15020 = ( n838 & ~n8281 ) | ( n838 & n15019 ) | ( ~n8281 & n15019 ) ;
  assign n15021 = n15020 ^ n11030 ^ 1'b0 ;
  assign n15022 = n15021 ^ n9354 ^ 1'b0 ;
  assign n15023 = n12196 ^ n8024 ^ n2965 ;
  assign n15024 = ( n8450 & n11545 ) | ( n8450 & ~n14722 ) | ( n11545 & ~n14722 ) ;
  assign n15025 = n3413 & ~n7712 ;
  assign n15026 = n15025 ^ n8949 ^ 1'b0 ;
  assign n15028 = ~n276 & n2020 ;
  assign n15029 = n15028 ^ n3312 ^ 1'b0 ;
  assign n15027 = n1819 & ~n7836 ;
  assign n15030 = n15029 ^ n15027 ^ 1'b0 ;
  assign n15031 = n15030 ^ n4442 ^ 1'b0 ;
  assign n15032 = n11936 ^ n10559 ^ n5891 ;
  assign n15033 = n1591 & n12121 ;
  assign n15034 = n11789 & n15033 ;
  assign n15035 = n3359 ^ n1276 ^ 1'b0 ;
  assign n15036 = n6325 & ~n15035 ;
  assign n15037 = n15036 ^ n13776 ^ n11022 ;
  assign n15038 = ( n3903 & ~n15034 ) | ( n3903 & n15037 ) | ( ~n15034 & n15037 ) ;
  assign n15039 = n15038 ^ n3585 ^ 1'b0 ;
  assign n15040 = ~n15032 & n15039 ;
  assign n15041 = n3858 ^ n2170 ^ 1'b0 ;
  assign n15042 = ( n5336 & n11132 ) | ( n5336 & ~n15041 ) | ( n11132 & ~n15041 ) ;
  assign n15043 = n362 | n9424 ;
  assign n15044 = n15043 ^ n11047 ^ 1'b0 ;
  assign n15045 = n6420 | n15044 ;
  assign n15046 = n15042 | n15045 ;
  assign n15047 = n15046 ^ n13605 ^ 1'b0 ;
  assign n15048 = n15047 ^ n13092 ^ 1'b0 ;
  assign n15049 = n2607 | n15048 ;
  assign n15050 = n10926 ^ n9387 ^ 1'b0 ;
  assign n15051 = ~n8945 & n15050 ;
  assign n15052 = n8219 ^ n7947 ^ n5088 ;
  assign n15053 = n15052 ^ n1348 ^ 1'b0 ;
  assign n15054 = ( ~n4583 & n4781 ) | ( ~n4583 & n6924 ) | ( n4781 & n6924 ) ;
  assign n15055 = n15053 | n15054 ;
  assign n15056 = n15055 ^ n4208 ^ 1'b0 ;
  assign n15057 = n3313 & n3790 ;
  assign n15058 = ( n5264 & n15056 ) | ( n5264 & ~n15057 ) | ( n15056 & ~n15057 ) ;
  assign n15059 = n11398 ^ n7108 ^ n317 ;
  assign n15060 = n14635 ^ n4865 ^ 1'b0 ;
  assign n15061 = n14703 & n15060 ;
  assign n15062 = n3771 | n5100 ;
  assign n15063 = n15062 ^ n586 ^ 1'b0 ;
  assign n15064 = ( n8725 & n12561 ) | ( n8725 & ~n15063 ) | ( n12561 & ~n15063 ) ;
  assign n15065 = ~n1130 & n15064 ;
  assign n15066 = n13141 ^ n5436 ^ 1'b0 ;
  assign n15067 = n15066 ^ n5545 ^ n4982 ;
  assign n15068 = n2602 ^ x93 ^ 1'b0 ;
  assign n15069 = n15068 ^ n4858 ^ x240 ;
  assign n15070 = n1917 & ~n15069 ;
  assign n15071 = ~n15067 & n15070 ;
  assign n15072 = ~n346 & n9014 ;
  assign n15073 = n2783 ^ n1932 ^ 1'b0 ;
  assign n15074 = n11420 | n15073 ;
  assign n15075 = n15074 ^ n11011 ^ n5427 ;
  assign n15076 = ~n726 & n7686 ;
  assign n15077 = n15076 ^ n1604 ^ 1'b0 ;
  assign n15078 = n1493 ^ n324 ^ 1'b0 ;
  assign n15079 = n15078 ^ n1050 ^ 1'b0 ;
  assign n15080 = n15077 & n15079 ;
  assign n15083 = x129 & ~n4284 ;
  assign n15084 = n2050 & n15083 ;
  assign n15081 = n1018 | n4849 ;
  assign n15082 = n2119 & n15081 ;
  assign n15085 = n15084 ^ n15082 ^ 1'b0 ;
  assign n15086 = ( n2724 & n7007 ) | ( n2724 & n12230 ) | ( n7007 & n12230 ) ;
  assign n15087 = ~n3994 & n4773 ;
  assign n15088 = ( x179 & ~n10422 ) | ( x179 & n15087 ) | ( ~n10422 & n15087 ) ;
  assign n15089 = n5567 ^ n3116 ^ 1'b0 ;
  assign n15093 = n5681 & n6759 ;
  assign n15090 = n4417 & n10038 ;
  assign n15091 = n15090 ^ n3453 ^ 1'b0 ;
  assign n15092 = n4065 & n15091 ;
  assign n15094 = n15093 ^ n15092 ^ 1'b0 ;
  assign n15095 = n13046 ^ n845 ^ 1'b0 ;
  assign n15096 = n10088 & ~n15095 ;
  assign n15097 = n2014 | n2463 ;
  assign n15098 = n15097 ^ n393 ^ 1'b0 ;
  assign n15099 = ~n7139 & n14411 ;
  assign n15100 = n10265 & n15099 ;
  assign n15101 = ( n11727 & n15098 ) | ( n11727 & n15100 ) | ( n15098 & n15100 ) ;
  assign n15102 = n12974 ^ n10463 ^ 1'b0 ;
  assign n15103 = ~n7283 & n15102 ;
  assign n15104 = ( n3441 & n6270 ) | ( n3441 & ~n7897 ) | ( n6270 & ~n7897 ) ;
  assign n15105 = ( n3578 & n11132 ) | ( n3578 & n15104 ) | ( n11132 & n15104 ) ;
  assign n15106 = n15105 ^ n6074 ^ 1'b0 ;
  assign n15107 = ~n7870 & n11505 ;
  assign n15108 = n4800 & ~n13599 ;
  assign n15109 = n15108 ^ n13359 ^ 1'b0 ;
  assign n15110 = n14097 ^ n8615 ^ 1'b0 ;
  assign n15111 = ~n12444 & n15110 ;
  assign n15117 = n1649 | n3682 ;
  assign n15118 = n15117 ^ x133 ^ 1'b0 ;
  assign n15116 = n14671 ^ n4410 ^ 1'b0 ;
  assign n15112 = n13693 ^ n6304 ^ n3237 ;
  assign n15113 = n5473 & n14377 ;
  assign n15114 = n12262 & ~n15113 ;
  assign n15115 = ~n15112 & n15114 ;
  assign n15119 = n15118 ^ n15116 ^ n15115 ;
  assign n15120 = n8376 ^ n1783 ^ n566 ;
  assign n15121 = n15120 ^ n8557 ^ 1'b0 ;
  assign n15125 = ( n4896 & n12344 ) | ( n4896 & ~n12814 ) | ( n12344 & ~n12814 ) ;
  assign n15122 = n7947 & n14262 ;
  assign n15123 = ~n2164 & n15122 ;
  assign n15124 = n6893 | n15123 ;
  assign n15126 = n15125 ^ n15124 ^ 1'b0 ;
  assign n15127 = n9756 | n12595 ;
  assign n15128 = ( n10186 & ~n10199 ) | ( n10186 & n13497 ) | ( ~n10199 & n13497 ) ;
  assign n15129 = n2270 & n6653 ;
  assign n15132 = n11503 ^ n10393 ^ n8779 ;
  assign n15130 = n7463 ^ n2732 ^ 1'b0 ;
  assign n15131 = n8296 & ~n15130 ;
  assign n15133 = n15132 ^ n15131 ^ 1'b0 ;
  assign n15134 = n2573 | n12278 ;
  assign n15135 = ~n9394 & n15134 ;
  assign n15136 = n8640 & n15135 ;
  assign n15137 = n15136 ^ n10158 ^ n1632 ;
  assign n15138 = ( n4996 & n15133 ) | ( n4996 & n15137 ) | ( n15133 & n15137 ) ;
  assign n15139 = n4711 & n10072 ;
  assign n15140 = n15139 ^ n1663 ^ 1'b0 ;
  assign n15141 = n1943 & n15140 ;
  assign n15142 = n11727 ^ n5775 ^ 1'b0 ;
  assign n15143 = n644 & n10268 ;
  assign n15144 = ( n14401 & n15142 ) | ( n14401 & ~n15143 ) | ( n15142 & ~n15143 ) ;
  assign n15145 = n3054 ^ n2436 ^ 1'b0 ;
  assign n15146 = n15144 | n15145 ;
  assign n15149 = ( n6511 & n11157 ) | ( n6511 & n12500 ) | ( n11157 & n12500 ) ;
  assign n15147 = x126 & n14568 ;
  assign n15148 = ( x7 & n2613 ) | ( x7 & n15147 ) | ( n2613 & n15147 ) ;
  assign n15150 = n15149 ^ n15148 ^ n4123 ;
  assign n15151 = ~n1619 & n4604 ;
  assign n15152 = ~n1395 & n15151 ;
  assign n15153 = n15152 ^ n10204 ^ n7217 ;
  assign n15154 = ~n10225 & n15153 ;
  assign n15155 = n10076 ^ n7846 ^ 1'b0 ;
  assign n15156 = n15155 ^ n11955 ^ n1029 ;
  assign n15157 = n12887 ^ n6718 ^ n4921 ;
  assign n15158 = n15157 ^ n2785 ^ 1'b0 ;
  assign n15159 = n15156 & n15158 ;
  assign n15160 = n6814 | n9500 ;
  assign n15161 = n12653 ^ n7481 ^ 1'b0 ;
  assign n15162 = ( n871 & ~n10191 ) | ( n871 & n15161 ) | ( ~n10191 & n15161 ) ;
  assign n15163 = n15162 ^ n8185 ^ n5712 ;
  assign n15167 = x121 & n2380 ;
  assign n15165 = n14792 ^ n4254 ^ 1'b0 ;
  assign n15166 = n10367 & n15165 ;
  assign n15164 = n261 | n2440 ;
  assign n15168 = n15167 ^ n15166 ^ n15164 ;
  assign n15169 = x114 & n6458 ;
  assign n15170 = n3026 & n15169 ;
  assign n15171 = n11231 ^ n8951 ^ 1'b0 ;
  assign n15172 = ~n15170 & n15171 ;
  assign n15173 = n8658 ^ n7211 ^ n1607 ;
  assign n15174 = x2 & ~n13718 ;
  assign n15175 = n2623 ^ n874 ^ 1'b0 ;
  assign n15176 = ~n10984 & n15175 ;
  assign n15177 = ~n15174 & n15176 ;
  assign n15178 = ( n14226 & ~n15173 ) | ( n14226 & n15177 ) | ( ~n15173 & n15177 ) ;
  assign n15179 = ~n9456 & n10659 ;
  assign n15180 = n7228 & n15179 ;
  assign n15181 = n15180 ^ n8619 ^ n6045 ;
  assign n15182 = n1285 ^ n482 ^ 1'b0 ;
  assign n15183 = n7314 & n15182 ;
  assign n15184 = ~x93 & n4530 ;
  assign n15185 = n15184 ^ n2310 ^ n1220 ;
  assign n15186 = n8977 & n15185 ;
  assign n15187 = ~n15183 & n15186 ;
  assign n15192 = n1953 | n7172 ;
  assign n15193 = n9765 & ~n15192 ;
  assign n15188 = ~n2704 & n5500 ;
  assign n15189 = n15188 ^ n13239 ^ 1'b0 ;
  assign n15190 = n681 | n15189 ;
  assign n15191 = n15190 ^ n11883 ^ 1'b0 ;
  assign n15194 = n15193 ^ n15191 ^ 1'b0 ;
  assign n15195 = n305 & n4895 ;
  assign n15196 = n15195 ^ n657 ^ 1'b0 ;
  assign n15197 = n15196 ^ n13309 ^ n9756 ;
  assign n15198 = ( n6037 & ~n8740 ) | ( n6037 & n13657 ) | ( ~n8740 & n13657 ) ;
  assign n15199 = n1068 | n6752 ;
  assign n15200 = n1986 ^ n1883 ^ n1277 ;
  assign n15201 = n3347 | n7538 ;
  assign n15202 = n2518 & ~n15201 ;
  assign n15203 = n15202 ^ n8613 ^ n1841 ;
  assign n15204 = n15203 ^ n14586 ^ 1'b0 ;
  assign n15205 = ~n15200 & n15204 ;
  assign n15206 = n1903 | n3933 ;
  assign n15207 = n11802 | n15206 ;
  assign n15208 = n15207 ^ n9195 ^ 1'b0 ;
  assign n15209 = n8231 ^ n7163 ^ n2726 ;
  assign n15217 = n7464 ^ n3728 ^ 1'b0 ;
  assign n15211 = n3617 ^ n3602 ^ 1'b0 ;
  assign n15212 = n892 & ~n15211 ;
  assign n15213 = ( n816 & n10210 ) | ( n816 & ~n15212 ) | ( n10210 & ~n15212 ) ;
  assign n15214 = n15213 ^ n7750 ^ n1981 ;
  assign n15210 = ~n4066 & n13516 ;
  assign n15215 = n15214 ^ n15210 ^ 1'b0 ;
  assign n15216 = n11564 | n15215 ;
  assign n15218 = n15217 ^ n15216 ^ 1'b0 ;
  assign n15219 = n6523 ^ n1180 ^ 1'b0 ;
  assign n15220 = n15219 ^ n6472 ^ 1'b0 ;
  assign n15221 = n9947 ^ n9260 ^ n6677 ;
  assign n15223 = ( n8969 & ~n13088 ) | ( n8969 & n14274 ) | ( ~n13088 & n14274 ) ;
  assign n15222 = n857 | n9697 ;
  assign n15224 = n15223 ^ n15222 ^ 1'b0 ;
  assign n15225 = ( n15220 & n15221 ) | ( n15220 & ~n15224 ) | ( n15221 & ~n15224 ) ;
  assign n15232 = ( ~x67 & n3463 ) | ( ~x67 & n6043 ) | ( n3463 & n6043 ) ;
  assign n15228 = n5637 ^ n5566 ^ n2878 ;
  assign n15226 = n2912 ^ n490 ^ 1'b0 ;
  assign n15227 = n3788 | n15226 ;
  assign n15229 = n15228 ^ n15227 ^ 1'b0 ;
  assign n15230 = n7176 | n15229 ;
  assign n15231 = n15230 ^ n9555 ^ n1720 ;
  assign n15233 = n15232 ^ n15231 ^ n13137 ;
  assign n15234 = n7369 ^ n2340 ^ 1'b0 ;
  assign n15235 = n9178 ^ n7879 ^ 1'b0 ;
  assign n15236 = n15234 | n15235 ;
  assign n15237 = ( n1734 & ~n4124 ) | ( n1734 & n5221 ) | ( ~n4124 & n5221 ) ;
  assign n15238 = n5514 ^ n1537 ^ x113 ;
  assign n15239 = n6199 | n15238 ;
  assign n15240 = n14435 & ~n15239 ;
  assign n15241 = n6705 | n15240 ;
  assign n15242 = n2719 | n15241 ;
  assign n15243 = n13994 ^ n3763 ^ 1'b0 ;
  assign n15244 = n374 & n15243 ;
  assign n15245 = n15244 ^ n11951 ^ n5284 ;
  assign n15246 = n448 | n1281 ;
  assign n15247 = n274 & ~n15246 ;
  assign n15248 = n3377 & ~n15247 ;
  assign n15249 = n15248 ^ n12728 ^ n4057 ;
  assign n15250 = ( n3298 & n11140 ) | ( n3298 & ~n15249 ) | ( n11140 & ~n15249 ) ;
  assign n15251 = n11321 ^ n7184 ^ n757 ;
  assign n15252 = n6597 | n15251 ;
  assign n15253 = n3129 ^ n2843 ^ 1'b0 ;
  assign n15254 = n4773 & ~n15253 ;
  assign n15255 = n15254 ^ n8735 ^ 1'b0 ;
  assign n15256 = n15252 & n15255 ;
  assign n15257 = ~n7616 & n10978 ;
  assign n15258 = n11768 & n15257 ;
  assign n15259 = ~n2899 & n3739 ;
  assign n15260 = n15259 ^ n6441 ^ 1'b0 ;
  assign n15261 = n12084 & ~n15260 ;
  assign n15262 = ~n13386 & n15261 ;
  assign n15263 = n15258 | n15262 ;
  assign n15264 = n15263 ^ n1703 ^ 1'b0 ;
  assign n15265 = n7685 | n11753 ;
  assign n15266 = n4712 | n15265 ;
  assign n15267 = n15266 ^ n376 ^ n352 ;
  assign n15272 = n8398 ^ n3496 ^ 1'b0 ;
  assign n15268 = n2256 & ~n3331 ;
  assign n15269 = ~n2083 & n15268 ;
  assign n15270 = n449 | n15269 ;
  assign n15271 = n15270 ^ n962 ^ 1'b0 ;
  assign n15273 = n15272 ^ n15271 ^ n4619 ;
  assign n15274 = n605 ^ x23 ^ 1'b0 ;
  assign n15275 = n15274 ^ n6246 ^ 1'b0 ;
  assign n15276 = ~n15273 & n15275 ;
  assign n15277 = n15276 ^ n13921 ^ n13890 ;
  assign n15278 = n6889 & ~n13019 ;
  assign n15281 = x138 & n2036 ;
  assign n15279 = n1776 & n9363 ;
  assign n15280 = ~n10538 & n15279 ;
  assign n15282 = n15281 ^ n15280 ^ n12622 ;
  assign n15283 = n11066 ^ n4797 ^ 1'b0 ;
  assign n15284 = n15283 ^ n14704 ^ n12459 ;
  assign n15285 = ( n904 & ~n1778 ) | ( n904 & n10079 ) | ( ~n1778 & n10079 ) ;
  assign n15286 = n3507 & n15285 ;
  assign n15287 = ~n1221 & n9316 ;
  assign n15288 = n518 & n15287 ;
  assign n15292 = n2968 & ~n6478 ;
  assign n15289 = ~n3851 & n12198 ;
  assign n15290 = ~n14690 & n15289 ;
  assign n15291 = ( n5849 & ~n9013 ) | ( n5849 & n15290 ) | ( ~n9013 & n15290 ) ;
  assign n15293 = n15292 ^ n15291 ^ n8885 ;
  assign n15294 = ( n3144 & n4280 ) | ( n3144 & ~n4316 ) | ( n4280 & ~n4316 ) ;
  assign n15295 = ~n1922 & n15294 ;
  assign n15296 = n15295 ^ n9904 ^ 1'b0 ;
  assign n15297 = n3083 | n15296 ;
  assign n15302 = n7836 ^ n5208 ^ 1'b0 ;
  assign n15303 = n4660 | n15302 ;
  assign n15304 = n15303 ^ n8625 ^ 1'b0 ;
  assign n15298 = ( ~n3111 & n4605 ) | ( ~n3111 & n5151 ) | ( n4605 & n5151 ) ;
  assign n15299 = x11 & ~x82 ;
  assign n15300 = ~n15298 & n15299 ;
  assign n15301 = n15300 ^ n867 ^ 1'b0 ;
  assign n15305 = n15304 ^ n15301 ^ n7153 ;
  assign n15306 = n7616 | n15305 ;
  assign n15307 = n15306 ^ n9665 ^ 1'b0 ;
  assign n15308 = ( n1573 & n2655 ) | ( n1573 & n4405 ) | ( n2655 & n4405 ) ;
  assign n15309 = n15308 ^ n6848 ^ n1281 ;
  assign n15310 = ~n14586 & n15309 ;
  assign n15311 = ~n3872 & n9658 ;
  assign n15312 = n15311 ^ n9377 ^ 1'b0 ;
  assign n15313 = n15312 ^ n5235 ^ n4306 ;
  assign n15314 = ~n843 & n3599 ;
  assign n15315 = n6876 ^ x42 ^ 1'b0 ;
  assign n15316 = n15315 ^ n12715 ^ 1'b0 ;
  assign n15317 = n15016 & n15316 ;
  assign n15318 = ( ~n15036 & n15314 ) | ( ~n15036 & n15317 ) | ( n15314 & n15317 ) ;
  assign n15319 = n7900 ^ n1581 ^ 1'b0 ;
  assign n15320 = ( n3796 & n11389 ) | ( n3796 & n15319 ) | ( n11389 & n15319 ) ;
  assign n15321 = ( ~n1451 & n6027 ) | ( ~n1451 & n12477 ) | ( n6027 & n12477 ) ;
  assign n15322 = n4329 ^ n2096 ^ x215 ;
  assign n15323 = n15322 ^ n6215 ^ 1'b0 ;
  assign n15324 = n15323 ^ n8741 ^ 1'b0 ;
  assign n15325 = n3144 & n15324 ;
  assign n15326 = ( ~n15320 & n15321 ) | ( ~n15320 & n15325 ) | ( n15321 & n15325 ) ;
  assign n15327 = ( ~n317 & n956 ) | ( ~n317 & n2657 ) | ( n956 & n2657 ) ;
  assign n15328 = ( n5710 & n9406 ) | ( n5710 & n15327 ) | ( n9406 & n15327 ) ;
  assign n15329 = n11327 & n11657 ;
  assign n15330 = ( n4459 & ~n5938 ) | ( n4459 & n11927 ) | ( ~n5938 & n11927 ) ;
  assign n15331 = n15330 ^ n7417 ^ 1'b0 ;
  assign n15332 = n6971 ^ n4484 ^ n2697 ;
  assign n15333 = n5257 ^ n1146 ^ n716 ;
  assign n15334 = ( n626 & n5416 ) | ( n626 & ~n5895 ) | ( n5416 & ~n5895 ) ;
  assign n15335 = ( ~n2639 & n13405 ) | ( ~n2639 & n15334 ) | ( n13405 & n15334 ) ;
  assign n15336 = n4826 & n15335 ;
  assign n15337 = n1598 & n8306 ;
  assign n15338 = n1837 & ~n8502 ;
  assign n15339 = ~n561 & n15338 ;
  assign n15340 = n5959 | n15339 ;
  assign n15341 = ( ~n15320 & n15337 ) | ( ~n15320 & n15340 ) | ( n15337 & n15340 ) ;
  assign n15342 = n10595 ^ n8298 ^ n3220 ;
  assign n15343 = n3530 ^ n1395 ^ 1'b0 ;
  assign n15344 = n11140 & ~n15343 ;
  assign n15345 = n15344 ^ n7735 ^ n6837 ;
  assign n15346 = n10848 ^ n6714 ^ 1'b0 ;
  assign n15347 = n2773 & n15346 ;
  assign n15348 = n2370 ^ x243 ^ 1'b0 ;
  assign n15349 = n15348 ^ n7406 ^ 1'b0 ;
  assign n15350 = n15347 & ~n15349 ;
  assign n15351 = n5819 & ~n15350 ;
  assign n15352 = ( n4341 & n15345 ) | ( n4341 & ~n15351 ) | ( n15345 & ~n15351 ) ;
  assign n15353 = n5438 | n15352 ;
  assign n15354 = ( ~n1607 & n7308 ) | ( ~n1607 & n14872 ) | ( n7308 & n14872 ) ;
  assign n15355 = ~n9808 & n15354 ;
  assign n15356 = n12045 ^ n7433 ^ 1'b0 ;
  assign n15357 = n3116 & n11925 ;
  assign n15358 = n836 | n5857 ;
  assign n15359 = n13303 | n15358 ;
  assign n15360 = n7746 & ~n15359 ;
  assign n15361 = ( n3177 & n15357 ) | ( n3177 & n15360 ) | ( n15357 & n15360 ) ;
  assign n15362 = ( ~n2343 & n3459 ) | ( ~n2343 & n4924 ) | ( n3459 & n4924 ) ;
  assign n15363 = n4327 ^ n2653 ^ 1'b0 ;
  assign n15364 = n15362 | n15363 ;
  assign n15365 = ~n2839 & n4698 ;
  assign n15366 = n11660 & ~n15365 ;
  assign n15367 = ~n1250 & n15366 ;
  assign n15368 = n15367 ^ n15168 ^ n8566 ;
  assign n15369 = n9921 ^ n1315 ^ 1'b0 ;
  assign n15370 = n15168 & n15369 ;
  assign n15372 = ( n6326 & n7784 ) | ( n6326 & n12921 ) | ( n7784 & n12921 ) ;
  assign n15371 = n12333 & ~n14205 ;
  assign n15373 = n15372 ^ n15371 ^ 1'b0 ;
  assign n15374 = n7211 & ~n7962 ;
  assign n15375 = n6653 & n15374 ;
  assign n15376 = n15375 ^ n5749 ^ 1'b0 ;
  assign n15377 = ~n3440 & n15376 ;
  assign n15378 = n15377 ^ n15258 ^ 1'b0 ;
  assign n15379 = n15378 ^ x140 ^ 1'b0 ;
  assign n15380 = n9549 ^ n9425 ^ 1'b0 ;
  assign n15385 = n3689 ^ n3034 ^ 1'b0 ;
  assign n15386 = n821 & ~n15385 ;
  assign n15381 = n5634 ^ n1351 ^ 1'b0 ;
  assign n15382 = ~n11253 & n15381 ;
  assign n15383 = n10909 ^ n2752 ^ 1'b0 ;
  assign n15384 = n15382 & ~n15383 ;
  assign n15387 = n15386 ^ n15384 ^ 1'b0 ;
  assign n15388 = ~n4382 & n15387 ;
  assign n15389 = ~n13226 & n15388 ;
  assign n15390 = ~n6725 & n13338 ;
  assign n15391 = n10663 ^ n3498 ^ 1'b0 ;
  assign n15392 = n15391 ^ n6079 ^ 1'b0 ;
  assign n15393 = n1062 & ~n8518 ;
  assign n15394 = n15393 ^ n4966 ^ 1'b0 ;
  assign n15395 = n15394 ^ n5236 ^ 1'b0 ;
  assign n15397 = n8790 ^ n4481 ^ 1'b0 ;
  assign n15396 = n5292 & ~n6956 ;
  assign n15398 = n15397 ^ n15396 ^ 1'b0 ;
  assign n15399 = n955 & n7519 ;
  assign n15400 = n1924 & n10829 ;
  assign n15401 = ~n15399 & n15400 ;
  assign n15402 = n558 & ~n6931 ;
  assign n15403 = n15402 ^ n3930 ^ 1'b0 ;
  assign n15404 = ( x115 & n2785 ) | ( x115 & n7589 ) | ( n2785 & n7589 ) ;
  assign n15405 = n8297 & ~n15404 ;
  assign n15406 = n15405 ^ n6277 ^ 1'b0 ;
  assign n15407 = n9717 & ~n12166 ;
  assign n15410 = n5326 ^ n1698 ^ 1'b0 ;
  assign n15408 = n8047 ^ n1805 ^ 1'b0 ;
  assign n15409 = n14140 | n15408 ;
  assign n15411 = n15410 ^ n15409 ^ n12697 ;
  assign n15412 = ~n2216 & n9812 ;
  assign n15413 = ~n6901 & n15412 ;
  assign n15414 = n11827 ^ n4306 ^ n576 ;
  assign n15415 = ( n2104 & n15413 ) | ( n2104 & n15414 ) | ( n15413 & n15414 ) ;
  assign n15417 = n2500 ^ n1199 ^ 1'b0 ;
  assign n15418 = n11173 & ~n15417 ;
  assign n15416 = n3739 & ~n14258 ;
  assign n15419 = n15418 ^ n15416 ^ 1'b0 ;
  assign n15420 = n10191 ^ n5622 ^ 1'b0 ;
  assign n15421 = ~n15419 & n15420 ;
  assign n15422 = n1164 & n12217 ;
  assign n15424 = n5332 ^ n4480 ^ n3374 ;
  assign n15425 = n15424 ^ n5974 ^ n3321 ;
  assign n15426 = ( n4806 & n15347 ) | ( n4806 & n15425 ) | ( n15347 & n15425 ) ;
  assign n15427 = n8142 & n15426 ;
  assign n15428 = n15427 ^ n10540 ^ 1'b0 ;
  assign n15429 = n2663 & ~n15428 ;
  assign n15430 = ~n5529 & n15429 ;
  assign n15431 = n7978 | n15430 ;
  assign n15432 = n3276 & ~n15431 ;
  assign n15423 = n6397 | n13339 ;
  assign n15433 = n15432 ^ n15423 ^ 1'b0 ;
  assign n15434 = n14633 ^ n8779 ^ 1'b0 ;
  assign n15435 = n11294 | n15434 ;
  assign n15436 = n15435 ^ n3954 ^ 1'b0 ;
  assign n15437 = n6781 & ~n11031 ;
  assign n15438 = n15436 & n15437 ;
  assign n15439 = ( ~n15422 & n15433 ) | ( ~n15422 & n15438 ) | ( n15433 & n15438 ) ;
  assign n15440 = ~n3748 & n10007 ;
  assign n15441 = n15440 ^ n1688 ^ 1'b0 ;
  assign n15443 = ( n4402 & n7043 ) | ( n4402 & ~n7293 ) | ( n7043 & ~n7293 ) ;
  assign n15442 = n809 & ~n6753 ;
  assign n15444 = n15443 ^ n15442 ^ 1'b0 ;
  assign n15445 = ~n3780 & n6329 ;
  assign n15446 = n5618 & n15445 ;
  assign n15447 = x82 & n12605 ;
  assign n15448 = ~n10559 & n15447 ;
  assign n15449 = n15448 ^ n8906 ^ 1'b0 ;
  assign n15450 = n15140 & ~n15449 ;
  assign n15451 = ( ~n14755 & n15446 ) | ( ~n14755 & n15450 ) | ( n15446 & n15450 ) ;
  assign n15452 = ( ~n3099 & n6430 ) | ( ~n3099 & n6683 ) | ( n6430 & n6683 ) ;
  assign n15453 = ( n4983 & n7223 ) | ( n4983 & n15452 ) | ( n7223 & n15452 ) ;
  assign n15454 = n5300 ^ n4624 ^ 1'b0 ;
  assign n15455 = n13467 ^ n9853 ^ 1'b0 ;
  assign n15456 = n11811 & ~n15455 ;
  assign n15457 = n15456 ^ n13957 ^ 1'b0 ;
  assign n15458 = ( x156 & n9788 ) | ( x156 & ~n14105 ) | ( n9788 & ~n14105 ) ;
  assign n15459 = n15458 ^ n6338 ^ 1'b0 ;
  assign n15460 = ( n1086 & n3745 ) | ( n1086 & n10846 ) | ( n3745 & n10846 ) ;
  assign n15461 = n3200 | n15460 ;
  assign n15462 = n8315 | n15461 ;
  assign n15463 = n15462 ^ n1367 ^ 1'b0 ;
  assign n15464 = n15463 ^ n9840 ^ n3991 ;
  assign n15465 = n4036 ^ n728 ^ x173 ;
  assign n15466 = n3527 ^ n2445 ^ n939 ;
  assign n15467 = n15466 ^ n7823 ^ 1'b0 ;
  assign n15468 = n12397 ^ n8247 ^ n3060 ;
  assign n15469 = n3568 ^ n982 ^ 1'b0 ;
  assign n15470 = n12803 & ~n15469 ;
  assign n15471 = n15470 ^ n5357 ^ 1'b0 ;
  assign n15472 = n1723 | n6362 ;
  assign n15473 = n15472 ^ n6402 ^ 1'b0 ;
  assign n15474 = ~n3930 & n14984 ;
  assign n15475 = ~n15473 & n15474 ;
  assign n15477 = n4136 ^ n3393 ^ n2171 ;
  assign n15478 = n15477 ^ n7044 ^ n449 ;
  assign n15476 = ( n3857 & ~n6142 ) | ( n3857 & n10615 ) | ( ~n6142 & n10615 ) ;
  assign n15479 = n15478 ^ n15476 ^ 1'b0 ;
  assign n15480 = n13718 & n15479 ;
  assign n15481 = n15480 ^ n13960 ^ n9109 ;
  assign n15482 = ~n585 & n2376 ;
  assign n15483 = n521 & ~n9576 ;
  assign n15484 = n3280 & n15483 ;
  assign n15485 = ( ~n10641 & n15482 ) | ( ~n10641 & n15484 ) | ( n15482 & n15484 ) ;
  assign n15486 = ( n1212 & ~n5513 ) | ( n1212 & n15485 ) | ( ~n5513 & n15485 ) ;
  assign n15487 = ( n8945 & n9044 ) | ( n8945 & n13927 ) | ( n9044 & n13927 ) ;
  assign n15488 = n995 | n3467 ;
  assign n15489 = n12388 | n15488 ;
  assign n15491 = ( n4048 & ~n4979 ) | ( n4048 & n8033 ) | ( ~n4979 & n8033 ) ;
  assign n15490 = n1676 & n5795 ;
  assign n15492 = n15491 ^ n15490 ^ 1'b0 ;
  assign n15493 = n3689 & n8950 ;
  assign n15494 = n15493 ^ n3502 ^ 1'b0 ;
  assign n15495 = n1735 & ~n5219 ;
  assign n15496 = n15495 ^ n12504 ^ 1'b0 ;
  assign n15497 = n4867 ^ n1801 ^ 1'b0 ;
  assign n15498 = n10895 | n15497 ;
  assign n15499 = n13306 | n15498 ;
  assign n15500 = ( ~n8271 & n12509 ) | ( ~n8271 & n12621 ) | ( n12509 & n12621 ) ;
  assign n15501 = n2453 | n7125 ;
  assign n15502 = n3096 | n15501 ;
  assign n15503 = n15502 ^ n13991 ^ 1'b0 ;
  assign n15504 = n3083 | n15503 ;
  assign n15509 = n3238 | n7143 ;
  assign n15510 = n15509 ^ n15273 ^ n11043 ;
  assign n15506 = ( x143 & n1260 ) | ( x143 & ~n3896 ) | ( n1260 & ~n3896 ) ;
  assign n15507 = n15506 ^ n9170 ^ n3118 ;
  assign n15508 = x205 & n15507 ;
  assign n15511 = n15510 ^ n15508 ^ 1'b0 ;
  assign n15505 = n4243 | n12042 ;
  assign n15512 = n15511 ^ n15505 ^ 1'b0 ;
  assign n15513 = ~n4619 & n9488 ;
  assign n15514 = n15513 ^ n4637 ^ 1'b0 ;
  assign n15520 = n8018 ^ n389 ^ x16 ;
  assign n15515 = n1477 | n8604 ;
  assign n15516 = n5775 | n15515 ;
  assign n15517 = n3608 ^ n3231 ^ 1'b0 ;
  assign n15518 = n6246 & n15517 ;
  assign n15519 = ( n10800 & n15516 ) | ( n10800 & ~n15518 ) | ( n15516 & ~n15518 ) ;
  assign n15521 = n15520 ^ n15519 ^ 1'b0 ;
  assign n15522 = n8133 | n15521 ;
  assign n15523 = ( ~n6320 & n6622 ) | ( ~n6320 & n12005 ) | ( n6622 & n12005 ) ;
  assign n15524 = n15523 ^ n4435 ^ 1'b0 ;
  assign n15525 = ~n7700 & n15524 ;
  assign n15526 = n6859 & ~n13826 ;
  assign n15527 = n13015 ^ n2604 ^ 1'b0 ;
  assign n15528 = n15526 & ~n15527 ;
  assign n15529 = n3066 ^ n1740 ^ 1'b0 ;
  assign n15530 = n4660 | n11903 ;
  assign n15531 = n14611 ^ n1483 ^ n1255 ;
  assign n15532 = ~n14502 & n15531 ;
  assign n15533 = n6716 & ~n15532 ;
  assign n15534 = n15533 ^ n4779 ^ 1'b0 ;
  assign n15535 = ( n15529 & n15530 ) | ( n15529 & ~n15534 ) | ( n15530 & ~n15534 ) ;
  assign n15536 = n6125 | n9034 ;
  assign n15537 = n15536 ^ n9691 ^ 1'b0 ;
  assign n15538 = ~n4469 & n14279 ;
  assign n15539 = n15538 ^ n2291 ^ 1'b0 ;
  assign n15540 = n6404 | n12186 ;
  assign n15541 = n15540 ^ n2925 ^ 1'b0 ;
  assign n15543 = n7812 ^ n3826 ^ n1789 ;
  assign n15542 = ~n7766 & n7987 ;
  assign n15544 = n15543 ^ n15542 ^ 1'b0 ;
  assign n15545 = n6238 | n15544 ;
  assign n15546 = n8798 & n11645 ;
  assign n15547 = n15546 ^ n10592 ^ 1'b0 ;
  assign n15548 = ( n779 & ~n10970 ) | ( n779 & n15547 ) | ( ~n10970 & n15547 ) ;
  assign n15552 = n5059 ^ n2937 ^ n2824 ;
  assign n15549 = n4352 ^ n2722 ^ 1'b0 ;
  assign n15550 = n3873 & n15549 ;
  assign n15551 = ~n10873 & n15550 ;
  assign n15553 = n15552 ^ n15551 ^ 1'b0 ;
  assign n15557 = n12319 ^ n7541 ^ 1'b0 ;
  assign n15558 = n10199 & n15557 ;
  assign n15554 = n5130 | n9473 ;
  assign n15555 = n13154 & ~n15554 ;
  assign n15556 = ( n3523 & n11789 ) | ( n3523 & n15555 ) | ( n11789 & n15555 ) ;
  assign n15559 = n15558 ^ n15556 ^ n5880 ;
  assign n15560 = n15138 ^ n2995 ^ 1'b0 ;
  assign n15561 = ~n15559 & n15560 ;
  assign n15562 = ( n7649 & ~n12326 ) | ( n7649 & n14632 ) | ( ~n12326 & n14632 ) ;
  assign n15563 = n4537 ^ n4490 ^ 1'b0 ;
  assign n15564 = n7582 & n15563 ;
  assign n15565 = n12813 & n15149 ;
  assign n15566 = ~n15564 & n15565 ;
  assign n15567 = n15566 ^ n11984 ^ 1'b0 ;
  assign n15568 = n11171 ^ n5276 ^ 1'b0 ;
  assign n15569 = n15568 ^ n2359 ^ n946 ;
  assign n15570 = ( n7470 & n12042 ) | ( n7470 & n15569 ) | ( n12042 & n15569 ) ;
  assign n15571 = n6199 ^ n5331 ^ 1'b0 ;
  assign n15572 = n11506 & n13433 ;
  assign n15573 = n15572 ^ n3754 ^ 1'b0 ;
  assign n15574 = n15573 ^ n6746 ^ 1'b0 ;
  assign n15575 = ~n15571 & n15574 ;
  assign n15576 = ( ~n3180 & n15570 ) | ( ~n3180 & n15575 ) | ( n15570 & n15575 ) ;
  assign n15577 = n872 & ~n3751 ;
  assign n15578 = n4416 & n15577 ;
  assign n15579 = n15578 ^ n6246 ^ n3917 ;
  assign n15580 = n4136 | n10160 ;
  assign n15581 = n15579 & ~n15580 ;
  assign n15582 = ~n7209 & n8872 ;
  assign n15587 = n11328 ^ n9252 ^ n4999 ;
  assign n15586 = n7686 ^ n5239 ^ x182 ;
  assign n15584 = n2489 & n3001 ;
  assign n15583 = n4190 & n8295 ;
  assign n15585 = n15584 ^ n15583 ^ n4847 ;
  assign n15588 = n15587 ^ n15586 ^ n15585 ;
  assign n15589 = n11556 & n15588 ;
  assign n15590 = ~n2519 & n3475 ;
  assign n15591 = n15590 ^ n10631 ^ n5299 ;
  assign n15592 = n2265 ^ n1305 ^ 1'b0 ;
  assign n15593 = n2272 & n15592 ;
  assign n15594 = n8227 ^ n2887 ^ x119 ;
  assign n15595 = n15594 ^ n4672 ^ 1'b0 ;
  assign n15596 = n15595 ^ n4833 ^ n642 ;
  assign n15597 = ( ~n10264 & n15593 ) | ( ~n10264 & n15596 ) | ( n15593 & n15596 ) ;
  assign n15598 = n10506 | n13651 ;
  assign n15599 = n10012 & ~n15598 ;
  assign n15602 = n9727 ^ n782 ^ 1'b0 ;
  assign n15603 = n5064 & ~n15602 ;
  assign n15600 = ( n597 & ~n1952 ) | ( n597 & n15123 ) | ( ~n1952 & n15123 ) ;
  assign n15601 = n9581 & n15600 ;
  assign n15604 = n15603 ^ n15601 ^ 1'b0 ;
  assign n15605 = n11965 ^ n10529 ^ n9499 ;
  assign n15608 = ( n3368 & n7190 ) | ( n3368 & n10791 ) | ( n7190 & n10791 ) ;
  assign n15606 = ~n7755 & n12438 ;
  assign n15607 = n15606 ^ n9874 ^ 1'b0 ;
  assign n15609 = n15608 ^ n15607 ^ 1'b0 ;
  assign n15610 = x156 & ~n15609 ;
  assign n15611 = n4379 & ~n12931 ;
  assign n15612 = n4178 ^ n285 ^ 1'b0 ;
  assign n15613 = n13729 & n15612 ;
  assign n15614 = ~n8962 & n12018 ;
  assign n15616 = n12287 ^ n764 ^ 1'b0 ;
  assign n15615 = n6901 ^ n2596 ^ n2140 ;
  assign n15617 = n15616 ^ n15615 ^ n12554 ;
  assign n15618 = n12551 & ~n14041 ;
  assign n15622 = n341 & ~n1805 ;
  assign n15623 = n15622 ^ x87 ^ 1'b0 ;
  assign n15619 = ~n5842 & n7972 ;
  assign n15620 = n15619 ^ n14270 ^ 1'b0 ;
  assign n15621 = n15620 ^ n764 ^ 1'b0 ;
  assign n15624 = n15623 ^ n15621 ^ n8870 ;
  assign n15625 = n14253 ^ n8172 ^ x203 ;
  assign n15626 = n15625 ^ n13252 ^ n4404 ;
  assign n15627 = n4604 & n12026 ;
  assign n15628 = n10605 | n15627 ;
  assign n15629 = n5679 ^ n2995 ^ 1'b0 ;
  assign n15630 = n681 | n15629 ;
  assign n15631 = ( n7272 & n8146 ) | ( n7272 & ~n15630 ) | ( n8146 & ~n15630 ) ;
  assign n15632 = n15631 ^ n7905 ^ 1'b0 ;
  assign n15633 = n12124 ^ n469 ^ 1'b0 ;
  assign n15634 = n15632 & ~n15633 ;
  assign n15635 = n4711 & n13369 ;
  assign n15636 = n15635 ^ n11962 ^ 1'b0 ;
  assign n15637 = n7783 & n15636 ;
  assign n15638 = ~n1811 & n15637 ;
  assign n15639 = n14012 | n15638 ;
  assign n15646 = ~n3930 & n12351 ;
  assign n15644 = ( n9304 & n9671 ) | ( n9304 & ~n11246 ) | ( n9671 & ~n11246 ) ;
  assign n15640 = n8660 | n14672 ;
  assign n15641 = n15640 ^ n12252 ^ 1'b0 ;
  assign n15642 = ~n12013 & n15641 ;
  assign n15643 = n15642 ^ n10325 ^ 1'b0 ;
  assign n15645 = n15644 ^ n15643 ^ 1'b0 ;
  assign n15647 = n15646 ^ n15645 ^ n13091 ;
  assign n15648 = n7414 & ~n7918 ;
  assign n15649 = n14775 & n15648 ;
  assign n15650 = x241 & ~n1926 ;
  assign n15651 = n15649 & n15650 ;
  assign n15652 = n5704 | n15651 ;
  assign n15653 = n15652 ^ n11678 ^ 1'b0 ;
  assign n15654 = ~n2514 & n12462 ;
  assign n15656 = n9043 ^ n7016 ^ n6411 ;
  assign n15657 = ( n7647 & n12353 ) | ( n7647 & n15656 ) | ( n12353 & n15656 ) ;
  assign n15658 = n15657 ^ n12013 ^ n1385 ;
  assign n15659 = n15658 ^ n6736 ^ 1'b0 ;
  assign n15655 = n1053 | n5680 ;
  assign n15660 = n15659 ^ n15655 ^ 1'b0 ;
  assign n15661 = n2438 & ~n4166 ;
  assign n15662 = n15661 ^ n6649 ^ n1782 ;
  assign n15663 = n15662 ^ n8332 ^ n3266 ;
  assign n15664 = n15553 ^ n9255 ^ n5388 ;
  assign n15665 = n2028 & n7477 ;
  assign n15666 = ( n626 & ~n2649 ) | ( n626 & n3377 ) | ( ~n2649 & n3377 ) ;
  assign n15667 = n15666 ^ n338 ^ 1'b0 ;
  assign n15668 = n6937 & n15667 ;
  assign n15669 = n1245 & ~n9794 ;
  assign n15670 = n15669 ^ n1671 ^ 1'b0 ;
  assign n15671 = n15670 ^ n807 ^ x99 ;
  assign n15672 = ( n5831 & ~n10549 ) | ( n5831 & n13527 ) | ( ~n10549 & n13527 ) ;
  assign n15678 = ~n581 & n1610 ;
  assign n15673 = n4714 ^ n1959 ^ n459 ;
  assign n15674 = n5415 ^ x135 ^ 1'b0 ;
  assign n15675 = ~n3200 & n15674 ;
  assign n15676 = n15675 ^ n8936 ^ 1'b0 ;
  assign n15677 = ( n317 & n15673 ) | ( n317 & n15676 ) | ( n15673 & n15676 ) ;
  assign n15679 = n15678 ^ n15677 ^ n4674 ;
  assign n15680 = ( n1607 & n3887 ) | ( n1607 & n12498 ) | ( n3887 & n12498 ) ;
  assign n15681 = n5567 & ~n8225 ;
  assign n15682 = n15681 ^ n10499 ^ n2402 ;
  assign n15683 = n6306 ^ n1455 ^ 1'b0 ;
  assign n15684 = n15683 ^ n5250 ^ n1442 ;
  assign n15685 = ( n8433 & n15682 ) | ( n8433 & ~n15684 ) | ( n15682 & ~n15684 ) ;
  assign n15686 = n15685 ^ n11177 ^ 1'b0 ;
  assign n15687 = n9503 ^ n2194 ^ 1'b0 ;
  assign n15688 = n15687 ^ n12035 ^ n11879 ;
  assign n15689 = n15686 & n15688 ;
  assign n15690 = ( ~n10573 & n15680 ) | ( ~n10573 & n15689 ) | ( n15680 & n15689 ) ;
  assign n15691 = ~n4396 & n11982 ;
  assign n15693 = ( n8279 & n8655 ) | ( n8279 & n9613 ) | ( n8655 & n9613 ) ;
  assign n15692 = n7173 ^ n3465 ^ 1'b0 ;
  assign n15694 = n15693 ^ n15692 ^ n9463 ;
  assign n15695 = n10139 & ~n12739 ;
  assign n15696 = n15695 ^ n9191 ^ 1'b0 ;
  assign n15697 = n4190 | n6215 ;
  assign n15698 = n15697 ^ n3276 ^ 1'b0 ;
  assign n15699 = n15698 ^ n7743 ^ n783 ;
  assign n15700 = n7613 & n7920 ;
  assign n15701 = ~n5662 & n15700 ;
  assign n15702 = n1948 & ~n15701 ;
  assign n15703 = n15699 & n15702 ;
  assign n15707 = n4224 & ~n6805 ;
  assign n15708 = n15707 ^ n7972 ^ 1'b0 ;
  assign n15709 = n15708 ^ n4287 ^ 1'b0 ;
  assign n15710 = n2261 & n15709 ;
  assign n15704 = n6911 ^ n4911 ^ n3775 ;
  assign n15705 = n10710 | n15704 ;
  assign n15706 = n15705 ^ n8787 ^ 1'b0 ;
  assign n15711 = n15710 ^ n15706 ^ n9384 ;
  assign n15712 = n2645 & ~n3732 ;
  assign n15713 = n15712 ^ n1383 ^ 1'b0 ;
  assign n15714 = n8795 ^ n4952 ^ 1'b0 ;
  assign n15715 = ( n10527 & n15713 ) | ( n10527 & ~n15714 ) | ( n15713 & ~n15714 ) ;
  assign n15716 = n2321 & ~n8217 ;
  assign n15717 = ~n7373 & n15716 ;
  assign n15718 = n15717 ^ n11407 ^ n10710 ;
  assign n15721 = ~n855 & n15683 ;
  assign n15722 = n688 & n15721 ;
  assign n15719 = n8574 & n9249 ;
  assign n15720 = ~n2544 & n15719 ;
  assign n15723 = n15722 ^ n15720 ^ n4671 ;
  assign n15724 = n7022 ^ n2834 ^ 1'b0 ;
  assign n15725 = n2638 & ~n4141 ;
  assign n15726 = x240 & n3085 ;
  assign n15727 = n15726 ^ n8307 ^ 1'b0 ;
  assign n15728 = ( ~x215 & n2154 ) | ( ~x215 & n2811 ) | ( n2154 & n2811 ) ;
  assign n15729 = n15728 ^ n4823 ^ 1'b0 ;
  assign n15730 = n1697 & n15729 ;
  assign n15731 = ( n1395 & ~n8929 ) | ( n1395 & n15730 ) | ( ~n8929 & n15730 ) ;
  assign n15732 = ~n4165 & n14311 ;
  assign n15733 = n15731 & ~n15732 ;
  assign n15734 = n3650 & n15733 ;
  assign n15735 = n15734 ^ n4156 ^ 1'b0 ;
  assign n15736 = n15727 | n15735 ;
  assign n15737 = n591 & ~n9430 ;
  assign n15738 = ( n728 & n12477 ) | ( n728 & n15737 ) | ( n12477 & n15737 ) ;
  assign n15739 = n7163 ^ n2890 ^ n1953 ;
  assign n15740 = n1586 | n12110 ;
  assign n15741 = n15740 ^ n8247 ^ 1'b0 ;
  assign n15742 = n15741 ^ n14290 ^ n13753 ;
  assign n15743 = ( n4446 & n5517 ) | ( n4446 & ~n15742 ) | ( n5517 & ~n15742 ) ;
  assign n15744 = ( ~n14852 & n15739 ) | ( ~n14852 & n15743 ) | ( n15739 & n15743 ) ;
  assign n15745 = n11725 ^ n10986 ^ n7128 ;
  assign n15746 = n12504 ^ n6529 ^ 1'b0 ;
  assign n15747 = n15746 ^ n2588 ^ n715 ;
  assign n15748 = n15747 ^ n1312 ^ 1'b0 ;
  assign n15749 = n5858 & n15748 ;
  assign n15750 = ( n10360 & n15745 ) | ( n10360 & n15749 ) | ( n15745 & n15749 ) ;
  assign n15751 = n15744 & n15750 ;
  assign n15752 = n3878 | n4337 ;
  assign n15755 = n9644 ^ n7490 ^ n6785 ;
  assign n15753 = ( x18 & n4467 ) | ( x18 & n6562 ) | ( n4467 & n6562 ) ;
  assign n15754 = n3327 | n15753 ;
  assign n15756 = n15755 ^ n15754 ^ 1'b0 ;
  assign n15757 = n15752 | n15756 ;
  assign n15758 = n13970 ^ n8515 ^ 1'b0 ;
  assign n15759 = n15758 ^ n15260 ^ 1'b0 ;
  assign n15760 = n290 & ~n15759 ;
  assign n15761 = n14807 ^ n8214 ^ 1'b0 ;
  assign n15762 = n11635 ^ n7185 ^ 1'b0 ;
  assign n15763 = n15762 ^ n12000 ^ n9884 ;
  assign n15764 = n14163 ^ n11084 ^ n6818 ;
  assign n15765 = n15119 ^ n7688 ^ 1'b0 ;
  assign n15766 = ~n3163 & n14778 ;
  assign n15767 = ~n5763 & n15766 ;
  assign n15768 = n9237 & ~n15767 ;
  assign n15769 = n5892 ^ n3166 ^ n2030 ;
  assign n15770 = n4499 | n10797 ;
  assign n15771 = n15770 ^ n13755 ^ 1'b0 ;
  assign n15772 = n15771 ^ n10251 ^ 1'b0 ;
  assign n15773 = ( n2336 & n4274 ) | ( n2336 & n15772 ) | ( n4274 & n15772 ) ;
  assign n15774 = n15773 ^ n5627 ^ 1'b0 ;
  assign n15775 = n7751 & ~n15774 ;
  assign n15776 = n7025 ^ n5918 ^ 1'b0 ;
  assign n15777 = ( n1062 & n5418 ) | ( n1062 & ~n15776 ) | ( n5418 & ~n15776 ) ;
  assign n15778 = n4238 ^ n3356 ^ 1'b0 ;
  assign n15779 = ~n11026 & n15778 ;
  assign n15780 = n10469 ^ n1714 ^ 1'b0 ;
  assign n15781 = ~n9578 & n15780 ;
  assign n15782 = n5291 ^ n1133 ^ 1'b0 ;
  assign n15783 = n11649 & n15782 ;
  assign n15784 = n15781 & ~n15783 ;
  assign n15785 = n3769 & ~n15784 ;
  assign n15786 = n15785 ^ n6514 ^ 1'b0 ;
  assign n15787 = n2707 & n5221 ;
  assign n15788 = n15787 ^ n7817 ^ 1'b0 ;
  assign n15789 = n391 & ~n9276 ;
  assign n15790 = n10010 & n15789 ;
  assign n15791 = n15790 ^ n2786 ^ 1'b0 ;
  assign n15792 = n15791 ^ n9608 ^ n9373 ;
  assign n15795 = ( ~n7125 & n10802 ) | ( ~n7125 & n11687 ) | ( n10802 & n11687 ) ;
  assign n15796 = ( n358 & n1299 ) | ( n358 & ~n3865 ) | ( n1299 & ~n3865 ) ;
  assign n15797 = n2443 & n15796 ;
  assign n15798 = ( n6218 & n8184 ) | ( n6218 & ~n14571 ) | ( n8184 & ~n14571 ) ;
  assign n15799 = ( n15795 & n15797 ) | ( n15795 & n15798 ) | ( n15797 & n15798 ) ;
  assign n15793 = n4889 & ~n9304 ;
  assign n15794 = n2093 & n15793 ;
  assign n15800 = n15799 ^ n15794 ^ 1'b0 ;
  assign n15801 = ~n9858 & n15800 ;
  assign n15802 = ~n605 & n15801 ;
  assign n15803 = n3463 ^ n1158 ^ 1'b0 ;
  assign n15804 = ~n2139 & n15803 ;
  assign n15805 = ~n420 & n15804 ;
  assign n15806 = n13039 & n15805 ;
  assign n15807 = ~n4235 & n6426 ;
  assign n15812 = n7910 ^ n480 ^ 1'b0 ;
  assign n15813 = ~n330 & n15812 ;
  assign n15808 = n976 | n5259 ;
  assign n15809 = n3833 & ~n15808 ;
  assign n15810 = ( n1359 & n8741 ) | ( n1359 & ~n15809 ) | ( n8741 & ~n15809 ) ;
  assign n15811 = ~n10222 & n15810 ;
  assign n15814 = n15813 ^ n15811 ^ 1'b0 ;
  assign n15815 = n15807 & n15814 ;
  assign n15816 = n2538 & n2796 ;
  assign n15817 = n15816 ^ n7708 ^ n6417 ;
  assign n15818 = n8196 ^ n1766 ^ 1'b0 ;
  assign n15819 = ~n15817 & n15818 ;
  assign n15820 = n14247 ^ n5193 ^ 1'b0 ;
  assign n15821 = n15820 ^ n10860 ^ n5992 ;
  assign n15822 = n11169 & n12418 ;
  assign n15823 = n2994 ^ n901 ^ 1'b0 ;
  assign n15824 = n8382 | n15823 ;
  assign n15825 = n8571 ^ n5873 ^ 1'b0 ;
  assign n15826 = ~n372 & n15825 ;
  assign n15827 = n2341 & ~n15826 ;
  assign n15828 = ( n6431 & n15824 ) | ( n6431 & ~n15827 ) | ( n15824 & ~n15827 ) ;
  assign n15829 = ( x148 & n707 ) | ( x148 & n1719 ) | ( n707 & n1719 ) ;
  assign n15830 = n15149 & ~n15829 ;
  assign n15831 = n12014 ^ n1886 ^ 1'b0 ;
  assign n15832 = n590 | n12060 ;
  assign n15833 = n15832 ^ n12351 ^ 1'b0 ;
  assign n15834 = n9473 ^ n2414 ^ 1'b0 ;
  assign n15835 = n4554 ^ n2329 ^ x124 ;
  assign n15836 = ~n386 & n15835 ;
  assign n15837 = ~n12817 & n15836 ;
  assign n15838 = n1520 ^ n1429 ^ n1251 ;
  assign n15839 = n5005 & ~n15838 ;
  assign n15840 = n2573 & n10721 ;
  assign n15841 = ~n3038 & n15840 ;
  assign n15842 = ( x212 & n1663 ) | ( x212 & ~n3670 ) | ( n1663 & ~n3670 ) ;
  assign n15843 = ( ~n4267 & n5408 ) | ( ~n4267 & n15842 ) | ( n5408 & n15842 ) ;
  assign n15844 = x21 & n6009 ;
  assign n15845 = n15844 ^ n6963 ^ 1'b0 ;
  assign n15846 = n15843 | n15845 ;
  assign n15847 = ~n2769 & n15846 ;
  assign n15848 = n15847 ^ n6215 ^ 1'b0 ;
  assign n15849 = n7685 ^ n6194 ^ 1'b0 ;
  assign n15850 = ~n14144 & n15849 ;
  assign n15851 = ( ~n2146 & n6222 ) | ( ~n2146 & n15850 ) | ( n6222 & n15850 ) ;
  assign n15852 = n1040 | n8859 ;
  assign n15853 = n12064 & ~n15852 ;
  assign n15856 = n3167 | n3254 ;
  assign n15857 = x109 | n15856 ;
  assign n15858 = ~n1174 & n15857 ;
  assign n15859 = n15858 ^ n2093 ^ 1'b0 ;
  assign n15860 = ( n8546 & ~n12756 ) | ( n8546 & n15859 ) | ( ~n12756 & n15859 ) ;
  assign n15854 = n9687 & n11008 ;
  assign n15855 = n15854 ^ n6345 ^ 1'b0 ;
  assign n15861 = n15860 ^ n15855 ^ 1'b0 ;
  assign n15862 = ~n3442 & n6796 ;
  assign n15871 = n7518 & n9586 ;
  assign n15868 = n2085 | n2432 ;
  assign n15869 = n15868 ^ n449 ^ 1'b0 ;
  assign n15863 = n5605 & ~n13480 ;
  assign n15864 = ~x181 & n15863 ;
  assign n15865 = ( ~n1700 & n4517 ) | ( ~n1700 & n6722 ) | ( n4517 & n6722 ) ;
  assign n15866 = n15865 ^ n9065 ^ 1'b0 ;
  assign n15867 = n15864 | n15866 ;
  assign n15870 = n15869 ^ n15867 ^ n3154 ;
  assign n15872 = n15871 ^ n15870 ^ n874 ;
  assign n15873 = n1108 | n1759 ;
  assign n15874 = n7394 ^ n1898 ^ 1'b0 ;
  assign n15875 = ~n6265 & n15874 ;
  assign n15876 = n15875 ^ n14803 ^ n1340 ;
  assign n15877 = n5682 & ~n10288 ;
  assign n15878 = ~n5526 & n15877 ;
  assign n15879 = n15878 ^ n7615 ^ n2415 ;
  assign n15880 = n15879 ^ n10852 ^ n7904 ;
  assign n15881 = n12576 & ~n15828 ;
  assign n15882 = n15414 & n15881 ;
  assign n15883 = n7304 ^ n4472 ^ n631 ;
  assign n15884 = ( ~n1873 & n7180 ) | ( ~n1873 & n10580 ) | ( n7180 & n10580 ) ;
  assign n15885 = n15883 & ~n15884 ;
  assign n15886 = n2087 & ~n10777 ;
  assign n15887 = n15886 ^ n14915 ^ 1'b0 ;
  assign n15888 = n4087 & ~n11515 ;
  assign n15889 = n6391 | n14148 ;
  assign n15890 = n2676 & ~n15889 ;
  assign n15891 = n8917 | n11775 ;
  assign n15892 = n15890 & ~n15891 ;
  assign n15893 = n15892 ^ n949 ^ 1'b0 ;
  assign n15894 = n5482 ^ n2362 ^ 1'b0 ;
  assign n15895 = ~n3366 & n15894 ;
  assign n15896 = n15895 ^ n15590 ^ n12276 ;
  assign n15897 = ( n5481 & ~n5714 ) | ( n5481 & n13609 ) | ( ~n5714 & n13609 ) ;
  assign n15898 = ( ~n3032 & n13925 ) | ( ~n3032 & n14413 ) | ( n13925 & n14413 ) ;
  assign n15899 = n3430 ^ n1673 ^ 1'b0 ;
  assign n15900 = ( n4019 & ~n7113 ) | ( n4019 & n15899 ) | ( ~n7113 & n15899 ) ;
  assign n15901 = n12696 ^ n5427 ^ 1'b0 ;
  assign n15902 = n12965 ^ n2333 ^ n1798 ;
  assign n15906 = n2937 | n3147 ;
  assign n15907 = ~n6118 & n15906 ;
  assign n15908 = n15907 ^ n4054 ^ 1'b0 ;
  assign n15903 = ~n1348 & n11173 ;
  assign n15904 = n15903 ^ n9749 ^ 1'b0 ;
  assign n15905 = n3013 | n15904 ;
  assign n15909 = n15908 ^ n15905 ^ 1'b0 ;
  assign n15910 = n14075 ^ n13957 ^ n2127 ;
  assign n15918 = n3401 & n5539 ;
  assign n15919 = n15918 ^ n2670 ^ 1'b0 ;
  assign n15911 = n3740 | n4632 ;
  assign n15912 = n15911 ^ n9576 ^ n4598 ;
  assign n15913 = n2896 | n8569 ;
  assign n15914 = n15913 ^ n4066 ^ 1'b0 ;
  assign n15915 = n4897 & n15914 ;
  assign n15916 = ~n15912 & n15915 ;
  assign n15917 = ~n2803 & n15916 ;
  assign n15920 = n15919 ^ n15917 ^ n1706 ;
  assign n15921 = n11866 ^ n8614 ^ n526 ;
  assign n15926 = n7461 ^ n7050 ^ n4669 ;
  assign n15927 = n3783 & n15926 ;
  assign n15925 = n3148 | n4924 ;
  assign n15922 = ( n675 & ~n1142 ) | ( n675 & n8200 ) | ( ~n1142 & n8200 ) ;
  assign n15923 = n6692 ^ n5123 ^ 1'b0 ;
  assign n15924 = n15922 | n15923 ;
  assign n15928 = n15927 ^ n15925 ^ n15924 ;
  assign n15929 = ~n5840 & n15928 ;
  assign n15930 = n373 | n2607 ;
  assign n15931 = n15930 ^ n8389 ^ 1'b0 ;
  assign n15932 = x57 & n9422 ;
  assign n15933 = ~n11366 & n15932 ;
  assign n15934 = n7614 ^ n3231 ^ 1'b0 ;
  assign n15935 = ~n3251 & n15934 ;
  assign n15936 = n633 & ~n1709 ;
  assign n15937 = ~n15935 & n15936 ;
  assign n15938 = n6030 ^ n3629 ^ n2353 ;
  assign n15939 = ( n3693 & n5209 ) | ( n3693 & n15938 ) | ( n5209 & n15938 ) ;
  assign n15940 = n2056 & ~n3954 ;
  assign n15941 = n15940 ^ x110 ^ 1'b0 ;
  assign n15942 = n1739 & ~n15941 ;
  assign n15943 = n4175 ^ n2927 ^ n1366 ;
  assign n15944 = n1737 | n15943 ;
  assign n15945 = ( n6338 & ~n7612 ) | ( n6338 & n15944 ) | ( ~n7612 & n15944 ) ;
  assign n15946 = ( ~n9799 & n15942 ) | ( ~n9799 & n15945 ) | ( n15942 & n15945 ) ;
  assign n15947 = n785 | n8159 ;
  assign n15948 = n14932 | n15947 ;
  assign n15949 = n15948 ^ n9311 ^ 1'b0 ;
  assign n15950 = n15949 ^ n4677 ^ 1'b0 ;
  assign n15951 = n9501 ^ n4809 ^ n4423 ;
  assign n15952 = ~n10496 & n15951 ;
  assign n15953 = ( ~x194 & n3769 ) | ( ~x194 & n6624 ) | ( n3769 & n6624 ) ;
  assign n15954 = n13899 & n15953 ;
  assign n15955 = n1854 & ~n11324 ;
  assign n15956 = n15955 ^ x197 ^ 1'b0 ;
  assign n15957 = n15292 & n15956 ;
  assign n15958 = n15957 ^ n12538 ^ 1'b0 ;
  assign n15959 = ~n2377 & n15958 ;
  assign n15960 = n1852 & n6647 ;
  assign n15961 = n15469 ^ n8128 ^ n4690 ;
  assign n15962 = n14830 & n15961 ;
  assign n15963 = n10549 ^ n7632 ^ 1'b0 ;
  assign n15964 = n3852 | n8367 ;
  assign n15965 = x98 | n15964 ;
  assign n15966 = n13241 ^ n8708 ^ 1'b0 ;
  assign n15967 = n11148 | n15966 ;
  assign n15968 = ( n4810 & ~n15965 ) | ( n4810 & n15967 ) | ( ~n15965 & n15967 ) ;
  assign n15969 = n7204 ^ n5725 ^ 1'b0 ;
  assign n15970 = n4636 ^ n3173 ^ 1'b0 ;
  assign n15971 = ( n9316 & n12415 ) | ( n9316 & ~n15851 ) | ( n12415 & ~n15851 ) ;
  assign n15972 = n9352 ^ n1807 ^ 1'b0 ;
  assign n15973 = ( n4494 & n8582 ) | ( n4494 & ~n8851 ) | ( n8582 & ~n8851 ) ;
  assign n15974 = ( n12269 & n15972 ) | ( n12269 & n15973 ) | ( n15972 & n15973 ) ;
  assign n15975 = n8552 ^ n2529 ^ n2427 ;
  assign n15976 = n15975 ^ n894 ^ 1'b0 ;
  assign n15977 = n10775 | n15976 ;
  assign n15978 = n3509 | n15977 ;
  assign n15979 = n3315 ^ n2191 ^ n1746 ;
  assign n15980 = ~n4904 & n15979 ;
  assign n15981 = ( n1016 & ~n6194 ) | ( n1016 & n13028 ) | ( ~n6194 & n13028 ) ;
  assign n15982 = n13121 ^ n12230 ^ 1'b0 ;
  assign n15983 = n15982 ^ n15061 ^ n12618 ;
  assign n15984 = n1902 & n7391 ;
  assign n15985 = n15984 ^ n3930 ^ 1'b0 ;
  assign n15986 = n15985 ^ n1708 ^ n326 ;
  assign n15987 = n6531 ^ n4874 ^ 1'b0 ;
  assign n15988 = n8513 & ~n15987 ;
  assign n15989 = n2686 ^ n2014 ^ n2001 ;
  assign n15990 = n15989 ^ n8959 ^ 1'b0 ;
  assign n15991 = n5111 ^ n3203 ^ 1'b0 ;
  assign n15992 = n3676 & n15991 ;
  assign n15993 = n15992 ^ n15312 ^ 1'b0 ;
  assign n15994 = ( x0 & n1873 ) | ( x0 & ~n3896 ) | ( n1873 & ~n3896 ) ;
  assign n15995 = n8243 & ~n8463 ;
  assign n15996 = ( n2948 & n4807 ) | ( n2948 & n15995 ) | ( n4807 & n15995 ) ;
  assign n15997 = n15996 ^ n10770 ^ 1'b0 ;
  assign n15998 = n2575 & ~n15997 ;
  assign n15999 = ( n334 & n15994 ) | ( n334 & n15998 ) | ( n15994 & n15998 ) ;
  assign n16000 = n9989 ^ n4147 ^ 1'b0 ;
  assign n16001 = n4444 & ~n16000 ;
  assign n16002 = n16001 ^ n11149 ^ n4760 ;
  assign n16003 = n10536 ^ n3027 ^ 1'b0 ;
  assign n16004 = n2479 & ~n10339 ;
  assign n16005 = n16004 ^ n15144 ^ n12970 ;
  assign n16006 = ( n8196 & n8347 ) | ( n8196 & n9809 ) | ( n8347 & n9809 ) ;
  assign n16007 = n950 | n4486 ;
  assign n16008 = ( x215 & n12462 ) | ( x215 & n16007 ) | ( n12462 & n16007 ) ;
  assign n16009 = n16008 ^ n10575 ^ 1'b0 ;
  assign n16010 = n11565 | n16009 ;
  assign n16011 = n9412 & ~n10297 ;
  assign n16012 = n16011 ^ n15247 ^ 1'b0 ;
  assign n16013 = ( ~n966 & n3673 ) | ( ~n966 & n6611 ) | ( n3673 & n6611 ) ;
  assign n16014 = n1241 | n16013 ;
  assign n16015 = n16014 ^ n7552 ^ 1'b0 ;
  assign n16016 = n15301 & ~n16015 ;
  assign n16017 = n3688 | n9146 ;
  assign n16018 = n16017 ^ n11821 ^ 1'b0 ;
  assign n16019 = ~n1045 & n2006 ;
  assign n16020 = n16019 ^ n13811 ^ 1'b0 ;
  assign n16021 = n10337 ^ n4479 ^ n3249 ;
  assign n16022 = n16021 ^ n10017 ^ 1'b0 ;
  assign n16023 = ( n4665 & n11440 ) | ( n4665 & n16022 ) | ( n11440 & n16022 ) ;
  assign n16026 = ~n1485 & n1542 ;
  assign n16027 = n482 & n4471 ;
  assign n16028 = n16027 ^ n540 ^ 1'b0 ;
  assign n16029 = n16026 | n16028 ;
  assign n16024 = n11594 ^ n4125 ^ n3788 ;
  assign n16025 = n16024 ^ n2987 ^ n416 ;
  assign n16030 = n16029 ^ n16025 ^ n12450 ;
  assign n16031 = ( n5338 & ~n8288 ) | ( n5338 & n16030 ) | ( ~n8288 & n16030 ) ;
  assign n16032 = n4356 ^ n738 ^ 1'b0 ;
  assign n16033 = n9016 & n16032 ;
  assign n16034 = n2236 ^ n668 ^ 1'b0 ;
  assign n16035 = n5315 ^ n4235 ^ 1'b0 ;
  assign n16036 = n2982 & n16035 ;
  assign n16037 = n16034 | n16036 ;
  assign n16038 = n16033 & ~n16037 ;
  assign n16039 = n5196 & n16038 ;
  assign n16040 = n272 | n4242 ;
  assign n16041 = n16040 ^ n13761 ^ 1'b0 ;
  assign n16042 = n2985 | n3765 ;
  assign n16043 = n10094 ^ n9165 ^ n5513 ;
  assign n16044 = n16043 ^ n8281 ^ 1'b0 ;
  assign n16045 = n16042 & ~n16044 ;
  assign n16046 = ~n16041 & n16045 ;
  assign n16047 = n5486 ^ x177 ^ 1'b0 ;
  assign n16048 = ( n6287 & n10963 ) | ( n6287 & n16047 ) | ( n10963 & n16047 ) ;
  assign n16049 = n16048 ^ n10759 ^ n4381 ;
  assign n16050 = n5820 | n11412 ;
  assign n16051 = n13441 ^ n12287 ^ n4373 ;
  assign n16052 = n16051 ^ n5574 ^ n5105 ;
  assign n16053 = n399 & n8297 ;
  assign n16054 = n7658 ^ n6670 ^ n4862 ;
  assign n16055 = n6324 | n16054 ;
  assign n16056 = n16053 & ~n16055 ;
  assign n16057 = n2337 ^ n1385 ^ 1'b0 ;
  assign n16058 = n13430 ^ n12273 ^ 1'b0 ;
  assign n16059 = n16058 ^ n8933 ^ 1'b0 ;
  assign n16060 = n2402 & ~n16059 ;
  assign n16061 = n1948 & n15307 ;
  assign n16062 = n16061 ^ n12815 ^ 1'b0 ;
  assign n16063 = ( n4014 & n5248 ) | ( n4014 & n11191 ) | ( n5248 & n11191 ) ;
  assign n16064 = ( n639 & ~n9075 ) | ( n639 & n13566 ) | ( ~n9075 & n13566 ) ;
  assign n16065 = ( n4611 & n16063 ) | ( n4611 & n16064 ) | ( n16063 & n16064 ) ;
  assign n16066 = ( n262 & ~n11685 ) | ( n262 & n12441 ) | ( ~n11685 & n12441 ) ;
  assign n16067 = n5034 ^ n2654 ^ 1'b0 ;
  assign n16068 = n16067 ^ n12655 ^ n11144 ;
  assign n16069 = n652 & ~n1317 ;
  assign n16070 = n16069 ^ n8127 ^ 1'b0 ;
  assign n16071 = n16070 ^ n9994 ^ 1'b0 ;
  assign n16075 = n3514 ^ n2825 ^ 1'b0 ;
  assign n16072 = ( n1398 & ~n8156 ) | ( n1398 & n14325 ) | ( ~n8156 & n14325 ) ;
  assign n16073 = ~n1475 & n16072 ;
  assign n16074 = ~n1173 & n16073 ;
  assign n16076 = n16075 ^ n16074 ^ 1'b0 ;
  assign n16077 = n9943 & n16076 ;
  assign n16078 = ( n1346 & n3338 ) | ( n1346 & n16077 ) | ( n3338 & n16077 ) ;
  assign n16079 = n16078 ^ n2369 ^ 1'b0 ;
  assign n16080 = n9999 ^ n7112 ^ 1'b0 ;
  assign n16081 = ~n7719 & n16080 ;
  assign n16082 = ~n7223 & n16081 ;
  assign n16083 = n16082 ^ n4837 ^ 1'b0 ;
  assign n16084 = ~n1903 & n7394 ;
  assign n16085 = ( ~n5461 & n6139 ) | ( ~n5461 & n12968 ) | ( n6139 & n12968 ) ;
  assign n16086 = ( n317 & n11987 ) | ( n317 & n16085 ) | ( n11987 & n16085 ) ;
  assign n16087 = n8779 & n10942 ;
  assign n16088 = n1233 ^ n1163 ^ n997 ;
  assign n16089 = n2081 | n6654 ;
  assign n16090 = n16089 ^ n7759 ^ n4104 ;
  assign n16091 = ( n1174 & n13516 ) | ( n1174 & ~n16090 ) | ( n13516 & ~n16090 ) ;
  assign n16092 = n1204 | n3276 ;
  assign n16094 = ~n284 & n8227 ;
  assign n16095 = n2643 & n16094 ;
  assign n16093 = n633 & n7085 ;
  assign n16096 = n16095 ^ n16093 ^ 1'b0 ;
  assign n16097 = n1201 & n5121 ;
  assign n16098 = ~n9174 & n16097 ;
  assign n16099 = n2945 & ~n16098 ;
  assign n16100 = ( n5718 & n6000 ) | ( n5718 & n7569 ) | ( n6000 & n7569 ) ;
  assign n16101 = n16100 ^ n3323 ^ 1'b0 ;
  assign n16102 = n16101 ^ n8513 ^ n6745 ;
  assign n16103 = n821 & ~n3847 ;
  assign n16104 = n16103 ^ n8704 ^ 1'b0 ;
  assign n16105 = ~n16102 & n16104 ;
  assign n16106 = ~n9211 & n16105 ;
  assign n16107 = ~n1130 & n7437 ;
  assign n16108 = ~n5332 & n16107 ;
  assign n16109 = n5755 | n16108 ;
  assign n16110 = ~n2461 & n3080 ;
  assign n16111 = n16110 ^ n1819 ^ 1'b0 ;
  assign n16112 = n15752 ^ n7479 ^ n1649 ;
  assign n16113 = n14577 & ~n16112 ;
  assign n16114 = ~n3223 & n16113 ;
  assign n16115 = n16114 ^ n12687 ^ n877 ;
  assign n16116 = n16115 ^ n12786 ^ 1'b0 ;
  assign n16117 = n5424 ^ n2136 ^ n634 ;
  assign n16118 = n16117 ^ n3650 ^ 1'b0 ;
  assign n16119 = n1381 & ~n16118 ;
  assign n16120 = n5456 & n7912 ;
  assign n16121 = n16120 ^ n10129 ^ 1'b0 ;
  assign n16125 = n4065 ^ n2482 ^ 1'b0 ;
  assign n16126 = n4148 & ~n16125 ;
  assign n16122 = n279 & ~n11990 ;
  assign n16123 = n3507 ^ n2234 ^ 1'b0 ;
  assign n16124 = n16122 & n16123 ;
  assign n16127 = n16126 ^ n16124 ^ n6642 ;
  assign n16128 = n12168 ^ n11614 ^ 1'b0 ;
  assign n16129 = n16128 ^ n13097 ^ n893 ;
  assign n16130 = n10684 ^ n3739 ^ 1'b0 ;
  assign n16131 = x133 & ~n16130 ;
  assign n16132 = ( n299 & ~n572 ) | ( n299 & n4759 ) | ( ~n572 & n4759 ) ;
  assign n16133 = ( n7551 & n13573 ) | ( n7551 & ~n16132 ) | ( n13573 & ~n16132 ) ;
  assign n16134 = ( n8678 & n16131 ) | ( n8678 & n16133 ) | ( n16131 & n16133 ) ;
  assign n16135 = n2753 & ~n3136 ;
  assign n16136 = n1834 & n16135 ;
  assign n16137 = n16136 ^ n12679 ^ n8131 ;
  assign n16138 = n1346 | n16137 ;
  assign n16139 = n8996 & ~n16138 ;
  assign n16140 = n5398 & ~n9197 ;
  assign n16141 = n4352 & n16140 ;
  assign n16145 = n13844 ^ n5968 ^ 1'b0 ;
  assign n16142 = n9798 ^ n926 ^ 1'b0 ;
  assign n16143 = n12479 | n16142 ;
  assign n16144 = ( ~n11532 & n14448 ) | ( ~n11532 & n16143 ) | ( n14448 & n16143 ) ;
  assign n16146 = n16145 ^ n16144 ^ n14274 ;
  assign n16147 = ~n16141 & n16146 ;
  assign n16148 = n11387 ^ n7377 ^ 1'b0 ;
  assign n16149 = n16148 ^ n11304 ^ 1'b0 ;
  assign n16150 = ( n2672 & n9016 ) | ( n2672 & ~n12069 ) | ( n9016 & ~n12069 ) ;
  assign n16151 = n16150 ^ n9265 ^ n5504 ;
  assign n16152 = n12056 ^ n5935 ^ 1'b0 ;
  assign n16158 = ( n881 & n1552 ) | ( n881 & n7965 ) | ( n1552 & n7965 ) ;
  assign n16156 = n12111 ^ n4745 ^ n4266 ;
  assign n16155 = n6967 ^ n3401 ^ n3032 ;
  assign n16153 = ( n2704 & ~n4332 ) | ( n2704 & n13810 ) | ( ~n4332 & n13810 ) ;
  assign n16154 = n12229 | n16153 ;
  assign n16157 = n16156 ^ n16155 ^ n16154 ;
  assign n16159 = n16158 ^ n16157 ^ n702 ;
  assign n16160 = n11190 ^ n3930 ^ n3528 ;
  assign n16161 = ~n3926 & n8291 ;
  assign n16162 = n16161 ^ n6742 ^ 1'b0 ;
  assign n16164 = ( n301 & ~n9139 ) | ( n301 & n14435 ) | ( ~n9139 & n14435 ) ;
  assign n16163 = n4393 ^ n1324 ^ n863 ;
  assign n16165 = n16164 ^ n16163 ^ 1'b0 ;
  assign n16166 = n3917 ^ n2966 ^ 1'b0 ;
  assign n16167 = ( n1742 & ~n2544 ) | ( n1742 & n4212 ) | ( ~n2544 & n4212 ) ;
  assign n16168 = n10863 | n16167 ;
  assign n16169 = n16168 ^ n13632 ^ 1'b0 ;
  assign n16170 = ( ~n3819 & n4711 ) | ( ~n3819 & n4854 ) | ( n4711 & n4854 ) ;
  assign n16171 = n16170 ^ n8000 ^ n6478 ;
  assign n16172 = n14890 ^ n8960 ^ 1'b0 ;
  assign n16173 = n11896 | n16172 ;
  assign n16174 = ( n3392 & n3397 ) | ( n3392 & n4741 ) | ( n3397 & n4741 ) ;
  assign n16175 = ~n689 & n16174 ;
  assign n16176 = n8484 ^ n8364 ^ n967 ;
  assign n16177 = n16176 ^ n10110 ^ n7800 ;
  assign n16185 = ( n3003 & n6758 ) | ( n3003 & ~n7310 ) | ( n6758 & ~n7310 ) ;
  assign n16178 = n15722 ^ n7007 ^ n4417 ;
  assign n16180 = ~n1979 & n12751 ;
  assign n16179 = n10951 ^ n9717 ^ n7101 ;
  assign n16181 = n16180 ^ n16179 ^ 1'b0 ;
  assign n16182 = ~n8607 & n16181 ;
  assign n16183 = ~n4895 & n16182 ;
  assign n16184 = n16178 | n16183 ;
  assign n16186 = n16185 ^ n16184 ^ 1'b0 ;
  assign n16187 = n12466 ^ n3867 ^ 1'b0 ;
  assign n16188 = n7240 ^ n6796 ^ x11 ;
  assign n16189 = n16188 ^ n13964 ^ n4989 ;
  assign n16190 = n5767 ^ n2175 ^ 1'b0 ;
  assign n16191 = n5012 | n16190 ;
  assign n16192 = n16191 ^ n11129 ^ 1'b0 ;
  assign n16193 = n8347 ^ n4749 ^ n686 ;
  assign n16194 = n3937 ^ n3843 ^ n3148 ;
  assign n16195 = n13211 ^ n4146 ^ n1173 ;
  assign n16196 = ~n2620 & n14870 ;
  assign n16197 = n16196 ^ n5051 ^ 1'b0 ;
  assign n16198 = n13372 & ~n16197 ;
  assign n16199 = ( n8502 & n16195 ) | ( n8502 & n16198 ) | ( n16195 & n16198 ) ;
  assign n16200 = n16199 ^ n11224 ^ n640 ;
  assign n16201 = n3760 ^ n3187 ^ 1'b0 ;
  assign n16202 = n6761 ^ n3748 ^ 1'b0 ;
  assign n16203 = n14159 & ~n14728 ;
  assign n16204 = n3781 ^ n3549 ^ n3543 ;
  assign n16205 = n4309 | n16204 ;
  assign n16206 = n1488 & ~n16205 ;
  assign n16207 = ~n3391 & n4281 ;
  assign n16208 = n16206 & n16207 ;
  assign n16209 = n5780 | n7285 ;
  assign n16210 = n1146 | n10930 ;
  assign n16211 = n8092 & ~n16210 ;
  assign n16213 = n9603 ^ n9080 ^ 1'b0 ;
  assign n16212 = ~n7914 & n12113 ;
  assign n16214 = n16213 ^ n16212 ^ 1'b0 ;
  assign n16215 = n9026 ^ n6132 ^ 1'b0 ;
  assign n16216 = n12573 & n16215 ;
  assign n16223 = n12306 & ~n13190 ;
  assign n16224 = n16223 ^ n2261 ^ 1'b0 ;
  assign n16222 = ( n4152 & ~n5233 ) | ( n4152 & n5833 ) | ( ~n5233 & n5833 ) ;
  assign n16225 = n16224 ^ n16222 ^ 1'b0 ;
  assign n16217 = n9903 ^ n5759 ^ 1'b0 ;
  assign n16218 = n10019 | n16217 ;
  assign n16219 = n16218 ^ n13250 ^ 1'b0 ;
  assign n16220 = n1168 | n16219 ;
  assign n16221 = n4694 & ~n16220 ;
  assign n16226 = n16225 ^ n16221 ^ 1'b0 ;
  assign n16238 = ~n4725 & n10914 ;
  assign n16235 = n6011 | n7953 ;
  assign n16236 = n16235 ^ n3233 ^ 1'b0 ;
  assign n16234 = n13635 ^ n964 ^ n350 ;
  assign n16237 = n16236 ^ n16234 ^ n4705 ;
  assign n16229 = n14418 ^ n5405 ^ 1'b0 ;
  assign n16230 = n2631 | n16229 ;
  assign n16227 = n5442 & ~n9839 ;
  assign n16228 = n7815 & n16227 ;
  assign n16231 = n16230 ^ n16228 ^ 1'b0 ;
  assign n16232 = ~n15687 & n16231 ;
  assign n16233 = ~n13687 & n16232 ;
  assign n16239 = n16238 ^ n16237 ^ n16233 ;
  assign n16240 = ~n1314 & n3320 ;
  assign n16241 = ~x45 & n16240 ;
  assign n16242 = n8757 ^ n8023 ^ 1'b0 ;
  assign n16243 = n4467 ^ n3676 ^ 1'b0 ;
  assign n16244 = n11498 | n16243 ;
  assign n16245 = ( n3006 & n3923 ) | ( n3006 & n16244 ) | ( n3923 & n16244 ) ;
  assign n16246 = n13487 ^ n10278 ^ 1'b0 ;
  assign n16247 = n8122 & n16246 ;
  assign n16248 = n5982 ^ n2791 ^ 1'b0 ;
  assign n16249 = n5044 ^ n3713 ^ n2326 ;
  assign n16250 = n16249 ^ n3974 ^ 1'b0 ;
  assign n16251 = ~n11175 & n11295 ;
  assign n16252 = ~n1819 & n16251 ;
  assign n16253 = ( n9981 & ~n16250 ) | ( n9981 & n16252 ) | ( ~n16250 & n16252 ) ;
  assign n16254 = ( n8253 & n16248 ) | ( n8253 & ~n16253 ) | ( n16248 & ~n16253 ) ;
  assign n16255 = n3984 & ~n8506 ;
  assign n16256 = n16255 ^ n14418 ^ n2634 ;
  assign n16257 = n2858 | n16256 ;
  assign n16258 = n1947 & ~n16257 ;
  assign n16259 = ( ~n1675 & n3049 ) | ( ~n1675 & n15443 ) | ( n3049 & n15443 ) ;
  assign n16260 = n15909 ^ n10274 ^ 1'b0 ;
  assign n16261 = n15422 ^ n13194 ^ 1'b0 ;
  assign n16262 = n7743 & n16261 ;
  assign n16264 = n11845 & n14141 ;
  assign n16265 = n16264 ^ n8591 ^ 1'b0 ;
  assign n16263 = n334 | n3563 ;
  assign n16266 = n16265 ^ n16263 ^ 1'b0 ;
  assign n16267 = n16266 ^ n2114 ^ 1'b0 ;
  assign n16270 = ( ~n5492 & n9872 ) | ( ~n5492 & n11503 ) | ( n9872 & n11503 ) ;
  assign n16268 = n3709 | n11767 ;
  assign n16269 = n9288 | n16268 ;
  assign n16271 = n16270 ^ n16269 ^ 1'b0 ;
  assign n16272 = n2828 | n5566 ;
  assign n16273 = ( n2573 & n6799 ) | ( n2573 & ~n16272 ) | ( n6799 & ~n16272 ) ;
  assign n16274 = n7142 & ~n16273 ;
  assign n16281 = n6329 ^ n3845 ^ 1'b0 ;
  assign n16282 = ( n486 & n3779 ) | ( n486 & ~n16281 ) | ( n3779 & ~n16281 ) ;
  assign n16283 = n16282 ^ n3335 ^ 1'b0 ;
  assign n16284 = ( n6423 & ~n10227 ) | ( n6423 & n16283 ) | ( ~n10227 & n16283 ) ;
  assign n16275 = ( n713 & ~n7533 ) | ( n713 & n11097 ) | ( ~n7533 & n11097 ) ;
  assign n16276 = n11324 ^ n7913 ^ n6479 ;
  assign n16277 = n16276 ^ n5479 ^ 1'b0 ;
  assign n16278 = ( n3335 & n16275 ) | ( n3335 & ~n16277 ) | ( n16275 & ~n16277 ) ;
  assign n16279 = n16278 ^ n9658 ^ 1'b0 ;
  assign n16280 = n11292 & ~n16279 ;
  assign n16285 = n16284 ^ n16280 ^ n14353 ;
  assign n16286 = ( n16271 & n16274 ) | ( n16271 & ~n16285 ) | ( n16274 & ~n16285 ) ;
  assign n16287 = ( n5772 & ~n10659 ) | ( n5772 & n15052 ) | ( ~n10659 & n15052 ) ;
  assign n16288 = ~n2554 & n6777 ;
  assign n16289 = n8726 & n16288 ;
  assign n16290 = n16289 ^ n16144 ^ 1'b0 ;
  assign n16291 = n11149 & ~n14462 ;
  assign n16292 = n11252 ^ n8357 ^ n5840 ;
  assign n16293 = n7254 ^ n5051 ^ 1'b0 ;
  assign n16294 = ( n4289 & ~n5523 ) | ( n4289 & n9706 ) | ( ~n5523 & n9706 ) ;
  assign n16295 = n4261 & ~n16294 ;
  assign n16296 = n16295 ^ n5544 ^ 1'b0 ;
  assign n16297 = n5371 & ~n16296 ;
  assign n16298 = n8809 & n16297 ;
  assign n16299 = n583 | n8757 ;
  assign n16300 = x21 | n16299 ;
  assign n16301 = n16300 ^ n5064 ^ n1452 ;
  assign n16302 = n16301 ^ n2113 ^ 1'b0 ;
  assign n16303 = ( n3248 & ~n15587 ) | ( n3248 & n16288 ) | ( ~n15587 & n16288 ) ;
  assign n16304 = n1342 & n4670 ;
  assign n16305 = ~n4670 & n16304 ;
  assign n16306 = n2860 | n16305 ;
  assign n16307 = ~n6103 & n16306 ;
  assign n16308 = ~n16306 & n16307 ;
  assign n16309 = n1452 ^ n561 ^ 1'b0 ;
  assign n16310 = n11192 & n16309 ;
  assign n16311 = ( ~n9794 & n9896 ) | ( ~n9794 & n16310 ) | ( n9896 & n16310 ) ;
  assign n16312 = n12685 ^ n11644 ^ 1'b0 ;
  assign n16313 = n1764 ^ n750 ^ 1'b0 ;
  assign n16314 = n16313 ^ n13241 ^ 1'b0 ;
  assign n16315 = n16314 ^ n10670 ^ 1'b0 ;
  assign n16316 = n16315 ^ n11553 ^ n4812 ;
  assign n16317 = n8619 & ~n16316 ;
  assign n16318 = n11143 ^ n6129 ^ 1'b0 ;
  assign n16319 = ~n5118 & n16318 ;
  assign n16320 = n3659 ^ x17 ^ 1'b0 ;
  assign n16321 = ~n15318 & n16320 ;
  assign n16322 = n6266 & ~n8667 ;
  assign n16323 = n9778 ^ n2515 ^ 1'b0 ;
  assign n16326 = n11587 ^ n4675 ^ 1'b0 ;
  assign n16324 = n12897 ^ n7252 ^ 1'b0 ;
  assign n16325 = n10765 & ~n16324 ;
  assign n16327 = n16326 ^ n16325 ^ n4587 ;
  assign n16328 = n4636 | n16327 ;
  assign n16329 = n8290 & ~n16328 ;
  assign n16330 = ~n8366 & n9366 ;
  assign n16331 = n16330 ^ n4524 ^ 1'b0 ;
  assign n16332 = n9919 & ~n16331 ;
  assign n16333 = n3510 | n14899 ;
  assign n16334 = ( n2807 & n7968 ) | ( n2807 & n16333 ) | ( n7968 & n16333 ) ;
  assign n16335 = n13306 ^ n2040 ^ 1'b0 ;
  assign n16336 = n7245 ^ n6260 ^ n1268 ;
  assign n16337 = n10020 | n16336 ;
  assign n16338 = n16337 ^ n5674 ^ 1'b0 ;
  assign n16339 = x240 & ~n2476 ;
  assign n16340 = n16339 ^ n3107 ^ 1'b0 ;
  assign n16341 = x140 & n16340 ;
  assign n16342 = n7558 & n16341 ;
  assign n16343 = ( n10002 & n12929 ) | ( n10002 & ~n16342 ) | ( n12929 & ~n16342 ) ;
  assign n16344 = n11982 ^ n10065 ^ 1'b0 ;
  assign n16345 = n3721 & ~n16344 ;
  assign n16346 = n16345 ^ n11840 ^ x50 ;
  assign n16348 = x84 & n1066 ;
  assign n16347 = n5281 | n14894 ;
  assign n16349 = n16348 ^ n16347 ^ 1'b0 ;
  assign n16350 = n1198 | n4900 ;
  assign n16351 = n12032 ^ n8786 ^ 1'b0 ;
  assign n16352 = n3849 & ~n16351 ;
  assign n16353 = n16350 & ~n16352 ;
  assign n16354 = n13859 ^ n7641 ^ 1'b0 ;
  assign n16355 = n416 | n16354 ;
  assign n16356 = n16355 ^ n4550 ^ 1'b0 ;
  assign n16357 = ~n9704 & n16356 ;
  assign n16358 = ( n2315 & n2534 ) | ( n2315 & n7331 ) | ( n2534 & n7331 ) ;
  assign n16359 = n350 & ~n2240 ;
  assign n16360 = n4550 | n16359 ;
  assign n16361 = n11770 | n16360 ;
  assign n16362 = n16361 ^ n7034 ^ n5838 ;
  assign n16363 = ( ~x79 & n10898 ) | ( ~x79 & n16362 ) | ( n10898 & n16362 ) ;
  assign n16364 = n16363 ^ n1379 ^ 1'b0 ;
  assign n16365 = n10432 & ~n16364 ;
  assign n16366 = ~n1405 & n16365 ;
  assign n16367 = ~n3091 & n16366 ;
  assign n16368 = n3770 | n4767 ;
  assign n16369 = n4670 ^ n3173 ^ n690 ;
  assign n16370 = n16369 ^ n285 ^ 1'b0 ;
  assign n16371 = n9732 & n16370 ;
  assign n16372 = n5882 & n16371 ;
  assign n16373 = ( n755 & ~n14639 ) | ( n755 & n15913 ) | ( ~n14639 & n15913 ) ;
  assign n16374 = n16292 ^ n8315 ^ n8010 ;
  assign n16376 = n2952 | n12417 ;
  assign n16377 = n6632 | n16376 ;
  assign n16378 = n16377 ^ n5954 ^ 1'b0 ;
  assign n16375 = ( ~n671 & n6222 ) | ( ~n671 & n9947 ) | ( n6222 & n9947 ) ;
  assign n16379 = n16378 ^ n16375 ^ 1'b0 ;
  assign n16380 = n2620 & n16379 ;
  assign n16381 = n16380 ^ n14499 ^ 1'b0 ;
  assign n16382 = n6326 & ~n15771 ;
  assign n16383 = n8337 & n16382 ;
  assign n16384 = n343 & ~n16383 ;
  assign n16385 = n14109 & n16384 ;
  assign n16386 = ~n3442 & n12391 ;
  assign n16387 = n16386 ^ n9526 ^ 1'b0 ;
  assign n16388 = n4833 & ~n6431 ;
  assign n16389 = ~n1524 & n16388 ;
  assign n16391 = n7485 ^ n5238 ^ 1'b0 ;
  assign n16392 = ~n7073 & n16391 ;
  assign n16393 = ~n15419 & n16392 ;
  assign n16394 = n4007 & n16393 ;
  assign n16390 = n10194 ^ n7391 ^ n2383 ;
  assign n16395 = n16394 ^ n16390 ^ 1'b0 ;
  assign n16396 = n10631 ^ n4230 ^ 1'b0 ;
  assign n16397 = ~x210 & n16396 ;
  assign n16398 = ( n11086 & n12484 ) | ( n11086 & ~n13873 ) | ( n12484 & ~n13873 ) ;
  assign n16399 = n6135 ^ n1818 ^ 1'b0 ;
  assign n16400 = n6875 | n8640 ;
  assign n16401 = n16116 ^ n15886 ^ 1'b0 ;
  assign n16402 = n7750 ^ n1629 ^ 1'b0 ;
  assign n16403 = n14758 ^ n9164 ^ n2638 ;
  assign n16404 = ~n4589 & n8533 ;
  assign n16405 = n16404 ^ n1680 ^ 1'b0 ;
  assign n16406 = n16405 ^ n9725 ^ n5537 ;
  assign n16407 = n3874 | n15594 ;
  assign n16408 = n16407 ^ n5954 ^ 1'b0 ;
  assign n16409 = n16406 & n16408 ;
  assign n16410 = n5405 & ~n8400 ;
  assign n16411 = ~n16409 & n16410 ;
  assign n16412 = ( ~n2233 & n3759 ) | ( ~n2233 & n4567 ) | ( n3759 & n4567 ) ;
  assign n16413 = ( x167 & n6803 ) | ( x167 & n16412 ) | ( n6803 & n16412 ) ;
  assign n16414 = n4728 ^ n284 ^ x36 ;
  assign n16415 = ( n9851 & ~n16413 ) | ( n9851 & n16414 ) | ( ~n16413 & n16414 ) ;
  assign n16416 = n11800 ^ n6318 ^ n4504 ;
  assign n16417 = n8535 ^ n4558 ^ n2971 ;
  assign n16418 = ~n16416 & n16417 ;
  assign n16419 = n16418 ^ n5510 ^ 1'b0 ;
  assign n16420 = n6501 | n7442 ;
  assign n16421 = n16420 ^ n9690 ^ 1'b0 ;
  assign n16422 = n2621 & n9655 ;
  assign n16423 = n13943 ^ n13396 ^ 1'b0 ;
  assign n16424 = n1775 | n16423 ;
  assign n16425 = n4949 | n9607 ;
  assign n16426 = n15347 | n16425 ;
  assign n16427 = ( n1868 & ~n12073 ) | ( n1868 & n16426 ) | ( ~n12073 & n16426 ) ;
  assign n16429 = ( x197 & n6001 ) | ( x197 & n7380 ) | ( n6001 & n7380 ) ;
  assign n16428 = n3159 | n15656 ;
  assign n16430 = n16429 ^ n16428 ^ 1'b0 ;
  assign n16431 = n16430 ^ n13203 ^ 1'b0 ;
  assign n16432 = n16431 ^ x241 ^ 1'b0 ;
  assign n16433 = ~n16427 & n16432 ;
  assign n16434 = n12234 ^ n12209 ^ n6205 ;
  assign n16435 = x119 & ~n3450 ;
  assign n16436 = n4110 & n16435 ;
  assign n16437 = ~n16434 & n16436 ;
  assign n16438 = ~n2808 & n6150 ;
  assign n16441 = n11186 ^ n9127 ^ n2725 ;
  assign n16439 = ( n1705 & n4016 ) | ( n1705 & ~n8739 ) | ( n4016 & ~n8739 ) ;
  assign n16440 = n2382 & n16439 ;
  assign n16442 = n16441 ^ n16440 ^ 1'b0 ;
  assign n16443 = n4520 ^ n764 ^ 1'b0 ;
  assign n16444 = n16442 & ~n16443 ;
  assign n16445 = n4300 & n16444 ;
  assign n16446 = ~n16438 & n16445 ;
  assign n16447 = n8715 ^ n1263 ^ 1'b0 ;
  assign n16448 = ( n461 & n5006 ) | ( n461 & ~n16447 ) | ( n5006 & ~n16447 ) ;
  assign n16449 = n9521 ^ n1858 ^ 1'b0 ;
  assign n16450 = n16449 ^ n4231 ^ 1'b0 ;
  assign n16451 = n15335 & ~n16450 ;
  assign n16452 = n16451 ^ n3619 ^ 1'b0 ;
  assign n16453 = n6538 & ~n16452 ;
  assign n16454 = n9252 ^ n4423 ^ n1414 ;
  assign n16455 = ( n466 & n4560 ) | ( n466 & ~n12219 ) | ( n4560 & ~n12219 ) ;
  assign n16456 = n16454 & ~n16455 ;
  assign n16458 = ~n5996 & n11171 ;
  assign n16457 = ~n4390 & n5978 ;
  assign n16459 = n16458 ^ n16457 ^ 1'b0 ;
  assign n16460 = n16310 & n16459 ;
  assign n16461 = ( ~n9002 & n14208 ) | ( ~n9002 & n15219 ) | ( n14208 & n15219 ) ;
  assign n16462 = n16461 ^ n9037 ^ 1'b0 ;
  assign n16463 = ~n3254 & n10259 ;
  assign n16464 = ~n8002 & n16463 ;
  assign n16470 = n10367 ^ n7223 ^ 1'b0 ;
  assign n16465 = n7824 | n8588 ;
  assign n16466 = n2924 & ~n16465 ;
  assign n16467 = n12306 ^ n1838 ^ 1'b0 ;
  assign n16468 = n11008 & n16467 ;
  assign n16469 = ~n16466 & n16468 ;
  assign n16471 = n16470 ^ n16469 ^ 1'b0 ;
  assign n16472 = n14658 ^ n1719 ^ 1'b0 ;
  assign n16473 = n13127 ^ n8379 ^ n7461 ;
  assign n16474 = n16473 ^ n9703 ^ 1'b0 ;
  assign n16475 = n16472 | n16474 ;
  assign n16476 = n13222 ^ n8608 ^ 1'b0 ;
  assign n16477 = n2532 & ~n16476 ;
  assign n16478 = ( n814 & n9064 ) | ( n814 & n10534 ) | ( n9064 & n10534 ) ;
  assign n16479 = n4066 & n16478 ;
  assign n16480 = n7751 ^ n6523 ^ 1'b0 ;
  assign n16481 = ~n16479 & n16480 ;
  assign n16482 = n4316 | n11127 ;
  assign n16483 = n16482 ^ n9378 ^ 1'b0 ;
  assign n16484 = n757 ^ n374 ^ 1'b0 ;
  assign n16485 = n16484 ^ n9904 ^ 1'b0 ;
  assign n16486 = ~n8384 & n16485 ;
  assign n16487 = n8840 ^ n3360 ^ 1'b0 ;
  assign n16488 = ~n4343 & n16487 ;
  assign n16489 = n16488 ^ x54 ^ 1'b0 ;
  assign n16490 = n2448 & ~n16489 ;
  assign n16491 = ( ~n5097 & n6166 ) | ( ~n5097 & n16490 ) | ( n6166 & n16490 ) ;
  assign n16492 = n9851 | n12960 ;
  assign n16493 = ( n1893 & n4987 ) | ( n1893 & n16001 ) | ( n4987 & n16001 ) ;
  assign n16494 = n829 & ~n1704 ;
  assign n16495 = ~x235 & n16494 ;
  assign n16496 = n16495 ^ n10514 ^ n5359 ;
  assign n16497 = n3060 & n7220 ;
  assign n16498 = x214 & ~n548 ;
  assign n16499 = ~n7782 & n16498 ;
  assign n16500 = ( x54 & n1795 ) | ( x54 & ~n3762 ) | ( n1795 & ~n3762 ) ;
  assign n16501 = n16500 ^ n10896 ^ 1'b0 ;
  assign n16502 = ~n16499 & n16501 ;
  assign n16503 = n16502 ^ n6858 ^ n3222 ;
  assign n16504 = n16503 ^ n3810 ^ 1'b0 ;
  assign n16505 = ~n3694 & n16198 ;
  assign n16506 = n16504 & n16505 ;
  assign n16507 = n11002 | n13582 ;
  assign n16508 = n5864 ^ n5070 ^ 1'b0 ;
  assign n16509 = n16508 ^ n2117 ^ 1'b0 ;
  assign n16510 = n4624 | n6665 ;
  assign n16511 = n16510 ^ n13681 ^ 1'b0 ;
  assign n16512 = ~n16509 & n16511 ;
  assign n16520 = ~n5744 & n5975 ;
  assign n16521 = n16520 ^ n6826 ^ 1'b0 ;
  assign n16522 = n9056 | n16521 ;
  assign n16523 = ( x59 & n5507 ) | ( x59 & ~n16522 ) | ( n5507 & ~n16522 ) ;
  assign n16519 = x140 & ~n3219 ;
  assign n16524 = n16523 ^ n16519 ^ 1'b0 ;
  assign n16516 = n12053 ^ n6253 ^ 1'b0 ;
  assign n16517 = ~n5825 & n16516 ;
  assign n16513 = n5390 & n9780 ;
  assign n16514 = ~n2380 & n16513 ;
  assign n16515 = n8988 | n16514 ;
  assign n16518 = n16517 ^ n16515 ^ 1'b0 ;
  assign n16525 = n16524 ^ n16518 ^ n16070 ;
  assign n16526 = n4118 ^ n1673 ^ n414 ;
  assign n16527 = n16526 ^ n4793 ^ n4190 ;
  assign n16528 = n16527 ^ n13491 ^ 1'b0 ;
  assign n16529 = n977 | n16528 ;
  assign n16530 = n16529 ^ n11678 ^ 1'b0 ;
  assign n16531 = n6703 ^ n1506 ^ n735 ;
  assign n16532 = n16531 ^ n6570 ^ 1'b0 ;
  assign n16533 = ~n3273 & n16532 ;
  assign n16534 = ( n1346 & ~n11005 ) | ( n1346 & n16533 ) | ( ~n11005 & n16533 ) ;
  assign n16535 = ( n14544 & ~n16530 ) | ( n14544 & n16534 ) | ( ~n16530 & n16534 ) ;
  assign n16536 = n14224 ^ n5253 ^ 1'b0 ;
  assign n16537 = n2719 & ~n16536 ;
  assign n16538 = ( n3580 & ~n5456 ) | ( n3580 & n16537 ) | ( ~n5456 & n16537 ) ;
  assign n16539 = n16101 ^ n11325 ^ 1'b0 ;
  assign n16540 = ( n7352 & n14075 ) | ( n7352 & ~n16539 ) | ( n14075 & ~n16539 ) ;
  assign n16541 = n15542 ^ n502 ^ 1'b0 ;
  assign n16542 = ( n9220 & ~n14952 ) | ( n9220 & n16541 ) | ( ~n14952 & n16541 ) ;
  assign n16543 = n4744 ^ n1556 ^ 1'b0 ;
  assign n16544 = n16542 & ~n16543 ;
  assign n16545 = n524 & ~n12613 ;
  assign n16546 = n16545 ^ n13901 ^ 1'b0 ;
  assign n16547 = ( n269 & n11330 ) | ( n269 & ~n13708 ) | ( n11330 & ~n13708 ) ;
  assign n16548 = n1930 | n4117 ;
  assign n16549 = n16548 ^ n3832 ^ 1'b0 ;
  assign n16550 = n3109 & n16549 ;
  assign n16551 = n16547 & n16550 ;
  assign n16552 = n10454 ^ n7615 ^ 1'b0 ;
  assign n16554 = n10820 ^ n7325 ^ n5292 ;
  assign n16553 = ~n1241 & n3463 ;
  assign n16555 = n16554 ^ n16553 ^ 1'b0 ;
  assign n16556 = ~n3690 & n16555 ;
  assign n16557 = ~n16552 & n16556 ;
  assign n16558 = n8169 & ~n16557 ;
  assign n16559 = ~n14536 & n16558 ;
  assign n16560 = n16559 ^ n10690 ^ n1850 ;
  assign n16561 = n702 | n2590 ;
  assign n16562 = n10024 ^ n5965 ^ n1397 ;
  assign n16563 = n12904 & ~n16562 ;
  assign n16564 = n11946 ^ n3675 ^ 1'b0 ;
  assign n16565 = n5573 & ~n16564 ;
  assign n16566 = n16565 ^ n16301 ^ n9481 ;
  assign n16572 = ~n859 & n8754 ;
  assign n16567 = n8953 ^ n7795 ^ 1'b0 ;
  assign n16568 = ~n7195 & n16567 ;
  assign n16569 = n7159 & n16568 ;
  assign n16570 = n16569 ^ n2782 ^ 1'b0 ;
  assign n16571 = n7322 & n16570 ;
  assign n16573 = n16572 ^ n16571 ^ 1'b0 ;
  assign n16574 = n11284 ^ n4535 ^ n2022 ;
  assign n16575 = n12080 ^ n7490 ^ 1'b0 ;
  assign n16576 = n10404 ^ n7102 ^ n5252 ;
  assign n16577 = n2638 & n16576 ;
  assign n16578 = n4322 & n16577 ;
  assign n16579 = n13218 ^ n2534 ^ 1'b0 ;
  assign n16580 = n2578 & n16579 ;
  assign n16581 = n13435 ^ n4226 ^ 1'b0 ;
  assign n16582 = n11676 ^ n2560 ^ 1'b0 ;
  assign n16583 = n7922 & ~n11676 ;
  assign n16584 = ~n1493 & n16583 ;
  assign n16585 = n898 | n6782 ;
  assign n16586 = ( n9039 & ~n16584 ) | ( n9039 & n16585 ) | ( ~n16584 & n16585 ) ;
  assign n16587 = n15365 ^ n7674 ^ 1'b0 ;
  assign n16588 = n1802 & ~n4053 ;
  assign n16589 = n2913 & n16588 ;
  assign n16590 = n15810 ^ n12783 ^ n12209 ;
  assign n16591 = n3817 ^ n2265 ^ 1'b0 ;
  assign n16592 = n8055 & n16591 ;
  assign n16593 = ( ~n6669 & n16590 ) | ( ~n6669 & n16592 ) | ( n16590 & n16592 ) ;
  assign n16594 = ~x165 & n8949 ;
  assign n16595 = ~n642 & n10388 ;
  assign n16596 = n16594 & n16595 ;
  assign n16597 = n7152 & ~n8907 ;
  assign n16598 = n16597 ^ n4815 ^ 1'b0 ;
  assign n16599 = ( n8291 & n11312 ) | ( n8291 & n16598 ) | ( n11312 & n16598 ) ;
  assign n16600 = n7331 & n16599 ;
  assign n16601 = ~n2139 & n6164 ;
  assign n16602 = ( n1884 & ~n5029 ) | ( n1884 & n6367 ) | ( ~n5029 & n6367 ) ;
  assign n16603 = n16602 ^ n4684 ^ n1496 ;
  assign n16604 = n5804 ^ n3133 ^ 1'b0 ;
  assign n16605 = n684 | n16604 ;
  assign n16606 = n16603 | n16605 ;
  assign n16607 = n16601 | n16606 ;
  assign n16610 = n1469 | n12429 ;
  assign n16611 = n16610 ^ n8426 ^ 1'b0 ;
  assign n16609 = n12423 ^ n11956 ^ n1604 ;
  assign n16608 = ~n1632 & n7762 ;
  assign n16612 = n16611 ^ n16609 ^ n16608 ;
  assign n16613 = n10104 | n10505 ;
  assign n16614 = n16613 ^ n7748 ^ 1'b0 ;
  assign n16615 = ~n3788 & n4759 ;
  assign n16616 = n2437 & n16615 ;
  assign n16617 = n4319 ^ n673 ^ 1'b0 ;
  assign n16618 = n6402 & n16617 ;
  assign n16619 = n16618 ^ n4842 ^ 1'b0 ;
  assign n16620 = ~n16616 & n16619 ;
  assign n16621 = n13521 ^ n317 ^ 1'b0 ;
  assign n16622 = n16620 & ~n16621 ;
  assign n16623 = n1735 & n1932 ;
  assign n16624 = n16623 ^ n16271 ^ n5500 ;
  assign n16625 = n3156 ^ n3004 ^ 1'b0 ;
  assign n16626 = ~n4243 & n16625 ;
  assign n16627 = n4575 & ~n9710 ;
  assign n16628 = ~n16626 & n16627 ;
  assign n16629 = n16628 ^ n7425 ^ 1'b0 ;
  assign n16630 = ~n7461 & n9015 ;
  assign n16631 = ( n5364 & ~n11088 ) | ( n5364 & n16630 ) | ( ~n11088 & n16630 ) ;
  assign n16632 = n13874 & ~n16631 ;
  assign n16633 = ~n10750 & n16632 ;
  assign n16634 = n1754 & ~n9504 ;
  assign n16635 = n15543 & n16634 ;
  assign n16636 = n10042 ^ n7750 ^ 1'b0 ;
  assign n16637 = n16289 | n16636 ;
  assign n16638 = ~n2066 & n7683 ;
  assign n16639 = n2398 ^ n758 ^ n633 ;
  assign n16640 = n5222 & n16639 ;
  assign n16641 = n5097 & n6045 ;
  assign n16642 = ( n13188 & n16640 ) | ( n13188 & n16641 ) | ( n16640 & n16641 ) ;
  assign n16643 = n7682 | n8548 ;
  assign n16644 = n16643 ^ n7788 ^ 1'b0 ;
  assign n16645 = n10952 ^ n4435 ^ 1'b0 ;
  assign n16646 = n6964 | n16645 ;
  assign n16652 = n4744 & ~n8022 ;
  assign n16649 = ( ~n2038 & n3805 ) | ( ~n2038 & n6872 ) | ( n3805 & n6872 ) ;
  assign n16650 = n3048 | n16649 ;
  assign n16651 = n16650 ^ n16145 ^ n908 ;
  assign n16647 = ( ~n996 & n5862 ) | ( ~n996 & n7484 ) | ( n5862 & n7484 ) ;
  assign n16648 = ~n3830 & n16647 ;
  assign n16653 = n16652 ^ n16651 ^ n16648 ;
  assign n16659 = ( n3285 & n8860 ) | ( n3285 & n8958 ) | ( n8860 & n8958 ) ;
  assign n16658 = n12381 ^ n9776 ^ n3549 ;
  assign n16654 = ( n4513 & n6520 ) | ( n4513 & ~n7254 ) | ( n6520 & ~n7254 ) ;
  assign n16655 = ( n3831 & n8930 ) | ( n3831 & n16654 ) | ( n8930 & n16654 ) ;
  assign n16656 = n16655 ^ n12406 ^ n4388 ;
  assign n16657 = ( n744 & ~n13583 ) | ( n744 & n16656 ) | ( ~n13583 & n16656 ) ;
  assign n16660 = n16659 ^ n16658 ^ n16657 ;
  assign n16661 = n3049 ^ n1591 ^ 1'b0 ;
  assign n16662 = ~n6866 & n16661 ;
  assign n16663 = n16662 ^ n9351 ^ 1'b0 ;
  assign n16664 = n13030 ^ n12262 ^ 1'b0 ;
  assign n16665 = ~n2089 & n16664 ;
  assign n16666 = n16663 & n16665 ;
  assign n16667 = n3625 & n16666 ;
  assign n16668 = n4570 & n16667 ;
  assign n16670 = n5811 ^ n637 ^ 1'b0 ;
  assign n16669 = ~n6393 & n8865 ;
  assign n16671 = n16670 ^ n16669 ^ 1'b0 ;
  assign n16672 = ~x29 & n3532 ;
  assign n16681 = n12232 ^ n8744 ^ n7761 ;
  assign n16682 = ~n1350 & n3752 ;
  assign n16683 = ~n16681 & n16682 ;
  assign n16673 = ~n3063 & n4556 ;
  assign n16674 = n16673 ^ n1593 ^ n1473 ;
  assign n16676 = ~n2319 & n2547 ;
  assign n16677 = n3474 & n16676 ;
  assign n16675 = n1898 ^ n586 ^ 1'b0 ;
  assign n16678 = n16677 ^ n16675 ^ 1'b0 ;
  assign n16679 = n16674 | n16678 ;
  assign n16680 = ~n12319 & n16679 ;
  assign n16684 = n16683 ^ n16680 ^ 1'b0 ;
  assign n16685 = ~n6372 & n16684 ;
  assign n16686 = n16685 ^ n9172 ^ n2125 ;
  assign n16687 = n11483 ^ n10386 ^ n1337 ;
  assign n16688 = n14817 ^ n10563 ^ 1'b0 ;
  assign n16689 = ( n388 & n1384 ) | ( n388 & ~n2646 ) | ( n1384 & ~n2646 ) ;
  assign n16690 = n16689 ^ n15038 ^ n9568 ;
  assign n16691 = n4682 | n5016 ;
  assign n16692 = ~n2093 & n10917 ;
  assign n16693 = n16692 ^ n12985 ^ 1'b0 ;
  assign n16694 = n16691 | n16693 ;
  assign n16695 = ( ~n5043 & n13518 ) | ( ~n5043 & n16694 ) | ( n13518 & n16694 ) ;
  assign n16696 = n5196 ^ n4068 ^ 1'b0 ;
  assign n16697 = n6398 & n16696 ;
  assign n16698 = ( ~n14284 & n15820 ) | ( ~n14284 & n16697 ) | ( n15820 & n16697 ) ;
  assign n16699 = n6081 & ~n7349 ;
  assign n16700 = n16699 ^ n13179 ^ n3095 ;
  assign n16703 = ~n1968 & n12266 ;
  assign n16704 = ~n5471 & n16703 ;
  assign n16705 = n16704 ^ n10458 ^ 1'b0 ;
  assign n16701 = ( n4924 & n9066 ) | ( n4924 & n9299 ) | ( n9066 & n9299 ) ;
  assign n16702 = n4156 & ~n16701 ;
  assign n16706 = n16705 ^ n16702 ^ 1'b0 ;
  assign n16707 = ~n16485 & n16706 ;
  assign n16708 = n12634 | n15576 ;
  assign n16709 = n16708 ^ n5777 ^ 1'b0 ;
  assign n16710 = n13204 ^ n4390 ^ 1'b0 ;
  assign n16711 = ~n2022 & n16710 ;
  assign n16712 = ~n11178 & n16711 ;
  assign n16713 = ~n9668 & n16712 ;
  assign n16714 = n1647 | n16713 ;
  assign n16715 = n16714 ^ n13745 ^ 1'b0 ;
  assign n16716 = n15879 ^ n11641 ^ n4779 ;
  assign n16717 = n8446 | n16716 ;
  assign n16718 = n16717 ^ n1359 ^ 1'b0 ;
  assign n16719 = ( ~n6809 & n7988 ) | ( ~n6809 & n12222 ) | ( n7988 & n12222 ) ;
  assign n16720 = n1331 & n4984 ;
  assign n16721 = n14717 & ~n16720 ;
  assign n16722 = n3459 ^ n2143 ^ n2116 ;
  assign n16723 = n4878 & ~n16722 ;
  assign n16724 = n16723 ^ n10240 ^ 1'b0 ;
  assign n16725 = n14477 ^ n3562 ^ n3016 ;
  assign n16726 = n1489 & ~n7248 ;
  assign n16727 = n16726 ^ n7057 ^ 1'b0 ;
  assign n16728 = n16727 ^ n16485 ^ 1'b0 ;
  assign n16729 = n9545 & n16728 ;
  assign n16730 = n13826 ^ n6171 ^ n4970 ;
  assign n16731 = n16730 ^ n1883 ^ 1'b0 ;
  assign n16732 = n7707 ^ n1075 ^ 1'b0 ;
  assign n16733 = n12059 ^ n1738 ^ 1'b0 ;
  assign n16734 = n16733 ^ n16670 ^ n9547 ;
  assign n16735 = n16734 ^ n15209 ^ 1'b0 ;
  assign n16736 = ~n16224 & n16735 ;
  assign n16737 = n5746 & ~n7817 ;
  assign n16738 = n16737 ^ n4712 ^ 1'b0 ;
  assign n16739 = n1508 | n16738 ;
  assign n16740 = n5309 & ~n16739 ;
  assign n16741 = n5094 ^ n2592 ^ 1'b0 ;
  assign n16742 = n16740 | n16741 ;
  assign n16743 = n3424 ^ n2260 ^ n593 ;
  assign n16744 = n16743 ^ n7731 ^ n2963 ;
  assign n16745 = n9901 & n16744 ;
  assign n16746 = ~n10791 & n16745 ;
  assign n16747 = ( ~n6666 & n7363 ) | ( ~n6666 & n16746 ) | ( n7363 & n16746 ) ;
  assign n16748 = ( ~n6821 & n7119 ) | ( ~n6821 & n11463 ) | ( n7119 & n11463 ) ;
  assign n16749 = ~n11007 & n15744 ;
  assign n16750 = ( n4740 & n16748 ) | ( n4740 & ~n16749 ) | ( n16748 & ~n16749 ) ;
  assign n16751 = n7637 ^ n6326 ^ 1'b0 ;
  assign n16752 = ~n687 & n16751 ;
  assign n16753 = ~n5470 & n16752 ;
  assign n16754 = ( n8359 & n12380 ) | ( n8359 & ~n12454 ) | ( n12380 & ~n12454 ) ;
  assign n16755 = ( ~n12692 & n16753 ) | ( ~n12692 & n16754 ) | ( n16753 & n16754 ) ;
  assign n16756 = n9234 & n15757 ;
  assign n16757 = ~n3750 & n16756 ;
  assign n16758 = n2430 & ~n8727 ;
  assign n16767 = ~n2767 & n7588 ;
  assign n16768 = n16767 ^ n10654 ^ 1'b0 ;
  assign n16759 = n6260 ^ n6085 ^ n2502 ;
  assign n16760 = ~n1252 & n16759 ;
  assign n16761 = n16760 ^ n7752 ^ n1663 ;
  assign n16762 = n3160 & n6299 ;
  assign n16763 = n16762 ^ n2606 ^ 1'b0 ;
  assign n16764 = ( ~n5223 & n8802 ) | ( ~n5223 & n16763 ) | ( n8802 & n16763 ) ;
  assign n16765 = n7014 | n16764 ;
  assign n16766 = ( n2265 & ~n16761 ) | ( n2265 & n16765 ) | ( ~n16761 & n16765 ) ;
  assign n16769 = n16768 ^ n16766 ^ n10122 ;
  assign n16770 = ( n6009 & n14492 ) | ( n6009 & n15398 ) | ( n14492 & n15398 ) ;
  assign n16772 = n4731 | n8145 ;
  assign n16771 = n8227 ^ n7089 ^ n6143 ;
  assign n16773 = n16772 ^ n16771 ^ 1'b0 ;
  assign n16774 = n6082 & n16773 ;
  assign n16775 = ( n2667 & n4763 ) | ( n2667 & n16774 ) | ( n4763 & n16774 ) ;
  assign n16776 = n10212 | n16775 ;
  assign n16777 = ~n10254 & n13279 ;
  assign n16778 = n16777 ^ n10572 ^ 1'b0 ;
  assign n16779 = ( n3996 & ~n11901 ) | ( n3996 & n16778 ) | ( ~n11901 & n16778 ) ;
  assign n16780 = ( ~n5954 & n6219 ) | ( ~n5954 & n13307 ) | ( n6219 & n13307 ) ;
  assign n16781 = n16780 ^ n7561 ^ 1'b0 ;
  assign n16782 = n6654 | n16781 ;
  assign n16784 = ( x109 & n750 ) | ( x109 & ~n2792 ) | ( n750 & ~n2792 ) ;
  assign n16785 = x216 & ~n11725 ;
  assign n16786 = n16785 ^ n4507 ^ 1'b0 ;
  assign n16787 = n16784 & ~n16786 ;
  assign n16788 = n7526 & n16787 ;
  assign n16783 = n7464 | n8933 ;
  assign n16789 = n16788 ^ n16783 ^ 1'b0 ;
  assign n16790 = n16789 ^ n9886 ^ 1'b0 ;
  assign n16791 = n3958 & ~n16790 ;
  assign n16792 = n8868 ^ n4703 ^ n1941 ;
  assign n16793 = ~n3643 & n9845 ;
  assign n16794 = n3942 & n16793 ;
  assign n16796 = n6216 ^ n3699 ^ 1'b0 ;
  assign n16797 = n5271 | n16796 ;
  assign n16795 = n7644 & ~n10549 ;
  assign n16798 = n16797 ^ n16795 ^ 1'b0 ;
  assign n16799 = n5681 | n8700 ;
  assign n16800 = n1099 | n16799 ;
  assign n16801 = n7753 & n16800 ;
  assign n16802 = n11021 ^ n5857 ^ x87 ;
  assign n16803 = n16802 ^ n11886 ^ 1'b0 ;
  assign n16804 = ( n9047 & n9568 ) | ( n9047 & ~n16803 ) | ( n9568 & ~n16803 ) ;
  assign n16805 = n4738 | n10569 ;
  assign n16806 = n16805 ^ n9237 ^ 1'b0 ;
  assign n16807 = n16806 ^ n10990 ^ n4847 ;
  assign n16808 = ( x221 & n13203 ) | ( x221 & ~n16807 ) | ( n13203 & ~n16807 ) ;
  assign n16809 = n7401 ^ n3257 ^ 1'b0 ;
  assign n16810 = n8433 ^ n4868 ^ n1051 ;
  assign n16811 = n14952 | n16810 ;
  assign n16812 = ( n2261 & n8398 ) | ( n2261 & n16811 ) | ( n8398 & n16811 ) ;
  assign n16813 = n10753 ^ n1564 ^ 1'b0 ;
  assign n16814 = n14735 ^ n9722 ^ 1'b0 ;
  assign n16815 = n12273 ^ n7304 ^ 1'b0 ;
  assign n16816 = ~n16814 & n16815 ;
  assign n16817 = x110 & n8116 ;
  assign n16818 = n16817 ^ n4741 ^ 1'b0 ;
  assign n16821 = ~n1325 & n2425 ;
  assign n16822 = ~n9735 & n16821 ;
  assign n16819 = n4852 & ~n6766 ;
  assign n16820 = n16819 ^ n366 ^ 1'b0 ;
  assign n16823 = n16822 ^ n16820 ^ 1'b0 ;
  assign n16824 = n16818 | n16823 ;
  assign n16825 = n481 & ~n6653 ;
  assign n16826 = n16825 ^ n2330 ^ 1'b0 ;
  assign n16827 = n16826 ^ n4935 ^ n2858 ;
  assign n16828 = n16827 ^ n11324 ^ n4185 ;
  assign n16829 = n16828 ^ n15827 ^ n7939 ;
  assign n16830 = n5444 ^ n1921 ^ 1'b0 ;
  assign n16831 = n8917 | n16830 ;
  assign n16832 = n16831 ^ n5369 ^ x183 ;
  assign n16833 = n11673 & n13032 ;
  assign n16834 = ~n8450 & n16833 ;
  assign n16835 = n9381 ^ n1030 ^ 1'b0 ;
  assign n16836 = n16834 | n16835 ;
  assign n16837 = n3018 | n4987 ;
  assign n16838 = n16837 ^ n2944 ^ 1'b0 ;
  assign n16839 = n12840 ^ n11349 ^ n7716 ;
  assign n16840 = ~n16838 & n16839 ;
  assign n16841 = ( n1333 & ~n7064 ) | ( n1333 & n7774 ) | ( ~n7064 & n7774 ) ;
  assign n16842 = ~n5137 & n7245 ;
  assign n16843 = ( n780 & n4793 ) | ( n780 & n16842 ) | ( n4793 & n16842 ) ;
  assign n16844 = n15513 & ~n16843 ;
  assign n16845 = ( n6190 & n16841 ) | ( n6190 & n16844 ) | ( n16841 & n16844 ) ;
  assign n16846 = n2944 & n4934 ;
  assign n16847 = n16846 ^ n5820 ^ n1660 ;
  assign n16848 = n16847 ^ n7288 ^ 1'b0 ;
  assign n16849 = n16848 ^ n16116 ^ 1'b0 ;
  assign n16850 = ~n3418 & n13715 ;
  assign n16851 = n16850 ^ n3787 ^ 1'b0 ;
  assign n16852 = ( n6625 & n7020 ) | ( n6625 & ~n16851 ) | ( n7020 & ~n16851 ) ;
  assign n16853 = n3122 | n4047 ;
  assign n16854 = n4786 & ~n16853 ;
  assign n16855 = ( x135 & n7643 ) | ( x135 & n13581 ) | ( n7643 & n13581 ) ;
  assign n16856 = n16854 | n16855 ;
  assign n16857 = n16852 | n16856 ;
  assign n16858 = ( ~n8864 & n9279 ) | ( ~n8864 & n11059 ) | ( n9279 & n11059 ) ;
  assign n16859 = n5785 & n16858 ;
  assign n16860 = n6125 & n16859 ;
  assign n16861 = n10216 ^ n7538 ^ n4866 ;
  assign n16862 = x108 & ~n16085 ;
  assign n16863 = n8303 & n16862 ;
  assign n16864 = n13632 ^ n4278 ^ 1'b0 ;
  assign n16865 = n9673 ^ n8295 ^ 1'b0 ;
  assign n16866 = n7676 & n16865 ;
  assign n16867 = n9664 & n13830 ;
  assign n16868 = n16867 ^ n5057 ^ n583 ;
  assign n16869 = n12162 ^ n958 ^ 1'b0 ;
  assign n16870 = n3858 & n16869 ;
  assign n16871 = n11838 ^ n5344 ^ n1952 ;
  assign n16872 = n13020 ^ n8706 ^ n2468 ;
  assign n16873 = ( x35 & n1868 ) | ( x35 & ~n3319 ) | ( n1868 & ~n3319 ) ;
  assign n16874 = n7216 & ~n16873 ;
  assign n16875 = ~n5666 & n16874 ;
  assign n16876 = n14365 | n16323 ;
  assign n16877 = n5836 & ~n16876 ;
  assign n16878 = n2796 & ~n8458 ;
  assign n16879 = n3945 & ~n15566 ;
  assign n16880 = ~n16878 & n16879 ;
  assign n16881 = n2464 ^ n1808 ^ 1'b0 ;
  assign n16882 = n10719 & ~n16881 ;
  assign n16883 = n4737 & n16882 ;
  assign n16884 = ( n13149 & ~n15464 ) | ( n13149 & n16883 ) | ( ~n15464 & n16883 ) ;
  assign n16885 = n5720 | n9237 ;
  assign n16886 = n394 & ~n4553 ;
  assign n16887 = n16886 ^ n9568 ^ 1'b0 ;
  assign n16888 = n16887 ^ n10053 ^ n732 ;
  assign n16889 = n5829 & n16888 ;
  assign n16890 = ~n9508 & n16889 ;
  assign n16891 = n4192 & n9315 ;
  assign n16892 = n16891 ^ n3767 ^ 1'b0 ;
  assign n16893 = n8508 & n16892 ;
  assign n16894 = n5050 ^ n2745 ^ n2276 ;
  assign n16895 = n7019 & n16894 ;
  assign n16896 = n16893 & ~n16895 ;
  assign n16897 = ( ~n684 & n12072 ) | ( ~n684 & n13291 ) | ( n12072 & n13291 ) ;
  assign n16903 = n2399 & ~n10887 ;
  assign n16899 = n474 | n14698 ;
  assign n16900 = n16899 ^ x154 ^ 1'b0 ;
  assign n16898 = ~n3008 & n13934 ;
  assign n16901 = n16900 ^ n16898 ^ 1'b0 ;
  assign n16902 = n2712 & n16901 ;
  assign n16904 = n16903 ^ n16902 ^ 1'b0 ;
  assign n16905 = n16904 ^ n15074 ^ n8525 ;
  assign n16908 = ~n1520 & n8940 ;
  assign n16909 = ( n3002 & ~n12536 ) | ( n3002 & n16908 ) | ( ~n12536 & n16908 ) ;
  assign n16906 = n7208 & ~n9585 ;
  assign n16907 = n16751 & ~n16906 ;
  assign n16910 = n16909 ^ n16907 ^ 1'b0 ;
  assign n16911 = n8375 | n16910 ;
  assign n16912 = ( n1920 & ~n15285 ) | ( n1920 & n15919 ) | ( ~n15285 & n15919 ) ;
  assign n16913 = n16912 ^ n15685 ^ 1'b0 ;
  assign n16916 = ~n6282 & n7802 ;
  assign n16917 = n16916 ^ n15680 ^ 1'b0 ;
  assign n16914 = n4254 & n4419 ;
  assign n16915 = n16914 ^ n5301 ^ n3995 ;
  assign n16918 = n16917 ^ n16915 ^ n1647 ;
  assign n16919 = ~n6088 & n14543 ;
  assign n16920 = n16919 ^ n16841 ^ 1'b0 ;
  assign n16926 = ( n8709 & ~n11296 ) | ( n8709 & n15337 ) | ( ~n11296 & n15337 ) ;
  assign n16927 = n16926 ^ n6451 ^ 1'b0 ;
  assign n16921 = n5038 ^ n1527 ^ 1'b0 ;
  assign n16922 = n2924 | n16921 ;
  assign n16923 = n7700 & n14197 ;
  assign n16924 = n16923 ^ n9644 ^ 1'b0 ;
  assign n16925 = ( ~n15644 & n16922 ) | ( ~n15644 & n16924 ) | ( n16922 & n16924 ) ;
  assign n16928 = n16927 ^ n16925 ^ n10865 ;
  assign n16929 = n3920 | n9196 ;
  assign n16930 = ( n4291 & n7465 ) | ( n4291 & ~n16929 ) | ( n7465 & ~n16929 ) ;
  assign n16931 = ( n16920 & n16928 ) | ( n16920 & n16930 ) | ( n16928 & n16930 ) ;
  assign n16932 = n1236 ^ n990 ^ x113 ;
  assign n16933 = n16932 ^ n4592 ^ 1'b0 ;
  assign n16934 = n1307 & n16933 ;
  assign n16935 = n16934 ^ n8817 ^ n6417 ;
  assign n16936 = n16935 ^ n1028 ^ 1'b0 ;
  assign n16937 = n6803 | n16936 ;
  assign n16938 = n6045 & ~n16937 ;
  assign n16939 = n16938 ^ n12708 ^ 1'b0 ;
  assign n16940 = n3325 ^ n540 ^ 1'b0 ;
  assign n16941 = n6175 ^ n3280 ^ 1'b0 ;
  assign n16942 = ~n16940 & n16941 ;
  assign n16943 = ~n15020 & n16194 ;
  assign n16944 = ~n16942 & n16943 ;
  assign n16945 = n2998 ^ n1969 ^ n1537 ;
  assign n16946 = ( n2554 & n15282 ) | ( n2554 & ~n16945 ) | ( n15282 & ~n16945 ) ;
  assign n16947 = n4360 & n9100 ;
  assign n16948 = n16947 ^ n8087 ^ 1'b0 ;
  assign n16949 = ~n2983 & n16134 ;
  assign n16950 = n16949 ^ n10425 ^ 1'b0 ;
  assign n16951 = n446 | n1494 ;
  assign n16952 = ( ~n7600 & n8227 ) | ( ~n7600 & n16951 ) | ( n8227 & n16951 ) ;
  assign n16953 = n16952 ^ n14594 ^ n8515 ;
  assign n16954 = n9865 ^ n8999 ^ 1'b0 ;
  assign n16955 = n6851 & ~n16954 ;
  assign n16956 = n16955 ^ n15930 ^ n562 ;
  assign n16957 = n9164 ^ n3429 ^ 1'b0 ;
  assign n16960 = n5540 ^ n452 ^ 1'b0 ;
  assign n16961 = ( n1576 & ~n4479 ) | ( n1576 & n16960 ) | ( ~n4479 & n16960 ) ;
  assign n16958 = ( ~n5716 & n6142 ) | ( ~n5716 & n11109 ) | ( n6142 & n11109 ) ;
  assign n16959 = ( n3598 & ~n8153 ) | ( n3598 & n16958 ) | ( ~n8153 & n16958 ) ;
  assign n16962 = n16961 ^ n16959 ^ x75 ;
  assign n16963 = n7318 | n8591 ;
  assign n16964 = n2244 & ~n16963 ;
  assign n16965 = n1643 | n16964 ;
  assign n16966 = n5384 | n16965 ;
  assign n16967 = n8905 & n16966 ;
  assign n16968 = n16967 ^ n3114 ^ 1'b0 ;
  assign n16969 = n16968 ^ n10016 ^ 1'b0 ;
  assign n16970 = n431 | n1113 ;
  assign n16971 = n16970 ^ n11924 ^ n9116 ;
  assign n16972 = n5455 | n16971 ;
  assign n16973 = n16972 ^ n2550 ^ 1'b0 ;
  assign n16974 = ( ~n8227 & n11699 ) | ( ~n8227 & n16973 ) | ( n11699 & n16973 ) ;
  assign n16975 = n10536 ^ n2369 ^ 1'b0 ;
  assign n16976 = n3382 | n16975 ;
  assign n16977 = n16974 | n16976 ;
  assign n16981 = ( n3927 & n4785 ) | ( n3927 & ~n10085 ) | ( n4785 & ~n10085 ) ;
  assign n16982 = n7709 & n16981 ;
  assign n16978 = ~n5249 & n8644 ;
  assign n16979 = ~n7796 & n8651 ;
  assign n16980 = n16978 | n16979 ;
  assign n16983 = n16982 ^ n16980 ^ n8477 ;
  assign n16984 = n16284 ^ n9757 ^ n6818 ;
  assign n16985 = n11986 ^ n1188 ^ 1'b0 ;
  assign n16986 = n16985 ^ n6061 ^ x218 ;
  assign n16987 = n1325 & n4533 ;
  assign n16988 = n16772 & ~n16987 ;
  assign n16989 = n4512 & n16988 ;
  assign n16990 = n11559 ^ n7633 ^ 1'b0 ;
  assign n16991 = n16990 ^ n6455 ^ 1'b0 ;
  assign n16992 = n16989 | n16991 ;
  assign n16993 = ( n2167 & n2944 ) | ( n2167 & n4386 ) | ( n2944 & n4386 ) ;
  assign n16994 = ( ~n2538 & n3824 ) | ( ~n2538 & n7250 ) | ( n3824 & n7250 ) ;
  assign n16995 = n16993 & ~n16994 ;
  assign n16996 = ~n780 & n9293 ;
  assign n16997 = ~n1158 & n16996 ;
  assign n16998 = n16997 ^ n7775 ^ 1'b0 ;
  assign n16999 = n16995 | n16998 ;
  assign n17005 = n7617 | n8529 ;
  assign n17006 = n4759 | n17005 ;
  assign n17003 = n2225 | n9526 ;
  assign n17004 = n5817 | n17003 ;
  assign n17000 = n6505 & n10745 ;
  assign n17001 = n17000 ^ n3033 ^ 1'b0 ;
  assign n17002 = n7108 & ~n17001 ;
  assign n17007 = n17006 ^ n17004 ^ n17002 ;
  assign n17008 = n3834 ^ n3711 ^ 1'b0 ;
  assign n17009 = ( ~n7382 & n8703 ) | ( ~n7382 & n12750 ) | ( n8703 & n12750 ) ;
  assign n17010 = n15906 ^ n7160 ^ n3457 ;
  assign n17014 = n10995 ^ n5773 ^ n4073 ;
  assign n17011 = n16231 ^ n8386 ^ n4713 ;
  assign n17012 = n17011 ^ n4856 ^ n2830 ;
  assign n17013 = n17012 ^ n12960 ^ n2159 ;
  assign n17015 = n17014 ^ n17013 ^ 1'b0 ;
  assign n17016 = n4266 | n9050 ;
  assign n17017 = n17016 ^ n8644 ^ 1'b0 ;
  assign n17018 = x61 & ~n17017 ;
  assign n17019 = ~n12205 & n14870 ;
  assign n17025 = n6388 ^ n2504 ^ 1'b0 ;
  assign n17026 = ( n3085 & n9865 ) | ( n3085 & n17025 ) | ( n9865 & n17025 ) ;
  assign n17027 = n17026 ^ n4396 ^ 1'b0 ;
  assign n17021 = ~n5984 & n14274 ;
  assign n17022 = n4466 & n17021 ;
  assign n17020 = n3687 & n7488 ;
  assign n17023 = n17022 ^ n17020 ^ 1'b0 ;
  assign n17024 = ~n8645 & n17023 ;
  assign n17028 = n17027 ^ n17024 ^ 1'b0 ;
  assign n17029 = ~n13840 & n16981 ;
  assign n17030 = n17029 ^ n12840 ^ 1'b0 ;
  assign n17031 = n16968 ^ n5492 ^ 1'b0 ;
  assign n17032 = n5662 & ~n17031 ;
  assign n17033 = n12873 & n17032 ;
  assign n17034 = n3711 & ~n7152 ;
  assign n17035 = n2184 | n7320 ;
  assign n17036 = n17035 ^ n10234 ^ n5530 ;
  assign n17037 = ( ~n1611 & n4077 ) | ( ~n1611 & n8364 ) | ( n4077 & n8364 ) ;
  assign n17038 = n17037 ^ x158 ^ 1'b0 ;
  assign n17039 = n6598 & ~n6649 ;
  assign n17040 = n587 & n17039 ;
  assign n17041 = ( n1052 & n9197 ) | ( n1052 & ~n17040 ) | ( n9197 & ~n17040 ) ;
  assign n17043 = n6178 | n11328 ;
  assign n17044 = n10433 & ~n17043 ;
  assign n17042 = ( n7871 & ~n10448 ) | ( n7871 & n15262 ) | ( ~n10448 & n15262 ) ;
  assign n17045 = n17044 ^ n17042 ^ 1'b0 ;
  assign n17046 = n11769 & n17045 ;
  assign n17047 = ( n1422 & n1961 ) | ( n1422 & ~n4996 ) | ( n1961 & ~n4996 ) ;
  assign n17048 = n13646 ^ n12101 ^ n5989 ;
  assign n17049 = ( n11264 & n17047 ) | ( n11264 & ~n17048 ) | ( n17047 & ~n17048 ) ;
  assign n17050 = n10601 & n17049 ;
  assign n17051 = n17050 ^ n12186 ^ 1'b0 ;
  assign n17052 = n17051 ^ n4585 ^ 1'b0 ;
  assign n17053 = n4871 | n10236 ;
  assign n17054 = n17053 ^ n4680 ^ 1'b0 ;
  assign n17055 = n2372 & n4555 ;
  assign n17056 = n17054 & n17055 ;
  assign n17057 = n7943 ^ n3214 ^ n3133 ;
  assign n17058 = ( ~n6047 & n6764 ) | ( ~n6047 & n17057 ) | ( n6764 & n17057 ) ;
  assign n17059 = n11027 | n17058 ;
  assign n17060 = n1738 & ~n17059 ;
  assign n17061 = n3562 | n17060 ;
  assign n17062 = n17061 ^ n13094 ^ 1'b0 ;
  assign n17064 = n10376 & ~n12026 ;
  assign n17063 = n12788 | n16974 ;
  assign n17065 = n17064 ^ n17063 ^ 1'b0 ;
  assign n17066 = ( n14614 & ~n17062 ) | ( n14614 & n17065 ) | ( ~n17062 & n17065 ) ;
  assign n17067 = n17066 ^ n13238 ^ 1'b0 ;
  assign n17068 = n6703 ^ n3600 ^ 1'b0 ;
  assign n17069 = n4260 & ~n17068 ;
  assign n17070 = n13995 ^ x36 ^ 1'b0 ;
  assign n17071 = ( n3097 & n5635 ) | ( n3097 & ~n9186 ) | ( n5635 & ~n9186 ) ;
  assign n17072 = n4066 | n17071 ;
  assign n17073 = n6430 & ~n17072 ;
  assign n17074 = n17070 | n17073 ;
  assign n17075 = ( n12360 & n17069 ) | ( n12360 & ~n17074 ) | ( n17069 & ~n17074 ) ;
  assign n17076 = n3565 ^ n3003 ^ n872 ;
  assign n17077 = ( n3926 & ~n8910 ) | ( n3926 & n17076 ) | ( ~n8910 & n17076 ) ;
  assign n17078 = n8818 ^ n2175 ^ 1'b0 ;
  assign n17079 = ( n871 & ~n10935 ) | ( n871 & n17078 ) | ( ~n10935 & n17078 ) ;
  assign n17080 = n17079 ^ n4987 ^ 1'b0 ;
  assign n17081 = ~n17077 & n17080 ;
  assign n17082 = ( n3991 & ~n6732 ) | ( n3991 & n13624 ) | ( ~n6732 & n13624 ) ;
  assign n17083 = n5538 & ~n15460 ;
  assign n17084 = x62 & ~n17083 ;
  assign n17085 = n17084 ^ n14111 ^ 1'b0 ;
  assign n17086 = n1742 | n17085 ;
  assign n17087 = n17086 ^ n12817 ^ n4061 ;
  assign n17088 = n8591 ^ n7145 ^ 1'b0 ;
  assign n17089 = ~n9067 & n17088 ;
  assign n17090 = n8430 ^ n3579 ^ 1'b0 ;
  assign n17091 = n2547 & ~n17090 ;
  assign n17096 = n5688 & n7732 ;
  assign n17097 = n17096 ^ n6307 ^ n5473 ;
  assign n17094 = n8594 | n8870 ;
  assign n17095 = n4620 | n17094 ;
  assign n17092 = n12798 ^ n825 ^ 1'b0 ;
  assign n17093 = n9008 & n17092 ;
  assign n17098 = n17097 ^ n17095 ^ n17093 ;
  assign n17099 = ( n7377 & n17091 ) | ( n7377 & n17098 ) | ( n17091 & n17098 ) ;
  assign n17104 = n4951 | n11120 ;
  assign n17105 = ( ~n1535 & n9125 ) | ( ~n1535 & n10001 ) | ( n9125 & n10001 ) ;
  assign n17106 = ( n6265 & ~n17104 ) | ( n6265 & n17105 ) | ( ~n17104 & n17105 ) ;
  assign n17101 = n6035 ^ n2952 ^ n602 ;
  assign n17100 = n1161 | n9564 ;
  assign n17102 = n17101 ^ n17100 ^ 1'b0 ;
  assign n17103 = ( ~n3347 & n9485 ) | ( ~n3347 & n17102 ) | ( n9485 & n17102 ) ;
  assign n17107 = n17106 ^ n17103 ^ 1'b0 ;
  assign n17114 = ( n2907 & n4567 ) | ( n2907 & ~n4925 ) | ( n4567 & ~n4925 ) ;
  assign n17108 = n14155 ^ n2215 ^ 1'b0 ;
  assign n17109 = n14318 & n17108 ;
  assign n17110 = n2500 & n2686 ;
  assign n17111 = n17110 ^ n2649 ^ 1'b0 ;
  assign n17112 = n3472 | n17111 ;
  assign n17113 = n17109 | n17112 ;
  assign n17115 = n17114 ^ n17113 ^ 1'b0 ;
  assign n17116 = n10214 ^ n2251 ^ 1'b0 ;
  assign n17117 = n3638 & ~n17116 ;
  assign n17122 = ( n898 & ~n1886 ) | ( n898 & n6021 ) | ( ~n1886 & n6021 ) ;
  assign n17118 = n6071 & n10638 ;
  assign n17119 = ~n12202 & n17118 ;
  assign n17120 = ( x221 & ~n6906 ) | ( x221 & n12708 ) | ( ~n6906 & n12708 ) ;
  assign n17121 = n17119 & n17120 ;
  assign n17123 = n17122 ^ n17121 ^ 1'b0 ;
  assign n17124 = n17123 ^ n9959 ^ 1'b0 ;
  assign n17125 = n17117 & n17124 ;
  assign n17126 = n16007 ^ n8249 ^ 1'b0 ;
  assign n17127 = n17125 & ~n17126 ;
  assign n17128 = ~n6440 & n8163 ;
  assign n17129 = n5091 | n12077 ;
  assign n17130 = n295 & ~n17129 ;
  assign n17131 = n3697 ^ n2844 ^ 1'b0 ;
  assign n17132 = n2001 | n17131 ;
  assign n17133 = n11050 | n17132 ;
  assign n17134 = n17133 ^ n8011 ^ 1'b0 ;
  assign n17135 = n2159 & ~n2737 ;
  assign n17136 = n17135 ^ n1778 ^ 1'b0 ;
  assign n17137 = n17136 ^ n7895 ^ n2121 ;
  assign n17138 = n17137 ^ n13317 ^ 1'b0 ;
  assign n17139 = n17134 & ~n17138 ;
  assign n17140 = n2391 | n5489 ;
  assign n17141 = ( ~n536 & n774 ) | ( ~n536 & n17140 ) | ( n774 & n17140 ) ;
  assign n17142 = n17141 ^ n12249 ^ 1'b0 ;
  assign n17143 = n8413 ^ n7358 ^ x169 ;
  assign n17144 = ( x242 & n13633 ) | ( x242 & ~n17143 ) | ( n13633 & ~n17143 ) ;
  assign n17145 = n8433 ^ n4835 ^ n4016 ;
  assign n17146 = n3503 & ~n3541 ;
  assign n17147 = n17146 ^ n11953 ^ 1'b0 ;
  assign n17148 = n17145 | n17147 ;
  assign n17149 = ( n5899 & n14137 ) | ( n5899 & ~n17148 ) | ( n14137 & ~n17148 ) ;
  assign n17150 = n11495 ^ n2178 ^ 1'b0 ;
  assign n17151 = n6406 & n6598 ;
  assign n17152 = n6809 & n17151 ;
  assign n17155 = n11419 ^ n10786 ^ n8480 ;
  assign n17153 = n1783 & n5968 ;
  assign n17154 = n11937 & n17153 ;
  assign n17156 = n17155 ^ n17154 ^ n14267 ;
  assign n17157 = n12345 | n13116 ;
  assign n17158 = ~n9861 & n15173 ;
  assign n17159 = ~n16928 & n17158 ;
  assign n17167 = n2367 ^ n2128 ^ 1'b0 ;
  assign n17168 = n15301 & ~n17167 ;
  assign n17169 = n17168 ^ n7949 ^ n4615 ;
  assign n17170 = n17169 ^ n12406 ^ 1'b0 ;
  assign n17171 = ~n14557 & n17170 ;
  assign n17160 = n7781 ^ n4053 ^ n259 ;
  assign n17161 = ( ~n13115 & n13439 ) | ( ~n13115 & n17160 ) | ( n13439 & n17160 ) ;
  assign n17162 = n17161 ^ n8780 ^ 1'b0 ;
  assign n17164 = n1405 & n5902 ;
  assign n17163 = n1179 & ~n2028 ;
  assign n17165 = n17164 ^ n17163 ^ 1'b0 ;
  assign n17166 = n17162 & n17165 ;
  assign n17172 = n17171 ^ n17166 ^ 1'b0 ;
  assign n17173 = n14573 ^ n14140 ^ 1'b0 ;
  assign n17174 = n6251 & n17173 ;
  assign n17175 = ( n11607 & n12143 ) | ( n11607 & n16526 ) | ( n12143 & n16526 ) ;
  assign n17178 = n4624 | n16987 ;
  assign n17179 = n4378 & ~n17178 ;
  assign n17176 = n11109 ^ n7898 ^ 1'b0 ;
  assign n17177 = ~n11570 & n17176 ;
  assign n17180 = n17179 ^ n17177 ^ 1'b0 ;
  assign n17183 = n9852 ^ n4662 ^ 1'b0 ;
  assign n17181 = n12217 ^ x78 ^ 1'b0 ;
  assign n17182 = n1475 & n17181 ;
  assign n17184 = n17183 ^ n17182 ^ 1'b0 ;
  assign n17188 = n7183 ^ n6159 ^ n926 ;
  assign n17186 = n6171 ^ n1738 ^ 1'b0 ;
  assign n17185 = n10043 & n12231 ;
  assign n17187 = n17186 ^ n17185 ^ 1'b0 ;
  assign n17189 = n17188 ^ n17187 ^ n5347 ;
  assign n17190 = ~n6227 & n13983 ;
  assign n17191 = n13059 & n17190 ;
  assign n17192 = n16733 ^ n5076 ^ n757 ;
  assign n17193 = ~n5556 & n17192 ;
  assign n17194 = n4131 & ~n17193 ;
  assign n17195 = n17194 ^ x194 ^ 1'b0 ;
  assign n17207 = n1188 & ~n9024 ;
  assign n17208 = n8555 & n17207 ;
  assign n17196 = n11620 ^ n410 ^ x109 ;
  assign n17197 = n4600 ^ x31 ^ 1'b0 ;
  assign n17198 = n4086 & ~n17197 ;
  assign n17199 = n1697 | n6999 ;
  assign n17200 = ( n4532 & n9247 ) | ( n4532 & n17199 ) | ( n9247 & n17199 ) ;
  assign n17201 = n5805 ^ n4419 ^ n1761 ;
  assign n17202 = n17201 ^ n10702 ^ 1'b0 ;
  assign n17203 = n17200 | n17202 ;
  assign n17204 = ( n8004 & ~n17198 ) | ( n8004 & n17203 ) | ( ~n17198 & n17203 ) ;
  assign n17205 = n17204 ^ n1570 ^ 1'b0 ;
  assign n17206 = n17196 & ~n17205 ;
  assign n17209 = n17208 ^ n17206 ^ 1'b0 ;
  assign n17210 = ( n14079 & n15214 ) | ( n14079 & ~n17029 ) | ( n15214 & ~n17029 ) ;
  assign n17211 = ~n989 & n15851 ;
  assign n17212 = n17211 ^ n7083 ^ 1'b0 ;
  assign n17213 = n11735 ^ n6103 ^ 1'b0 ;
  assign n17214 = n8070 & ~n17213 ;
  assign n17215 = n6893 ^ n2221 ^ 1'b0 ;
  assign n17216 = n17214 & n17215 ;
  assign n17217 = n8387 & n17216 ;
  assign n17218 = n17217 ^ n11966 ^ 1'b0 ;
  assign n17219 = n11177 ^ n2588 ^ x137 ;
  assign n17220 = ( ~n4118 & n7717 ) | ( ~n4118 & n17219 ) | ( n7717 & n17219 ) ;
  assign n17221 = ( n4394 & n17218 ) | ( n4394 & n17220 ) | ( n17218 & n17220 ) ;
  assign n17222 = ~n8964 & n12469 ;
  assign n17223 = n17222 ^ n8931 ^ 1'b0 ;
  assign n17224 = n7902 ^ n4740 ^ 1'b0 ;
  assign n17225 = n9134 ^ n2125 ^ n1543 ;
  assign n17226 = n17225 ^ n7143 ^ n3073 ;
  assign n17227 = n324 | n17226 ;
  assign n17228 = n17224 & ~n17227 ;
  assign n17229 = n17228 ^ n13948 ^ 1'b0 ;
  assign n17230 = n17223 | n17229 ;
  assign n17231 = n4239 & n7472 ;
  assign n17232 = n17231 ^ n14290 ^ 1'b0 ;
  assign n17233 = n17232 ^ n14267 ^ 1'b0 ;
  assign n17234 = n12447 & n17233 ;
  assign n17236 = n5235 ^ n1246 ^ 1'b0 ;
  assign n17237 = n4294 & n17236 ;
  assign n17235 = n4904 | n14184 ;
  assign n17238 = n17237 ^ n17235 ^ 1'b0 ;
  assign n17239 = n4811 ^ n4156 ^ 1'b0 ;
  assign n17240 = ( ~n5839 & n6281 ) | ( ~n5839 & n7826 ) | ( n6281 & n7826 ) ;
  assign n17241 = ( n336 & ~n17239 ) | ( n336 & n17240 ) | ( ~n17239 & n17240 ) ;
  assign n17245 = n6191 ^ n3395 ^ 1'b0 ;
  assign n17246 = ~n1964 & n17245 ;
  assign n17247 = n10688 | n17246 ;
  assign n17248 = x151 | n17247 ;
  assign n17242 = n2458 & n11165 ;
  assign n17243 = n17242 ^ n7762 ^ n4749 ;
  assign n17244 = n14715 & n17243 ;
  assign n17249 = n17248 ^ n17244 ^ n6662 ;
  assign n17250 = n17249 ^ n13335 ^ n2758 ;
  assign n17251 = n15228 ^ n4110 ^ 1'b0 ;
  assign n17252 = n4066 & n17251 ;
  assign n17253 = ~n3896 & n17252 ;
  assign n17254 = n17253 ^ n5388 ^ 1'b0 ;
  assign n17257 = n14402 ^ n10840 ^ n2635 ;
  assign n17255 = n3845 ^ n1307 ^ n1294 ;
  assign n17256 = ( ~n7733 & n11318 ) | ( ~n7733 & n17255 ) | ( n11318 & n17255 ) ;
  assign n17258 = n17257 ^ n17256 ^ n11563 ;
  assign n17259 = n6174 ^ n4040 ^ n1090 ;
  assign n17260 = ~n2575 & n17259 ;
  assign n17261 = n7688 & ~n11955 ;
  assign n17262 = n10370 & n10961 ;
  assign n17263 = n17262 ^ n8374 ^ 1'b0 ;
  assign n17264 = n17145 ^ n7595 ^ 1'b0 ;
  assign n17265 = n13354 & ~n17264 ;
  assign n17266 = n17265 ^ n11801 ^ 1'b0 ;
  assign n17267 = n12171 ^ n11376 ^ n2145 ;
  assign n17268 = n11476 ^ n3488 ^ n881 ;
  assign n17269 = ~n11781 & n17268 ;
  assign n17274 = n9034 ^ n4819 ^ 1'b0 ;
  assign n17275 = n15473 & ~n17274 ;
  assign n17270 = n15926 ^ n1578 ^ n578 ;
  assign n17271 = ( n2592 & ~n11727 ) | ( n2592 & n16499 ) | ( ~n11727 & n16499 ) ;
  assign n17272 = n13760 & ~n17271 ;
  assign n17273 = ( n10389 & n17270 ) | ( n10389 & n17272 ) | ( n17270 & n17272 ) ;
  assign n17276 = n17275 ^ n17273 ^ n6228 ;
  assign n17277 = x52 & ~n3482 ;
  assign n17278 = ~n3924 & n17277 ;
  assign n17279 = n7230 ^ n1308 ^ 1'b0 ;
  assign n17281 = x107 & n1681 ;
  assign n17282 = n17281 ^ n1218 ^ 1'b0 ;
  assign n17283 = n15543 | n17282 ;
  assign n17280 = n13488 | n15019 ;
  assign n17284 = n17283 ^ n17280 ^ 1'b0 ;
  assign n17290 = n5455 | n8662 ;
  assign n17288 = ~n1674 & n10645 ;
  assign n17289 = n1701 & n17288 ;
  assign n17285 = n5295 & ~n11789 ;
  assign n17286 = n17285 ^ n2362 ^ 1'b0 ;
  assign n17287 = n17286 ^ n6622 ^ 1'b0 ;
  assign n17291 = n17290 ^ n17289 ^ n17287 ;
  assign n17294 = n2423 & ~n2760 ;
  assign n17292 = n7688 & ~n10377 ;
  assign n17293 = n8660 & n17292 ;
  assign n17295 = n17294 ^ n17293 ^ n15594 ;
  assign n17296 = n6473 & n8647 ;
  assign n17297 = n7112 ^ n2397 ^ 1'b0 ;
  assign n17298 = n17297 ^ n7013 ^ 1'b0 ;
  assign n17299 = n6071 ^ n4690 ^ 1'b0 ;
  assign n17300 = n3906 | n17299 ;
  assign n17301 = n17300 ^ n9519 ^ n4045 ;
  assign n17302 = n8295 ^ n1969 ^ 1'b0 ;
  assign n17303 = n16927 | n17302 ;
  assign n17306 = n14212 ^ n7685 ^ 1'b0 ;
  assign n17304 = n1370 & n3858 ;
  assign n17305 = n17304 ^ n9987 ^ 1'b0 ;
  assign n17307 = n17306 ^ n17305 ^ 1'b0 ;
  assign n17311 = n9203 & n12245 ;
  assign n17312 = n17311 ^ n12359 ^ 1'b0 ;
  assign n17313 = n5439 ^ n1742 ^ 1'b0 ;
  assign n17314 = n7805 & ~n17313 ;
  assign n17315 = n9646 & n17314 ;
  assign n17316 = n4328 & n5126 ;
  assign n17317 = ( n17312 & n17315 ) | ( n17312 & ~n17316 ) | ( n17315 & ~n17316 ) ;
  assign n17308 = ( n1325 & n8660 ) | ( n1325 & n10017 ) | ( n8660 & n10017 ) ;
  assign n17309 = n17308 ^ n1284 ^ 1'b0 ;
  assign n17310 = ~n6721 & n17309 ;
  assign n17318 = n17317 ^ n17310 ^ n8869 ;
  assign n17319 = n15231 ^ n14298 ^ n7991 ;
  assign n17321 = n4725 ^ n2559 ^ 1'b0 ;
  assign n17320 = n12369 ^ n6241 ^ n6035 ;
  assign n17322 = n17321 ^ n17320 ^ 1'b0 ;
  assign n17330 = n5137 ^ n1311 ^ n665 ;
  assign n17323 = n7973 | n12151 ;
  assign n17324 = n7752 ^ n5259 ^ 1'b0 ;
  assign n17325 = n3004 & n17324 ;
  assign n17326 = n3868 & n9019 ;
  assign n17327 = n17326 ^ n7070 ^ 1'b0 ;
  assign n17328 = n17325 & n17327 ;
  assign n17329 = n17323 & n17328 ;
  assign n17331 = n17330 ^ n17329 ^ 1'b0 ;
  assign n17332 = n17322 & ~n17331 ;
  assign n17333 = ~n8560 & n17332 ;
  assign n17334 = n17333 ^ n2815 ^ 1'b0 ;
  assign n17340 = ~n2333 & n13141 ;
  assign n17341 = n17340 ^ n16272 ^ 1'b0 ;
  assign n17342 = ~n13561 & n17341 ;
  assign n17335 = ~n8528 & n10004 ;
  assign n17336 = n5324 & n17335 ;
  assign n17337 = ~n14600 & n17336 ;
  assign n17338 = n17337 ^ x60 ^ 1'b0 ;
  assign n17339 = n10252 | n17338 ;
  assign n17343 = n17342 ^ n17339 ^ 1'b0 ;
  assign n17344 = n9660 & ~n17343 ;
  assign n17345 = n7613 ^ n4501 ^ n3331 ;
  assign n17346 = n14175 ^ n3823 ^ 1'b0 ;
  assign n17347 = n2512 & ~n17346 ;
  assign n17348 = n6739 & n17347 ;
  assign n17349 = ~n17345 & n17348 ;
  assign n17350 = n13122 ^ n5444 ^ n4639 ;
  assign n17351 = n17350 ^ n10325 ^ n5381 ;
  assign n17352 = n17351 ^ n9201 ^ n3527 ;
  assign n17353 = n8662 | n17352 ;
  assign n17354 = ( ~n4158 & n14769 ) | ( ~n4158 & n16177 ) | ( n14769 & n16177 ) ;
  assign n17355 = n9779 ^ n8365 ^ n3214 ;
  assign n17356 = n14691 & ~n17355 ;
  assign n17357 = n17356 ^ n14981 ^ 1'b0 ;
  assign n17358 = n5460 ^ n1558 ^ 1'b0 ;
  assign n17359 = n17358 ^ n4833 ^ n4553 ;
  assign n17360 = n17359 ^ n7403 ^ 1'b0 ;
  assign n17361 = x140 & n17360 ;
  assign n17362 = n8618 ^ n2094 ^ 1'b0 ;
  assign n17363 = n2380 & n17362 ;
  assign n17364 = ~n477 & n17363 ;
  assign n17365 = ~n13356 & n17364 ;
  assign n17366 = ~n893 & n4595 ;
  assign n17367 = ~n17365 & n17366 ;
  assign n17368 = ~x108 & n11627 ;
  assign n17369 = n4080 ^ n3035 ^ 1'b0 ;
  assign n17370 = n7830 | n17369 ;
  assign n17371 = n17370 ^ n7090 ^ 1'b0 ;
  assign n17372 = n16329 ^ n7890 ^ n3523 ;
  assign n17373 = n4734 & n6743 ;
  assign n17374 = n17373 ^ n3647 ^ 1'b0 ;
  assign n17375 = n17374 ^ x218 ^ 1'b0 ;
  assign n17376 = ( n14802 & n16124 ) | ( n14802 & ~n17375 ) | ( n16124 & ~n17375 ) ;
  assign n17377 = n17376 ^ n9137 ^ 1'b0 ;
  assign n17378 = n4691 & ~n9843 ;
  assign n17379 = ( n1839 & n14787 ) | ( n1839 & n17378 ) | ( n14787 & n17378 ) ;
  assign n17380 = ( n2918 & n3601 ) | ( n2918 & ~n17379 ) | ( n3601 & ~n17379 ) ;
  assign n17381 = n17380 ^ n6310 ^ n2124 ;
  assign n17382 = n17381 ^ n2747 ^ 1'b0 ;
  assign n17383 = ( n1104 & n2841 ) | ( n1104 & ~n5155 ) | ( n2841 & ~n5155 ) ;
  assign n17384 = n3639 & n17383 ;
  assign n17385 = n2192 | n17384 ;
  assign n17386 = n17385 ^ n3526 ^ n3004 ;
  assign n17387 = n9361 ^ n8070 ^ n4762 ;
  assign n17388 = n17387 ^ n13295 ^ 1'b0 ;
  assign n17389 = n17386 | n17388 ;
  assign n17399 = n17286 ^ n7260 ^ 1'b0 ;
  assign n17396 = ( n2250 & n3830 ) | ( n2250 & ~n12342 ) | ( n3830 & ~n12342 ) ;
  assign n17397 = n17396 ^ n14411 ^ n1437 ;
  assign n17390 = n11037 ^ n469 ^ 1'b0 ;
  assign n17391 = ~n4995 & n17390 ;
  assign n17392 = n3832 & n17391 ;
  assign n17393 = n17392 ^ n5125 ^ 1'b0 ;
  assign n17394 = n15152 | n17393 ;
  assign n17395 = n7841 & ~n17394 ;
  assign n17398 = n17397 ^ n17395 ^ 1'b0 ;
  assign n17400 = n17399 ^ n17398 ^ n5160 ;
  assign n17401 = ~n7447 & n17355 ;
  assign n17402 = n3340 | n4432 ;
  assign n17403 = n6699 | n17402 ;
  assign n17404 = n17403 ^ n2795 ^ 1'b0 ;
  assign n17405 = n11873 | n17404 ;
  assign n17406 = n17405 ^ n3585 ^ 1'b0 ;
  assign n17407 = ( n1784 & ~n2262 ) | ( n1784 & n9124 ) | ( ~n2262 & n9124 ) ;
  assign n17411 = n1819 ^ x209 ^ 1'b0 ;
  assign n17412 = ( n8452 & n15730 ) | ( n8452 & n17411 ) | ( n15730 & n17411 ) ;
  assign n17409 = x12 & n5839 ;
  assign n17410 = n17409 ^ n5062 ^ 1'b0 ;
  assign n17408 = n11504 ^ n4789 ^ n1508 ;
  assign n17413 = n17412 ^ n17410 ^ n17408 ;
  assign n17414 = ( n3026 & ~n17407 ) | ( n3026 & n17413 ) | ( ~n17407 & n17413 ) ;
  assign n17415 = n17414 ^ n2769 ^ 1'b0 ;
  assign n17416 = n7589 | n11151 ;
  assign n17417 = n6560 & ~n17416 ;
  assign n17418 = n10907 ^ n8706 ^ 1'b0 ;
  assign n17419 = n2479 & ~n17418 ;
  assign n17420 = n17419 ^ n12110 ^ n12045 ;
  assign n17421 = n5789 ^ n4790 ^ 1'b0 ;
  assign n17422 = n17420 & ~n17421 ;
  assign n17423 = ( n1964 & ~n5053 ) | ( n1964 & n7752 ) | ( ~n5053 & n7752 ) ;
  assign n17424 = n2338 & ~n17423 ;
  assign n17425 = n7318 ^ n2388 ^ 1'b0 ;
  assign n17426 = n2547 & n8317 ;
  assign n17427 = n10655 & n17426 ;
  assign n17428 = n17427 ^ n6381 ^ 1'b0 ;
  assign n17429 = n17428 ^ n14956 ^ n7040 ;
  assign n17430 = n17429 ^ n16507 ^ n10819 ;
  assign n17431 = n3313 & n6874 ;
  assign n17432 = ( n2547 & ~n12143 ) | ( n2547 & n17431 ) | ( ~n12143 & n17431 ) ;
  assign n17434 = n13857 ^ n6899 ^ n4813 ;
  assign n17433 = n14148 ^ x21 ^ 1'b0 ;
  assign n17435 = n17434 ^ n17433 ^ 1'b0 ;
  assign n17436 = n13305 & ~n17435 ;
  assign n17437 = n9554 | n10699 ;
  assign n17438 = n1485 & ~n17437 ;
  assign n17439 = n11384 & ~n14524 ;
  assign n17440 = ( n7630 & ~n12746 ) | ( n7630 & n13187 ) | ( ~n12746 & n13187 ) ;
  assign n17442 = n1522 & n8165 ;
  assign n17441 = n1766 ^ x27 ^ 1'b0 ;
  assign n17443 = n17442 ^ n17441 ^ 1'b0 ;
  assign n17444 = n14259 | n17443 ;
  assign n17446 = n4717 ^ n3906 ^ n1352 ;
  assign n17445 = ( ~n2308 & n3587 ) | ( ~n2308 & n15594 ) | ( n3587 & n15594 ) ;
  assign n17447 = n17446 ^ n17445 ^ n3003 ;
  assign n17448 = n8905 ^ n6856 ^ 1'b0 ;
  assign n17449 = ~n9987 & n17448 ;
  assign n17450 = n17449 ^ x151 ^ 1'b0 ;
  assign n17451 = ~n7143 & n7742 ;
  assign n17452 = n16446 & n17451 ;
  assign n17453 = ( ~n3368 & n9974 ) | ( ~n3368 & n17452 ) | ( n9974 & n17452 ) ;
  assign n17454 = n3740 & n7014 ;
  assign n17455 = n17454 ^ n2567 ^ 1'b0 ;
  assign n17456 = n9991 ^ n3917 ^ 1'b0 ;
  assign n17457 = n9938 ^ n6685 ^ 1'b0 ;
  assign n17458 = n14832 ^ n10842 ^ n6527 ;
  assign n17460 = n8366 ^ n5240 ^ 1'b0 ;
  assign n17461 = ~n7568 & n17460 ;
  assign n17459 = ~n7127 & n17392 ;
  assign n17462 = n17461 ^ n17459 ^ 1'b0 ;
  assign n17463 = ( x132 & n426 ) | ( x132 & ~n3770 ) | ( n426 & ~n3770 ) ;
  assign n17467 = n11536 ^ n429 ^ 1'b0 ;
  assign n17465 = n13023 ^ n8314 ^ n2510 ;
  assign n17464 = n6792 | n10332 ;
  assign n17466 = n17465 ^ n17464 ^ 1'b0 ;
  assign n17468 = n17467 ^ n17466 ^ 1'b0 ;
  assign n17469 = n1680 ^ n1292 ^ 1'b0 ;
  assign n17470 = ~n420 & n17469 ;
  assign n17471 = n17467 ^ n8315 ^ 1'b0 ;
  assign n17472 = n17470 & ~n17471 ;
  assign n17473 = n6621 & ~n6735 ;
  assign n17474 = ~n17472 & n17473 ;
  assign n17475 = n3683 ^ n2486 ^ n919 ;
  assign n17476 = n9570 ^ n8700 ^ 1'b0 ;
  assign n17477 = ( n3632 & n5443 ) | ( n3632 & n17476 ) | ( n5443 & n17476 ) ;
  assign n17478 = n17475 & n17477 ;
  assign n17479 = n17478 ^ n8504 ^ 1'b0 ;
  assign n17480 = n13039 ^ n6204 ^ 1'b0 ;
  assign n17481 = n2477 | n17480 ;
  assign n17482 = n16775 & ~n17481 ;
  assign n17483 = ~n17479 & n17482 ;
  assign n17484 = ( ~n2002 & n10282 ) | ( ~n2002 & n11156 ) | ( n10282 & n11156 ) ;
  assign n17485 = n5042 ^ n1026 ^ 1'b0 ;
  assign n17486 = n17485 ^ n4840 ^ 1'b0 ;
  assign n17487 = n4386 ^ n2455 ^ 1'b0 ;
  assign n17488 = n16095 | n17487 ;
  assign n17489 = n4917 ^ n3146 ^ n448 ;
  assign n17490 = ~n3945 & n17489 ;
  assign n17491 = n14524 ^ n6653 ^ n2927 ;
  assign n17492 = n5167 & n7453 ;
  assign n17493 = n4700 ^ n870 ^ n868 ;
  assign n17494 = n17493 ^ n4977 ^ 1'b0 ;
  assign n17495 = ~n284 & n17494 ;
  assign n17496 = x251 & ~n3849 ;
  assign n17497 = n17496 ^ x72 ^ 1'b0 ;
  assign n17498 = n7748 & ~n17497 ;
  assign n17499 = n17498 ^ n2692 ^ n1778 ;
  assign n17500 = n11722 ^ n4946 ^ n3280 ;
  assign n17501 = ( n1943 & ~n17499 ) | ( n1943 & n17500 ) | ( ~n17499 & n17500 ) ;
  assign n17504 = n2978 & ~n11564 ;
  assign n17505 = n8366 & n17504 ;
  assign n17506 = n17505 ^ n10531 ^ 1'b0 ;
  assign n17507 = n14578 & ~n17506 ;
  assign n17502 = n12906 & ~n14620 ;
  assign n17503 = n10873 & ~n17502 ;
  assign n17508 = n17507 ^ n17503 ^ 1'b0 ;
  assign n17509 = n15425 ^ n8235 ^ 1'b0 ;
  assign n17510 = n4154 & ~n15390 ;
  assign n17511 = n14117 ^ n10156 ^ 1'b0 ;
  assign n17512 = ~n16234 & n17511 ;
  assign n17513 = n17512 ^ n7383 ^ 1'b0 ;
  assign n17517 = n8108 | n13418 ;
  assign n17518 = n17517 ^ n1771 ^ 1'b0 ;
  assign n17519 = n583 | n17518 ;
  assign n17514 = n15875 ^ n11484 ^ 1'b0 ;
  assign n17515 = n5440 | n17514 ;
  assign n17516 = n5646 | n17515 ;
  assign n17520 = n17519 ^ n17516 ^ n9408 ;
  assign n17521 = ~n1709 & n4756 ;
  assign n17522 = ~n335 & n17521 ;
  assign n17523 = n17522 ^ n1125 ^ 1'b0 ;
  assign n17524 = ~n8369 & n17523 ;
  assign n17525 = n17524 ^ n9960 ^ 1'b0 ;
  assign n17526 = n8120 ^ n327 ^ 1'b0 ;
  assign n17527 = n17525 | n17526 ;
  assign n17528 = n17527 ^ n14111 ^ 1'b0 ;
  assign n17529 = n16701 ^ n7673 ^ n3385 ;
  assign n17530 = n13939 ^ n10553 ^ 1'b0 ;
  assign n17531 = n17529 & n17530 ;
  assign n17532 = ~n4037 & n6615 ;
  assign n17533 = n5025 & ~n16195 ;
  assign n17534 = n13672 ^ n2569 ^ n1247 ;
  assign n17535 = n5009 | n17534 ;
  assign n17536 = n17535 ^ n7217 ^ 1'b0 ;
  assign n17537 = n3530 & ~n12967 ;
  assign n17538 = ~n9106 & n9903 ;
  assign n17544 = n12462 ^ n5393 ^ 1'b0 ;
  assign n17539 = n11899 ^ n7301 ^ n4552 ;
  assign n17540 = ~n16037 & n17539 ;
  assign n17541 = n14101 & n17540 ;
  assign n17542 = n6406 ^ n4453 ^ 1'b0 ;
  assign n17543 = ~n17541 & n17542 ;
  assign n17545 = n17544 ^ n17543 ^ 1'b0 ;
  assign n17546 = n17538 | n17545 ;
  assign n17547 = n3980 & n16508 ;
  assign n17548 = ~n665 & n17547 ;
  assign n17549 = ( n5694 & n8375 ) | ( n5694 & n17548 ) | ( n8375 & n17548 ) ;
  assign n17550 = ~n5757 & n7238 ;
  assign n17551 = n14686 ^ n614 ^ 1'b0 ;
  assign n17552 = n4378 ^ n3809 ^ 1'b0 ;
  assign n17553 = ~n13368 & n17552 ;
  assign n17554 = n17553 ^ n11403 ^ n5529 ;
  assign n17555 = n12232 & ~n17554 ;
  assign n17556 = ~n2707 & n6353 ;
  assign n17557 = ( ~n14064 & n15593 ) | ( ~n14064 & n17556 ) | ( n15593 & n17556 ) ;
  assign n17559 = n9781 ^ n1838 ^ 1'b0 ;
  assign n17558 = n2828 & ~n9377 ;
  assign n17560 = n17559 ^ n17558 ^ 1'b0 ;
  assign n17561 = ( ~n4439 & n5336 ) | ( ~n4439 & n17560 ) | ( n5336 & n17560 ) ;
  assign n17562 = ( n8802 & n9061 ) | ( n8802 & n17561 ) | ( n9061 & n17561 ) ;
  assign n17563 = n400 | n1183 ;
  assign n17564 = ( ~n4686 & n7051 ) | ( ~n4686 & n17563 ) | ( n7051 & n17563 ) ;
  assign n17565 = ( ~n503 & n1843 ) | ( ~n503 & n5059 ) | ( n1843 & n5059 ) ;
  assign n17566 = n17565 ^ n11021 ^ n1582 ;
  assign n17567 = n17566 ^ n10014 ^ 1'b0 ;
  assign n17568 = n3319 & n17567 ;
  assign n17569 = n11968 | n17568 ;
  assign n17573 = n10898 ^ n10078 ^ 1'b0 ;
  assign n17570 = n6856 & ~n8333 ;
  assign n17571 = n17570 ^ n15212 ^ 1'b0 ;
  assign n17572 = n17571 ^ n1189 ^ 1'b0 ;
  assign n17574 = n17573 ^ n17572 ^ 1'b0 ;
  assign n17575 = n783 | n7235 ;
  assign n17576 = n13785 ^ n12483 ^ 1'b0 ;
  assign n17577 = n2033 & ~n17576 ;
  assign n17578 = ~n4908 & n17577 ;
  assign n17579 = n6804 | n16599 ;
  assign n17580 = n7653 & ~n15058 ;
  assign n17581 = n13000 ^ n6750 ^ 1'b0 ;
  assign n17589 = ~n3424 & n15252 ;
  assign n17587 = n2427 ^ x85 ^ 1'b0 ;
  assign n17588 = ( n4167 & ~n7300 ) | ( n4167 & n17587 ) | ( ~n7300 & n17587 ) ;
  assign n17582 = n875 & ~n1272 ;
  assign n17583 = n17582 ^ n6752 ^ 1'b0 ;
  assign n17584 = n1007 & n17583 ;
  assign n17585 = ~n15335 & n17584 ;
  assign n17586 = n17585 ^ n13388 ^ n6397 ;
  assign n17590 = n17589 ^ n17588 ^ n17586 ;
  assign n17591 = n5300 & ~n15704 ;
  assign n17592 = n17591 ^ n3225 ^ 1'b0 ;
  assign n17593 = n17592 ^ n7577 ^ n6372 ;
  assign n17594 = n16121 ^ n9522 ^ 1'b0 ;
  assign n17595 = n17593 & n17594 ;
  assign n17596 = n10170 ^ n7463 ^ 1'b0 ;
  assign n17597 = ( n9260 & n11348 ) | ( n9260 & ~n17596 ) | ( n11348 & ~n17596 ) ;
  assign n17598 = n1372 & ~n5984 ;
  assign n17599 = ~n13469 & n17598 ;
  assign n17600 = n4308 | n5157 ;
  assign n17601 = n14857 ^ n12794 ^ n8409 ;
  assign n17602 = ( ~n6960 & n17430 ) | ( ~n6960 & n17601 ) | ( n17430 & n17601 ) ;
  assign n17603 = n6205 ^ n4142 ^ 1'b0 ;
  assign n17604 = ~n13950 & n17603 ;
  assign n17605 = n11673 ^ n7058 ^ 1'b0 ;
  assign n17606 = n11384 & ~n17605 ;
  assign n17607 = ( n3126 & ~n13675 ) | ( n3126 & n17606 ) | ( ~n13675 & n17606 ) ;
  assign n17608 = n16775 ^ n9405 ^ 1'b0 ;
  assign n17609 = ~n16509 & n17608 ;
  assign n17610 = n17609 ^ n13544 ^ 1'b0 ;
  assign n17611 = n704 & n17610 ;
  assign n17612 = ~n7920 & n17611 ;
  assign n17613 = ~n12137 & n17612 ;
  assign n17625 = n9551 ^ n436 ^ 1'b0 ;
  assign n17626 = n8372 | n17625 ;
  assign n17614 = n6201 & ~n7461 ;
  assign n17615 = n17614 ^ n9795 ^ 1'b0 ;
  assign n17618 = n7534 ^ n7429 ^ n428 ;
  assign n17616 = n438 & ~n1283 ;
  assign n17617 = n17616 ^ n2399 ^ 1'b0 ;
  assign n17619 = n17618 ^ n17617 ^ 1'b0 ;
  assign n17620 = n8514 & n17619 ;
  assign n17621 = n17620 ^ n2169 ^ 1'b0 ;
  assign n17622 = ~n8289 & n17621 ;
  assign n17623 = n841 & n17622 ;
  assign n17624 = ( n8423 & n17615 ) | ( n8423 & ~n17623 ) | ( n17615 & ~n17623 ) ;
  assign n17627 = n17626 ^ n17624 ^ n1173 ;
  assign n17630 = n2950 & n17294 ;
  assign n17631 = n17630 ^ n6887 ^ 1'b0 ;
  assign n17632 = ~n7748 & n17631 ;
  assign n17628 = n9789 ^ n6995 ^ n3970 ;
  assign n17629 = n17628 ^ n11252 ^ 1'b0 ;
  assign n17633 = n17632 ^ n17629 ^ n16946 ;
  assign n17634 = n12027 ^ n11291 ^ 1'b0 ;
  assign n17635 = ~n5132 & n17634 ;
  assign n17636 = n17635 ^ n15200 ^ 1'b0 ;
  assign n17637 = n16703 ^ n7366 ^ 1'b0 ;
  assign n17638 = n17636 | n17637 ;
  assign n17639 = n10875 ^ n3173 ^ n408 ;
  assign n17640 = n17639 ^ n11808 ^ n5151 ;
  assign n17641 = ( n14555 & n15728 ) | ( n14555 & ~n17640 ) | ( n15728 & ~n17640 ) ;
  assign n17642 = n9311 ^ x89 ^ 1'b0 ;
  assign n17643 = n1346 | n17642 ;
  assign n17644 = n4976 | n17643 ;
  assign n17645 = n2763 & ~n17644 ;
  assign n17646 = n15519 ^ n12811 ^ 1'b0 ;
  assign n17647 = ( ~n2530 & n4916 ) | ( ~n2530 & n7664 ) | ( n4916 & n7664 ) ;
  assign n17648 = n3621 & n17647 ;
  assign n17649 = n5889 & n7734 ;
  assign n17654 = n8545 & ~n11212 ;
  assign n17655 = n1894 & n17654 ;
  assign n17653 = ~n11784 & n14374 ;
  assign n17650 = n3159 | n3840 ;
  assign n17651 = n17650 ^ n6495 ^ 1'b0 ;
  assign n17652 = n17651 ^ n12168 ^ n2859 ;
  assign n17656 = n17655 ^ n17653 ^ n17652 ;
  assign n17659 = n6387 | n14600 ;
  assign n17657 = ~n9009 & n16955 ;
  assign n17658 = ~n12783 & n17657 ;
  assign n17660 = n17659 ^ n17658 ^ 1'b0 ;
  assign n17661 = ~n12363 & n14336 ;
  assign n17662 = n17661 ^ n13660 ^ 1'b0 ;
  assign n17663 = n3269 & ~n4968 ;
  assign n17664 = n17663 ^ n8546 ^ 1'b0 ;
  assign n17665 = n17664 ^ n6521 ^ 1'b0 ;
  assign n17666 = n348 & n17665 ;
  assign n17667 = n12477 ^ n11136 ^ n4911 ;
  assign n17668 = n17667 ^ n10696 ^ 1'b0 ;
  assign n17673 = n16196 ^ n2686 ^ 1'b0 ;
  assign n17674 = n14467 ^ n13544 ^ 1'b0 ;
  assign n17675 = n11278 | n17674 ;
  assign n17676 = n17673 & ~n17675 ;
  assign n17669 = ( n1451 & ~n4958 ) | ( n1451 & n7576 ) | ( ~n4958 & n7576 ) ;
  assign n17670 = n13204 ^ n5650 ^ 1'b0 ;
  assign n17671 = n13127 & ~n17670 ;
  assign n17672 = n17669 | n17671 ;
  assign n17677 = n17676 ^ n17672 ^ n4315 ;
  assign n17678 = n11929 ^ n5843 ^ 1'b0 ;
  assign n17679 = ( ~n989 & n7903 ) | ( ~n989 & n17678 ) | ( n7903 & n17678 ) ;
  assign n17680 = n17679 ^ n8935 ^ 1'b0 ;
  assign n17681 = n321 & ~n17680 ;
  assign n17682 = n16477 ^ n6637 ^ n1591 ;
  assign n17683 = ~n3771 & n17682 ;
  assign n17684 = n12454 ^ n10214 ^ 1'b0 ;
  assign n17685 = n8336 & n17684 ;
  assign n17686 = ~n17289 & n17685 ;
  assign n17687 = n8367 & n17686 ;
  assign n17688 = n13025 ^ n4588 ^ 1'b0 ;
  assign n17689 = ~n17687 & n17688 ;
  assign n17690 = ( n1350 & n7787 ) | ( n1350 & ~n13319 ) | ( n7787 & ~n13319 ) ;
  assign n17691 = n17690 ^ n11612 ^ 1'b0 ;
  assign n17692 = n6368 | n17691 ;
  assign n17693 = ( ~n280 & n4989 ) | ( ~n280 & n16775 ) | ( n4989 & n16775 ) ;
  assign n17694 = n16238 ^ n6643 ^ 1'b0 ;
  assign n17695 = n2744 & ~n17694 ;
  assign n17696 = n17695 ^ n15181 ^ n1971 ;
  assign n17697 = ~n10394 & n12369 ;
  assign n17698 = n17697 ^ n4472 ^ n2414 ;
  assign n17699 = ~n6705 & n16490 ;
  assign n17700 = n17699 ^ n11246 ^ 1'b0 ;
  assign n17701 = n17700 ^ n8503 ^ n5259 ;
  assign n17702 = ~n1429 & n12081 ;
  assign n17703 = n17702 ^ n16112 ^ 1'b0 ;
  assign n17704 = n17703 ^ n12393 ^ 1'b0 ;
  assign n17705 = n3222 & n17051 ;
  assign n17706 = n6073 & n17705 ;
  assign n17709 = n4698 & n11689 ;
  assign n17710 = n6921 & n17709 ;
  assign n17707 = ( n853 & n1994 ) | ( n853 & n7641 ) | ( n1994 & n7641 ) ;
  assign n17708 = ( n4064 & n9175 ) | ( n4064 & ~n17707 ) | ( n9175 & ~n17707 ) ;
  assign n17711 = n17710 ^ n17708 ^ n8393 ;
  assign n17721 = n10288 ^ n5133 ^ 1'b0 ;
  assign n17717 = n9827 ^ n1589 ^ 1'b0 ;
  assign n17718 = ~n14192 & n17717 ;
  assign n17716 = ~n3433 & n6396 ;
  assign n17719 = n17718 ^ n17716 ^ 1'b0 ;
  assign n17712 = n3719 & ~n9463 ;
  assign n17713 = n8196 & n17712 ;
  assign n17714 = n12547 ^ n11261 ^ 1'b0 ;
  assign n17715 = ~n17713 & n17714 ;
  assign n17720 = n17719 ^ n17715 ^ n12560 ;
  assign n17722 = n17721 ^ n17720 ^ 1'b0 ;
  assign n17723 = n11916 ^ n4363 ^ n2782 ;
  assign n17724 = x242 & ~n17723 ;
  assign n17725 = n17724 ^ n3803 ^ 1'b0 ;
  assign n17726 = ( n6536 & n13108 ) | ( n6536 & n17725 ) | ( n13108 & n17725 ) ;
  assign n17727 = n17726 ^ n14318 ^ 1'b0 ;
  assign n17728 = ( n3075 & ~n5242 ) | ( n3075 & n17543 ) | ( ~n5242 & n17543 ) ;
  assign n17733 = n4826 ^ n3619 ^ n1392 ;
  assign n17734 = n17733 ^ n3508 ^ n1284 ;
  assign n17729 = ( ~n730 & n3721 ) | ( ~n730 & n13497 ) | ( n3721 & n13497 ) ;
  assign n17730 = x37 & n17729 ;
  assign n17731 = n17730 ^ n5612 ^ 1'b0 ;
  assign n17732 = ( n4108 & n7355 ) | ( n4108 & n17731 ) | ( n7355 & n17731 ) ;
  assign n17735 = n17734 ^ n17732 ^ 1'b0 ;
  assign n17736 = n11825 | n11832 ;
  assign n17737 = n11116 | n17736 ;
  assign n17738 = n11938 ^ n7371 ^ 1'b0 ;
  assign n17739 = x45 & n17738 ;
  assign n17740 = n17739 ^ n16491 ^ 1'b0 ;
  assign n17741 = n5608 & n17740 ;
  assign n17742 = n16145 ^ n8635 ^ 1'b0 ;
  assign n17743 = n3690 | n5990 ;
  assign n17744 = n17743 ^ n285 ^ 1'b0 ;
  assign n17745 = n16447 | n17744 ;
  assign n17746 = n17745 ^ n5559 ^ 1'b0 ;
  assign n17747 = n3786 & ~n11645 ;
  assign n17748 = n17747 ^ n4796 ^ 1'b0 ;
  assign n17750 = n3360 | n16191 ;
  assign n17751 = n17750 ^ n7121 ^ 1'b0 ;
  assign n17752 = n17751 ^ n1269 ^ 1'b0 ;
  assign n17753 = n10729 & ~n17752 ;
  assign n17749 = n9002 | n10679 ;
  assign n17754 = n17753 ^ n17749 ^ 1'b0 ;
  assign n17755 = ( n1294 & ~n9252 ) | ( n1294 & n17754 ) | ( ~n9252 & n17754 ) ;
  assign n17756 = n2541 | n9246 ;
  assign n17757 = n17756 ^ n3126 ^ 1'b0 ;
  assign n17758 = n14688 ^ n14382 ^ n3148 ;
  assign n17759 = n17758 ^ n3015 ^ 1'b0 ;
  assign n17760 = n3917 & n4240 ;
  assign n17761 = ~n5405 & n17760 ;
  assign n17762 = ( ~x103 & n14675 ) | ( ~x103 & n17761 ) | ( n14675 & n17761 ) ;
  assign n17763 = ( x32 & n3496 ) | ( x32 & n8537 ) | ( n3496 & n8537 ) ;
  assign n17764 = n17763 ^ n7000 ^ n4986 ;
  assign n17765 = n9087 ^ x107 ^ 1'b0 ;
  assign n17766 = n17764 | n17765 ;
  assign n17770 = n10552 ^ n7929 ^ 1'b0 ;
  assign n17771 = n4914 | n17770 ;
  assign n17767 = n6419 ^ n3115 ^ 1'b0 ;
  assign n17768 = n1504 & n17767 ;
  assign n17769 = ~n17733 & n17768 ;
  assign n17772 = n17771 ^ n17769 ^ 1'b0 ;
  assign n17773 = n16512 | n17772 ;
  assign n17774 = n2461 | n11134 ;
  assign n17775 = n17774 ^ n14843 ^ 1'b0 ;
  assign n17776 = n6708 & n14012 ;
  assign n17777 = ~n3771 & n17776 ;
  assign n17778 = n17775 & n17777 ;
  assign n17779 = n12146 ^ n4682 ^ 1'b0 ;
  assign n17780 = n17779 ^ n3616 ^ 1'b0 ;
  assign n17781 = n3985 ^ n3852 ^ 1'b0 ;
  assign n17782 = ~n3478 & n17781 ;
  assign n17783 = ~n14897 & n17782 ;
  assign n17784 = n9405 ^ n4056 ^ 1'b0 ;
  assign n17785 = ~n6241 & n17784 ;
  assign n17786 = n3711 ^ n3129 ^ n1108 ;
  assign n17787 = n17786 ^ n642 ^ n479 ;
  assign n17788 = ( ~n10597 & n11295 ) | ( ~n10597 & n17787 ) | ( n11295 & n17787 ) ;
  assign n17789 = ~n2960 & n17788 ;
  assign n17790 = n8868 & ~n17789 ;
  assign n17791 = ( n1051 & n11235 ) | ( n1051 & n12101 ) | ( n11235 & n12101 ) ;
  assign n17792 = n12071 ^ n3999 ^ 1'b0 ;
  assign n17793 = n14849 | n17792 ;
  assign n17794 = ~n8915 & n17793 ;
  assign n17795 = n3517 & ~n4146 ;
  assign n17796 = ~n12381 & n17795 ;
  assign n17797 = n7015 & n14636 ;
  assign n17800 = n13439 ^ n12914 ^ 1'b0 ;
  assign n17798 = n17327 ^ n4013 ^ 1'b0 ;
  assign n17799 = n16294 | n17798 ;
  assign n17801 = n17800 ^ n17799 ^ 1'b0 ;
  assign n17802 = n6451 ^ n2869 ^ n2825 ;
  assign n17805 = n5532 ^ n5116 ^ 1'b0 ;
  assign n17806 = n4803 & ~n17805 ;
  assign n17807 = ( ~n5447 & n10204 ) | ( ~n5447 & n17806 ) | ( n10204 & n17806 ) ;
  assign n17808 = n17807 ^ n15518 ^ n7787 ;
  assign n17803 = n14621 ^ n11270 ^ n6203 ;
  assign n17804 = n1199 | n17803 ;
  assign n17809 = n17808 ^ n17804 ^ 1'b0 ;
  assign n17810 = n5585 ^ n3702 ^ 1'b0 ;
  assign n17811 = n11782 ^ n8811 ^ 1'b0 ;
  assign n17812 = n17810 & ~n17811 ;
  assign n17813 = n17812 ^ n3521 ^ n861 ;
  assign n17814 = ~n907 & n12126 ;
  assign n17815 = n17814 ^ n9975 ^ 1'b0 ;
  assign n17816 = n17441 ^ n2860 ^ 1'b0 ;
  assign n17817 = ( ~n7289 & n17815 ) | ( ~n7289 & n17816 ) | ( n17815 & n17816 ) ;
  assign n17818 = n8477 ^ n8333 ^ 1'b0 ;
  assign n17819 = n17818 ^ n2745 ^ 1'b0 ;
  assign n17820 = ~n9779 & n14344 ;
  assign n17821 = ( n1593 & ~n7950 ) | ( n1593 & n17820 ) | ( ~n7950 & n17820 ) ;
  assign n17822 = n17821 ^ n16964 ^ n3285 ;
  assign n17823 = ( n998 & ~n3580 ) | ( n998 & n4933 ) | ( ~n3580 & n4933 ) ;
  assign n17824 = n17823 ^ n16132 ^ n3863 ;
  assign n17825 = n11398 & n17824 ;
  assign n17826 = n10958 ^ n8122 ^ n6658 ;
  assign n17827 = ( n1311 & n4935 ) | ( n1311 & n7782 ) | ( n4935 & n7782 ) ;
  assign n17828 = n17827 ^ n6168 ^ n2436 ;
  assign n17829 = n10514 ^ n7223 ^ 1'b0 ;
  assign n17830 = n17423 & n17829 ;
  assign n17831 = ~n8699 & n17830 ;
  assign n17832 = n17828 & n17831 ;
  assign n17833 = n12060 & n17516 ;
  assign n17834 = n3951 ^ n874 ^ 1'b0 ;
  assign n17835 = n5025 ^ n1045 ^ 1'b0 ;
  assign n17836 = n17834 | n17835 ;
  assign n17837 = n4287 ^ n3269 ^ n1372 ;
  assign n17838 = n17837 ^ n7950 ^ n6212 ;
  assign n17839 = n17836 | n17838 ;
  assign n17840 = n17839 ^ n4956 ^ 1'b0 ;
  assign n17841 = n8014 ^ n6382 ^ 1'b0 ;
  assign n17842 = n16981 ^ n2934 ^ 1'b0 ;
  assign n17843 = n6258 & n8005 ;
  assign n17844 = n17843 ^ n6481 ^ 1'b0 ;
  assign n17845 = n12207 & ~n17844 ;
  assign n17846 = n17845 ^ n8195 ^ 1'b0 ;
  assign n17847 = ( ~n3471 & n17842 ) | ( ~n3471 & n17846 ) | ( n17842 & n17846 ) ;
  assign n17848 = n1522 & ~n9989 ;
  assign n17865 = n4813 & ~n8614 ;
  assign n17866 = n2319 & n17865 ;
  assign n17849 = ~n7168 & n8878 ;
  assign n17850 = n17849 ^ n4445 ^ 1'b0 ;
  assign n17852 = n12541 ^ n5524 ^ n3368 ;
  assign n17851 = ( n1934 & n2388 ) | ( n1934 & ~n10028 ) | ( n2388 & ~n10028 ) ;
  assign n17853 = n17852 ^ n17851 ^ 1'b0 ;
  assign n17854 = n3074 & n17853 ;
  assign n17855 = n9611 ^ n9174 ^ 1'b0 ;
  assign n17856 = n17854 & n17855 ;
  assign n17857 = ~n7029 & n7414 ;
  assign n17858 = n2016 & n17857 ;
  assign n17859 = ( n2169 & n14515 ) | ( n2169 & n17858 ) | ( n14515 & n17858 ) ;
  assign n17860 = n17859 ^ n8977 ^ 1'b0 ;
  assign n17861 = n521 & ~n17860 ;
  assign n17862 = n8494 | n17861 ;
  assign n17863 = ( n17850 & ~n17856 ) | ( n17850 & n17862 ) | ( ~n17856 & n17862 ) ;
  assign n17864 = n2983 | n17863 ;
  assign n17867 = n17866 ^ n17864 ^ 1'b0 ;
  assign n17868 = ( n11862 & ~n17848 ) | ( n11862 & n17867 ) | ( ~n17848 & n17867 ) ;
  assign n17869 = n7538 ^ n6673 ^ 1'b0 ;
  assign n17870 = n10249 | n17869 ;
  assign n17871 = ~n8539 & n17870 ;
  assign n17872 = n6033 & ~n10710 ;
  assign n17873 = ( n5082 & n13814 ) | ( n5082 & ~n17872 ) | ( n13814 & ~n17872 ) ;
  assign n17874 = n14340 ^ n11722 ^ 1'b0 ;
  assign n17875 = n5263 ^ n3491 ^ n2450 ;
  assign n17876 = n17875 ^ n4723 ^ 1'b0 ;
  assign n17877 = n16348 ^ n3285 ^ 1'b0 ;
  assign n17878 = n17877 ^ n2400 ^ 1'b0 ;
  assign n17881 = ( n870 & n3599 ) | ( n870 & n4432 ) | ( n3599 & n4432 ) ;
  assign n17879 = ~n7734 & n9724 ;
  assign n17880 = n17879 ^ n13282 ^ 1'b0 ;
  assign n17882 = n17881 ^ n17880 ^ 1'b0 ;
  assign n17883 = n3995 & n17882 ;
  assign n17884 = ~n4055 & n17883 ;
  assign n17885 = n4662 ^ n1112 ^ 1'b0 ;
  assign n17886 = n15816 ^ n8768 ^ n3436 ;
  assign n17887 = n17886 ^ n6022 ^ n5117 ;
  assign n17888 = n13760 & ~n17887 ;
  assign n17895 = n7011 ^ n6398 ^ 1'b0 ;
  assign n17896 = n4659 & n17895 ;
  assign n17897 = ( n5506 & n7200 ) | ( n5506 & ~n17896 ) | ( n7200 & ~n17896 ) ;
  assign n17894 = n7574 | n13818 ;
  assign n17889 = n4081 & n9589 ;
  assign n17890 = n17889 ^ n10369 ^ 1'b0 ;
  assign n17891 = n11321 ^ n9607 ^ n7785 ;
  assign n17892 = ( n6240 & n17890 ) | ( n6240 & n17891 ) | ( n17890 & n17891 ) ;
  assign n17893 = n17892 ^ n10755 ^ n1785 ;
  assign n17898 = n17897 ^ n17894 ^ n17893 ;
  assign n17899 = n10057 ^ n8644 ^ 1'b0 ;
  assign n17900 = n10156 | n13155 ;
  assign n17901 = n17900 ^ n6160 ^ 1'b0 ;
  assign n17902 = n17901 ^ n10020 ^ n8977 ;
  assign n17903 = ( n1137 & ~n3872 ) | ( n1137 & n11519 ) | ( ~n3872 & n11519 ) ;
  assign n17904 = ( n457 & ~n1569 ) | ( n457 & n4281 ) | ( ~n1569 & n4281 ) ;
  assign n17905 = ~n17903 & n17904 ;
  assign n17906 = x244 & ~n5784 ;
  assign n17907 = n8125 & n17906 ;
  assign n17908 = n17907 ^ n10849 ^ 1'b0 ;
  assign n17909 = n11281 ^ n8306 ^ 1'b0 ;
  assign n17910 = n17908 | n17909 ;
  assign n17911 = n4790 ^ n1472 ^ 1'b0 ;
  assign n17912 = ~n3450 & n17911 ;
  assign n17913 = n17912 ^ n9049 ^ 1'b0 ;
  assign n17914 = n17910 | n17913 ;
  assign n17915 = n17914 ^ n4289 ^ 1'b0 ;
  assign n17916 = n7349 | n8614 ;
  assign n17917 = n17916 ^ x73 ^ 1'b0 ;
  assign n17918 = n4390 | n13251 ;
  assign n17919 = n17917 | n17918 ;
  assign n17920 = n17919 ^ n9480 ^ n4257 ;
  assign n17921 = n16072 ^ n6453 ^ n5385 ;
  assign n17922 = n17921 ^ n15080 ^ n5780 ;
  assign n17923 = n14379 ^ n4066 ^ 1'b0 ;
  assign n17924 = n1464 | n17923 ;
  assign n17925 = n17924 ^ n2232 ^ n2191 ;
  assign n17932 = n1311 & ~n4540 ;
  assign n17933 = n17932 ^ n6341 ^ n4596 ;
  assign n17934 = n4183 | n10430 ;
  assign n17935 = ( ~n8217 & n11185 ) | ( ~n8217 & n17934 ) | ( n11185 & n17934 ) ;
  assign n17936 = ( n11336 & ~n17933 ) | ( n11336 & n17935 ) | ( ~n17933 & n17935 ) ;
  assign n17926 = n12694 ^ n5386 ^ 1'b0 ;
  assign n17927 = n4840 & n17926 ;
  assign n17928 = ( n2666 & ~n3585 ) | ( n2666 & n6270 ) | ( ~n3585 & n6270 ) ;
  assign n17929 = ( n4440 & n11323 ) | ( n4440 & ~n17928 ) | ( n11323 & ~n17928 ) ;
  assign n17930 = n10872 & ~n17929 ;
  assign n17931 = ~n17927 & n17930 ;
  assign n17937 = n17936 ^ n17931 ^ n11801 ;
  assign n17938 = ( n556 & n1958 ) | ( n556 & ~n17937 ) | ( n1958 & ~n17937 ) ;
  assign n17939 = n7625 | n17048 ;
  assign n17940 = n17939 ^ n1236 ^ 1'b0 ;
  assign n17941 = n4758 & n10199 ;
  assign n17942 = n17941 ^ n10137 ^ 1'b0 ;
  assign n17943 = n11272 ^ n10474 ^ 1'b0 ;
  assign n17944 = ( n4501 & n12698 ) | ( n4501 & ~n17943 ) | ( n12698 & ~n17943 ) ;
  assign n17945 = n12532 ^ n11795 ^ 1'b0 ;
  assign n17946 = n8817 & n17945 ;
  assign n17947 = n17946 ^ n11250 ^ 1'b0 ;
  assign n17948 = ( n8253 & n10514 ) | ( n8253 & ~n12199 ) | ( n10514 & ~n12199 ) ;
  assign n17949 = n15977 & n17948 ;
  assign n17950 = n1542 & n17949 ;
  assign n17954 = n5602 ^ n3239 ^ n1868 ;
  assign n17955 = x9 & ~n17954 ;
  assign n17956 = n7759 & n17955 ;
  assign n17957 = n2201 & ~n17956 ;
  assign n17958 = n17957 ^ n4412 ^ 1'b0 ;
  assign n17951 = ~n3496 & n11546 ;
  assign n17952 = ~n12785 & n17951 ;
  assign n17953 = n17952 ^ n16004 ^ n14796 ;
  assign n17959 = n17958 ^ n17953 ^ n12767 ;
  assign n17960 = n14377 ^ n8184 ^ n1112 ;
  assign n17961 = n17960 ^ n11658 ^ n7236 ;
  assign n17962 = n5567 & ~n17961 ;
  assign n17963 = n17721 & ~n17962 ;
  assign n17964 = n17963 ^ n6621 ^ 1'b0 ;
  assign n17965 = n6696 & n11815 ;
  assign n17966 = ~n5449 & n17965 ;
  assign n17967 = n2545 | n17966 ;
  assign n17968 = n2140 & ~n16709 ;
  assign n17969 = n12748 & ~n17051 ;
  assign n17970 = ( ~n2465 & n10485 ) | ( ~n2465 & n13054 ) | ( n10485 & n13054 ) ;
  assign n17979 = ( ~x73 & n2132 ) | ( ~x73 & n7105 ) | ( n2132 & n7105 ) ;
  assign n17980 = n2716 | n17979 ;
  assign n17975 = n5073 & ~n5796 ;
  assign n17976 = n6737 & n17975 ;
  assign n17972 = n3565 | n11373 ;
  assign n17973 = n17972 ^ n2503 ^ 1'b0 ;
  assign n17974 = n17973 ^ n7770 ^ n735 ;
  assign n17977 = n17976 ^ n17974 ^ n8976 ;
  assign n17971 = ( n747 & ~n1610 ) | ( n747 & n6391 ) | ( ~n1610 & n6391 ) ;
  assign n17978 = n17977 ^ n17971 ^ n13650 ;
  assign n17981 = n17980 ^ n17978 ^ n3366 ;
  assign n17982 = ~n2673 & n6352 ;
  assign n17983 = ( n16766 & n17981 ) | ( n16766 & ~n17982 ) | ( n17981 & ~n17982 ) ;
  assign n17984 = n733 ^ n537 ^ x174 ;
  assign n17985 = n4571 & ~n17984 ;
  assign n17986 = n9455 ^ n5639 ^ n3694 ;
  assign n17987 = ( n3488 & n7806 ) | ( n3488 & ~n17986 ) | ( n7806 & ~n17986 ) ;
  assign n17988 = n13655 & ~n17987 ;
  assign n17989 = n7501 & n17988 ;
  assign n17990 = n14073 ^ n13508 ^ n8133 ;
  assign n17991 = n15598 ^ n8964 ^ 1'b0 ;
  assign n17992 = n7499 & n17991 ;
  assign n17993 = ~n11958 & n15552 ;
  assign n17994 = n17993 ^ n5445 ^ 1'b0 ;
  assign n17995 = ( ~n10214 & n13541 ) | ( ~n10214 & n17994 ) | ( n13541 & n17994 ) ;
  assign n17996 = n4593 ^ n716 ^ 1'b0 ;
  assign n17997 = n3782 & ~n17996 ;
  assign n17998 = n6053 & n17997 ;
  assign n17999 = n8396 & n17998 ;
  assign n18000 = ( n6507 & ~n17062 ) | ( n6507 & n17999 ) | ( ~n17062 & n17999 ) ;
  assign n18001 = ~n3845 & n18000 ;
  assign n18002 = n5545 ^ n3523 ^ n1049 ;
  assign n18003 = ( n2741 & n6990 ) | ( n2741 & n18002 ) | ( n6990 & n18002 ) ;
  assign n18004 = n17629 ^ n7414 ^ n6935 ;
  assign n18005 = n7673 ^ n2663 ^ 1'b0 ;
  assign n18006 = n18005 ^ n3671 ^ n3233 ;
  assign n18007 = n5529 | n6541 ;
  assign n18008 = n18007 ^ n6753 ^ 1'b0 ;
  assign n18009 = n3736 & n8977 ;
  assign n18010 = n18009 ^ n6092 ^ 1'b0 ;
  assign n18011 = n3225 | n18010 ;
  assign n18012 = n18008 | n18011 ;
  assign n18013 = n3172 | n12465 ;
  assign n18016 = n6642 & n14690 ;
  assign n18017 = n18016 ^ n7103 ^ 1'b0 ;
  assign n18014 = n11298 | n11687 ;
  assign n18015 = n6129 | n18014 ;
  assign n18018 = n18017 ^ n18015 ^ 1'b0 ;
  assign n18019 = ~n4369 & n18018 ;
  assign n18020 = n14718 ^ n7326 ^ n6458 ;
  assign n18021 = n7860 ^ n7184 ^ n4471 ;
  assign n18022 = n1415 & n16758 ;
  assign n18023 = n18021 & n18022 ;
  assign n18024 = ~n8937 & n18023 ;
  assign n18025 = n5638 ^ n4240 ^ n1503 ;
  assign n18026 = n18025 ^ n10024 ^ n2709 ;
  assign n18027 = n11227 & ~n18026 ;
  assign n18028 = n8508 ^ n3986 ^ 1'b0 ;
  assign n18029 = n18028 ^ n5733 ^ 1'b0 ;
  assign n18030 = n18029 ^ n5820 ^ 1'b0 ;
  assign n18031 = ~n9216 & n18030 ;
  assign n18032 = n3173 & n5707 ;
  assign n18033 = n14008 ^ n4244 ^ 1'b0 ;
  assign n18034 = n18032 & n18033 ;
  assign n18035 = n10684 ^ n4585 ^ n1936 ;
  assign n18036 = ~n790 & n18035 ;
  assign n18037 = n3888 | n10027 ;
  assign n18038 = n18036 & n18037 ;
  assign n18039 = n2065 & ~n5948 ;
  assign n18040 = n18039 ^ n2229 ^ 1'b0 ;
  assign n18041 = n8172 ^ n3261 ^ 1'b0 ;
  assign n18042 = ~n3165 & n18041 ;
  assign n18043 = n9660 ^ n3746 ^ n1597 ;
  assign n18044 = n18042 & ~n18043 ;
  assign n18045 = n18044 ^ n1884 ^ 1'b0 ;
  assign n18046 = ( n5422 & n18040 ) | ( n5422 & ~n18045 ) | ( n18040 & ~n18045 ) ;
  assign n18047 = n5573 & ~n6950 ;
  assign n18048 = n18047 ^ x154 ^ 1'b0 ;
  assign n18049 = n18048 ^ n8754 ^ n6639 ;
  assign n18050 = n10648 & n18049 ;
  assign n18051 = ( n6991 & n7588 ) | ( n6991 & ~n17883 ) | ( n7588 & ~n17883 ) ;
  assign n18052 = n8518 ^ n6852 ^ 1'b0 ;
  assign n18053 = n18052 ^ n14563 ^ 1'b0 ;
  assign n18054 = n17559 ^ n15616 ^ n13335 ;
  assign n18055 = n6205 & ~n18054 ;
  assign n18056 = n18055 ^ n5566 ^ 1'b0 ;
  assign n18063 = ( n516 & n4622 ) | ( n516 & ~n7581 ) | ( n4622 & ~n7581 ) ;
  assign n18057 = n9901 ^ n7672 ^ n5795 ;
  assign n18058 = n409 & ~n18057 ;
  assign n18059 = n18058 ^ n690 ^ 1'b0 ;
  assign n18060 = ~n11623 & n14030 ;
  assign n18061 = ~n338 & n18060 ;
  assign n18062 = n18059 & ~n18061 ;
  assign n18064 = n18063 ^ n18062 ^ 1'b0 ;
  assign n18065 = ( n1537 & ~n3335 ) | ( n1537 & n15055 ) | ( ~n3335 & n15055 ) ;
  assign n18066 = ~x10 & n12834 ;
  assign n18067 = n18065 & n18066 ;
  assign n18068 = ( n611 & n1594 ) | ( n611 & n5741 ) | ( n1594 & n5741 ) ;
  assign n18069 = ( n5092 & n13993 ) | ( n5092 & n18068 ) | ( n13993 & n18068 ) ;
  assign n18070 = n7413 ^ n6030 ^ n5928 ;
  assign n18071 = ~n10185 & n13295 ;
  assign n18072 = ~n2793 & n13582 ;
  assign n18073 = ~n18071 & n18072 ;
  assign n18074 = n18073 ^ n6596 ^ 1'b0 ;
  assign n18075 = n5116 & n18074 ;
  assign n18076 = ( n5359 & n11565 ) | ( n5359 & ~n18075 ) | ( n11565 & ~n18075 ) ;
  assign n18077 = n410 & n6530 ;
  assign n18078 = ( ~n3243 & n4180 ) | ( ~n3243 & n10364 ) | ( n4180 & n10364 ) ;
  assign n18079 = n18078 ^ n16608 ^ n6468 ;
  assign n18080 = n4327 & n18079 ;
  assign n18081 = n9451 & n18080 ;
  assign n18082 = n18003 ^ n7790 ^ 1'b0 ;
  assign n18083 = ( n10509 & n13363 ) | ( n10509 & ~n14251 ) | ( n13363 & ~n14251 ) ;
  assign n18084 = n9622 & ~n18083 ;
  assign n18085 = n13724 ^ n12750 ^ 1'b0 ;
  assign n18086 = ( ~n6247 & n18084 ) | ( ~n6247 & n18085 ) | ( n18084 & n18085 ) ;
  assign n18087 = n2251 & n11661 ;
  assign n18088 = n3353 & n16670 ;
  assign n18089 = ~n13439 & n18088 ;
  assign n18090 = n9779 | n12599 ;
  assign n18091 = n18089 | n18090 ;
  assign n18092 = n18091 ^ n7366 ^ 1'b0 ;
  assign n18093 = ( ~n10735 & n11796 ) | ( ~n10735 & n14695 ) | ( n11796 & n14695 ) ;
  assign n18094 = ( n2119 & n2179 ) | ( n2119 & ~n4517 ) | ( n2179 & ~n4517 ) ;
  assign n18095 = n9970 | n13260 ;
  assign n18096 = n18095 ^ n1839 ^ 1'b0 ;
  assign n18097 = n818 & n10914 ;
  assign n18098 = ( n3909 & n7554 ) | ( n3909 & ~n7683 ) | ( n7554 & ~n7683 ) ;
  assign n18099 = n18098 ^ n10846 ^ 1'b0 ;
  assign n18100 = n18097 & ~n18099 ;
  assign n18106 = ~n3301 & n4199 ;
  assign n18101 = n4514 ^ n3021 ^ n1678 ;
  assign n18102 = n13282 & ~n18101 ;
  assign n18103 = n18102 ^ n8552 ^ 1'b0 ;
  assign n18104 = ( n756 & ~n1806 ) | ( n756 & n3907 ) | ( ~n1806 & n3907 ) ;
  assign n18105 = ( n5457 & n18103 ) | ( n5457 & n18104 ) | ( n18103 & n18104 ) ;
  assign n18107 = n18106 ^ n18105 ^ n6518 ;
  assign n18108 = n7477 ^ n2865 ^ n1159 ;
  assign n18109 = n18108 ^ n8438 ^ 1'b0 ;
  assign n18110 = n14373 ^ n12163 ^ n8559 ;
  assign n18111 = ~n4251 & n8624 ;
  assign n18112 = n18111 ^ n9658 ^ n3238 ;
  assign n18113 = n7441 | n18112 ;
  assign n18114 = n18113 ^ n3190 ^ 1'b0 ;
  assign n18115 = n8638 & ~n18114 ;
  assign n18116 = ( n5160 & n9663 ) | ( n5160 & ~n18115 ) | ( n9663 & ~n18115 ) ;
  assign n18117 = ~n1425 & n18116 ;
  assign n18125 = n2175 & n7163 ;
  assign n18126 = ~n16961 & n18125 ;
  assign n18120 = ( ~n2100 & n8676 ) | ( ~n2100 & n12113 ) | ( n8676 & n12113 ) ;
  assign n18121 = n18120 ^ n3792 ^ 1'b0 ;
  assign n18122 = n18121 ^ n400 ^ 1'b0 ;
  assign n18123 = n11302 ^ n6744 ^ 1'b0 ;
  assign n18124 = n18122 & n18123 ;
  assign n18118 = n14817 ^ n2994 ^ 1'b0 ;
  assign n18119 = n5222 | n18118 ;
  assign n18127 = n18126 ^ n18124 ^ n18119 ;
  assign n18128 = n405 & n11896 ;
  assign n18129 = n18128 ^ n15548 ^ n2845 ;
  assign n18131 = n9213 ^ n6455 ^ 1'b0 ;
  assign n18132 = n444 & n18131 ;
  assign n18130 = n3578 | n16836 ;
  assign n18133 = n18132 ^ n18130 ^ 1'b0 ;
  assign n18134 = n7664 ^ n4937 ^ 1'b0 ;
  assign n18135 = ( ~n798 & n6829 ) | ( ~n798 & n16822 ) | ( n6829 & n16822 ) ;
  assign n18136 = n18135 ^ n15019 ^ 1'b0 ;
  assign n18137 = n18134 & n18136 ;
  assign n18138 = n17887 ^ n16584 ^ 1'b0 ;
  assign n18139 = n1444 | n18138 ;
  assign n18140 = n17850 ^ n3186 ^ 1'b0 ;
  assign n18141 = n18140 ^ n16713 ^ 1'b0 ;
  assign n18142 = n2243 & ~n6111 ;
  assign n18143 = n18142 ^ n5418 ^ 1'b0 ;
  assign n18144 = ( n5402 & n17800 ) | ( n5402 & ~n18143 ) | ( n17800 & ~n18143 ) ;
  assign n18145 = n18144 ^ n11681 ^ 1'b0 ;
  assign n18146 = ~n7993 & n18145 ;
  assign n18147 = n7388 & ~n11244 ;
  assign n18148 = ( n5544 & ~n10030 ) | ( n5544 & n18010 ) | ( ~n10030 & n18010 ) ;
  assign n18149 = ( ~n10496 & n14406 ) | ( ~n10496 & n18148 ) | ( n14406 & n18148 ) ;
  assign n18150 = n14821 ^ n9897 ^ 1'b0 ;
  assign n18151 = n4826 | n18150 ;
  assign n18152 = n18151 ^ n17351 ^ n4151 ;
  assign n18153 = n8631 ^ n6795 ^ n3407 ;
  assign n18154 = n18153 ^ n13744 ^ 1'b0 ;
  assign n18155 = n6629 ^ n3420 ^ n3331 ;
  assign n18156 = ( n2121 & ~n3075 ) | ( n2121 & n18155 ) | ( ~n3075 & n18155 ) ;
  assign n18157 = n18156 ^ n17657 ^ 1'b0 ;
  assign n18158 = n10715 ^ n1665 ^ 1'b0 ;
  assign n18159 = n18157 & n18158 ;
  assign n18160 = n1173 | n8192 ;
  assign n18161 = n18160 ^ n7924 ^ 1'b0 ;
  assign n18162 = ~n1379 & n2464 ;
  assign n18163 = n18161 & n18162 ;
  assign n18164 = n18163 ^ n17445 ^ 1'b0 ;
  assign n18165 = n2081 & n4522 ;
  assign n18166 = n8838 & ~n15719 ;
  assign n18167 = ( n8606 & ~n18165 ) | ( n8606 & n18166 ) | ( ~n18165 & n18166 ) ;
  assign n18168 = ( n3617 & n12070 ) | ( n3617 & n18167 ) | ( n12070 & n18167 ) ;
  assign n18172 = n6064 | n14091 ;
  assign n18169 = ( n493 & n1601 ) | ( n493 & n2540 ) | ( n1601 & n2540 ) ;
  assign n18170 = n5397 ^ n3115 ^ 1'b0 ;
  assign n18171 = n18169 | n18170 ;
  assign n18173 = n18172 ^ n18171 ^ n8681 ;
  assign n18174 = n6252 & n9423 ;
  assign n18175 = n18174 ^ n15845 ^ n6693 ;
  assign n18176 = ~n7165 & n7410 ;
  assign n18177 = n18176 ^ n16826 ^ 1'b0 ;
  assign n18178 = n5135 ^ n5008 ^ n2631 ;
  assign n18179 = n18178 ^ n12521 ^ 1'b0 ;
  assign n18180 = ~n4968 & n18179 ;
  assign n18183 = n5554 ^ n1908 ^ 1'b0 ;
  assign n18184 = n3289 & n18183 ;
  assign n18185 = n18184 ^ n17366 ^ n1095 ;
  assign n18181 = ~n3032 & n14929 ;
  assign n18182 = n10057 | n18181 ;
  assign n18186 = n18185 ^ n18182 ^ 1'b0 ;
  assign n18187 = ( x188 & n9150 ) | ( x188 & ~n14489 ) | ( n9150 & ~n14489 ) ;
  assign n18188 = ( ~n1133 & n8304 ) | ( ~n1133 & n18187 ) | ( n8304 & n18187 ) ;
  assign n18192 = ~n5612 & n15183 ;
  assign n18193 = ~n10423 & n18192 ;
  assign n18194 = n18193 ^ n9064 ^ 1'b0 ;
  assign n18195 = n3907 & ~n18194 ;
  assign n18189 = n15949 ^ n5523 ^ n1949 ;
  assign n18190 = ~n5433 & n18189 ;
  assign n18191 = n18190 ^ n17522 ^ 1'b0 ;
  assign n18196 = n18195 ^ n18191 ^ n9124 ;
  assign n18197 = n12558 ^ n3427 ^ n966 ;
  assign n18198 = n3248 & n9825 ;
  assign n18199 = n18198 ^ n17384 ^ 1'b0 ;
  assign n18200 = n18199 ^ n2227 ^ n1723 ;
  assign n18201 = n1594 & ~n12919 ;
  assign n18202 = n8910 & ~n18201 ;
  assign n18203 = n18202 ^ n9610 ^ 1'b0 ;
  assign n18204 = n12806 & ~n18203 ;
  assign n18205 = n18200 & n18204 ;
  assign n18206 = x83 & n18205 ;
  assign n18207 = ~n13328 & n18206 ;
  assign n18208 = n18207 ^ n1795 ^ 1'b0 ;
  assign n18209 = ( n3060 & n9083 ) | ( n3060 & n12590 ) | ( n9083 & n12590 ) ;
  assign n18210 = ( n5809 & ~n6096 ) | ( n5809 & n9411 ) | ( ~n6096 & n9411 ) ;
  assign n18211 = n1146 & n18210 ;
  assign n18212 = ~n18209 & n18211 ;
  assign n18214 = ( x230 & n7796 ) | ( x230 & n11760 ) | ( n7796 & n11760 ) ;
  assign n18213 = n10427 | n10608 ;
  assign n18215 = n18214 ^ n18213 ^ 1'b0 ;
  assign n18216 = n4669 & n10509 ;
  assign n18217 = ( n12348 & ~n15783 ) | ( n12348 & n18216 ) | ( ~n15783 & n18216 ) ;
  assign n18221 = n3099 ^ n595 ^ 1'b0 ;
  assign n18222 = n9619 | n18221 ;
  assign n18223 = ( n3006 & n3623 ) | ( n3006 & ~n18222 ) | ( n3623 & ~n18222 ) ;
  assign n18218 = n2436 & n5461 ;
  assign n18219 = ~x82 & n9572 ;
  assign n18220 = n18218 & n18219 ;
  assign n18224 = n18223 ^ n18220 ^ n13645 ;
  assign n18225 = n18217 | n18224 ;
  assign n18226 = n7108 | n18225 ;
  assign n18227 = n8769 | n10460 ;
  assign n18228 = n18227 ^ n2525 ^ 1'b0 ;
  assign n18232 = ( ~n3240 & n3924 ) | ( ~n3240 & n9417 ) | ( n3924 & n9417 ) ;
  assign n18233 = n6089 & n18232 ;
  assign n18234 = n2458 & n18233 ;
  assign n18229 = n3841 ^ n593 ^ 1'b0 ;
  assign n18230 = ( ~n1146 & n3549 ) | ( ~n1146 & n13408 ) | ( n3549 & n13408 ) ;
  assign n18231 = ( n1726 & ~n18229 ) | ( n1726 & n18230 ) | ( ~n18229 & n18230 ) ;
  assign n18235 = n18234 ^ n18231 ^ 1'b0 ;
  assign n18238 = n7043 ^ n825 ^ 1'b0 ;
  assign n18239 = n2020 & n18238 ;
  assign n18236 = n8620 & n9735 ;
  assign n18237 = n18236 ^ n13089 ^ n7069 ;
  assign n18240 = n18239 ^ n18237 ^ n9851 ;
  assign n18244 = ( ~n1539 & n3441 ) | ( ~n1539 & n4272 ) | ( n3441 & n4272 ) ;
  assign n18241 = n12527 ^ n2657 ^ 1'b0 ;
  assign n18242 = n8429 & ~n18241 ;
  assign n18243 = ( x102 & n5891 ) | ( x102 & n18242 ) | ( n5891 & n18242 ) ;
  assign n18245 = n18244 ^ n18243 ^ 1'b0 ;
  assign n18247 = ~n8622 & n10287 ;
  assign n18246 = ( n652 & ~n3425 ) | ( n652 & n7236 ) | ( ~n3425 & n7236 ) ;
  assign n18248 = n18247 ^ n18246 ^ n1494 ;
  assign n18249 = n18248 ^ n16670 ^ n13687 ;
  assign n18250 = n4548 & ~n18249 ;
  assign n18251 = n8802 | n18250 ;
  assign n18252 = n18245 & ~n18251 ;
  assign n18254 = n16533 ^ n8122 ^ n3927 ;
  assign n18253 = n17000 ^ n7856 ^ n4041 ;
  assign n18255 = n18254 ^ n18253 ^ 1'b0 ;
  assign n18256 = n18255 ^ n3167 ^ n2960 ;
  assign n18257 = n2722 & n18256 ;
  assign n18258 = ( n1380 & ~n7826 ) | ( n1380 & n9902 ) | ( ~n7826 & n9902 ) ;
  assign n18259 = n10009 ^ n4238 ^ n3759 ;
  assign n18260 = ( n8062 & n11031 ) | ( n8062 & ~n18259 ) | ( n11031 & ~n18259 ) ;
  assign n18261 = n9247 ^ n8531 ^ n8350 ;
  assign n18262 = n9628 ^ n6611 ^ n3499 ;
  assign n18263 = n18262 ^ n9067 ^ 1'b0 ;
  assign n18264 = n7593 & n18263 ;
  assign n18265 = n12046 ^ n6923 ^ n2139 ;
  assign n18266 = n693 & ~n18265 ;
  assign n18267 = n18266 ^ n17433 ^ 1'b0 ;
  assign n18268 = n18264 & ~n18267 ;
  assign n18269 = ~n2518 & n18268 ;
  assign n18270 = n18261 & n18269 ;
  assign n18287 = n11907 | n11961 ;
  assign n18288 = n18287 ^ n2954 ^ 1'b0 ;
  assign n18289 = ( x199 & n4109 ) | ( x199 & n7790 ) | ( n4109 & n7790 ) ;
  assign n18290 = n3406 | n8331 ;
  assign n18291 = n18290 ^ n2169 ^ 1'b0 ;
  assign n18292 = n18291 ^ n7511 ^ n496 ;
  assign n18293 = n18289 & n18292 ;
  assign n18294 = n18288 & n18293 ;
  assign n18295 = n18294 ^ n10123 ^ 1'b0 ;
  assign n18271 = n7332 ^ n2139 ^ n936 ;
  assign n18272 = n6148 & n8495 ;
  assign n18273 = n18272 ^ n5439 ^ 1'b0 ;
  assign n18274 = n7673 ^ n1932 ^ 1'b0 ;
  assign n18275 = n18273 | n18274 ;
  assign n18276 = n4098 & ~n18275 ;
  assign n18277 = n5512 & n18276 ;
  assign n18278 = n18277 ^ n7558 ^ 1'b0 ;
  assign n18279 = n7425 & n18278 ;
  assign n18280 = n4644 ^ n3587 ^ 1'b0 ;
  assign n18281 = x222 & ~n18280 ;
  assign n18282 = n18281 ^ n7363 ^ n2021 ;
  assign n18283 = ~n11255 & n18282 ;
  assign n18284 = ~n11006 & n18283 ;
  assign n18285 = ( n11447 & n18279 ) | ( n11447 & n18284 ) | ( n18279 & n18284 ) ;
  assign n18286 = n18271 & n18285 ;
  assign n18296 = n18295 ^ n18286 ^ 1'b0 ;
  assign n18297 = n5737 & n11171 ;
  assign n18298 = n6822 & n18297 ;
  assign n18299 = n18298 ^ n12070 ^ n1840 ;
  assign n18300 = n4393 ^ n1920 ^ 1'b0 ;
  assign n18301 = n4217 & ~n18300 ;
  assign n18302 = ~n585 & n18301 ;
  assign n18303 = n5086 & n18302 ;
  assign n18304 = n4340 & n18303 ;
  assign n18305 = n9814 & n13228 ;
  assign n18306 = ~n18304 & n18305 ;
  assign n18310 = ( n5781 & n6607 ) | ( n5781 & ~n17732 ) | ( n6607 & ~n17732 ) ;
  assign n18307 = n4639 ^ n3178 ^ 1'b0 ;
  assign n18308 = ~n3390 & n18307 ;
  assign n18309 = ~n15899 & n18308 ;
  assign n18311 = n18310 ^ n18309 ^ 1'b0 ;
  assign n18312 = n12038 | n18311 ;
  assign n18313 = n1935 | n4393 ;
  assign n18314 = n4898 | n18313 ;
  assign n18315 = n10077 & n18314 ;
  assign n18316 = n13772 ^ n3330 ^ 1'b0 ;
  assign n18317 = n18315 & n18316 ;
  assign n18318 = n18317 ^ n6960 ^ 1'b0 ;
  assign n18319 = n18318 ^ n9340 ^ 1'b0 ;
  assign n18320 = n17265 ^ n16720 ^ n4902 ;
  assign n18321 = n16665 & n18320 ;
  assign n18322 = n16312 ^ n12333 ^ n4781 ;
  assign n18323 = n13107 ^ n5112 ^ n2522 ;
  assign n18324 = n3418 | n18323 ;
  assign n18326 = n7595 ^ n4932 ^ n681 ;
  assign n18327 = ( n2629 & ~n6316 ) | ( n2629 & n18326 ) | ( ~n6316 & n18326 ) ;
  assign n18325 = n5760 & n14875 ;
  assign n18328 = n18327 ^ n18325 ^ 1'b0 ;
  assign n18329 = n18324 | n18328 ;
  assign n18331 = x82 & ~n6260 ;
  assign n18330 = n1919 | n10657 ;
  assign n18332 = n18331 ^ n18330 ^ n9775 ;
  assign n18333 = n5507 ^ n1077 ^ 1'b0 ;
  assign n18334 = ~n4025 & n18333 ;
  assign n18335 = ( n8149 & n14942 ) | ( n8149 & ~n18334 ) | ( n14942 & ~n18334 ) ;
  assign n18336 = n18335 ^ n750 ^ 1'b0 ;
  assign n18337 = n488 ^ x187 ^ 1'b0 ;
  assign n18338 = n18337 ^ n5793 ^ n5368 ;
  assign n18339 = n18338 ^ n7790 ^ 1'b0 ;
  assign n18340 = n18339 ^ n10274 ^ 1'b0 ;
  assign n18347 = ~n3427 & n3507 ;
  assign n18348 = n18347 ^ n7158 ^ 1'b0 ;
  assign n18349 = n18348 ^ n1894 ^ 1'b0 ;
  assign n18345 = n7936 ^ n3915 ^ n1591 ;
  assign n18342 = n12150 | n17499 ;
  assign n18343 = n14210 & ~n18342 ;
  assign n18344 = n8617 | n18343 ;
  assign n18346 = n18345 ^ n18344 ^ 1'b0 ;
  assign n18341 = n17655 ^ n5307 ^ 1'b0 ;
  assign n18350 = n18349 ^ n18346 ^ n18341 ;
  assign n18351 = n3203 | n8091 ;
  assign n18352 = ( n367 & n14868 ) | ( n367 & n18351 ) | ( n14868 & n18351 ) ;
  assign n18353 = n5233 ^ n2412 ^ 1'b0 ;
  assign n18354 = n5451 & ~n18353 ;
  assign n18355 = n18354 ^ n6913 ^ n6326 ;
  assign n18356 = ( n17999 & n18352 ) | ( n17999 & n18355 ) | ( n18352 & n18355 ) ;
  assign n18357 = ~n17687 & n18356 ;
  assign n18358 = n11345 & n11492 ;
  assign n18359 = n18358 ^ n16638 ^ 1'b0 ;
  assign n18360 = n4813 ^ n3707 ^ 1'b0 ;
  assign n18361 = ( ~x5 & n1959 ) | ( ~x5 & n11157 ) | ( n1959 & n11157 ) ;
  assign n18362 = n18361 ^ n9927 ^ 1'b0 ;
  assign n18363 = n8800 | n18362 ;
  assign n18364 = ~n12291 & n18363 ;
  assign n18365 = n4581 | n15830 ;
  assign n18366 = n2442 | n15636 ;
  assign n18367 = n6689 ^ x129 ^ 1'b0 ;
  assign n18368 = n611 | n18367 ;
  assign n18369 = n18366 | n18368 ;
  assign n18374 = n5683 ^ n954 ^ 1'b0 ;
  assign n18370 = ( n1775 & n4811 ) | ( n1775 & ~n7577 ) | ( n4811 & ~n7577 ) ;
  assign n18371 = ( n7058 & n10376 ) | ( n7058 & n18370 ) | ( n10376 & n18370 ) ;
  assign n18372 = n1961 ^ x10 ^ 1'b0 ;
  assign n18373 = n18371 & ~n18372 ;
  assign n18375 = n18374 ^ n18373 ^ n3031 ;
  assign n18376 = n2796 | n18375 ;
  assign n18377 = n18376 ^ n6462 ^ 1'b0 ;
  assign n18378 = n7217 & n8818 ;
  assign n18379 = n18378 ^ n9974 ^ 1'b0 ;
  assign n18380 = n6075 ^ n5567 ^ n1706 ;
  assign n18381 = n6788 | n18380 ;
  assign n18382 = n2029 | n6815 ;
  assign n18383 = n5219 ^ n1785 ^ 1'b0 ;
  assign n18384 = n9605 | n18383 ;
  assign n18385 = ( ~n5214 & n12950 ) | ( ~n5214 & n18384 ) | ( n12950 & n18384 ) ;
  assign n18386 = ( x144 & n18382 ) | ( x144 & n18385 ) | ( n18382 & n18385 ) ;
  assign n18387 = ~n1701 & n18386 ;
  assign n18388 = n18387 ^ n6497 ^ 1'b0 ;
  assign n18389 = n13438 ^ n13246 ^ 1'b0 ;
  assign n18392 = n9562 ^ n8280 ^ 1'b0 ;
  assign n18393 = ~n3298 & n18392 ;
  assign n18390 = ~n6193 & n7154 ;
  assign n18391 = n18214 & ~n18390 ;
  assign n18394 = n18393 ^ n18391 ^ 1'b0 ;
  assign n18395 = n8203 ^ n5878 ^ 1'b0 ;
  assign n18396 = n2026 | n5848 ;
  assign n18397 = ( ~n12137 & n18395 ) | ( ~n12137 & n18396 ) | ( n18395 & n18396 ) ;
  assign n18398 = ~n6689 & n10428 ;
  assign n18399 = ~n4484 & n9040 ;
  assign n18401 = n1233 ^ n757 ^ 1'b0 ;
  assign n18402 = n5340 | n18401 ;
  assign n18403 = ( n4382 & ~n8290 ) | ( n4382 & n18402 ) | ( ~n8290 & n18402 ) ;
  assign n18400 = n3520 | n8982 ;
  assign n18404 = n18403 ^ n18400 ^ 1'b0 ;
  assign n18405 = n18404 ^ x188 ^ 1'b0 ;
  assign n18406 = n18399 & ~n18405 ;
  assign n18407 = ( ~n1383 & n1848 ) | ( ~n1383 & n6307 ) | ( n1848 & n6307 ) ;
  assign n18408 = n11976 & n16435 ;
  assign n18409 = n18408 ^ n13415 ^ 1'b0 ;
  assign n18410 = n6982 & ~n18409 ;
  assign n18411 = ~n9915 & n18410 ;
  assign n18412 = n18407 & n18411 ;
  assign n18413 = n3080 | n5381 ;
  assign n18414 = n2130 & ~n18413 ;
  assign n18415 = n5601 ^ n676 ^ 1'b0 ;
  assign n18416 = ~n6005 & n12233 ;
  assign n18417 = n17870 & n18416 ;
  assign n18418 = n18415 & ~n18417 ;
  assign n18419 = n18414 & n18418 ;
  assign n18420 = n2819 | n6295 ;
  assign n18421 = x153 & n18420 ;
  assign n18422 = n13856 ^ n1317 ^ 1'b0 ;
  assign n18423 = n12359 & ~n18422 ;
  assign n18424 = n15556 & n18423 ;
  assign n18425 = ( ~n4057 & n18421 ) | ( ~n4057 & n18424 ) | ( n18421 & n18424 ) ;
  assign n18426 = n10524 & n12630 ;
  assign n18427 = n18426 ^ n7228 ^ 1'b0 ;
  assign n18428 = n16493 ^ n7152 ^ 1'b0 ;
  assign n18429 = n9191 & ~n18428 ;
  assign n18430 = n9309 & ~n15424 ;
  assign n18431 = n18430 ^ n313 ^ 1'b0 ;
  assign n18433 = n8200 | n14502 ;
  assign n18434 = n18433 ^ n12509 ^ 1'b0 ;
  assign n18432 = n2063 | n6282 ;
  assign n18435 = n18434 ^ n18432 ^ 1'b0 ;
  assign n18436 = ( n15523 & n18431 ) | ( n15523 & ~n18435 ) | ( n18431 & ~n18435 ) ;
  assign n18437 = n3584 & ~n18436 ;
  assign n18438 = n18437 ^ n9334 ^ 1'b0 ;
  assign n18441 = ( ~n4114 & n5112 ) | ( ~n4114 & n9625 ) | ( n5112 & n9625 ) ;
  assign n18439 = n894 | n947 ;
  assign n18440 = n18439 ^ n2737 ^ 1'b0 ;
  assign n18442 = n18441 ^ n18440 ^ 1'b0 ;
  assign n18443 = n4163 & ~n4881 ;
  assign n18444 = n18443 ^ n8658 ^ 1'b0 ;
  assign n18445 = n12733 & n18444 ;
  assign n18446 = ( n593 & n3792 ) | ( n593 & n8019 ) | ( n3792 & n8019 ) ;
  assign n18447 = n18446 ^ n16412 ^ n7138 ;
  assign n18448 = ~n3397 & n15683 ;
  assign n18449 = ~n18447 & n18448 ;
  assign n18450 = ( ~n1928 & n3310 ) | ( ~n1928 & n4304 ) | ( n3310 & n4304 ) ;
  assign n18451 = ~n15315 & n18450 ;
  assign n18452 = x27 & n18451 ;
  assign n18453 = n18449 & n18452 ;
  assign n18454 = n11043 & n16803 ;
  assign n18457 = n367 & n1209 ;
  assign n18458 = n9678 ^ n9120 ^ 1'b0 ;
  assign n18459 = n18457 | n18458 ;
  assign n18455 = ~n1654 & n2574 ;
  assign n18456 = n18455 ^ n9853 ^ 1'b0 ;
  assign n18460 = n18459 ^ n18456 ^ n12393 ;
  assign n18461 = n18460 ^ n8321 ^ n6272 ;
  assign n18462 = ( n4946 & n4978 ) | ( n4946 & ~n9759 ) | ( n4978 & ~n9759 ) ;
  assign n18463 = ( n3070 & n13799 ) | ( n3070 & n16765 ) | ( n13799 & n16765 ) ;
  assign n18464 = ( n3496 & ~n18462 ) | ( n3496 & n18463 ) | ( ~n18462 & n18463 ) ;
  assign n18465 = ~n4622 & n6160 ;
  assign n18466 = n18465 ^ n1810 ^ 1'b0 ;
  assign n18467 = n6033 & n18466 ;
  assign n18468 = n3336 & ~n18467 ;
  assign n18469 = n18468 ^ n10949 ^ 1'b0 ;
  assign n18470 = ( n11009 & n12098 ) | ( n11009 & ~n15644 ) | ( n12098 & ~n15644 ) ;
  assign n18471 = n18470 ^ n8230 ^ n3487 ;
  assign n18472 = n18471 ^ n11294 ^ 1'b0 ;
  assign n18473 = ( ~n8056 & n14972 ) | ( ~n8056 & n15672 ) | ( n14972 & n15672 ) ;
  assign n18474 = n13127 ^ n542 ^ 1'b0 ;
  assign n18475 = n541 & n18474 ;
  assign n18476 = ~n1837 & n18475 ;
  assign n18477 = ~n284 & n7752 ;
  assign n18478 = n10571 ^ n2441 ^ 1'b0 ;
  assign n18483 = ( n4315 & n9865 ) | ( n4315 & n13828 ) | ( n9865 & n13828 ) ;
  assign n18484 = ( n2812 & ~n4740 ) | ( n2812 & n18483 ) | ( ~n4740 & n18483 ) ;
  assign n18479 = ~n5137 & n9655 ;
  assign n18480 = n7356 ^ n2791 ^ 1'b0 ;
  assign n18481 = n18479 | n18480 ;
  assign n18482 = n18481 ^ n15843 ^ n15649 ;
  assign n18485 = n18484 ^ n18482 ^ n7494 ;
  assign n18486 = n8243 ^ n6374 ^ 1'b0 ;
  assign n18487 = n11810 ^ n3088 ^ 1'b0 ;
  assign n18488 = n9305 ^ n9109 ^ 1'b0 ;
  assign n18489 = n1435 & ~n4386 ;
  assign n18490 = n4619 & n18489 ;
  assign n18491 = ( ~n1556 & n18488 ) | ( ~n1556 & n18490 ) | ( n18488 & n18490 ) ;
  assign n18494 = n1208 & n6251 ;
  assign n18495 = ~n7012 & n18494 ;
  assign n18492 = n6612 | n7172 ;
  assign n18493 = n18492 ^ n13749 ^ n10076 ;
  assign n18496 = n18495 ^ n18493 ^ 1'b0 ;
  assign n18497 = n7925 & n16095 ;
  assign n18498 = ~n15234 & n18497 ;
  assign n18499 = ( n1944 & n12061 ) | ( n1944 & ~n18498 ) | ( n12061 & ~n18498 ) ;
  assign n18500 = ( n3018 & n7865 ) | ( n3018 & n8273 ) | ( n7865 & n8273 ) ;
  assign n18501 = ~n11936 & n18500 ;
  assign n18502 = n18501 ^ n3780 ^ 1'b0 ;
  assign n18503 = ( n3745 & ~n4048 ) | ( n3745 & n6739 ) | ( ~n4048 & n6739 ) ;
  assign n18504 = n11115 | n18503 ;
  assign n18505 = ( ~n6070 & n6481 ) | ( ~n6070 & n8781 ) | ( n6481 & n8781 ) ;
  assign n18506 = ~x153 & n4442 ;
  assign n18507 = n758 & ~n18506 ;
  assign n18508 = n18505 & n18507 ;
  assign n18509 = x81 & n8357 ;
  assign n18511 = x158 & ~n1164 ;
  assign n18512 = n18511 ^ n1854 ^ 1'b0 ;
  assign n18510 = n13037 ^ n10114 ^ n2211 ;
  assign n18513 = n18512 ^ n18510 ^ n5650 ;
  assign n18514 = n15456 ^ n14958 ^ n321 ;
  assign n18515 = n6465 | n9295 ;
  assign n18516 = n6488 & n17120 ;
  assign n18517 = n18516 ^ n16824 ^ 1'b0 ;
  assign n18518 = n17651 ^ n14193 ^ 1'b0 ;
  assign n18519 = n6863 | n10838 ;
  assign n18520 = ( n8894 & ~n18518 ) | ( n8894 & n18519 ) | ( ~n18518 & n18519 ) ;
  assign n18521 = n12837 ^ n10707 ^ 1'b0 ;
  assign n18522 = ( n2128 & ~n6064 ) | ( n2128 & n18521 ) | ( ~n6064 & n18521 ) ;
  assign n18523 = n1311 ^ n564 ^ 1'b0 ;
  assign n18524 = n816 & n16350 ;
  assign n18525 = n18524 ^ n6784 ^ 1'b0 ;
  assign n18526 = n14155 ^ n2553 ^ x11 ;
  assign n18527 = ( n9160 & n13017 ) | ( n9160 & n18526 ) | ( n13017 & n18526 ) ;
  assign n18528 = n10546 | n16230 ;
  assign n18529 = n18527 & ~n18528 ;
  assign n18530 = n8053 ^ n4717 ^ n1654 ;
  assign n18531 = n5907 | n5980 ;
  assign n18532 = n2946 | n18531 ;
  assign n18533 = n16768 & ~n18532 ;
  assign n18534 = n18533 ^ n14072 ^ n3586 ;
  assign n18535 = ( n1454 & n6449 ) | ( n1454 & ~n18534 ) | ( n6449 & ~n18534 ) ;
  assign n18536 = n675 | n18535 ;
  assign n18537 = ( n16195 & n18530 ) | ( n16195 & n18536 ) | ( n18530 & n18536 ) ;
  assign n18538 = n14433 ^ n13459 ^ n7373 ;
  assign n18539 = n18317 & ~n18538 ;
  assign n18540 = n18539 ^ n12059 ^ 1'b0 ;
  assign n18541 = ~n6247 & n7460 ;
  assign n18542 = n18541 ^ n14829 ^ 1'b0 ;
  assign n18543 = n2340 & ~n18542 ;
  assign n18544 = n4087 & n18543 ;
  assign n18545 = n18544 ^ n15919 ^ 1'b0 ;
  assign n18546 = n13161 ^ n9142 ^ 1'b0 ;
  assign n18547 = n10251 & n18546 ;
  assign n18548 = n13213 ^ n11246 ^ 1'b0 ;
  assign n18549 = n13160 | n18548 ;
  assign n18550 = n2008 | n18549 ;
  assign n18551 = n7750 | n18550 ;
  assign n18554 = x217 & ~n10728 ;
  assign n18555 = ~n3074 & n18554 ;
  assign n18552 = n11439 ^ n4329 ^ 1'b0 ;
  assign n18553 = n9119 & n18552 ;
  assign n18556 = n18555 ^ n18553 ^ 1'b0 ;
  assign n18557 = ( n8548 & ~n11192 ) | ( n8548 & n18556 ) | ( ~n11192 & n18556 ) ;
  assign n18558 = ~n5248 & n8780 ;
  assign n18559 = n18220 & n18558 ;
  assign n18560 = ~n4260 & n6930 ;
  assign n18561 = n18559 & n18560 ;
  assign n18562 = n3375 ^ n3114 ^ 1'b0 ;
  assign n18563 = ~n5053 & n18562 ;
  assign n18564 = n12893 & n18563 ;
  assign n18565 = ~n3712 & n18564 ;
  assign n18566 = n18565 ^ n2963 ^ 1'b0 ;
  assign n18567 = n7756 ^ n4745 ^ 1'b0 ;
  assign n18568 = ( n885 & n2654 ) | ( n885 & n8533 ) | ( n2654 & n8533 ) ;
  assign n18569 = n18568 ^ n17884 ^ 1'b0 ;
  assign n18570 = n8453 ^ n633 ^ 1'b0 ;
  assign n18571 = n12247 ^ n6360 ^ n3598 ;
  assign n18572 = n1220 & n9654 ;
  assign n18573 = n18572 ^ n3919 ^ 1'b0 ;
  assign n18574 = n18573 ^ n16917 ^ n4497 ;
  assign n18575 = ( n1336 & ~n6270 ) | ( n1336 & n13039 ) | ( ~n6270 & n13039 ) ;
  assign n18576 = n18575 ^ n17997 ^ n6347 ;
  assign n18577 = ( n6928 & n18574 ) | ( n6928 & ~n18576 ) | ( n18574 & ~n18576 ) ;
  assign n18578 = n13718 ^ n2160 ^ n855 ;
  assign n18579 = n10873 ^ n10248 ^ n3091 ;
  assign n18580 = n12546 ^ n737 ^ 1'b0 ;
  assign n18581 = x92 & ~n18580 ;
  assign n18582 = n6420 & n18581 ;
  assign n18583 = n18582 ^ n9616 ^ 1'b0 ;
  assign n18585 = ( n10034 & n15784 ) | ( n10034 & ~n18352 ) | ( n15784 & ~n18352 ) ;
  assign n18584 = n8858 | n9087 ;
  assign n18586 = n18585 ^ n18584 ^ 1'b0 ;
  assign n18587 = n8895 ^ n3724 ^ n500 ;
  assign n18588 = n9030 & ~n10416 ;
  assign n18589 = n1024 & ~n18588 ;
  assign n18590 = n18589 ^ n926 ^ 1'b0 ;
  assign n18591 = n4002 & n12726 ;
  assign n18592 = n18591 ^ n14056 ^ n7291 ;
  assign n18593 = n11245 ^ n930 ^ 1'b0 ;
  assign n18599 = n3225 & n8424 ;
  assign n18600 = n1121 & n18599 ;
  assign n18601 = ~n964 & n7108 ;
  assign n18602 = n18601 ^ n12522 ^ 1'b0 ;
  assign n18603 = ( ~n12682 & n18600 ) | ( ~n12682 & n18602 ) | ( n18600 & n18602 ) ;
  assign n18594 = n1629 & n11235 ;
  assign n18595 = n18594 ^ n15930 ^ 1'b0 ;
  assign n18596 = n3382 ^ n2909 ^ n1640 ;
  assign n18597 = n18595 & ~n18596 ;
  assign n18598 = ~n1631 & n18597 ;
  assign n18604 = n18603 ^ n18598 ^ n10053 ;
  assign n18605 = n4548 & n12462 ;
  assign n18606 = ~n6125 & n6735 ;
  assign n18607 = n18606 ^ n4059 ^ 1'b0 ;
  assign n18608 = n13554 | n18607 ;
  assign n18609 = n17489 ^ n17472 ^ n6114 ;
  assign n18610 = n4187 & ~n6276 ;
  assign n18611 = n18610 ^ n11418 ^ 1'b0 ;
  assign n18612 = ~n3502 & n18611 ;
  assign n18615 = ( n2074 & n4799 ) | ( n2074 & n8008 ) | ( n4799 & n8008 ) ;
  assign n18616 = n3071 | n18615 ;
  assign n18613 = n11001 ^ n7962 ^ 1'b0 ;
  assign n18614 = n6033 | n18613 ;
  assign n18617 = n18616 ^ n18614 ^ 1'b0 ;
  assign n18618 = ( ~n15528 & n18612 ) | ( ~n15528 & n18617 ) | ( n18612 & n18617 ) ;
  assign n18619 = x79 & ~n2049 ;
  assign n18620 = n18619 ^ n9765 ^ n9691 ;
  assign n18621 = n7721 ^ n6584 ^ 1'b0 ;
  assign n18622 = n3979 & n18621 ;
  assign n18623 = n9446 & ~n18622 ;
  assign n18624 = ( n13664 & n18620 ) | ( n13664 & n18623 ) | ( n18620 & n18623 ) ;
  assign n18625 = ( n4044 & n5462 ) | ( n4044 & n14024 ) | ( n5462 & n14024 ) ;
  assign n18626 = n18625 ^ n14839 ^ 1'b0 ;
  assign n18627 = n18624 | n18626 ;
  assign n18629 = ~n1261 & n7846 ;
  assign n18630 = n6402 & ~n18629 ;
  assign n18631 = n9592 & n18630 ;
  assign n18628 = n3839 & ~n12613 ;
  assign n18632 = n18631 ^ n18628 ^ 1'b0 ;
  assign n18633 = n18632 ^ n3019 ^ 1'b0 ;
  assign n18634 = n14051 | n18633 ;
  assign n18641 = n5825 ^ n316 ^ x166 ;
  assign n18642 = n18641 ^ n18040 ^ n8087 ;
  assign n18643 = n9564 | n18642 ;
  assign n18635 = ~n3521 & n6249 ;
  assign n18636 = n18635 ^ n5369 ^ 1'b0 ;
  assign n18637 = n8149 | n18431 ;
  assign n18638 = n18637 ^ n7047 ^ 1'b0 ;
  assign n18639 = ( n11777 & n18636 ) | ( n11777 & n18638 ) | ( n18636 & n18638 ) ;
  assign n18640 = n18639 ^ n11764 ^ n1348 ;
  assign n18644 = n18643 ^ n18640 ^ n5521 ;
  assign n18645 = n7146 ^ n4239 ^ 1'b0 ;
  assign n18646 = ~n12426 & n14745 ;
  assign n18647 = ( n459 & n7881 ) | ( n459 & n11595 ) | ( n7881 & n11595 ) ;
  assign n18648 = n1802 & n9205 ;
  assign n18649 = n18648 ^ n4240 ^ 1'b0 ;
  assign n18650 = ( n10687 & n18647 ) | ( n10687 & ~n18649 ) | ( n18647 & ~n18649 ) ;
  assign n18651 = n10714 ^ n3778 ^ n2963 ;
  assign n18652 = n4626 & n18651 ;
  assign n18653 = n11649 & ~n17585 ;
  assign n18654 = n18652 & n18653 ;
  assign n18655 = n9641 | n11996 ;
  assign n18656 = n2458 & n8624 ;
  assign n18657 = ~n4292 & n18656 ;
  assign n18658 = ( n10680 & ~n17347 ) | ( n10680 & n18657 ) | ( ~n17347 & n18657 ) ;
  assign n18659 = n18658 ^ n16761 ^ 1'b0 ;
  assign n18660 = n18659 ^ n462 ^ 1'b0 ;
  assign n18661 = n9285 | n17391 ;
  assign n18662 = ~n5521 & n18661 ;
  assign n18663 = n5144 & ~n10792 ;
  assign n18665 = n11453 ^ n9581 ^ n7364 ;
  assign n18664 = n13864 ^ n8621 ^ n7474 ;
  assign n18666 = n18665 ^ n18664 ^ n3941 ;
  assign n18667 = ( n16244 & n18663 ) | ( n16244 & ~n18666 ) | ( n18663 & ~n18666 ) ;
  assign n18668 = n11419 ^ n2041 ^ 1'b0 ;
  assign n18669 = ~n9164 & n13066 ;
  assign n18670 = n18669 ^ n1934 ^ 1'b0 ;
  assign n18671 = ( n13191 & ~n18668 ) | ( n13191 & n18670 ) | ( ~n18668 & n18670 ) ;
  assign n18676 = n9726 ^ n4714 ^ n2241 ;
  assign n18677 = n5868 & ~n13061 ;
  assign n18678 = n18676 & n18677 ;
  assign n18679 = n18678 ^ n15466 ^ 1'b0 ;
  assign n18680 = n9089 | n18679 ;
  assign n18672 = ( n7199 & n9534 ) | ( n7199 & n10448 ) | ( n9534 & n10448 ) ;
  assign n18673 = n4978 ^ n3452 ^ 1'b0 ;
  assign n18674 = n18673 ^ n13349 ^ 1'b0 ;
  assign n18675 = n18672 | n18674 ;
  assign n18681 = n18680 ^ n18675 ^ n9966 ;
  assign n18686 = x80 & n6862 ;
  assign n18687 = n14402 & n18686 ;
  assign n18688 = n18687 ^ n10288 ^ n9585 ;
  assign n18682 = ( n1564 & n5592 ) | ( n1564 & ~n6420 ) | ( n5592 & ~n6420 ) ;
  assign n18683 = ~n18402 & n18682 ;
  assign n18684 = n18683 ^ n11825 ^ n9652 ;
  assign n18685 = n10631 & n18684 ;
  assign n18689 = n18688 ^ n18685 ^ 1'b0 ;
  assign n18690 = n17904 & n18331 ;
  assign n18691 = n15531 & n18690 ;
  assign n18692 = n5762 | n18691 ;
  assign n18693 = n18692 ^ n11457 ^ 1'b0 ;
  assign n18694 = n4436 & n18693 ;
  assign n18695 = n2481 | n6152 ;
  assign n18696 = n4338 | n18695 ;
  assign n18697 = n18696 ^ n999 ^ 1'b0 ;
  assign n18698 = n17111 ^ n16570 ^ 1'b0 ;
  assign n18699 = n5217 ^ n3923 ^ x106 ;
  assign n18700 = n6428 | n8760 ;
  assign n18701 = n18699 | n18700 ;
  assign n18702 = n11064 | n18701 ;
  assign n18706 = ~n8880 & n16665 ;
  assign n18707 = n18706 ^ n12244 ^ 1'b0 ;
  assign n18708 = n18707 ^ n11550 ^ 1'b0 ;
  assign n18703 = n11866 ^ n8880 ^ n1941 ;
  assign n18704 = n16115 ^ n8036 ^ 1'b0 ;
  assign n18705 = n18703 & ~n18704 ;
  assign n18709 = n18708 ^ n18705 ^ n996 ;
  assign n18710 = n2035 & n8231 ;
  assign n18711 = n18710 ^ n10507 ^ 1'b0 ;
  assign n18712 = n949 | n18711 ;
  assign n18713 = n2870 ^ n704 ^ 1'b0 ;
  assign n18714 = n18201 | n18713 ;
  assign n18715 = n4465 | n5486 ;
  assign n18716 = n10379 ^ n2492 ^ 1'b0 ;
  assign n18717 = n11551 & ~n18716 ;
  assign n18718 = ~n13717 & n18717 ;
  assign n18719 = n13577 ^ n11300 ^ n7727 ;
  assign n18720 = n5407 ^ n1700 ^ n524 ;
  assign n18721 = n11689 & ~n18720 ;
  assign n18722 = n18721 ^ n3585 ^ 1'b0 ;
  assign n18723 = n18722 ^ n11638 ^ n1188 ;
  assign n18724 = n2854 ^ n468 ^ 1'b0 ;
  assign n18725 = n6092 & n18724 ;
  assign n18726 = ~n2850 & n6540 ;
  assign n18727 = ~n14588 & n18726 ;
  assign n18728 = ( n18279 & n18725 ) | ( n18279 & ~n18727 ) | ( n18725 & ~n18727 ) ;
  assign n18729 = n6066 ^ n5941 ^ 1'b0 ;
  assign n18730 = ( n7263 & n13831 ) | ( n7263 & n18729 ) | ( n13831 & n18729 ) ;
  assign n18731 = n8939 ^ n1912 ^ 1'b0 ;
  assign n18732 = n898 & n3857 ;
  assign n18733 = n18732 ^ n9953 ^ 1'b0 ;
  assign n18734 = n282 & ~n8025 ;
  assign n18735 = ( n18151 & n18733 ) | ( n18151 & n18734 ) | ( n18733 & n18734 ) ;
  assign n18736 = n766 & n10151 ;
  assign n18737 = ~n13237 & n18736 ;
  assign n18738 = n4341 ^ n1568 ^ 1'b0 ;
  assign n18739 = n16852 | n18738 ;
  assign n18740 = n3322 | n7574 ;
  assign n18741 = n18739 | n18740 ;
  assign n18742 = n3664 ^ n2694 ^ 1'b0 ;
  assign n18743 = n17074 ^ n16537 ^ n15771 ;
  assign n18744 = n17223 ^ n8506 ^ n7976 ;
  assign n18745 = ( n3009 & n15841 ) | ( n3009 & n18744 ) | ( n15841 & n18744 ) ;
  assign n18746 = n14852 ^ n7963 ^ n477 ;
  assign n18747 = n18746 ^ n3555 ^ 1'b0 ;
  assign n18748 = n5646 ^ n4733 ^ n4240 ;
  assign n18749 = n15240 & ~n18748 ;
  assign n18751 = n14945 ^ n10079 ^ n9285 ;
  assign n18750 = n10763 ^ n10498 ^ 1'b0 ;
  assign n18752 = n18751 ^ n18750 ^ 1'b0 ;
  assign n18753 = ~n4626 & n18752 ;
  assign n18754 = n18753 ^ n18741 ^ n13819 ;
  assign n18755 = n14906 ^ n12244 ^ 1'b0 ;
  assign n18756 = n14159 | n18755 ;
  assign n18757 = n13257 & ~n18756 ;
  assign n18758 = ~n4047 & n18757 ;
  assign n18759 = n15579 ^ n12658 ^ n7662 ;
  assign n18760 = n18759 ^ n13178 ^ n767 ;
  assign n18761 = n4513 ^ n1997 ^ n861 ;
  assign n18762 = n18703 & n18761 ;
  assign n18763 = n18762 ^ n14091 ^ 1'b0 ;
  assign n18764 = ~n1099 & n3645 ;
  assign n18765 = n2254 & ~n18764 ;
  assign n18766 = ( n1037 & n7752 ) | ( n1037 & ~n18765 ) | ( n7752 & ~n18765 ) ;
  assign n18767 = n13028 & ~n16860 ;
  assign n18768 = ( n15730 & n18766 ) | ( n15730 & ~n18767 ) | ( n18766 & ~n18767 ) ;
  assign n18770 = ( n1624 & n3353 ) | ( n1624 & ~n4027 ) | ( n3353 & ~n4027 ) ;
  assign n18771 = ( n1014 & ~n15623 ) | ( n1014 & n18770 ) | ( ~n15623 & n18770 ) ;
  assign n18769 = ~n3140 & n12210 ;
  assign n18772 = n18771 ^ n18769 ^ n9927 ;
  assign n18773 = n13573 ^ n944 ^ 1'b0 ;
  assign n18779 = n3254 & ~n5602 ;
  assign n18777 = n3387 ^ n2482 ^ n2040 ;
  assign n18778 = n18777 ^ n9369 ^ 1'b0 ;
  assign n18780 = n18779 ^ n18778 ^ n17171 ;
  assign n18781 = n18780 ^ n9018 ^ 1'b0 ;
  assign n18774 = n5368 ^ n317 ^ 1'b0 ;
  assign n18775 = n871 | n5270 ;
  assign n18776 = n18774 | n18775 ;
  assign n18782 = n18781 ^ n18776 ^ 1'b0 ;
  assign n18783 = ~n18773 & n18782 ;
  assign n18784 = n8763 & ~n10854 ;
  assign n18785 = n2961 & n18784 ;
  assign n18786 = ( n393 & n5299 ) | ( n393 & ~n18785 ) | ( n5299 & ~n18785 ) ;
  assign n18787 = ( ~n1545 & n15199 ) | ( ~n1545 & n18786 ) | ( n15199 & n18786 ) ;
  assign n18790 = n5228 ^ n1246 ^ 1'b0 ;
  assign n18788 = ~n8839 & n11087 ;
  assign n18789 = n18788 ^ n4555 ^ 1'b0 ;
  assign n18791 = n18790 ^ n18789 ^ n10757 ;
  assign n18796 = n4455 ^ n3000 ^ n2941 ;
  assign n18792 = n1323 ^ x200 ^ 1'b0 ;
  assign n18793 = n3665 & n18792 ;
  assign n18794 = n18793 ^ n8475 ^ 1'b0 ;
  assign n18795 = n3459 | n18794 ;
  assign n18797 = n18796 ^ n18795 ^ n10699 ;
  assign n18798 = n18797 ^ n17934 ^ 1'b0 ;
  assign n18799 = n6831 & ~n15956 ;
  assign n18800 = n9137 & n18799 ;
  assign n18801 = ( ~n3314 & n3651 ) | ( ~n3314 & n18800 ) | ( n3651 & n18800 ) ;
  assign n18802 = n967 | n6974 ;
  assign n18803 = n18801 & ~n18802 ;
  assign n18804 = n416 | n15351 ;
  assign n18805 = n18804 ^ n3301 ^ 1'b0 ;
  assign n18806 = n13491 ^ n1482 ^ 1'b0 ;
  assign n18807 = n3672 | n18806 ;
  assign n18808 = n18805 | n18807 ;
  assign n18809 = n6832 & ~n12399 ;
  assign n18810 = n18809 ^ n6240 ^ 1'b0 ;
  assign n18811 = n18810 ^ n11591 ^ n10743 ;
  assign n18812 = n10389 & n12474 ;
  assign n18813 = ~n6449 & n18474 ;
  assign n18814 = n18813 ^ n258 ^ 1'b0 ;
  assign n18815 = ( ~n8483 & n14628 ) | ( ~n8483 & n18814 ) | ( n14628 & n18814 ) ;
  assign n18816 = ( ~n4093 & n6690 ) | ( ~n4093 & n18815 ) | ( n6690 & n18815 ) ;
  assign n18817 = n18526 ^ n14787 ^ n2560 ;
  assign n18822 = n3644 & ~n17226 ;
  assign n18823 = n18822 ^ n4733 ^ 1'b0 ;
  assign n18820 = n2106 & n12456 ;
  assign n18821 = ~n7361 & n18820 ;
  assign n18818 = n1136 | n5276 ;
  assign n18819 = n2782 & ~n18818 ;
  assign n18824 = n18823 ^ n18821 ^ n18819 ;
  assign n18825 = ( n6518 & ~n9746 ) | ( n6518 & n12721 ) | ( ~n9746 & n12721 ) ;
  assign n18826 = ( n3171 & n6273 ) | ( n3171 & ~n18825 ) | ( n6273 & ~n18825 ) ;
  assign n18827 = n3983 & ~n14563 ;
  assign n18828 = ( n2441 & n14611 ) | ( n2441 & ~n17325 ) | ( n14611 & ~n17325 ) ;
  assign n18829 = ( n2453 & n12443 ) | ( n2453 & ~n18828 ) | ( n12443 & ~n18828 ) ;
  assign n18830 = n4152 & ~n18829 ;
  assign n18831 = ~n13220 & n18830 ;
  assign n18832 = ( n6800 & n13904 ) | ( n6800 & ~n18767 ) | ( n13904 & ~n18767 ) ;
  assign n18833 = n15298 ^ n8335 ^ n3303 ;
  assign n18834 = n10521 & ~n18833 ;
  assign n18835 = x19 & n5214 ;
  assign n18838 = ( x132 & n2722 ) | ( x132 & ~n3428 ) | ( n2722 & ~n3428 ) ;
  assign n18836 = n2341 ^ x5 ^ 1'b0 ;
  assign n18837 = n12531 | n18836 ;
  assign n18839 = n18838 ^ n18837 ^ 1'b0 ;
  assign n18840 = ( ~n3496 & n8240 ) | ( ~n3496 & n18839 ) | ( n8240 & n18839 ) ;
  assign n18844 = n9042 ^ n6451 ^ 1'b0 ;
  assign n18845 = n18844 ^ n7913 ^ 1'b0 ;
  assign n18841 = n10027 ^ n9877 ^ n5735 ;
  assign n18842 = n8614 ^ n7932 ^ n5791 ;
  assign n18843 = n18841 & n18842 ;
  assign n18846 = n18845 ^ n18843 ^ 1'b0 ;
  assign n18852 = n4612 ^ n3530 ^ n2180 ;
  assign n18853 = n18852 ^ n4862 ^ 1'b0 ;
  assign n18854 = n18853 ^ n9852 ^ n5003 ;
  assign n18847 = ( n2553 & n9632 ) | ( n2553 & ~n10139 ) | ( n9632 & ~n10139 ) ;
  assign n18848 = n8495 ^ n3032 ^ n2106 ;
  assign n18849 = ~n789 & n18848 ;
  assign n18850 = n18849 ^ n4390 ^ 1'b0 ;
  assign n18851 = n18847 & n18850 ;
  assign n18855 = n18854 ^ n18851 ^ 1'b0 ;
  assign n18856 = ( ~n2103 & n18652 ) | ( ~n2103 & n18855 ) | ( n18652 & n18855 ) ;
  assign n18857 = n10436 | n18856 ;
  assign n18858 = n2468 & ~n18857 ;
  assign n18859 = n14381 & ~n16250 ;
  assign n18860 = n16932 ^ n10448 ^ 1'b0 ;
  assign n18861 = n11512 & n18860 ;
  assign n18862 = n3857 | n16221 ;
  assign n18863 = n18861 & ~n18862 ;
  assign n18864 = ~n6897 & n10793 ;
  assign n18865 = ~n18863 & n18864 ;
  assign n18866 = ( n2281 & n3240 ) | ( n2281 & ~n6699 ) | ( n3240 & ~n6699 ) ;
  assign n18867 = n18866 ^ n11840 ^ 1'b0 ;
  assign n18868 = n5037 | n18867 ;
  assign n18869 = x54 & ~n11055 ;
  assign n18872 = n748 & n13421 ;
  assign n18870 = n9102 & ~n18374 ;
  assign n18871 = ~n8011 & n18870 ;
  assign n18873 = n18872 ^ n18871 ^ n11546 ;
  assign n18874 = ( n306 & ~n2066 ) | ( n306 & n7517 ) | ( ~n2066 & n7517 ) ;
  assign n18875 = n13496 ^ n287 ^ 1'b0 ;
  assign n18876 = n18874 | n18875 ;
  assign n18877 = n4417 ^ n711 ^ 1'b0 ;
  assign n18878 = ~n2669 & n18877 ;
  assign n18879 = ( n14439 & ~n18122 ) | ( n14439 & n18878 ) | ( ~n18122 & n18878 ) ;
  assign n18880 = n17498 ^ n7170 ^ 1'b0 ;
  assign n18881 = n18880 ^ n13604 ^ n4544 ;
  assign n18882 = n3665 & ~n7957 ;
  assign n18883 = n15799 ^ n15641 ^ 1'b0 ;
  assign n18884 = n18883 ^ n759 ^ n749 ;
  assign n18885 = n8421 ^ n1883 ^ 1'b0 ;
  assign n18886 = n17679 | n18885 ;
  assign n18887 = n9997 ^ n9463 ^ n5851 ;
  assign n18888 = ( ~n18417 & n18886 ) | ( ~n18417 & n18887 ) | ( n18886 & n18887 ) ;
  assign n18890 = n4497 & ~n10529 ;
  assign n18891 = n18890 ^ n1853 ^ 1'b0 ;
  assign n18892 = n18891 ^ n5015 ^ n1567 ;
  assign n18889 = n3772 | n18239 ;
  assign n18893 = n18892 ^ n18889 ^ n6757 ;
  assign n18894 = n8861 ^ n2087 ^ 1'b0 ;
  assign n18895 = n18495 | n18894 ;
  assign n18896 = n18895 ^ n2297 ^ 1'b0 ;
  assign n18897 = n7742 ^ n5129 ^ 1'b0 ;
  assign n18898 = n1697 & ~n4455 ;
  assign n18899 = n1896 & n18898 ;
  assign n18900 = n2508 & n7166 ;
  assign n18901 = n5949 & n11341 ;
  assign n18902 = n18900 & n18901 ;
  assign n18903 = n18902 ^ n4424 ^ 1'b0 ;
  assign n18904 = ~n18899 & n18903 ;
  assign n18905 = n2823 & ~n9373 ;
  assign n18906 = n18905 ^ n3395 ^ 1'b0 ;
  assign n18907 = ( n5512 & n9922 ) | ( n5512 & ~n18906 ) | ( n9922 & ~n18906 ) ;
  assign n18908 = n756 | n6639 ;
  assign n18909 = n9056 & ~n18908 ;
  assign n18910 = n1586 | n18909 ;
  assign n18911 = n18910 ^ n10090 ^ 1'b0 ;
  assign n18912 = n17286 ^ n6216 ^ 1'b0 ;
  assign n18913 = n18911 & n18912 ;
  assign n18914 = n9568 ^ n7288 ^ 1'b0 ;
  assign n18915 = ~n1742 & n18914 ;
  assign n18916 = n13461 ^ n5647 ^ 1'b0 ;
  assign n18917 = n12109 | n13901 ;
  assign n18918 = n6453 ^ n2395 ^ n1684 ;
  assign n18919 = n18918 ^ n10687 ^ 1'b0 ;
  assign n18928 = n7024 ^ n6374 ^ n3397 ;
  assign n18929 = n18928 ^ n11171 ^ 1'b0 ;
  assign n18930 = n18929 ^ n15734 ^ 1'b0 ;
  assign n18931 = ~n11148 & n18930 ;
  assign n18932 = ( n8059 & n9295 ) | ( n8059 & n18931 ) | ( n9295 & n18931 ) ;
  assign n18921 = n18668 ^ n3430 ^ n1775 ;
  assign n18922 = ( n4413 & n5316 ) | ( n4413 & n18921 ) | ( n5316 & n18921 ) ;
  assign n18923 = n5542 & ~n18922 ;
  assign n18924 = ~n17186 & n18923 ;
  assign n18925 = n18924 ^ n793 ^ 1'b0 ;
  assign n18926 = ~n11853 & n18925 ;
  assign n18920 = n2075 & ~n16416 ;
  assign n18927 = n18926 ^ n18920 ^ n1776 ;
  assign n18933 = n18932 ^ n18927 ^ n17349 ;
  assign n18934 = ~n573 & n9381 ;
  assign n18935 = n18934 ^ n11363 ^ 1'b0 ;
  assign n18936 = n18935 ^ n12063 ^ n11374 ;
  assign n18937 = n18936 ^ n12191 ^ n1205 ;
  assign n18938 = ~n8768 & n17992 ;
  assign n18939 = n18938 ^ n15397 ^ 1'b0 ;
  assign n18940 = ( n2265 & n6771 ) | ( n2265 & ~n16585 ) | ( n6771 & ~n16585 ) ;
  assign n18941 = ~n2986 & n4728 ;
  assign n18942 = n18941 ^ n2696 ^ 1'b0 ;
  assign n18943 = n9070 | n18942 ;
  assign n18944 = n14090 & ~n18943 ;
  assign n18945 = ( n6554 & n15238 ) | ( n6554 & n18944 ) | ( n15238 & n18944 ) ;
  assign n18946 = n7679 ^ n7321 ^ 1'b0 ;
  assign n18947 = n9789 ^ n4639 ^ n2929 ;
  assign n18948 = n18947 ^ n11207 ^ 1'b0 ;
  assign n18949 = n10367 & ~n18948 ;
  assign n18950 = ~n9107 & n11357 ;
  assign n18951 = n1450 & n2825 ;
  assign n18952 = ~n13428 & n13987 ;
  assign n18953 = n18951 & n18952 ;
  assign n18954 = ~n7341 & n11594 ;
  assign n18955 = n11623 & n18954 ;
  assign n18956 = ( ~n9322 & n10419 ) | ( ~n9322 & n18955 ) | ( n10419 & n18955 ) ;
  assign n18957 = n15555 & n16852 ;
  assign n18958 = n3437 | n5458 ;
  assign n18959 = n18958 ^ n4866 ^ 1'b0 ;
  assign n18960 = ( n4907 & n14664 ) | ( n4907 & n18959 ) | ( n14664 & n18959 ) ;
  assign n18961 = n18960 ^ n15851 ^ 1'b0 ;
  assign n18962 = n6332 ^ n4594 ^ n3678 ;
  assign n18963 = n3110 ^ n915 ^ 1'b0 ;
  assign n18964 = ~n2071 & n9648 ;
  assign n18965 = n18964 ^ x153 ^ 1'b0 ;
  assign n18966 = n333 & ~n2781 ;
  assign n18967 = n18965 & n18966 ;
  assign n18968 = n18967 ^ n3303 ^ 1'b0 ;
  assign n18969 = n18963 & n18968 ;
  assign n18970 = n18969 ^ n13869 ^ 1'b0 ;
  assign n18971 = ( n12422 & ~n16683 ) | ( n12422 & n16860 ) | ( ~n16683 & n16860 ) ;
  assign n18972 = n18153 ^ n15846 ^ n15469 ;
  assign n18973 = n1664 & ~n16649 ;
  assign n18974 = n11051 & n18973 ;
  assign n18975 = n16768 & n18974 ;
  assign n18976 = n18975 ^ n6169 ^ n3499 ;
  assign n18977 = n18976 ^ n18161 ^ n10529 ;
  assign n18991 = n284 | n9361 ;
  assign n18992 = n4300 | n18991 ;
  assign n18988 = n1958 & n7140 ;
  assign n18989 = ~n6852 & n18988 ;
  assign n18990 = n18989 ^ n1894 ^ 1'b0 ;
  assign n18983 = n11352 ^ n1525 ^ 1'b0 ;
  assign n18984 = n2106 & n18983 ;
  assign n18978 = n6408 ^ n2249 ^ x152 ;
  assign n18979 = n18978 ^ n16970 ^ 1'b0 ;
  assign n18980 = n13708 & n16901 ;
  assign n18981 = n13561 & n18980 ;
  assign n18982 = n18979 & ~n18981 ;
  assign n18985 = n18984 ^ n18982 ^ 1'b0 ;
  assign n18986 = n6113 | n18985 ;
  assign n18987 = n18986 ^ n17152 ^ 1'b0 ;
  assign n18993 = n18992 ^ n18990 ^ n18987 ;
  assign n18994 = n2340 | n7090 ;
  assign n18995 = n17827 ^ n12317 ^ 1'b0 ;
  assign n18996 = n18994 & ~n18995 ;
  assign n18997 = n18996 ^ n7783 ^ 1'b0 ;
  assign n18998 = ( x102 & ~n10936 ) | ( x102 & n18997 ) | ( ~n10936 & n18997 ) ;
  assign n19000 = n3072 ^ n1943 ^ 1'b0 ;
  assign n18999 = n18162 ^ n16973 ^ n6659 ;
  assign n19001 = n19000 ^ n18999 ^ 1'b0 ;
  assign n19002 = n18998 | n19001 ;
  assign n19005 = n13905 ^ n7282 ^ 1'b0 ;
  assign n19006 = n19005 ^ n11352 ^ 1'b0 ;
  assign n19007 = n19006 ^ n12024 ^ 1'b0 ;
  assign n19003 = n17875 ^ n14266 ^ n8644 ;
  assign n19004 = ~n15909 & n19003 ;
  assign n19008 = n19007 ^ n19004 ^ 1'b0 ;
  assign n19009 = ( n3781 & ~n4928 ) | ( n3781 & n13655 ) | ( ~n4928 & n13655 ) ;
  assign n19010 = n14808 ^ n11303 ^ 1'b0 ;
  assign n19011 = n19009 & n19010 ;
  assign n19012 = n19011 ^ n16697 ^ n8480 ;
  assign n19013 = n19012 ^ n11505 ^ 1'b0 ;
  assign n19014 = n7112 ^ n776 ^ 1'b0 ;
  assign n19015 = n16472 ^ n14267 ^ 1'b0 ;
  assign n19016 = n6821 & n12122 ;
  assign n19017 = n19016 ^ n14916 ^ 1'b0 ;
  assign n19018 = n13909 ^ n2529 ^ n2514 ;
  assign n19019 = n3348 & n9521 ;
  assign n19020 = n19019 ^ n2100 ^ 1'b0 ;
  assign n19021 = n19020 ^ n3075 ^ 1'b0 ;
  assign n19022 = n19018 | n19021 ;
  assign n19023 = ~n1226 & n3917 ;
  assign n19024 = n7395 & n19023 ;
  assign n19025 = n17216 ^ n1916 ^ 1'b0 ;
  assign n19026 = n19024 | n19025 ;
  assign n19027 = n8955 ^ n8397 ^ 1'b0 ;
  assign n19028 = n3701 | n9973 ;
  assign n19029 = ~n19027 & n19028 ;
  assign n19030 = n19029 ^ n2405 ^ 1'b0 ;
  assign n19031 = n19030 ^ n6097 ^ n2620 ;
  assign n19032 = n2139 ^ n2050 ^ 1'b0 ;
  assign n19033 = ( n10464 & n10474 ) | ( n10464 & ~n13717 ) | ( n10474 & ~n13717 ) ;
  assign n19034 = n12834 ^ n6111 ^ n3372 ;
  assign n19035 = ~n12867 & n14749 ;
  assign n19036 = ~n4700 & n12997 ;
  assign n19037 = ~n4139 & n19036 ;
  assign n19038 = n3126 ^ n806 ^ 1'b0 ;
  assign n19039 = n19038 ^ n11029 ^ 1'b0 ;
  assign n19040 = n4816 & ~n10009 ;
  assign n19041 = ( n6222 & n8550 ) | ( n6222 & ~n14603 ) | ( n8550 & ~n14603 ) ;
  assign n19042 = n2916 & n18814 ;
  assign n19043 = n19042 ^ n10585 ^ n4226 ;
  assign n19044 = n626 & ~n16410 ;
  assign n19045 = ~n3765 & n8225 ;
  assign n19046 = ( ~n3509 & n9851 ) | ( ~n3509 & n13260 ) | ( n9851 & n13260 ) ;
  assign n19047 = n4021 & n19046 ;
  assign n19048 = n16208 ^ n7123 ^ 1'b0 ;
  assign n19049 = n8281 | n19048 ;
  assign n19050 = n12344 ^ n7930 ^ n681 ;
  assign n19051 = ( ~n1091 & n12472 ) | ( ~n1091 & n19050 ) | ( n12472 & n19050 ) ;
  assign n19052 = n8935 ^ n4147 ^ 1'b0 ;
  assign n19053 = n2042 & ~n19052 ;
  assign n19054 = ( n13852 & n17413 ) | ( n13852 & n19053 ) | ( n17413 & n19053 ) ;
  assign n19055 = n15348 ^ n5008 ^ 1'b0 ;
  assign n19056 = n4141 | n16124 ;
  assign n19057 = n18842 ^ n4757 ^ 1'b0 ;
  assign n19058 = n17701 & ~n19057 ;
  assign n19060 = n8779 & n18619 ;
  assign n19061 = n941 & n4828 ;
  assign n19062 = n19060 & n19061 ;
  assign n19059 = n2933 & ~n8411 ;
  assign n19063 = n19062 ^ n19059 ^ 1'b0 ;
  assign n19064 = n2445 | n2695 ;
  assign n19065 = n1345 & ~n19064 ;
  assign n19066 = n19065 ^ n2564 ^ 1'b0 ;
  assign n19067 = n1854 & n19066 ;
  assign n19068 = n19067 ^ n829 ^ 1'b0 ;
  assign n19069 = n5678 | n8217 ;
  assign n19070 = n19069 ^ n17171 ^ n6270 ;
  assign n19071 = n5975 | n10612 ;
  assign n19072 = n7428 & n8500 ;
  assign n19073 = n19072 ^ n2841 ^ 1'b0 ;
  assign n19074 = n19073 ^ n454 ^ 1'b0 ;
  assign n19075 = n9695 & ~n19074 ;
  assign n19076 = ( n2928 & ~n19071 ) | ( n2928 & n19075 ) | ( ~n19071 & n19075 ) ;
  assign n19079 = n3043 | n9659 ;
  assign n19080 = n19079 ^ n9762 ^ 1'b0 ;
  assign n19077 = ~n6977 & n10919 ;
  assign n19078 = ( n7300 & n17077 ) | ( n7300 & ~n19077 ) | ( n17077 & ~n19077 ) ;
  assign n19081 = n19080 ^ n19078 ^ 1'b0 ;
  assign n19086 = ( ~n299 & n1053 ) | ( ~n299 & n13991 ) | ( n1053 & n13991 ) ;
  assign n19083 = ~n7566 & n12483 ;
  assign n19084 = n4052 & n19083 ;
  assign n19082 = n9884 & n10724 ;
  assign n19085 = n19084 ^ n19082 ^ 1'b0 ;
  assign n19087 = n19086 ^ n19085 ^ n6608 ;
  assign n19088 = ( n10223 & ~n13575 ) | ( n10223 & n18909 ) | ( ~n13575 & n18909 ) ;
  assign n19089 = n12538 & ~n14258 ;
  assign n19090 = n1220 & n5918 ;
  assign n19091 = n19090 ^ n13074 ^ n3251 ;
  assign n19092 = n19091 ^ n13394 ^ 1'b0 ;
  assign n19093 = n5136 & n19092 ;
  assign n19094 = ( n10427 & n15991 ) | ( n10427 & n19093 ) | ( n15991 & n19093 ) ;
  assign n19095 = n3302 & n18220 ;
  assign n19096 = ~n8333 & n9521 ;
  assign n19097 = n19096 ^ n8896 ^ 1'b0 ;
  assign n19098 = n19097 ^ n14533 ^ n4364 ;
  assign n19099 = ~n16980 & n19098 ;
  assign n19100 = n8747 | n15747 ;
  assign n19101 = n19099 | n19100 ;
  assign n19102 = ~n5762 & n19101 ;
  assign n19103 = n19095 & n19102 ;
  assign n19107 = n2781 | n2862 ;
  assign n19108 = n19107 ^ n4156 ^ n4121 ;
  assign n19104 = n19097 ^ n9886 ^ 1'b0 ;
  assign n19105 = n4373 & ~n19104 ;
  assign n19106 = ( n8530 & ~n11347 ) | ( n8530 & n19105 ) | ( ~n11347 & n19105 ) ;
  assign n19109 = n19108 ^ n19106 ^ n1045 ;
  assign n19110 = n14956 ^ n12550 ^ n1578 ;
  assign n19111 = ~n4334 & n7149 ;
  assign n19112 = n1225 & n19111 ;
  assign n19113 = n19112 ^ n7641 ^ 1'b0 ;
  assign n19114 = n19113 ^ n18268 ^ n12096 ;
  assign n19115 = n1474 | n6168 ;
  assign n19116 = n4382 & ~n19115 ;
  assign n19117 = n1930 | n19116 ;
  assign n19118 = n19117 ^ n18396 ^ 1'b0 ;
  assign n19119 = n9438 ^ n3247 ^ 1'b0 ;
  assign n19120 = ~n9742 & n19119 ;
  assign n19121 = n2819 & n19120 ;
  assign n19122 = n6591 & ~n7302 ;
  assign n19123 = n19121 & n19122 ;
  assign n19124 = ( n1736 & n9816 ) | ( n1736 & ~n14132 ) | ( n9816 & ~n14132 ) ;
  assign n19125 = n19124 ^ n3891 ^ 1'b0 ;
  assign n19126 = n12293 ^ n1411 ^ 1'b0 ;
  assign n19127 = n13875 ^ n8635 ^ 1'b0 ;
  assign n19128 = n5912 & ~n19127 ;
  assign n19129 = n19128 ^ n12077 ^ 1'b0 ;
  assign n19130 = n9126 & n15237 ;
  assign n19131 = n19129 & ~n19130 ;
  assign n19134 = ( ~n1799 & n2669 ) | ( ~n1799 & n8918 ) | ( n2669 & n8918 ) ;
  assign n19135 = n12915 & ~n19134 ;
  assign n19136 = n19135 ^ n10994 ^ 1'b0 ;
  assign n19132 = ( n11929 & n12000 ) | ( n11929 & ~n17201 ) | ( n12000 & ~n17201 ) ;
  assign n19133 = n19132 ^ n14302 ^ n8210 ;
  assign n19137 = n19136 ^ n19133 ^ n8612 ;
  assign n19138 = n15487 ^ n12894 ^ n4153 ;
  assign n19139 = n4373 & n10423 ;
  assign n19140 = n3491 & n19139 ;
  assign n19141 = n9461 & n16518 ;
  assign n19142 = n2113 & n19141 ;
  assign n19143 = n8400 ^ n1046 ^ 1'b0 ;
  assign n19144 = n19143 ^ n4051 ^ 1'b0 ;
  assign n19145 = n6607 ^ n4837 ^ 1'b0 ;
  assign n19146 = ~n1113 & n19145 ;
  assign n19147 = ~n10561 & n19146 ;
  assign n19149 = n2986 ^ n1083 ^ 1'b0 ;
  assign n19148 = n12999 ^ n6027 ^ 1'b0 ;
  assign n19150 = n19149 ^ n19148 ^ n11872 ;
  assign n19151 = n780 | n825 ;
  assign n19152 = n767 & ~n19151 ;
  assign n19153 = n19152 ^ n9700 ^ n3683 ;
  assign n19154 = ~n6173 & n19153 ;
  assign n19155 = ~n3656 & n13544 ;
  assign n19156 = ~n8910 & n19155 ;
  assign n19157 = n19156 ^ n18294 ^ n14207 ;
  assign n19158 = n19154 | n19157 ;
  assign n19159 = n19158 ^ n14513 ^ 1'b0 ;
  assign n19160 = n3425 & n13379 ;
  assign n19161 = n4079 | n19160 ;
  assign n19162 = n3238 ^ n3015 ^ 1'b0 ;
  assign n19163 = n6938 | n19162 ;
  assign n19164 = n19163 ^ n11253 ^ 1'b0 ;
  assign n19165 = n19164 ^ n6390 ^ n5500 ;
  assign n19166 = ~n7165 & n12409 ;
  assign n19167 = ~n19165 & n19166 ;
  assign n19168 = n11581 | n19167 ;
  assign n19169 = n19168 ^ n4281 ^ 1'b0 ;
  assign n19170 = n770 & ~n14543 ;
  assign n19171 = n2906 | n6218 ;
  assign n19172 = ( n957 & n13794 ) | ( n957 & n19171 ) | ( n13794 & n19171 ) ;
  assign n19173 = n19172 ^ n10069 ^ n6404 ;
  assign n19174 = n617 | n17439 ;
  assign n19175 = n6316 ^ n4168 ^ 1'b0 ;
  assign n19176 = n17934 ^ n11049 ^ 1'b0 ;
  assign n19177 = n19175 | n19176 ;
  assign n19178 = n19177 ^ n10085 ^ 1'b0 ;
  assign n19179 = n4961 ^ n4281 ^ 1'b0 ;
  assign n19180 = ( ~n1533 & n19178 ) | ( ~n1533 & n19179 ) | ( n19178 & n19179 ) ;
  assign n19181 = n4684 ^ n4118 ^ 1'b0 ;
  assign n19182 = n15020 | n19181 ;
  assign n19183 = n7200 & ~n13755 ;
  assign n19184 = ~n8513 & n19183 ;
  assign n19185 = n2934 | n19184 ;
  assign n19186 = n19182 & ~n19185 ;
  assign n19187 = n9003 & ~n19186 ;
  assign n19194 = n5930 & n7252 ;
  assign n19195 = n19194 ^ n10239 ^ 1'b0 ;
  assign n19192 = n4393 & n4505 ;
  assign n19193 = n19192 ^ n12028 ^ n8450 ;
  assign n19196 = n19195 ^ n19193 ^ n7628 ;
  assign n19197 = n19196 ^ n11438 ^ n950 ;
  assign n19188 = n14341 ^ n2119 ^ 1'b0 ;
  assign n19189 = n15473 & ~n19188 ;
  assign n19190 = ( n3629 & ~n15066 ) | ( n3629 & n19189 ) | ( ~n15066 & n19189 ) ;
  assign n19191 = n11042 & n19190 ;
  assign n19198 = n19197 ^ n19191 ^ 1'b0 ;
  assign n19199 = ( ~n4832 & n8494 ) | ( ~n4832 & n19198 ) | ( n8494 & n19198 ) ;
  assign n19200 = ~n8586 & n10370 ;
  assign n19201 = n5240 & n19200 ;
  assign n19202 = x153 & n5462 ;
  assign n19203 = n19201 & n19202 ;
  assign n19204 = n11907 ^ n11524 ^ n6658 ;
  assign n19209 = ~n3713 & n6862 ;
  assign n19208 = n6788 & n7212 ;
  assign n19210 = n19209 ^ n19208 ^ 1'b0 ;
  assign n19207 = n2779 | n3107 ;
  assign n19205 = ~n9699 & n12409 ;
  assign n19206 = n13480 & ~n19205 ;
  assign n19211 = n19210 ^ n19207 ^ n19206 ;
  assign n19212 = n19211 ^ n16266 ^ n6237 ;
  assign n19213 = ( n1365 & ~n4615 ) | ( n1365 & n7060 ) | ( ~n4615 & n7060 ) ;
  assign n19214 = ( n4046 & n6593 ) | ( n4046 & n19213 ) | ( n6593 & n19213 ) ;
  assign n19215 = n11685 ^ n3986 ^ 1'b0 ;
  assign n19216 = n1975 & n19215 ;
  assign n19217 = n3668 ^ x5 ^ 1'b0 ;
  assign n19218 = n19216 & n19217 ;
  assign n19219 = ~n8598 & n19218 ;
  assign n19220 = ~n19214 & n19219 ;
  assign n19221 = n9149 ^ n8778 ^ 1'b0 ;
  assign n19222 = n2024 & n19221 ;
  assign n19223 = ~n13722 & n19222 ;
  assign n19224 = n19223 ^ n5681 ^ 1'b0 ;
  assign n19225 = n11559 ^ n6213 ^ 1'b0 ;
  assign n19226 = ( ~n5036 & n17276 ) | ( ~n5036 & n19225 ) | ( n17276 & n19225 ) ;
  assign n19227 = n16154 ^ n15558 ^ 1'b0 ;
  assign n19228 = n3109 & ~n5853 ;
  assign n19229 = n19228 ^ n9390 ^ n8488 ;
  assign n19230 = ( n3832 & n6680 ) | ( n3832 & ~n19229 ) | ( n6680 & ~n19229 ) ;
  assign n19231 = n15926 ^ n6043 ^ n4080 ;
  assign n19232 = ~n8314 & n19231 ;
  assign n19233 = n19232 ^ n9704 ^ 1'b0 ;
  assign n19234 = n10312 ^ n6089 ^ n5979 ;
  assign n19235 = n19233 & ~n19234 ;
  assign n19237 = ~n5171 & n5234 ;
  assign n19238 = n10926 & n19237 ;
  assign n19239 = ( ~n5168 & n9540 ) | ( ~n5168 & n19238 ) | ( n9540 & n19238 ) ;
  assign n19240 = n19239 ^ n5618 ^ 1'b0 ;
  assign n19241 = n17321 & n19240 ;
  assign n19236 = n7140 & ~n10930 ;
  assign n19242 = n19241 ^ n19236 ^ n13147 ;
  assign n19243 = n14857 ^ n12871 ^ n8292 ;
  assign n19244 = n14907 ^ n7659 ^ n4340 ;
  assign n19245 = n19244 ^ n15240 ^ n1769 ;
  assign n19246 = n17544 ^ n15424 ^ 1'b0 ;
  assign n19247 = n4902 & n19246 ;
  assign n19248 = n19247 ^ n3085 ^ 1'b0 ;
  assign n19249 = n8149 ^ n739 ^ 1'b0 ;
  assign n19250 = n1569 | n19249 ;
  assign n19251 = n19250 ^ n10791 ^ n5050 ;
  assign n19252 = n11866 ^ n7878 ^ n555 ;
  assign n19261 = ( n1743 & ~n4328 ) | ( n1743 & n5096 ) | ( ~n4328 & n5096 ) ;
  assign n19262 = n19261 ^ n11778 ^ 1'b0 ;
  assign n19263 = ( n8632 & n12191 ) | ( n8632 & n19262 ) | ( n12191 & n19262 ) ;
  assign n19253 = ( n5877 & ~n12596 ) | ( n5877 & n14686 ) | ( ~n12596 & n14686 ) ;
  assign n19256 = n9930 ^ n8358 ^ 1'b0 ;
  assign n19255 = n10723 | n12270 ;
  assign n19257 = n19256 ^ n19255 ^ n2647 ;
  assign n19258 = n19257 ^ n10745 ^ n1226 ;
  assign n19254 = n13605 & n18173 ;
  assign n19259 = n19258 ^ n19254 ^ 1'b0 ;
  assign n19260 = n19253 & ~n19259 ;
  assign n19264 = n19263 ^ n19260 ^ 1'b0 ;
  assign n19265 = n7563 ^ n2192 ^ n765 ;
  assign n19266 = n11683 | n19265 ;
  assign n19267 = n19266 ^ n13778 ^ 1'b0 ;
  assign n19268 = ( n14255 & ~n14691 ) | ( n14255 & n19267 ) | ( ~n14691 & n19267 ) ;
  assign n19269 = n9190 & ~n17817 ;
  assign n19270 = ~n3281 & n9610 ;
  assign n19271 = ~n3159 & n8059 ;
  assign n19272 = ~n19270 & n19271 ;
  assign n19277 = n1887 & ~n4527 ;
  assign n19278 = ~n1101 & n19277 ;
  assign n19273 = n577 | n5604 ;
  assign n19274 = n19273 ^ n9610 ^ 1'b0 ;
  assign n19275 = ( n1390 & n3438 ) | ( n1390 & ~n19274 ) | ( n3438 & ~n19274 ) ;
  assign n19276 = ( ~n4465 & n15868 ) | ( ~n4465 & n19275 ) | ( n15868 & n19275 ) ;
  assign n19279 = n19278 ^ n19276 ^ n1318 ;
  assign n19280 = ( ~n6939 & n11324 ) | ( ~n6939 & n12014 ) | ( n11324 & n12014 ) ;
  assign n19281 = n19280 ^ n3512 ^ n2260 ;
  assign n19283 = n13785 ^ n8981 ^ n6337 ;
  assign n19282 = n18079 ^ n10022 ^ n1173 ;
  assign n19284 = n19283 ^ n19282 ^ 1'b0 ;
  assign n19285 = n19281 & n19284 ;
  assign n19286 = n2592 | n5938 ;
  assign n19287 = n10109 | n19286 ;
  assign n19288 = n5729 & ~n17522 ;
  assign n19289 = ~n8663 & n19288 ;
  assign n19290 = n19289 ^ n3775 ^ 1'b0 ;
  assign n19291 = n12776 & n19290 ;
  assign n19293 = n5324 ^ n2909 ^ 1'b0 ;
  assign n19294 = n19293 ^ n12255 ^ 1'b0 ;
  assign n19295 = n8632 | n19294 ;
  assign n19292 = n2267 | n3133 ;
  assign n19296 = n19295 ^ n19292 ^ 1'b0 ;
  assign n19306 = ~n734 & n16003 ;
  assign n19307 = ( n6092 & ~n8930 ) | ( n6092 & n19306 ) | ( ~n8930 & n19306 ) ;
  assign n19301 = n1128 | n4201 ;
  assign n19302 = n1064 & ~n19301 ;
  assign n19303 = ( ~n5762 & n17423 ) | ( ~n5762 & n19302 ) | ( n17423 & n19302 ) ;
  assign n19304 = n19303 ^ n16958 ^ n1357 ;
  assign n19305 = n4635 & ~n19304 ;
  assign n19308 = n19307 ^ n19305 ^ 1'b0 ;
  assign n19300 = ( n8301 & ~n14019 ) | ( n8301 & n19250 ) | ( ~n14019 & n19250 ) ;
  assign n19297 = ( x190 & ~n7478 ) | ( x190 & n18770 ) | ( ~n7478 & n18770 ) ;
  assign n19298 = n19297 ^ n9466 ^ n3133 ;
  assign n19299 = n19298 ^ n5338 ^ n5059 ;
  assign n19309 = n19308 ^ n19300 ^ n19299 ;
  assign n19310 = n13822 ^ n12991 ^ 1'b0 ;
  assign n19311 = n5730 | n19310 ;
  assign n19312 = n19311 ^ n13317 ^ 1'b0 ;
  assign n19313 = n9659 ^ n6021 ^ n2299 ;
  assign n19314 = n19313 ^ n5328 ^ 1'b0 ;
  assign n19315 = ~n15899 & n19314 ;
  assign n19316 = ~n4156 & n19315 ;
  assign n19317 = n19316 ^ n16686 ^ n9976 ;
  assign n19318 = n15251 ^ n13112 ^ n9865 ;
  assign n19319 = n16255 ^ x231 ^ 1'b0 ;
  assign n19320 = n1362 | n19319 ;
  assign n19321 = n19320 ^ n2208 ^ 1'b0 ;
  assign n19322 = n2704 ^ n1004 ^ 1'b0 ;
  assign n19323 = ~n1665 & n3320 ;
  assign n19324 = n19323 ^ n2883 ^ 1'b0 ;
  assign n19325 = n16689 ^ n3037 ^ 1'b0 ;
  assign n19326 = ~n16958 & n19325 ;
  assign n19327 = ( ~n10490 & n19324 ) | ( ~n10490 & n19326 ) | ( n19324 & n19326 ) ;
  assign n19328 = x76 & ~n372 ;
  assign n19329 = ~x76 & n19328 ;
  assign n19330 = n782 & ~n1861 ;
  assign n19331 = n19329 & n19330 ;
  assign n19332 = ~n1123 & n19331 ;
  assign n19333 = ( x79 & n1218 ) | ( x79 & n2014 ) | ( n1218 & n2014 ) ;
  assign n19334 = n10300 & n19333 ;
  assign n19335 = n19332 & n19334 ;
  assign n19336 = n5635 ^ n2558 ^ n798 ;
  assign n19337 = ~n19335 & n19336 ;
  assign n19338 = n19335 & n19337 ;
  assign n19339 = n5735 & ~n5928 ;
  assign n19340 = ~n5735 & n19339 ;
  assign n19341 = n19338 | n19340 ;
  assign n19342 = n19338 & ~n19341 ;
  assign n19343 = n2758 & ~n9787 ;
  assign n19344 = ~n2758 & n19343 ;
  assign n19345 = n19342 | n19344 ;
  assign n19346 = n19342 & ~n19345 ;
  assign n19347 = n9732 ^ n4464 ^ n4300 ;
  assign n19348 = n12387 & ~n18304 ;
  assign n19349 = n19347 & n19348 ;
  assign n19350 = n19346 | n19349 ;
  assign n19351 = n19350 ^ n15593 ^ 1'b0 ;
  assign n19352 = n8849 ^ n5753 ^ n2726 ;
  assign n19353 = n17911 ^ n4381 ^ 1'b0 ;
  assign n19354 = n19352 & ~n19353 ;
  assign n19356 = ( x159 & ~n5595 ) | ( x159 & n12491 ) | ( ~n5595 & n12491 ) ;
  assign n19355 = n11766 ^ n9161 ^ 1'b0 ;
  assign n19357 = n19356 ^ n19355 ^ n9086 ;
  assign n19358 = ~n15279 & n19357 ;
  assign n19359 = n12783 | n18664 ;
  assign n19360 = ( n14168 & n15034 ) | ( n14168 & ~n19359 ) | ( n15034 & ~n19359 ) ;
  assign n19362 = n4671 ^ n516 ^ 1'b0 ;
  assign n19363 = ~n1396 & n19362 ;
  assign n19361 = ~n6985 & n12267 ;
  assign n19364 = n19363 ^ n19361 ^ 1'b0 ;
  assign n19365 = n11161 ^ n7689 ^ 1'b0 ;
  assign n19366 = n15683 ^ n5664 ^ n3927 ;
  assign n19367 = n19366 ^ n822 ^ 1'b0 ;
  assign n19368 = n4570 & ~n19367 ;
  assign n19369 = n5954 | n19368 ;
  assign n19370 = n19369 ^ n9102 ^ n2781 ;
  assign n19378 = ~n660 & n4224 ;
  assign n19379 = ( n503 & n18253 ) | ( n503 & ~n19378 ) | ( n18253 & ~n19378 ) ;
  assign n19371 = ( x217 & n2722 ) | ( x217 & n13019 ) | ( n2722 & n13019 ) ;
  assign n19372 = n4110 & n8911 ;
  assign n19373 = n19372 ^ n1735 ^ 1'b0 ;
  assign n19374 = n19373 ^ x189 ^ 1'b0 ;
  assign n19375 = n19371 & ~n19374 ;
  assign n19376 = n19375 ^ n14779 ^ 1'b0 ;
  assign n19377 = ~n1305 & n19376 ;
  assign n19380 = n19379 ^ n19377 ^ 1'b0 ;
  assign n19381 = ~n16836 & n19380 ;
  assign n19382 = n16760 ^ n11387 ^ 1'b0 ;
  assign n19383 = n13966 & n19382 ;
  assign n19384 = n1489 & n4131 ;
  assign n19385 = ~n19383 & n19384 ;
  assign n19386 = ( ~n679 & n1735 ) | ( ~n679 & n14573 ) | ( n1735 & n14573 ) ;
  assign n19387 = n14762 ^ n8579 ^ 1'b0 ;
  assign n19388 = n17595 & ~n19387 ;
  assign n19389 = n1272 | n3299 ;
  assign n19390 = n19389 ^ n10225 ^ 1'b0 ;
  assign n19391 = n10938 ^ n3680 ^ 1'b0 ;
  assign n19392 = n19391 ^ n19223 ^ 1'b0 ;
  assign n19393 = n632 | n19392 ;
  assign n19394 = n19393 ^ n6556 ^ 1'b0 ;
  assign n19395 = ( ~n1321 & n12598 ) | ( ~n1321 & n18717 ) | ( n12598 & n18717 ) ;
  assign n19396 = n4261 & n6381 ;
  assign n19397 = n19396 ^ n9598 ^ 1'b0 ;
  assign n19398 = n19397 ^ n3387 ^ x75 ;
  assign n19399 = n5800 ^ n1998 ^ n1045 ;
  assign n19400 = n15929 & ~n19399 ;
  assign n19402 = n5272 & n8186 ;
  assign n19401 = n732 | n3769 ;
  assign n19403 = n19402 ^ n19401 ^ n1107 ;
  assign n19404 = n6423 ^ n4388 ^ n2517 ;
  assign n19405 = n12333 ^ n10656 ^ 1'b0 ;
  assign n19406 = n19404 | n19405 ;
  assign n19407 = n7034 ^ n2599 ^ n554 ;
  assign n19408 = n19407 ^ n15167 ^ n10450 ;
  assign n19409 = n5264 ^ n3065 ^ n2132 ;
  assign n19410 = n1600 ^ n969 ^ 1'b0 ;
  assign n19411 = n7428 & n19410 ;
  assign n19412 = ( n12338 & ~n19409 ) | ( n12338 & n19411 ) | ( ~n19409 & n19411 ) ;
  assign n19413 = n8008 & n15683 ;
  assign n19414 = n1542 & n19413 ;
  assign n19415 = ( n4183 & n12891 ) | ( n4183 & ~n19414 ) | ( n12891 & ~n19414 ) ;
  assign n19416 = n19415 ^ n8729 ^ 1'b0 ;
  assign n19417 = n12883 ^ n7105 ^ 1'b0 ;
  assign n19418 = ~n6737 & n6889 ;
  assign n19419 = n19418 ^ n8235 ^ 1'b0 ;
  assign n19420 = ( n13160 & ~n19417 ) | ( n13160 & n19419 ) | ( ~n19417 & n19419 ) ;
  assign n19421 = ( ~n3385 & n13729 ) | ( ~n3385 & n19420 ) | ( n13729 & n19420 ) ;
  assign n19422 = ~n8588 & n19421 ;
  assign n19423 = ~n4604 & n19422 ;
  assign n19425 = ( n1219 & n6246 ) | ( n1219 & ~n9767 ) | ( n6246 & ~n9767 ) ;
  assign n19424 = n3790 ^ n544 ^ 1'b0 ;
  assign n19426 = n19425 ^ n19424 ^ n18311 ;
  assign n19427 = n15304 ^ n2236 ^ 1'b0 ;
  assign n19428 = n13967 ^ n3383 ^ 1'b0 ;
  assign n19429 = n8726 ^ n7698 ^ n2947 ;
  assign n19430 = n7226 ^ n6368 ^ 1'b0 ;
  assign n19431 = ~n9900 & n19430 ;
  assign n19432 = ( ~n2210 & n18120 ) | ( ~n2210 & n19431 ) | ( n18120 & n19431 ) ;
  assign n19433 = ( n266 & n19429 ) | ( n266 & n19432 ) | ( n19429 & n19432 ) ;
  assign n19434 = n550 & n4054 ;
  assign n19435 = n8411 ^ x158 ^ 1'b0 ;
  assign n19436 = ( n15068 & n19434 ) | ( n15068 & n19435 ) | ( n19434 & n19435 ) ;
  assign n19440 = n7741 & ~n14129 ;
  assign n19441 = n19440 ^ n7700 ^ 1'b0 ;
  assign n19442 = ~n259 & n19441 ;
  assign n19443 = n19442 ^ n3322 ^ 1'b0 ;
  assign n19437 = n11055 & ~n14249 ;
  assign n19438 = n19437 ^ n18800 ^ 1'b0 ;
  assign n19439 = ~n15570 & n19438 ;
  assign n19444 = n19443 ^ n19439 ^ 1'b0 ;
  assign n19445 = ( n9531 & ~n11946 ) | ( n9531 & n18035 ) | ( ~n11946 & n18035 ) ;
  assign n19446 = ( n2608 & n4455 ) | ( n2608 & n19445 ) | ( n4455 & n19445 ) ;
  assign n19447 = n1475 | n3075 ;
  assign n19448 = n19447 ^ n6495 ^ 1'b0 ;
  assign n19449 = n4240 ^ n890 ^ 1'b0 ;
  assign n19450 = n7334 & n19449 ;
  assign n19451 = n19450 ^ n12793 ^ 1'b0 ;
  assign n19452 = ~n19448 & n19451 ;
  assign n19453 = n18063 ^ n7190 ^ x101 ;
  assign n19454 = ( x3 & n7177 ) | ( x3 & n19453 ) | ( n7177 & n19453 ) ;
  assign n19455 = ~n1052 & n19454 ;
  assign n19456 = n1783 & ~n9321 ;
  assign n19457 = n11391 & ~n19456 ;
  assign n19458 = n13191 & n17376 ;
  assign n19459 = n19458 ^ n3238 ^ 1'b0 ;
  assign n19460 = ~n19457 & n19459 ;
  assign n19461 = n6737 ^ n1372 ^ n284 ;
  assign n19462 = n7135 ^ n362 ^ x97 ;
  assign n19463 = ~n5947 & n11006 ;
  assign n19464 = n938 ^ x20 ^ 1'b0 ;
  assign n19465 = n19464 ^ n5204 ^ n2382 ;
  assign n19466 = n19465 ^ n6878 ^ 1'b0 ;
  assign n19467 = n19463 & n19466 ;
  assign n19468 = ( n19461 & n19462 ) | ( n19461 & ~n19467 ) | ( n19462 & ~n19467 ) ;
  assign n19469 = n14677 ^ n5359 ^ 1'b0 ;
  assign n19470 = n12120 & ~n19469 ;
  assign n19471 = n6155 ^ n5299 ^ 1'b0 ;
  assign n19472 = n19470 & ~n19471 ;
  assign n19473 = ( ~n4434 & n10327 ) | ( ~n4434 & n18178 ) | ( n10327 & n18178 ) ;
  assign n19474 = ( n7664 & n9049 ) | ( n7664 & n19473 ) | ( n9049 & n19473 ) ;
  assign n19475 = n4045 | n19474 ;
  assign n19476 = n12847 ^ n9570 ^ 1'b0 ;
  assign n19477 = ( n11550 & ~n16863 ) | ( n11550 & n19476 ) | ( ~n16863 & n19476 ) ;
  assign n19478 = ( n9289 & n10546 ) | ( n9289 & n18301 ) | ( n10546 & n18301 ) ;
  assign n19479 = n1465 & ~n5754 ;
  assign n19480 = n19479 ^ n9804 ^ 1'b0 ;
  assign n19481 = n6173 ^ n3753 ^ 1'b0 ;
  assign n19482 = ( n19478 & n19480 ) | ( n19478 & n19481 ) | ( n19480 & n19481 ) ;
  assign n19483 = ( n3369 & n6658 ) | ( n3369 & ~n8154 ) | ( n6658 & ~n8154 ) ;
  assign n19484 = ~n13685 & n14539 ;
  assign n19485 = ~n19483 & n19484 ;
  assign n19486 = n19485 ^ n2167 ^ 1'b0 ;
  assign n19487 = n18015 ^ n1601 ^ 1'b0 ;
  assign n19488 = n12767 & n19487 ;
  assign n19489 = n15302 ^ n10174 ^ n7404 ;
  assign n19490 = n15528 ^ n7447 ^ 1'b0 ;
  assign n19491 = n8397 & ~n19490 ;
  assign n19492 = n19311 ^ n4497 ^ 1'b0 ;
  assign n19493 = n14704 ^ n2272 ^ 1'b0 ;
  assign n19494 = n16210 & ~n19493 ;
  assign n19495 = n19492 & n19494 ;
  assign n19496 = n7192 ^ n6205 ^ n5191 ;
  assign n19497 = n19496 ^ n18861 ^ 1'b0 ;
  assign n19498 = n19495 | n19497 ;
  assign n19499 = n2291 ^ n1886 ^ 1'b0 ;
  assign n19500 = n19499 ^ n9916 ^ 1'b0 ;
  assign n19501 = n1630 & n8872 ;
  assign n19502 = n19501 ^ n3665 ^ 1'b0 ;
  assign n19503 = n9585 & ~n19502 ;
  assign n19504 = ~n7026 & n19503 ;
  assign n19505 = n11427 | n19504 ;
  assign n19506 = ~n3816 & n8261 ;
  assign n19507 = ~n9495 & n19506 ;
  assign n19508 = n19507 ^ n8117 ^ 1'b0 ;
  assign n19509 = n19508 ^ n6730 ^ 1'b0 ;
  assign n19510 = n17493 | n19509 ;
  assign n19513 = n17751 ^ n602 ^ 1'b0 ;
  assign n19514 = n1928 & n19513 ;
  assign n19511 = n10186 ^ n8239 ^ n5799 ;
  assign n19512 = n19511 ^ n18776 ^ n15795 ;
  assign n19515 = n19514 ^ n19512 ^ n11849 ;
  assign n19516 = ~n4449 & n10300 ;
  assign n19517 = n8352 & n19516 ;
  assign n19518 = n19517 ^ n18978 ^ 1'b0 ;
  assign n19519 = n13951 ^ n11801 ^ n11024 ;
  assign n19520 = ~n10149 & n19519 ;
  assign n19521 = n13706 ^ n6991 ^ x156 ;
  assign n19522 = n12030 | n19521 ;
  assign n19523 = n11055 ^ n4777 ^ 1'b0 ;
  assign n19524 = n8927 | n19523 ;
  assign n19525 = n19524 ^ n2934 ^ 1'b0 ;
  assign n19526 = n4770 ^ n1879 ^ n374 ;
  assign n19527 = n19526 ^ n12003 ^ n4067 ;
  assign n19528 = ( n13687 & n19525 ) | ( n13687 & n19527 ) | ( n19525 & n19527 ) ;
  assign n19530 = n8541 ^ n6611 ^ 1'b0 ;
  assign n19529 = n1455 | n15657 ;
  assign n19531 = n19530 ^ n19529 ^ 1'b0 ;
  assign n19532 = n6455 & ~n12446 ;
  assign n19533 = ~n19531 & n19532 ;
  assign n19534 = n13464 & ~n15494 ;
  assign n19535 = n12179 ^ n2774 ^ 1'b0 ;
  assign n19536 = n6917 ^ n3148 ^ 1'b0 ;
  assign n19537 = n2229 & ~n19536 ;
  assign n19538 = n19537 ^ n18770 ^ n8822 ;
  assign n19539 = n9366 ^ n4874 ^ 1'b0 ;
  assign n19540 = ( n5012 & n12485 ) | ( n5012 & n19539 ) | ( n12485 & n19539 ) ;
  assign n19541 = n7930 & ~n19540 ;
  assign n19542 = n17952 | n19541 ;
  assign n19543 = n19542 ^ n5823 ^ 1'b0 ;
  assign n19544 = n7941 ^ n1638 ^ 1'b0 ;
  assign n19545 = n5042 | n19544 ;
  assign n19546 = n1278 | n14051 ;
  assign n19547 = n5953 | n19546 ;
  assign n19548 = n6889 & n13213 ;
  assign n19549 = ~n19547 & n19548 ;
  assign n19550 = n2394 | n19549 ;
  assign n19551 = n13927 | n19550 ;
  assign n19552 = n8042 & ~n13600 ;
  assign n19553 = n19552 ^ n4417 ^ 1'b0 ;
  assign n19554 = ( n7983 & ~n10850 ) | ( n7983 & n19553 ) | ( ~n10850 & n19553 ) ;
  assign n19555 = n3448 & n15274 ;
  assign n19556 = n19555 ^ n644 ^ 1'b0 ;
  assign n19557 = ( n6531 & n11179 ) | ( n6531 & ~n19556 ) | ( n11179 & ~n19556 ) ;
  assign n19558 = n12887 & n15822 ;
  assign n19559 = n19209 ^ n10080 ^ 1'b0 ;
  assign n19560 = ~n10096 & n19559 ;
  assign n19561 = n19560 ^ n14853 ^ n9492 ;
  assign n19562 = n3452 ^ n3292 ^ n2427 ;
  assign n19563 = n19278 ^ n12121 ^ 1'b0 ;
  assign n19564 = n5990 & ~n19563 ;
  assign n19565 = n7878 ^ n4823 ^ 1'b0 ;
  assign n19566 = n13125 | n15850 ;
  assign n19567 = ( n13589 & ~n19565 ) | ( n13589 & n19566 ) | ( ~n19565 & n19566 ) ;
  assign n19572 = n7191 ^ n4761 ^ 1'b0 ;
  assign n19573 = n18629 | n19572 ;
  assign n19568 = n5373 & n7050 ;
  assign n19569 = ~n14658 & n19568 ;
  assign n19570 = n19569 ^ n2683 ^ 1'b0 ;
  assign n19571 = n5687 & n19570 ;
  assign n19574 = n19573 ^ n19571 ^ x154 ;
  assign n19575 = n5329 ^ n2406 ^ 1'b0 ;
  assign n19576 = n9332 | n19575 ;
  assign n19577 = n9093 | n19576 ;
  assign n19578 = ~n12500 & n18916 ;
  assign n19579 = n860 ^ n631 ^ n264 ;
  assign n19580 = n19579 ^ n16008 ^ n14818 ;
  assign n19581 = n19580 ^ n8896 ^ 1'b0 ;
  assign n19582 = n10387 | n16195 ;
  assign n19583 = n15693 ^ n5686 ^ 1'b0 ;
  assign n19584 = n19583 ^ n2156 ^ 1'b0 ;
  assign n19585 = n277 & ~n8919 ;
  assign n19586 = ~n13111 & n19585 ;
  assign n19587 = ( n4769 & n9174 ) | ( n4769 & n10860 ) | ( n9174 & n10860 ) ;
  assign n19588 = ~n13518 & n19587 ;
  assign n19589 = n19588 ^ n3305 ^ 1'b0 ;
  assign n19590 = n12917 | n18624 ;
  assign n19591 = n1719 | n7779 ;
  assign n19592 = n19591 ^ n19163 ^ 1'b0 ;
  assign n19593 = n18003 | n19592 ;
  assign n19594 = n6361 ^ n2995 ^ 1'b0 ;
  assign n19595 = ~n735 & n1876 ;
  assign n19596 = n19595 ^ n11150 ^ n2502 ;
  assign n19598 = n4912 ^ n3520 ^ 1'b0 ;
  assign n19597 = n10976 & ~n12384 ;
  assign n19599 = n19598 ^ n19597 ^ 1'b0 ;
  assign n19600 = n8858 | n10325 ;
  assign n19601 = n7173 | n19600 ;
  assign n19602 = ~n2502 & n6129 ;
  assign n19603 = n19602 ^ n11587 ^ 1'b0 ;
  assign n19604 = n19601 & n19603 ;
  assign n19605 = n19604 ^ n16222 ^ n6390 ;
  assign n19606 = n5866 ^ n4419 ^ n1029 ;
  assign n19607 = ( n4893 & n13899 ) | ( n4893 & n19606 ) | ( n13899 & n19606 ) ;
  assign n19608 = n19605 & ~n19607 ;
  assign n19618 = n13040 ^ n12426 ^ 1'b0 ;
  assign n19619 = n1566 & ~n19618 ;
  assign n19609 = n4030 ^ n3996 ^ 1'b0 ;
  assign n19610 = ( n1385 & n10239 ) | ( n1385 & n19609 ) | ( n10239 & n19609 ) ;
  assign n19611 = n1037 & ~n19610 ;
  assign n19612 = n19611 ^ n12393 ^ 1'b0 ;
  assign n19614 = ~n6586 & n12333 ;
  assign n19613 = n8063 & n13056 ;
  assign n19615 = n19614 ^ n19613 ^ 1'b0 ;
  assign n19616 = n19615 ^ n14794 ^ x212 ;
  assign n19617 = ( ~n11165 & n19612 ) | ( ~n11165 & n19616 ) | ( n19612 & n19616 ) ;
  assign n19620 = n19619 ^ n19617 ^ n15152 ;
  assign n19622 = n10454 & ~n16831 ;
  assign n19623 = ~n7919 & n19622 ;
  assign n19621 = n4021 & n7565 ;
  assign n19624 = n19623 ^ n19621 ^ 1'b0 ;
  assign n19625 = n868 | n8802 ;
  assign n19626 = n19625 ^ n14307 ^ 1'b0 ;
  assign n19627 = n18337 ^ n15112 ^ 1'b0 ;
  assign n19632 = n6270 ^ n3088 ^ 1'b0 ;
  assign n19628 = ( n426 & n643 ) | ( n426 & n1554 ) | ( n643 & n1554 ) ;
  assign n19629 = n6022 ^ n5751 ^ 1'b0 ;
  assign n19630 = ( n15712 & n16228 ) | ( n15712 & ~n19629 ) | ( n16228 & ~n19629 ) ;
  assign n19631 = n19628 & n19630 ;
  assign n19633 = n19632 ^ n19631 ^ 1'b0 ;
  assign n19634 = n14296 ^ n7968 ^ n7060 ;
  assign n19635 = n19634 ^ n2925 ^ n1272 ;
  assign n19636 = ( n7576 & ~n19633 ) | ( n7576 & n19635 ) | ( ~n19633 & n19635 ) ;
  assign n19638 = n7748 ^ n2042 ^ 1'b0 ;
  assign n19639 = n5064 & ~n19638 ;
  assign n19637 = ~n10615 & n13822 ;
  assign n19640 = n19639 ^ n19637 ^ 1'b0 ;
  assign n19641 = n13910 & ~n19640 ;
  assign n19642 = ~n6269 & n19641 ;
  assign n19643 = ( ~n2536 & n9137 ) | ( ~n2536 & n19642 ) | ( n9137 & n19642 ) ;
  assign n19644 = n9417 ^ n3639 ^ 1'b0 ;
  assign n19645 = n19643 | n19644 ;
  assign n19646 = ( n10406 & n12767 ) | ( n10406 & ~n19645 ) | ( n12767 & ~n19645 ) ;
  assign n19651 = ~n1452 & n3369 ;
  assign n19650 = ( n879 & n1345 ) | ( n879 & ~n5965 ) | ( n1345 & ~n5965 ) ;
  assign n19652 = n19651 ^ n19650 ^ 1'b0 ;
  assign n19653 = n9056 | n19652 ;
  assign n19654 = n19653 ^ n9293 ^ 1'b0 ;
  assign n19655 = n14899 & ~n19654 ;
  assign n19647 = n2374 ^ n1635 ^ n633 ;
  assign n19648 = ( ~n789 & n17199 ) | ( ~n789 & n19647 ) | ( n17199 & n19647 ) ;
  assign n19649 = n19648 ^ n11725 ^ 1'b0 ;
  assign n19656 = n19655 ^ n19649 ^ n13848 ;
  assign n19657 = n8834 ^ n6037 ^ n605 ;
  assign n19658 = n19657 ^ n15787 ^ 1'b0 ;
  assign n19659 = n14627 & ~n19658 ;
  assign n19660 = n19659 ^ n12418 ^ 1'b0 ;
  assign n19661 = n19660 ^ n18881 ^ 1'b0 ;
  assign n19662 = n19656 & n19661 ;
  assign n19663 = n19545 ^ n15175 ^ n7786 ;
  assign n19664 = n765 & n2793 ;
  assign n19665 = n19664 ^ n7981 ^ n1513 ;
  assign n19666 = ( x170 & n17057 ) | ( x170 & n19665 ) | ( n17057 & n19665 ) ;
  assign n19667 = n19666 ^ n17647 ^ n14147 ;
  assign n19668 = ~n4223 & n15224 ;
  assign n19669 = n16838 ^ n604 ^ 1'b0 ;
  assign n19670 = n4866 | n19669 ;
  assign n19674 = n8497 ^ n6648 ^ n5027 ;
  assign n19675 = ( n13942 & n14954 ) | ( n13942 & n19674 ) | ( n14954 & n19674 ) ;
  assign n19671 = n1684 ^ n1511 ^ 1'b0 ;
  assign n19672 = n5532 | n19671 ;
  assign n19673 = n12215 & ~n19672 ;
  assign n19676 = n19675 ^ n19673 ^ n5405 ;
  assign n19677 = n6349 & n9931 ;
  assign n19678 = n845 | n7238 ;
  assign n19679 = n19677 & ~n19678 ;
  assign n19680 = ( n4789 & n5196 ) | ( n4789 & ~n19679 ) | ( n5196 & ~n19679 ) ;
  assign n19681 = n16056 & ~n19680 ;
  assign n19682 = n18071 ^ n13046 ^ n11378 ;
  assign n19683 = ~n867 & n1360 ;
  assign n19684 = n8970 & n19683 ;
  assign n19685 = x194 & n7897 ;
  assign n19686 = n19685 ^ n10377 ^ 1'b0 ;
  assign n19687 = n3828 & ~n19686 ;
  assign n19691 = ~n6912 & n18828 ;
  assign n19688 = ~n3970 & n14396 ;
  assign n19689 = n19688 ^ n17006 ^ n1438 ;
  assign n19690 = n12343 | n19689 ;
  assign n19692 = n19691 ^ n19690 ^ 1'b0 ;
  assign n19693 = n15308 ^ n9708 ^ 1'b0 ;
  assign n19694 = n19692 & ~n19693 ;
  assign n19695 = n10694 ^ n3828 ^ n3499 ;
  assign n19696 = ( n6683 & n11612 ) | ( n6683 & n19695 ) | ( n11612 & n19695 ) ;
  assign n19697 = n11498 ^ n5880 ^ 1'b0 ;
  assign n19698 = ~n18887 & n19697 ;
  assign n19699 = n7540 ^ n1455 ^ 1'b0 ;
  assign n19700 = ( n15688 & n17386 ) | ( n15688 & n19699 ) | ( n17386 & n19699 ) ;
  assign n19701 = n7192 | n13614 ;
  assign n19702 = n8873 | n19701 ;
  assign n19703 = n19702 ^ n8343 ^ 1'b0 ;
  assign n19704 = ( ~n676 & n4097 ) | ( ~n676 & n19703 ) | ( n4097 & n19703 ) ;
  assign n19705 = n19704 ^ n10179 ^ 1'b0 ;
  assign n19706 = ~n4531 & n19705 ;
  assign n19707 = n19706 ^ n14595 ^ 1'b0 ;
  assign n19708 = ( ~n1106 & n3091 ) | ( ~n1106 & n12910 ) | ( n3091 & n12910 ) ;
  assign n19709 = ( n8915 & ~n13175 ) | ( n8915 & n19708 ) | ( ~n13175 & n19708 ) ;
  assign n19710 = n19709 ^ n14958 ^ x198 ;
  assign n19711 = n12835 ^ n10268 ^ x144 ;
  assign n19712 = n19711 ^ n10138 ^ 1'b0 ;
  assign n19713 = n10030 ^ n496 ^ 1'b0 ;
  assign n19714 = n19712 & ~n19713 ;
  assign n19716 = n6249 & ~n11287 ;
  assign n19717 = n16377 & ~n19595 ;
  assign n19718 = ~n3962 & n19717 ;
  assign n19719 = n4558 ^ n1175 ^ 1'b0 ;
  assign n19720 = ~n3892 & n19719 ;
  assign n19721 = n19718 & n19720 ;
  assign n19722 = n19716 & ~n19721 ;
  assign n19715 = n4300 & n16468 ;
  assign n19723 = n19722 ^ n19715 ^ 1'b0 ;
  assign n19724 = n8145 ^ n6657 ^ n2113 ;
  assign n19725 = n19724 ^ n2575 ^ n600 ;
  assign n19726 = n9758 | n12029 ;
  assign n19727 = n9073 | n19726 ;
  assign n19728 = n19725 & ~n19727 ;
  assign n19729 = n7697 ^ n4329 ^ n1859 ;
  assign n19730 = n5395 & n19729 ;
  assign n19731 = n19730 ^ n12837 ^ 1'b0 ;
  assign n19732 = n4506 & n19731 ;
  assign n19733 = n19732 ^ n9882 ^ 1'b0 ;
  assign n19734 = n19733 ^ n3843 ^ n2519 ;
  assign n19735 = n10961 ^ n3973 ^ 1'b0 ;
  assign n19736 = n10163 & n19735 ;
  assign n19737 = ~n5061 & n14896 ;
  assign n19738 = ~n1706 & n19737 ;
  assign n19739 = n19738 ^ n5372 ^ n3172 ;
  assign n19740 = ( n17971 & n19736 ) | ( n17971 & n19739 ) | ( n19736 & n19739 ) ;
  assign n19741 = n15686 | n19740 ;
  assign n19742 = n4249 & n8219 ;
  assign n19743 = n19742 ^ n337 ^ 1'b0 ;
  assign n19744 = n3101 | n19743 ;
  assign n19745 = n13055 | n18796 ;
  assign n19746 = n19261 ^ n3186 ^ 1'b0 ;
  assign n19747 = n11174 & n19746 ;
  assign n19748 = ~n5649 & n18979 ;
  assign n19749 = n8219 & ~n10722 ;
  assign n19750 = n19749 ^ n13534 ^ 1'b0 ;
  assign n19751 = n19750 ^ n9767 ^ n1735 ;
  assign n19752 = n11859 & ~n15842 ;
  assign n19753 = ( n6897 & ~n16423 ) | ( n6897 & n19752 ) | ( ~n16423 & n19752 ) ;
  assign n19754 = n13616 ^ n7421 ^ 1'b0 ;
  assign n19755 = n9328 | n9463 ;
  assign n19756 = n19755 ^ n3116 ^ 1'b0 ;
  assign n19757 = n19756 ^ n11024 ^ 1'b0 ;
  assign n19761 = ~n2965 & n12406 ;
  assign n19762 = ~n9162 & n19761 ;
  assign n19763 = ~n8947 & n19762 ;
  assign n19758 = n6173 | n10165 ;
  assign n19759 = n10599 | n13554 ;
  assign n19760 = ( n6421 & n19758 ) | ( n6421 & n19759 ) | ( n19758 & n19759 ) ;
  assign n19764 = n19763 ^ n19760 ^ n8768 ;
  assign n19766 = n10456 ^ n5322 ^ 1'b0 ;
  assign n19767 = n1039 | n19766 ;
  assign n19765 = n16378 ^ n5896 ^ 1'b0 ;
  assign n19768 = n19767 ^ n19765 ^ n3260 ;
  assign n19769 = n12155 ^ n11498 ^ n1414 ;
  assign n19770 = n16818 ^ n10509 ^ 1'b0 ;
  assign n19771 = n19499 & ~n19770 ;
  assign n19772 = n14053 & n19771 ;
  assign n19773 = n2052 & n2335 ;
  assign n19774 = n2872 | n19773 ;
  assign n19775 = n2405 & ~n19774 ;
  assign n19776 = n19775 ^ n19012 ^ 1'b0 ;
  assign n19777 = n556 | n9258 ;
  assign n19778 = n7555 ^ n7029 ^ 1'b0 ;
  assign n19779 = ( n2749 & n2994 ) | ( n2749 & ~n19778 ) | ( n2994 & ~n19778 ) ;
  assign n19780 = ~n13431 & n19779 ;
  assign n19781 = n19780 ^ n6776 ^ 1'b0 ;
  assign n19786 = ( x64 & ~x101 ) | ( x64 & n7049 ) | ( ~x101 & n7049 ) ;
  assign n19782 = n11698 ^ n6804 ^ 1'b0 ;
  assign n19783 = n15208 & n19782 ;
  assign n19784 = n19783 ^ n14461 ^ 1'b0 ;
  assign n19785 = n508 & ~n19784 ;
  assign n19787 = n19786 ^ n19785 ^ n8731 ;
  assign n19788 = ( ~n6475 & n12381 ) | ( ~n6475 & n16618 ) | ( n12381 & n16618 ) ;
  assign n19789 = n1834 | n5513 ;
  assign n19790 = n19789 ^ n5454 ^ 1'b0 ;
  assign n19791 = n19790 ^ n9148 ^ 1'b0 ;
  assign n19792 = n17681 ^ n13262 ^ 1'b0 ;
  assign n19793 = n3883 ^ n3553 ^ 1'b0 ;
  assign n19794 = n19793 ^ n2247 ^ 1'b0 ;
  assign n19795 = n17631 & ~n19794 ;
  assign n19796 = ( n15375 & n19656 ) | ( n15375 & n19795 ) | ( n19656 & n19795 ) ;
  assign n19797 = n6716 ^ n3462 ^ 1'b0 ;
  assign n19798 = ( ~n9852 & n10895 ) | ( ~n9852 & n19797 ) | ( n10895 & n19797 ) ;
  assign n19799 = n1717 | n13248 ;
  assign n19800 = ~n1932 & n13589 ;
  assign n19801 = ~n19799 & n19800 ;
  assign n19802 = ( ~n15163 & n18709 ) | ( ~n15163 & n19801 ) | ( n18709 & n19801 ) ;
  assign n19803 = n17796 ^ n10416 ^ n6500 ;
  assign n19804 = n7643 | n11486 ;
  assign n19805 = n9347 & ~n19804 ;
  assign n19806 = n1654 ^ n1367 ^ n938 ;
  assign n19807 = n19806 ^ n8971 ^ 1'b0 ;
  assign n19808 = ~n19805 & n19807 ;
  assign n19809 = n9807 ^ n2887 ^ 1'b0 ;
  assign n19810 = n17854 & ~n19809 ;
  assign n19811 = ~n5615 & n8717 ;
  assign n19812 = n19811 ^ n1367 ^ 1'b0 ;
  assign n19813 = n19810 & n19812 ;
  assign n19814 = n477 & ~n19813 ;
  assign n19815 = ~n1442 & n1603 ;
  assign n19816 = ( n1206 & n8209 ) | ( n1206 & ~n15842 ) | ( n8209 & ~n15842 ) ;
  assign n19817 = ~n583 & n14197 ;
  assign n19818 = ~n19816 & n19817 ;
  assign n19819 = n19818 ^ n6178 ^ n3071 ;
  assign n19820 = ( n19814 & n19815 ) | ( n19814 & ~n19819 ) | ( n19815 & ~n19819 ) ;
  assign n19822 = ( n2760 & n6317 ) | ( n2760 & ~n13704 ) | ( n6317 & ~n13704 ) ;
  assign n19821 = n2930 | n13118 ;
  assign n19823 = n19822 ^ n19821 ^ 1'b0 ;
  assign n19824 = ( ~x34 & n2574 ) | ( ~x34 & n11715 ) | ( n2574 & n11715 ) ;
  assign n19825 = n10911 | n19824 ;
  assign n19826 = n6580 ^ n5907 ^ 1'b0 ;
  assign n19827 = ~n18942 & n19826 ;
  assign n19828 = ~n18201 & n19827 ;
  assign n19829 = n916 ^ x176 ^ 1'b0 ;
  assign n19830 = n19829 ^ n5197 ^ n2191 ;
  assign n19831 = n10155 ^ n4285 ^ n389 ;
  assign n19832 = n19831 ^ n13342 ^ n6543 ;
  assign n19833 = ~n272 & n1798 ;
  assign n19834 = ~n2083 & n19833 ;
  assign n19835 = ( n2927 & ~n2965 ) | ( n2927 & n19834 ) | ( ~n2965 & n19834 ) ;
  assign n19836 = n19835 ^ n2986 ^ 1'b0 ;
  assign n19837 = ( ~n8503 & n19266 ) | ( ~n8503 & n19836 ) | ( n19266 & n19836 ) ;
  assign n19838 = n14565 & ~n19837 ;
  assign n19839 = n7105 & ~n16199 ;
  assign n19840 = n11150 & n19839 ;
  assign n19841 = n19840 ^ n19030 ^ 1'b0 ;
  assign n19842 = ~n7748 & n11009 ;
  assign n19843 = n13554 & n19842 ;
  assign n19846 = ~n2258 & n12280 ;
  assign n19847 = n19846 ^ n8398 ^ 1'b0 ;
  assign n19848 = n7838 ^ n5641 ^ 1'b0 ;
  assign n19849 = ( n5222 & n19847 ) | ( n5222 & ~n19848 ) | ( n19847 & ~n19848 ) ;
  assign n19850 = n19849 ^ n12083 ^ 1'b0 ;
  assign n19851 = n2803 & n19850 ;
  assign n19844 = n19233 ^ n13030 ^ 1'b0 ;
  assign n19845 = n19844 ^ n3596 ^ n2376 ;
  assign n19852 = n19851 ^ n19845 ^ n4536 ;
  assign n19853 = n11987 ^ n5171 ^ n3395 ;
  assign n19854 = n19853 ^ n16686 ^ 1'b0 ;
  assign n19855 = n1814 | n19854 ;
  assign n19856 = n1878 | n4588 ;
  assign n19857 = n2971 & ~n3577 ;
  assign n19858 = ( n2692 & n9905 ) | ( n2692 & n11343 ) | ( n9905 & n11343 ) ;
  assign n19859 = ( n17232 & ~n19857 ) | ( n17232 & n19858 ) | ( ~n19857 & n19858 ) ;
  assign n19860 = ( n10450 & n14172 ) | ( n10450 & n19859 ) | ( n14172 & n19859 ) ;
  assign n19861 = n19860 ^ n9758 ^ 1'b0 ;
  assign n19863 = n2134 & ~n4837 ;
  assign n19862 = n16701 ^ n6178 ^ 1'b0 ;
  assign n19864 = n19863 ^ n19862 ^ 1'b0 ;
  assign n19865 = n8357 | n12130 ;
  assign n19866 = n6071 ^ n5513 ^ 1'b0 ;
  assign n19867 = n16156 | n19866 ;
  assign n19868 = n19867 ^ n15315 ^ n6449 ;
  assign n19869 = n12794 & n19868 ;
  assign n19870 = ~n17245 & n19869 ;
  assign n19871 = n19870 ^ n13851 ^ n9701 ;
  assign n19872 = n19871 ^ n5201 ^ n3585 ;
  assign n19873 = ( n8564 & n19865 ) | ( n8564 & n19872 ) | ( n19865 & n19872 ) ;
  assign n19874 = n11318 ^ n890 ^ x223 ;
  assign n19875 = ( n1908 & ~n7308 ) | ( n1908 & n19874 ) | ( ~n7308 & n19874 ) ;
  assign n19876 = n19875 ^ n2850 ^ n594 ;
  assign n19877 = n1415 & ~n8493 ;
  assign n19878 = n16565 ^ n3365 ^ 1'b0 ;
  assign n19879 = n4989 | n19878 ;
  assign n19880 = n19877 & ~n19879 ;
  assign n19881 = n10337 & n19880 ;
  assign n19882 = n19881 ^ n7044 ^ 1'b0 ;
  assign n19883 = n13891 ^ n7449 ^ 1'b0 ;
  assign n19884 = ~n3906 & n19883 ;
  assign n19885 = n466 & n19884 ;
  assign n19886 = ~n19882 & n19885 ;
  assign n19887 = n16605 ^ n6212 ^ n5968 ;
  assign n19888 = ( ~n700 & n12586 ) | ( ~n700 & n19887 ) | ( n12586 & n19887 ) ;
  assign n19889 = n12298 & ~n19888 ;
  assign n19890 = n15558 ^ n4427 ^ 1'b0 ;
  assign n19891 = n8554 & ~n19890 ;
  assign n19892 = n19891 ^ n12114 ^ 1'b0 ;
  assign n19893 = ~n4141 & n19892 ;
  assign n19894 = n19893 ^ n2194 ^ 1'b0 ;
  assign n19896 = ( n758 & n3322 ) | ( n758 & ~n10997 ) | ( n3322 & ~n10997 ) ;
  assign n19895 = n10615 ^ n8215 ^ n3352 ;
  assign n19897 = n19896 ^ n19895 ^ n6527 ;
  assign n19898 = n9581 ^ n9240 ^ 1'b0 ;
  assign n19899 = n963 | n10281 ;
  assign n19900 = n19899 ^ n19716 ^ 1'b0 ;
  assign n19901 = n19900 ^ n18291 ^ n849 ;
  assign n19902 = n13178 ^ n12157 ^ 1'b0 ;
  assign n19903 = ( n15696 & ~n16930 ) | ( n15696 & n19902 ) | ( ~n16930 & n19902 ) ;
  assign n19904 = ( n736 & ~n8169 ) | ( n736 & n12125 ) | ( ~n8169 & n12125 ) ;
  assign n19905 = n6798 ^ n3193 ^ n534 ;
  assign n19906 = ~n3432 & n19905 ;
  assign n19907 = n17710 & n19906 ;
  assign n19909 = n3483 & n9904 ;
  assign n19910 = ~n3348 & n19909 ;
  assign n19911 = n19910 ^ n5669 ^ n2916 ;
  assign n19908 = n14891 | n17971 ;
  assign n19912 = n19911 ^ n19908 ^ 1'b0 ;
  assign n19913 = n15491 ^ n10701 ^ 1'b0 ;
  assign n19914 = ( n10249 & n17585 ) | ( n10249 & n19913 ) | ( n17585 & n19913 ) ;
  assign n19915 = n8279 ^ n4997 ^ 1'b0 ;
  assign n19916 = n18090 ^ n11048 ^ n10851 ;
  assign n19917 = n16468 ^ n14776 ^ n4567 ;
  assign n19918 = ( n17979 & n18531 ) | ( n17979 & n19352 ) | ( n18531 & n19352 ) ;
  assign n19919 = n12357 & ~n19918 ;
  assign n19920 = ~n19917 & n19919 ;
  assign n19921 = ~n4060 & n11858 ;
  assign n19922 = ~n3362 & n19921 ;
  assign n19923 = n9360 ^ n5868 ^ 1'b0 ;
  assign n19924 = ( n3465 & ~n7837 ) | ( n3465 & n10786 ) | ( ~n7837 & n10786 ) ;
  assign n19925 = ( ~n809 & n8595 ) | ( ~n809 & n19924 ) | ( n8595 & n19924 ) ;
  assign n19926 = n7349 & ~n10772 ;
  assign n19927 = n19925 | n19926 ;
  assign n19928 = n5380 | n10672 ;
  assign n19929 = n19928 ^ n8612 ^ n6530 ;
  assign n19930 = ~n4634 & n12826 ;
  assign n19931 = n19930 ^ n13616 ^ n9972 ;
  assign n19932 = n4977 & ~n19931 ;
  assign n19933 = n19932 ^ n2945 ^ 1'b0 ;
  assign n19934 = n19929 & n19933 ;
  assign n19935 = ~n14969 & n19934 ;
  assign n19937 = n8930 ^ n7732 ^ n2013 ;
  assign n19936 = n5322 | n15390 ;
  assign n19938 = n19937 ^ n19936 ^ 1'b0 ;
  assign n19939 = x156 | n1317 ;
  assign n19940 = n19939 ^ n6475 ^ 1'b0 ;
  assign n19941 = n642 | n12170 ;
  assign n19942 = n19940 | n19941 ;
  assign n19943 = ~n9342 & n19942 ;
  assign n19944 = n13312 & n19943 ;
  assign n19945 = ~n5979 & n9347 ;
  assign n19946 = n2363 | n19945 ;
  assign n19947 = n2211 | n19946 ;
  assign n19948 = n8008 & n12665 ;
  assign n19950 = n11632 ^ n6566 ^ 1'b0 ;
  assign n19951 = n19950 ^ n14270 ^ n9551 ;
  assign n19952 = n7327 | n19951 ;
  assign n19953 = n19952 ^ n3906 ^ 1'b0 ;
  assign n19949 = n5085 & n17671 ;
  assign n19954 = n19953 ^ n19949 ^ 1'b0 ;
  assign n19955 = ~n2117 & n15796 ;
  assign n19956 = n19955 ^ n7107 ^ 1'b0 ;
  assign n19957 = n19956 ^ n17737 ^ 1'b0 ;
  assign n19958 = ( n5990 & n7761 ) | ( n5990 & ~n19957 ) | ( n7761 & ~n19957 ) ;
  assign n19959 = n6664 ^ n2668 ^ n2036 ;
  assign n19960 = ( n4997 & n11212 ) | ( n4997 & ~n19959 ) | ( n11212 & ~n19959 ) ;
  assign n19961 = ( n937 & n1666 ) | ( n937 & n5090 ) | ( n1666 & n5090 ) ;
  assign n19962 = ( n10654 & ~n14717 ) | ( n10654 & n19961 ) | ( ~n14717 & n19961 ) ;
  assign n19963 = ( x71 & n3456 ) | ( x71 & ~n7484 ) | ( n3456 & ~n7484 ) ;
  assign n19964 = n19963 ^ n4521 ^ 1'b0 ;
  assign n19965 = n693 | n2582 ;
  assign n19966 = ( n1806 & ~n7181 ) | ( n1806 & n19965 ) | ( ~n7181 & n19965 ) ;
  assign n19967 = n6466 | n19966 ;
  assign n19968 = n19967 ^ n12444 ^ n5992 ;
  assign n19969 = n19968 ^ n2595 ^ 1'b0 ;
  assign n19970 = ~n17226 & n19969 ;
  assign n19972 = n2792 ^ n980 ^ 1'b0 ;
  assign n19973 = n8092 & n19972 ;
  assign n19971 = n8557 & ~n13787 ;
  assign n19974 = n19973 ^ n19971 ^ 1'b0 ;
  assign n19975 = ( ~n10391 & n10789 ) | ( ~n10391 & n19974 ) | ( n10789 & n19974 ) ;
  assign n19976 = ( n10951 & n16413 ) | ( n10951 & ~n19105 ) | ( n16413 & ~n19105 ) ;
  assign n19977 = n11789 & n19976 ;
  assign n19978 = ( n2822 & n2958 ) | ( n2822 & ~n4247 ) | ( n2958 & ~n4247 ) ;
  assign n19979 = n19978 ^ n11231 ^ 1'b0 ;
  assign n19980 = n7812 | n19979 ;
  assign n19981 = ( ~x111 & x215 ) | ( ~x111 & n19980 ) | ( x215 & n19980 ) ;
  assign n19982 = n8201 & n19981 ;
  assign n19983 = n10533 ^ n598 ^ 1'b0 ;
  assign n19984 = n16412 ^ n3535 ^ 1'b0 ;
  assign n19985 = ( n7507 & n19983 ) | ( n7507 & ~n19984 ) | ( n19983 & ~n19984 ) ;
  assign n19986 = n11058 | n19985 ;
  assign n19987 = n19986 ^ n13593 ^ 1'b0 ;
  assign n19988 = n11427 & ~n18028 ;
  assign n19989 = n19988 ^ x10 ^ 1'b0 ;
  assign n19990 = n4652 | n19989 ;
  assign n19991 = n15194 & ~n19184 ;
  assign n19992 = ~n19990 & n19991 ;
  assign n19993 = ( n937 & ~n11253 ) | ( n937 & n16997 ) | ( ~n11253 & n16997 ) ;
  assign n19994 = n11286 ^ n2197 ^ n1524 ;
  assign n19995 = ( n19959 & n19993 ) | ( n19959 & n19994 ) | ( n19993 & n19994 ) ;
  assign n19996 = n17474 | n19992 ;
  assign n19997 = n15321 ^ n9876 ^ 1'b0 ;
  assign n19998 = n9589 & ~n19997 ;
  assign n19999 = n4196 ^ n3071 ^ n1662 ;
  assign n20000 = n14675 & ~n19999 ;
  assign n20001 = n20000 ^ n14725 ^ 1'b0 ;
  assign n20002 = n20001 ^ n13970 ^ 1'b0 ;
  assign n20003 = n8159 & ~n20002 ;
  assign n20004 = n5649 | n7061 ;
  assign n20005 = n5027 & ~n20004 ;
  assign n20006 = n13915 | n20005 ;
  assign n20007 = n5891 & ~n20006 ;
  assign n20008 = n1108 & ~n20007 ;
  assign n20009 = n20008 ^ n7540 ^ 1'b0 ;
  assign n20010 = n19359 ^ n18725 ^ n5413 ;
  assign n20011 = n17412 ^ n2864 ^ 1'b0 ;
  assign n20012 = n19270 & ~n20011 ;
  assign n20013 = ~n15842 & n20012 ;
  assign n20014 = n10280 & n20013 ;
  assign n20015 = ( n8854 & n9150 ) | ( n8854 & ~n19303 ) | ( n9150 & ~n19303 ) ;
  assign n20016 = n20015 ^ n12586 ^ 1'b0 ;
  assign n20017 = n7113 ^ n5372 ^ n262 ;
  assign n20018 = ( n3955 & ~n5447 ) | ( n3955 & n19146 ) | ( ~n5447 & n19146 ) ;
  assign n20019 = n11730 & ~n20018 ;
  assign n20020 = n20017 & ~n20019 ;
  assign n20021 = ( n5571 & n10228 ) | ( n5571 & n10973 ) | ( n10228 & n10973 ) ;
  assign n20022 = n12480 | n15816 ;
  assign n20023 = n20021 | n20022 ;
  assign n20024 = n20023 ^ n5942 ^ 1'b0 ;
  assign n20025 = n5639 & n15510 ;
  assign n20026 = ( x74 & x82 ) | ( x74 & ~n3813 ) | ( x82 & ~n3813 ) ;
  assign n20027 = n2989 & ~n3009 ;
  assign n20028 = n20026 & n20027 ;
  assign n20029 = n8677 | n20028 ;
  assign n20030 = n18187 ^ n12599 ^ 1'b0 ;
  assign n20031 = n14297 | n20030 ;
  assign n20032 = n10448 ^ n6739 ^ n1037 ;
  assign n20033 = n20032 ^ n6081 ^ 1'b0 ;
  assign n20034 = n6130 & n20033 ;
  assign n20035 = n5774 | n8294 ;
  assign n20036 = x44 & n20035 ;
  assign n20037 = n2039 ^ n293 ^ 1'b0 ;
  assign n20038 = n3516 & ~n20037 ;
  assign n20039 = n15084 & n20038 ;
  assign n20040 = ~n8549 & n10556 ;
  assign n20041 = n20040 ^ n9314 ^ 1'b0 ;
  assign n20042 = ( n5733 & n10557 ) | ( n5733 & n12033 ) | ( n10557 & n12033 ) ;
  assign n20043 = ( ~n432 & n20041 ) | ( ~n432 & n20042 ) | ( n20041 & n20042 ) ;
  assign n20044 = n13317 & ~n13950 ;
  assign n20045 = n16034 & n20044 ;
  assign n20046 = n884 & ~n5568 ;
  assign n20047 = n20046 ^ n14575 ^ n1877 ;
  assign n20048 = ~n16763 & n20047 ;
  assign n20049 = n20048 ^ n19419 ^ 1'b0 ;
  assign n20050 = ( ~n3052 & n7367 ) | ( ~n3052 & n19675 ) | ( n7367 & n19675 ) ;
  assign n20051 = n8977 | n20050 ;
  assign n20052 = n15333 | n16126 ;
  assign n20053 = n18921 ^ n6658 ^ 1'b0 ;
  assign n20054 = n814 | n20053 ;
  assign n20055 = n20054 ^ n12033 ^ 1'b0 ;
  assign n20056 = n4763 & ~n20055 ;
  assign n20057 = ~n13932 & n20056 ;
  assign n20058 = ( ~n9451 & n18304 ) | ( ~n9451 & n20057 ) | ( n18304 & n20057 ) ;
  assign n20059 = ~n2737 & n10518 ;
  assign n20060 = n20059 ^ n2402 ^ 1'b0 ;
  assign n20061 = n20060 ^ n15790 ^ 1'b0 ;
  assign n20062 = ~n1342 & n10547 ;
  assign n20063 = n9586 & n20062 ;
  assign n20064 = ( n6641 & n8013 ) | ( n6641 & n20063 ) | ( n8013 & n20063 ) ;
  assign n20065 = n20064 ^ n14583 ^ 1'b0 ;
  assign n20068 = ~n6689 & n11801 ;
  assign n20069 = n20068 ^ n3345 ^ 1'b0 ;
  assign n20066 = n6895 ^ n2834 ^ 1'b0 ;
  assign n20067 = n11565 & n20066 ;
  assign n20070 = n20069 ^ n20067 ^ n8651 ;
  assign n20071 = n9632 ^ n5125 ^ 1'b0 ;
  assign n20072 = ~n3377 & n20071 ;
  assign n20073 = ( n12538 & n13252 ) | ( n12538 & n19214 ) | ( n13252 & n19214 ) ;
  assign n20074 = n12539 ^ n2453 ^ n1365 ;
  assign n20075 = n4208 ^ n1827 ^ 1'b0 ;
  assign n20076 = ~n12764 & n20075 ;
  assign n20077 = n20076 ^ n4268 ^ 1'b0 ;
  assign n20078 = n20077 ^ n17095 ^ 1'b0 ;
  assign n20079 = n20074 & n20078 ;
  assign n20080 = n3120 & ~n10027 ;
  assign n20081 = n20080 ^ n19870 ^ 1'b0 ;
  assign n20082 = ~n8254 & n20081 ;
  assign n20083 = ( ~n7321 & n12624 ) | ( ~n7321 & n16362 ) | ( n12624 & n16362 ) ;
  assign n20086 = ~n1304 & n16478 ;
  assign n20087 = n20086 ^ n2815 ^ 1'b0 ;
  assign n20088 = n10761 & ~n20087 ;
  assign n20084 = n1666 & ~n3655 ;
  assign n20085 = n5948 & n20084 ;
  assign n20089 = n20088 ^ n20085 ^ n6642 ;
  assign n20090 = n20089 ^ n11820 ^ 1'b0 ;
  assign n20091 = n16353 ^ n15094 ^ n9570 ;
  assign n20092 = n7080 ^ n6566 ^ n3425 ;
  assign n20094 = n10966 ^ n6245 ^ 1'b0 ;
  assign n20093 = ( n4381 & n6267 ) | ( n4381 & n11685 ) | ( n6267 & n11685 ) ;
  assign n20095 = n20094 ^ n20093 ^ 1'b0 ;
  assign n20096 = ( n4189 & ~n20092 ) | ( n4189 & n20095 ) | ( ~n20092 & n20095 ) ;
  assign n20097 = ~n2917 & n5685 ;
  assign n20098 = n16854 ^ n14899 ^ n1671 ;
  assign n20099 = n14218 ^ n9755 ^ 1'b0 ;
  assign n20100 = n20098 | n20099 ;
  assign n20101 = ( n16178 & ~n20097 ) | ( n16178 & n20100 ) | ( ~n20097 & n20100 ) ;
  assign n20102 = ( n1607 & ~n14156 ) | ( n1607 & n15273 ) | ( ~n14156 & n15273 ) ;
  assign n20103 = n15835 & ~n20102 ;
  assign n20104 = ~n2080 & n5427 ;
  assign n20105 = ( n5954 & n10034 ) | ( n5954 & ~n20104 ) | ( n10034 & ~n20104 ) ;
  assign n20106 = ~n5514 & n20105 ;
  assign n20107 = ~n18587 & n20106 ;
  assign n20108 = n20107 ^ n3769 ^ 1'b0 ;
  assign n20109 = n5807 & ~n11785 ;
  assign n20110 = ~n19233 & n20109 ;
  assign n20111 = ( ~n1556 & n13125 ) | ( ~n1556 & n20110 ) | ( n13125 & n20110 ) ;
  assign n20112 = n9295 ^ n643 ^ 1'b0 ;
  assign n20113 = n20112 ^ n9033 ^ 1'b0 ;
  assign n20114 = n11234 & n20113 ;
  assign n20115 = n18934 ^ n14027 ^ n6858 ;
  assign n20116 = n13873 & ~n20115 ;
  assign n20117 = n20116 ^ n2221 ^ 1'b0 ;
  assign n20118 = n7191 | n12788 ;
  assign n20119 = n15632 & ~n20118 ;
  assign n20120 = n20119 ^ n7801 ^ 1'b0 ;
  assign n20121 = n20120 ^ n10826 ^ 1'b0 ;
  assign n20122 = n18021 | n20121 ;
  assign n20123 = n7369 ^ n3817 ^ n1744 ;
  assign n20124 = n20123 ^ n1910 ^ 1'b0 ;
  assign n20125 = n4942 & ~n10018 ;
  assign n20126 = n20125 ^ n18338 ^ n3739 ;
  assign n20127 = ~n8399 & n20104 ;
  assign n20128 = n6294 & n20127 ;
  assign n20129 = ( n2466 & ~n3713 ) | ( n2466 & n20128 ) | ( ~n3713 & n20128 ) ;
  assign n20130 = n3160 ^ n929 ^ 1'b0 ;
  assign n20131 = n5529 ^ n4510 ^ n3501 ;
  assign n20132 = ( ~n8907 & n13316 ) | ( ~n8907 & n20131 ) | ( n13316 & n20131 ) ;
  assign n20133 = n9997 | n15638 ;
  assign n20134 = n20132 | n20133 ;
  assign n20135 = ( n13479 & n20130 ) | ( n13479 & ~n20134 ) | ( n20130 & ~n20134 ) ;
  assign n20136 = n3425 & n11051 ;
  assign n20137 = n3640 & n14448 ;
  assign n20138 = n19930 ^ n1867 ^ 1'b0 ;
  assign n20139 = ~n2344 & n20138 ;
  assign n20140 = n10078 & n20139 ;
  assign n20141 = n13502 & n20140 ;
  assign n20142 = ( ~n8723 & n20137 ) | ( ~n8723 & n20141 ) | ( n20137 & n20141 ) ;
  assign n20143 = n13873 ^ n1475 ^ 1'b0 ;
  assign n20144 = n20143 ^ n8731 ^ 1'b0 ;
  assign n20145 = ~n6848 & n8452 ;
  assign n20146 = n20145 ^ n15753 ^ n3091 ;
  assign n20147 = n8286 | n20146 ;
  assign n20148 = n20144 & ~n20147 ;
  assign n20149 = ~n2653 & n16292 ;
  assign n20150 = n20148 & n20149 ;
  assign n20151 = n340 & ~n19526 ;
  assign n20152 = n1594 | n1879 ;
  assign n20153 = n20152 ^ n19615 ^ 1'b0 ;
  assign n20154 = n17926 ^ n2030 ^ 1'b0 ;
  assign n20155 = n20154 ^ n15193 ^ n3465 ;
  assign n20156 = n20155 ^ n17008 ^ n2382 ;
  assign n20157 = ~n4823 & n17739 ;
  assign n20158 = ~x207 & n20157 ;
  assign n20159 = n1811 & ~n4405 ;
  assign n20160 = n20159 ^ n3372 ^ 1'b0 ;
  assign n20161 = ~n20158 & n20160 ;
  assign n20162 = ( ~n4470 & n8952 ) | ( ~n4470 & n15600 ) | ( n8952 & n15600 ) ;
  assign n20163 = n12126 ^ n9612 ^ n5800 ;
  assign n20166 = n17664 ^ n15439 ^ 1'b0 ;
  assign n20167 = n12908 & ~n20166 ;
  assign n20164 = n2755 | n15244 ;
  assign n20165 = n4624 & n20164 ;
  assign n20168 = n20167 ^ n20165 ^ 1'b0 ;
  assign n20169 = ~n2728 & n11803 ;
  assign n20170 = n5910 | n16724 ;
  assign n20171 = n2816 & n8098 ;
  assign n20172 = n20171 ^ n3515 ^ 1'b0 ;
  assign n20173 = n20172 ^ n4596 ^ n3553 ;
  assign n20174 = n20173 ^ n8506 ^ n1578 ;
  assign n20175 = n20174 ^ n12269 ^ n8059 ;
  assign n20176 = n4440 ^ n3362 ^ 1'b0 ;
  assign n20177 = n20175 & ~n20176 ;
  assign n20179 = n4813 ^ n2460 ^ n1852 ;
  assign n20178 = n3050 & ~n11623 ;
  assign n20180 = n20179 ^ n20178 ^ n2321 ;
  assign n20181 = n6658 ^ n3397 ^ 1'b0 ;
  assign n20182 = n4934 & ~n20181 ;
  assign n20183 = ~n9552 & n20182 ;
  assign n20184 = n20183 ^ n18535 ^ 1'b0 ;
  assign n20185 = n18624 ^ n780 ^ n345 ;
  assign n20186 = ~n6906 & n15927 ;
  assign n20187 = n3513 & n20186 ;
  assign n20188 = n20187 ^ n3402 ^ 1'b0 ;
  assign n20189 = n9519 & n20188 ;
  assign n20190 = n15590 ^ n773 ^ 1'b0 ;
  assign n20191 = ~n2344 & n20190 ;
  assign n20192 = n13274 | n20191 ;
  assign n20193 = ( ~x73 & n1953 ) | ( ~x73 & n20192 ) | ( n1953 & n20192 ) ;
  assign n20195 = n3542 & ~n3599 ;
  assign n20196 = ~n2073 & n20195 ;
  assign n20194 = n13213 ^ n12580 ^ n10376 ;
  assign n20197 = n20196 ^ n20194 ^ 1'b0 ;
  assign n20198 = n16769 ^ n6426 ^ 1'b0 ;
  assign n20199 = n17983 ^ n9228 ^ 1'b0 ;
  assign n20200 = n12965 | n20199 ;
  assign n20201 = ~n8610 & n10777 ;
  assign n20202 = n20201 ^ n18115 ^ 1'b0 ;
  assign n20204 = ( ~n3063 & n4350 ) | ( ~n3063 & n5992 ) | ( n4350 & n5992 ) ;
  assign n20203 = n8044 | n17203 ;
  assign n20205 = n20204 ^ n20203 ^ n12135 ;
  assign n20206 = n10063 ^ n5902 ^ n1843 ;
  assign n20207 = ( n6939 & ~n10329 ) | ( n6939 & n20206 ) | ( ~n10329 & n20206 ) ;
  assign n20208 = ( n1557 & ~n8019 ) | ( n1557 & n11683 ) | ( ~n8019 & n11683 ) ;
  assign n20209 = n3476 | n12312 ;
  assign n20210 = ( ~n1934 & n3801 ) | ( ~n1934 & n20209 ) | ( n3801 & n20209 ) ;
  assign n20211 = n20208 & ~n20210 ;
  assign n20212 = n20207 & n20211 ;
  assign n20213 = n11892 ^ n2541 ^ 1'b0 ;
  assign n20214 = ~n3502 & n3805 ;
  assign n20215 = ~n968 & n1292 ;
  assign n20216 = n20215 ^ n19739 ^ 1'b0 ;
  assign n20217 = n16162 ^ n12622 ^ 1'b0 ;
  assign n20218 = n5827 & n20217 ;
  assign n20219 = n20218 ^ n18214 ^ n13733 ;
  assign n20226 = ~n6959 & n7163 ;
  assign n20224 = ~n16405 & n17017 ;
  assign n20225 = n20224 ^ n10660 ^ 1'b0 ;
  assign n20227 = n20226 ^ n20225 ^ n13664 ;
  assign n20228 = ~n1304 & n11858 ;
  assign n20229 = n20228 ^ x246 ^ 1'b0 ;
  assign n20230 = n20227 & ~n20229 ;
  assign n20220 = n3690 & n5038 ;
  assign n20221 = n3465 | n20220 ;
  assign n20222 = n12917 & ~n20221 ;
  assign n20223 = n2100 | n20222 ;
  assign n20231 = n20230 ^ n20223 ^ 1'b0 ;
  assign n20232 = n12593 ^ n3771 ^ 1'b0 ;
  assign n20233 = n11891 & ~n20232 ;
  assign n20234 = n15203 ^ n2759 ^ n899 ;
  assign n20235 = n8593 ^ n7452 ^ n5090 ;
  assign n20236 = n10382 | n15380 ;
  assign n20237 = ~n20235 & n20236 ;
  assign n20238 = n20234 & ~n20237 ;
  assign n20239 = n6047 & n20238 ;
  assign n20240 = ~n5057 & n6901 ;
  assign n20241 = n20240 ^ n284 ^ 1'b0 ;
  assign n20242 = ( n11275 & ~n19143 ) | ( n11275 & n20241 ) | ( ~n19143 & n20241 ) ;
  assign n20243 = x142 & ~n15005 ;
  assign n20244 = n11487 & n20243 ;
  assign n20245 = ~n13014 & n13213 ;
  assign n20247 = n6863 ^ n6110 ^ n2684 ;
  assign n20246 = ~n1752 & n17539 ;
  assign n20248 = n20247 ^ n20246 ^ 1'b0 ;
  assign n20249 = ( n8362 & n15579 ) | ( n8362 & n16669 ) | ( n15579 & n16669 ) ;
  assign n20253 = ( n2108 & n2967 ) | ( n2108 & n8730 ) | ( n2967 & n8730 ) ;
  assign n20250 = n3512 & n18071 ;
  assign n20251 = n1921 & ~n20250 ;
  assign n20252 = n10229 & n20251 ;
  assign n20254 = n20253 ^ n20252 ^ 1'b0 ;
  assign n20259 = n18116 ^ n7686 ^ n6061 ;
  assign n20255 = ~n1411 & n11009 ;
  assign n20256 = n20255 ^ n19228 ^ 1'b0 ;
  assign n20257 = n20256 ^ n8895 ^ n2180 ;
  assign n20258 = n16813 & ~n20257 ;
  assign n20260 = n20259 ^ n20258 ^ 1'b0 ;
  assign n20261 = n20254 | n20260 ;
  assign n20262 = n20261 ^ n19132 ^ 1'b0 ;
  assign n20263 = ~n11570 & n20262 ;
  assign n20264 = n7280 & n20263 ;
  assign n20265 = ~n261 & n18339 ;
  assign n20272 = n2262 & ~n5944 ;
  assign n20270 = ( n9257 & ~n13474 ) | ( n9257 & n15180 ) | ( ~n13474 & n15180 ) ;
  assign n20266 = n15646 ^ x17 ^ 1'b0 ;
  assign n20267 = n10113 ^ n4423 ^ 1'b0 ;
  assign n20268 = n20266 | n20267 ;
  assign n20269 = n20268 ^ n19492 ^ n16230 ;
  assign n20271 = n20270 ^ n20269 ^ 1'b0 ;
  assign n20273 = n20272 ^ n20271 ^ 1'b0 ;
  assign n20274 = ~n17009 & n20273 ;
  assign n20275 = n9309 & n9924 ;
  assign n20276 = n20275 ^ n10342 ^ 1'b0 ;
  assign n20277 = ( n14474 & ~n14520 ) | ( n14474 & n20276 ) | ( ~n14520 & n20276 ) ;
  assign n20278 = n20277 ^ n12494 ^ 1'b0 ;
  assign n20279 = ~n15922 & n20278 ;
  assign n20280 = n7383 & ~n16934 ;
  assign n20281 = n20280 ^ n3703 ^ 1'b0 ;
  assign n20282 = ( n2075 & n7304 ) | ( n2075 & ~n11578 ) | ( n7304 & ~n11578 ) ;
  assign n20283 = n1191 & ~n1684 ;
  assign n20284 = n2825 & ~n20283 ;
  assign n20285 = n15921 & ~n20284 ;
  assign n20286 = ( n15994 & ~n20282 ) | ( n15994 & n20285 ) | ( ~n20282 & n20285 ) ;
  assign n20287 = n20281 & ~n20286 ;
  assign n20288 = n20287 ^ n14638 ^ 1'b0 ;
  assign n20289 = ~n6311 & n13054 ;
  assign n20290 = n13758 ^ n5075 ^ n3771 ;
  assign n20291 = ( n2177 & n5494 ) | ( n2177 & ~n20290 ) | ( n5494 & ~n20290 ) ;
  assign n20292 = ~n1757 & n4268 ;
  assign n20293 = ~n7046 & n20292 ;
  assign n20294 = ( n3248 & n4905 ) | ( n3248 & ~n18500 ) | ( n4905 & ~n18500 ) ;
  assign n20295 = n20294 ^ n4935 ^ 1'b0 ;
  assign n20296 = n6670 & n13173 ;
  assign n20297 = x169 & ~n3196 ;
  assign n20298 = n20297 ^ n20179 ^ 1'b0 ;
  assign n20299 = x168 & n20298 ;
  assign n20300 = ( ~n3845 & n20296 ) | ( ~n3845 & n20299 ) | ( n20296 & n20299 ) ;
  assign n20301 = n5649 | n20300 ;
  assign n20302 = n11912 ^ n354 ^ 1'b0 ;
  assign n20303 = n20302 ^ n19266 ^ 1'b0 ;
  assign n20304 = n18942 ^ n3208 ^ 1'b0 ;
  assign n20305 = ~n4008 & n20304 ;
  assign n20306 = ( ~n8291 & n13508 ) | ( ~n8291 & n20305 ) | ( n13508 & n20305 ) ;
  assign n20307 = n20306 ^ n4311 ^ 1'b0 ;
  assign n20308 = n20303 | n20307 ;
  assign n20309 = ~n2322 & n12563 ;
  assign n20310 = n14843 & n20309 ;
  assign n20311 = n20310 ^ n11565 ^ 1'b0 ;
  assign n20312 = n20311 ^ n10557 ^ n8306 ;
  assign n20313 = ( n15526 & n16241 ) | ( n15526 & ~n20312 ) | ( n16241 & ~n20312 ) ;
  assign n20314 = n16926 ^ n2569 ^ 1'b0 ;
  assign n20315 = ~n11021 & n20314 ;
  assign n20316 = ~n19455 & n20315 ;
  assign n20317 = n9853 ^ n4118 ^ 1'b0 ;
  assign n20318 = n1542 | n16355 ;
  assign n20319 = n20318 ^ n5680 ^ 1'b0 ;
  assign n20320 = n18606 ^ n8977 ^ 1'b0 ;
  assign n20321 = ~n20319 & n20320 ;
  assign n20322 = n11352 ^ n1516 ^ 1'b0 ;
  assign n20323 = ~n9840 & n20322 ;
  assign n20324 = ~n7871 & n20323 ;
  assign n20325 = n20324 ^ n11544 ^ 1'b0 ;
  assign n20326 = n8210 ^ n3509 ^ n617 ;
  assign n20327 = n19450 ^ n14963 ^ 1'b0 ;
  assign n20328 = n20326 | n20327 ;
  assign n20334 = ( n4179 & n6025 ) | ( n4179 & n19163 ) | ( n6025 & n19163 ) ;
  assign n20335 = n3227 | n5325 ;
  assign n20336 = n20334 | n20335 ;
  assign n20329 = n2721 | n17502 ;
  assign n20330 = n7686 & ~n20329 ;
  assign n20331 = n20330 ^ n2649 ^ 1'b0 ;
  assign n20332 = n20331 ^ n12033 ^ n3955 ;
  assign n20333 = ( n14643 & n15368 ) | ( n14643 & ~n20332 ) | ( n15368 & ~n20332 ) ;
  assign n20337 = n20336 ^ n20333 ^ 1'b0 ;
  assign n20338 = n20328 | n20337 ;
  assign n20339 = n16500 ^ n13373 ^ n8468 ;
  assign n20340 = n15771 ^ n10869 ^ 1'b0 ;
  assign n20341 = ~n20339 & n20340 ;
  assign n20342 = ( n19947 & n20338 ) | ( n19947 & ~n20341 ) | ( n20338 & ~n20341 ) ;
  assign n20343 = n10538 ^ n7633 ^ n2045 ;
  assign n20344 = ( n2633 & n10535 ) | ( n2633 & ~n20343 ) | ( n10535 & ~n20343 ) ;
  assign n20345 = n17058 ^ n5864 ^ 1'b0 ;
  assign n20346 = n4490 ^ n3816 ^ n2547 ;
  assign n20347 = ( x14 & n9273 ) | ( x14 & n20346 ) | ( n9273 & n20346 ) ;
  assign n20348 = n1548 & n5605 ;
  assign n20349 = n20348 ^ n7062 ^ 1'b0 ;
  assign n20350 = n20349 ^ n7481 ^ n7024 ;
  assign n20351 = n20350 ^ n14680 ^ n5526 ;
  assign n20352 = n20351 ^ n2720 ^ n1370 ;
  assign n20353 = n17239 ^ n17176 ^ 1'b0 ;
  assign n20354 = n3737 & n4595 ;
  assign n20355 = n20354 ^ n16217 ^ 1'b0 ;
  assign n20356 = ( n774 & ~n20353 ) | ( n774 & n20355 ) | ( ~n20353 & n20355 ) ;
  assign n20357 = n20352 | n20356 ;
  assign n20358 = n7484 ^ n2045 ^ 1'b0 ;
  assign n20359 = n20358 ^ n12064 ^ 1'b0 ;
  assign n20360 = n11215 ^ n2502 ^ 1'b0 ;
  assign n20361 = n20359 & ~n20360 ;
  assign n20362 = n20361 ^ n15008 ^ n10104 ;
  assign n20363 = n6008 | n16995 ;
  assign n20364 = n7410 | n20363 ;
  assign n20365 = n2332 & n15172 ;
  assign n20366 = n20365 ^ n7116 ^ 1'b0 ;
  assign n20367 = n8440 ^ n3037 ^ 1'b0 ;
  assign n20368 = ( n11078 & n15362 ) | ( n11078 & n18725 ) | ( n15362 & n18725 ) ;
  assign n20369 = n7203 & ~n7990 ;
  assign n20370 = n20369 ^ n4732 ^ 1'b0 ;
  assign n20371 = n8284 ^ n3517 ^ 1'b0 ;
  assign n20372 = n2588 & ~n5596 ;
  assign n20373 = ~n18738 & n20372 ;
  assign n20374 = ( ~n8737 & n20371 ) | ( ~n8737 & n20373 ) | ( n20371 & n20373 ) ;
  assign n20375 = n20374 ^ n18746 ^ n11671 ;
  assign n20376 = n1841 ^ x82 ^ 1'b0 ;
  assign n20377 = n20376 ^ n8772 ^ 1'b0 ;
  assign n20378 = n20377 ^ n15319 ^ 1'b0 ;
  assign n20379 = n6331 & ~n20378 ;
  assign n20380 = n20379 ^ n18596 ^ n5231 ;
  assign n20381 = n12713 & ~n20380 ;
  assign n20382 = n20381 ^ n8240 ^ 1'b0 ;
  assign n20385 = n756 & n12795 ;
  assign n20386 = n20385 ^ n739 ^ 1'b0 ;
  assign n20384 = ( ~n4934 & n7119 ) | ( ~n4934 & n10418 ) | ( n7119 & n10418 ) ;
  assign n20383 = ~n11396 & n16029 ;
  assign n20387 = n20386 ^ n20384 ^ n20383 ;
  assign n20391 = n9916 & ~n12823 ;
  assign n20392 = n12960 & n20391 ;
  assign n20388 = ~n5592 & n7382 ;
  assign n20389 = ~n13750 & n20388 ;
  assign n20390 = n20389 ^ n14934 ^ n9670 ;
  assign n20393 = n20392 ^ n20390 ^ 1'b0 ;
  assign n20394 = n14244 ^ n8409 ^ 1'b0 ;
  assign n20395 = n18288 | n20394 ;
  assign n20396 = n1676 & ~n20395 ;
  assign n20397 = ~n16951 & n20396 ;
  assign n20398 = ( n8581 & n9188 ) | ( n8581 & ~n20397 ) | ( n9188 & ~n20397 ) ;
  assign n20399 = n3844 | n11677 ;
  assign n20400 = n8689 & ~n20399 ;
  assign n20401 = n10178 ^ n6344 ^ 1'b0 ;
  assign n20402 = ~n20400 & n20401 ;
  assign n20403 = ~n9359 & n15598 ;
  assign n20404 = ( n16504 & n18977 ) | ( n16504 & ~n20403 ) | ( n18977 & ~n20403 ) ;
  assign n20405 = n2643 | n20404 ;
  assign n20406 = n20405 ^ n10637 ^ 1'b0 ;
  assign n20407 = x54 & n6666 ;
  assign n20408 = n20407 ^ n5444 ^ 1'b0 ;
  assign n20409 = n11283 ^ x149 ^ 1'b0 ;
  assign n20410 = ( n3759 & n14064 ) | ( n3759 & n20409 ) | ( n14064 & n20409 ) ;
  assign n20411 = ~n18848 & n20410 ;
  assign n20414 = n18374 ^ n1334 ^ 1'b0 ;
  assign n20415 = ~n2728 & n20414 ;
  assign n20412 = ~n1075 & n5026 ;
  assign n20413 = n8933 & n20412 ;
  assign n20416 = n20415 ^ n20413 ^ 1'b0 ;
  assign n20417 = n769 & n5087 ;
  assign n20419 = n9110 ^ x127 ^ 1'b0 ;
  assign n20420 = n18351 & ~n20419 ;
  assign n20418 = n2101 & ~n4998 ;
  assign n20421 = n20420 ^ n20418 ^ 1'b0 ;
  assign n20422 = n7902 ^ n5524 ^ 1'b0 ;
  assign n20423 = n20421 | n20422 ;
  assign n20424 = ( n1385 & n2722 ) | ( n1385 & ~n7281 ) | ( n2722 & ~n7281 ) ;
  assign n20425 = n20423 | n20424 ;
  assign n20426 = n20417 | n20425 ;
  assign n20427 = n20426 ^ n9004 ^ 1'b0 ;
  assign n20428 = n4220 & ~n20427 ;
  assign n20429 = ~n5015 & n11327 ;
  assign n20430 = n20429 ^ n12239 ^ 1'b0 ;
  assign n20431 = n20430 ^ n20346 ^ n9205 ;
  assign n20432 = ( n11859 & ~n12585 ) | ( n11859 & n20431 ) | ( ~n12585 & n20431 ) ;
  assign n20433 = n1773 ^ n1317 ^ n393 ;
  assign n20434 = n20433 ^ n7702 ^ 1'b0 ;
  assign n20435 = n20434 ^ n17635 ^ n1474 ;
  assign n20436 = ( n5195 & n7200 ) | ( n5195 & n8848 ) | ( n7200 & n8848 ) ;
  assign n20437 = n20436 ^ n14180 ^ n2559 ;
  assign n20438 = n16652 & n20437 ;
  assign n20439 = ~n14452 & n20438 ;
  assign n20440 = n20439 ^ n6937 ^ 1'b0 ;
  assign n20441 = n16534 ^ x116 ^ 1'b0 ;
  assign n20442 = n15380 ^ n13934 ^ n322 ;
  assign n20443 = n1434 & n6579 ;
  assign n20444 = n20443 ^ n7711 ^ 1'b0 ;
  assign n20445 = n13686 ^ n7198 ^ 1'b0 ;
  assign n20446 = ( ~n6124 & n20444 ) | ( ~n6124 & n20445 ) | ( n20444 & n20445 ) ;
  assign n20447 = n20446 ^ n12622 ^ n745 ;
  assign n20448 = n20442 | n20447 ;
  assign n20449 = n20441 | n20448 ;
  assign n20450 = n20449 ^ n17306 ^ 1'b0 ;
  assign n20451 = ~n2279 & n13220 ;
  assign n20452 = n20451 ^ n1922 ^ 1'b0 ;
  assign n20453 = n1608 & n16847 ;
  assign n20454 = n20452 & ~n20453 ;
  assign n20455 = n20454 ^ n17256 ^ 1'b0 ;
  assign n20456 = n3942 & ~n20455 ;
  assign n20457 = ( n8326 & ~n14373 ) | ( n8326 & n20456 ) | ( ~n14373 & n20456 ) ;
  assign n20458 = ( ~x157 & n284 ) | ( ~x157 & n20457 ) | ( n284 & n20457 ) ;
  assign n20459 = n12322 ^ n10349 ^ n609 ;
  assign n20468 = n10478 ^ n2597 ^ 1'b0 ;
  assign n20460 = n716 & n2594 ;
  assign n20461 = n20460 ^ n4054 ^ n1958 ;
  assign n20462 = ( n7824 & ~n8566 ) | ( n7824 & n20461 ) | ( ~n8566 & n20461 ) ;
  assign n20463 = n2498 & n14290 ;
  assign n20464 = n3378 | n20463 ;
  assign n20465 = n20464 ^ n7034 ^ 1'b0 ;
  assign n20466 = n20462 | n20465 ;
  assign n20467 = n20466 ^ n12088 ^ 1'b0 ;
  assign n20469 = n20468 ^ n20467 ^ 1'b0 ;
  assign n20470 = n15312 ^ n9126 ^ 1'b0 ;
  assign n20471 = n6865 & ~n20470 ;
  assign n20472 = ~n4860 & n20471 ;
  assign n20473 = n20472 ^ n11679 ^ 1'b0 ;
  assign n20474 = n16626 & n20473 ;
  assign n20475 = n8809 & n20474 ;
  assign n20476 = ( n1744 & n8233 ) | ( n1744 & ~n12992 ) | ( n8233 & ~n12992 ) ;
  assign n20477 = n20476 ^ n14293 ^ 1'b0 ;
  assign n20478 = n5356 & n8911 ;
  assign n20479 = n20478 ^ n5613 ^ 1'b0 ;
  assign n20480 = n14349 & ~n20479 ;
  assign n20481 = n20480 ^ n16570 ^ 1'b0 ;
  assign n20482 = n7021 ^ n4279 ^ n633 ;
  assign n20483 = n13708 ^ n3032 ^ n268 ;
  assign n20487 = n5592 | n7136 ;
  assign n20484 = n10517 ^ n8745 ^ n2930 ;
  assign n20485 = n8557 & n20484 ;
  assign n20486 = n19373 & n20485 ;
  assign n20488 = n20487 ^ n20486 ^ 1'b0 ;
  assign n20489 = n10404 | n20488 ;
  assign n20490 = n3995 & ~n8098 ;
  assign n20492 = n5444 ^ n3813 ^ 1'b0 ;
  assign n20493 = n8400 | n20492 ;
  assign n20491 = ~n5081 & n7377 ;
  assign n20494 = n20493 ^ n20491 ^ 1'b0 ;
  assign n20495 = n20490 | n20494 ;
  assign n20496 = n15378 | n18456 ;
  assign n20497 = n18604 & ~n20496 ;
  assign n20498 = n20352 ^ n16648 ^ n13347 ;
  assign n20499 = n10674 ^ n6420 ^ n399 ;
  assign n20500 = ~n5665 & n20499 ;
  assign n20501 = n6368 & n20500 ;
  assign n20502 = n20501 ^ n15406 ^ n4301 ;
  assign n20503 = n14313 ^ n3395 ^ 1'b0 ;
  assign n20504 = n15153 ^ n6244 ^ n5736 ;
  assign n20505 = ~n7970 & n9732 ;
  assign n20506 = n20505 ^ n11209 ^ 1'b0 ;
  assign n20507 = n20504 | n20506 ;
  assign n20508 = n17157 ^ n4852 ^ 1'b0 ;
  assign n20509 = n20508 ^ n19894 ^ n16665 ;
  assign n20510 = n9109 & n13326 ;
  assign n20511 = ~n2965 & n20510 ;
  assign n20512 = n19161 ^ n16421 ^ n8554 ;
  assign n20516 = n4139 & n7586 ;
  assign n20513 = n6311 ^ n5759 ^ 1'b0 ;
  assign n20514 = n6566 & ~n20513 ;
  assign n20515 = n14677 & n20514 ;
  assign n20517 = n20516 ^ n20515 ^ 1'b0 ;
  assign n20518 = ( n17176 & ~n20454 ) | ( n17176 & n20517 ) | ( ~n20454 & n20517 ) ;
  assign n20519 = n2663 & ~n13748 ;
  assign n20520 = n20519 ^ n9845 ^ n5091 ;
  assign n20521 = n3902 & ~n9024 ;
  assign n20522 = n20521 ^ n5409 ^ 1'b0 ;
  assign n20523 = n6442 & n12024 ;
  assign n20524 = ~n11670 & n20523 ;
  assign n20525 = n7968 ^ n7380 ^ 1'b0 ;
  assign n20526 = ( n17314 & n20524 ) | ( n17314 & ~n20525 ) | ( n20524 & ~n20525 ) ;
  assign n20527 = n11445 | n20349 ;
  assign n20528 = n20527 ^ n11079 ^ 1'b0 ;
  assign n20529 = n7401 ^ n2016 ^ x152 ;
  assign n20530 = ( n15021 & ~n18850 ) | ( n15021 & n20529 ) | ( ~n18850 & n20529 ) ;
  assign n20537 = n16155 | n19836 ;
  assign n20538 = n20537 ^ n8070 ^ 1'b0 ;
  assign n20535 = ~x159 & n6846 ;
  assign n20536 = ~n5584 & n20535 ;
  assign n20533 = ( ~n3260 & n3947 ) | ( ~n3260 & n6292 ) | ( n3947 & n6292 ) ;
  assign n20531 = n13094 ^ n8399 ^ 1'b0 ;
  assign n20532 = n20531 ^ n16503 ^ n10102 ;
  assign n20534 = n20533 ^ n20532 ^ 1'b0 ;
  assign n20539 = n20538 ^ n20536 ^ n20534 ;
  assign n20540 = ( ~n12309 & n13176 ) | ( ~n12309 & n14070 ) | ( n13176 & n14070 ) ;
  assign n20541 = n9769 ^ x100 ^ 1'b0 ;
  assign n20542 = n8174 & n20541 ;
  assign n20543 = n9315 & ~n10502 ;
  assign n20544 = ~n20542 & n20543 ;
  assign n20545 = n10732 ^ n1520 ^ 1'b0 ;
  assign n20546 = ( n770 & n1947 ) | ( n770 & ~n5115 ) | ( n1947 & ~n5115 ) ;
  assign n20547 = n5851 & n20546 ;
  assign n20548 = ~n20545 & n20547 ;
  assign n20549 = n8903 & ~n11476 ;
  assign n20550 = n20549 ^ n8808 ^ 1'b0 ;
  assign n20551 = ( n8139 & n20548 ) | ( n8139 & n20550 ) | ( n20548 & n20550 ) ;
  assign n20552 = n20551 ^ n693 ^ 1'b0 ;
  assign n20553 = n10731 & n20552 ;
  assign n20554 = n16911 & n20553 ;
  assign n20555 = n16170 ^ n1705 ^ 1'b0 ;
  assign n20556 = n8348 | n20555 ;
  assign n20557 = n20556 ^ n4021 ^ 1'b0 ;
  assign n20558 = ~n713 & n5571 ;
  assign n20559 = n20558 ^ n10509 ^ 1'b0 ;
  assign n20560 = n16774 ^ n4053 ^ 1'b0 ;
  assign n20561 = n13545 ^ n13388 ^ n1268 ;
  assign n20562 = n20561 ^ n7494 ^ x140 ;
  assign n20563 = n4064 & ~n6019 ;
  assign n20564 = ~n17232 & n19011 ;
  assign n20565 = n20564 ^ n20482 ^ 1'b0 ;
  assign n20566 = n7905 ^ n1020 ^ 1'b0 ;
  assign n20567 = n8306 & n20566 ;
  assign n20568 = ( n5424 & n11089 ) | ( n5424 & ~n11898 ) | ( n11089 & ~n11898 ) ;
  assign n20569 = ( n5376 & ~n20567 ) | ( n5376 & n20568 ) | ( ~n20567 & n20568 ) ;
  assign n20570 = ( n1363 & n8868 ) | ( n1363 & ~n20569 ) | ( n8868 & ~n20569 ) ;
  assign n20571 = n15421 ^ n13289 ^ 1'b0 ;
  assign n20572 = n20571 ^ n13462 ^ 1'b0 ;
  assign n20574 = n13813 | n18243 ;
  assign n20575 = x173 & n20574 ;
  assign n20573 = n6334 ^ n2021 ^ 1'b0 ;
  assign n20576 = n20575 ^ n20573 ^ n11907 ;
  assign n20577 = ( n388 & n12715 ) | ( n388 & ~n15772 ) | ( n12715 & ~n15772 ) ;
  assign n20583 = n1091 & n13646 ;
  assign n20578 = n1610 ^ n753 ^ 1'b0 ;
  assign n20579 = n9268 & n20578 ;
  assign n20580 = ~n4589 & n4851 ;
  assign n20581 = n20580 ^ n1871 ^ 1'b0 ;
  assign n20582 = ( n9286 & n20579 ) | ( n9286 & n20581 ) | ( n20579 & n20581 ) ;
  assign n20584 = n20583 ^ n20582 ^ n10921 ;
  assign n20585 = n12487 ^ n940 ^ 1'b0 ;
  assign n20586 = ~n9039 & n20585 ;
  assign n20587 = ~n586 & n8946 ;
  assign n20588 = n5302 ^ n1737 ^ 1'b0 ;
  assign n20589 = n12348 & n20588 ;
  assign n20590 = n1059 | n6958 ;
  assign n20591 = n2414 & ~n20590 ;
  assign n20592 = ( ~n8200 & n9658 ) | ( ~n8200 & n20591 ) | ( n9658 & n20591 ) ;
  assign n20593 = n20592 ^ n15692 ^ n2234 ;
  assign n20594 = ~n16089 & n20516 ;
  assign n20595 = ~n829 & n20594 ;
  assign n20596 = n3913 & ~n9714 ;
  assign n20597 = n4105 & ~n10728 ;
  assign n20598 = n20597 ^ n2607 ^ 1'b0 ;
  assign n20599 = ~n13578 & n20598 ;
  assign n20600 = n17719 & n20599 ;
  assign n20601 = n12873 ^ n10102 ^ n7669 ;
  assign n20602 = n20601 ^ n19605 ^ n7752 ;
  assign n20609 = n10284 ^ n6826 ^ n2451 ;
  assign n20603 = x167 & x222 ;
  assign n20604 = n737 & n20603 ;
  assign n20605 = n20604 ^ n7969 ^ 1'b0 ;
  assign n20606 = ( ~n1434 & n4805 ) | ( ~n1434 & n7687 ) | ( n4805 & n7687 ) ;
  assign n20607 = n13633 | n20606 ;
  assign n20608 = ( ~n10628 & n20605 ) | ( ~n10628 & n20607 ) | ( n20605 & n20607 ) ;
  assign n20610 = n20609 ^ n20608 ^ n12470 ;
  assign n20611 = n19453 ^ n6819 ^ n511 ;
  assign n20612 = n6969 | n7261 ;
  assign n20613 = n20612 ^ n5347 ^ 1'b0 ;
  assign n20614 = ( n10220 & ~n18963 ) | ( n10220 & n20613 ) | ( ~n18963 & n20613 ) ;
  assign n20618 = n890 & ~n12166 ;
  assign n20619 = n17751 & n20618 ;
  assign n20620 = n9093 & ~n20619 ;
  assign n20615 = n7254 ^ n6048 ^ 1'b0 ;
  assign n20616 = n20615 ^ n1783 ^ 1'b0 ;
  assign n20617 = ( n10307 & n12101 ) | ( n10307 & ~n20616 ) | ( n12101 & ~n20616 ) ;
  assign n20621 = n20620 ^ n20617 ^ x195 ;
  assign n20622 = n20614 | n20621 ;
  assign n20623 = n15061 | n20622 ;
  assign n20624 = n17483 ^ n16675 ^ 1'b0 ;
  assign n20625 = n12766 ^ n3186 ^ 1'b0 ;
  assign n20626 = n6891 ^ n1470 ^ 1'b0 ;
  assign n20627 = ~n7131 & n11579 ;
  assign n20628 = n20627 ^ n4930 ^ 1'b0 ;
  assign n20629 = ~n9626 & n20628 ;
  assign n20630 = ( n5921 & n15414 ) | ( n5921 & n20629 ) | ( n15414 & n20629 ) ;
  assign n20631 = ( n20625 & n20626 ) | ( n20625 & ~n20630 ) | ( n20626 & ~n20630 ) ;
  assign n20632 = ~n7440 & n13294 ;
  assign n20633 = n11564 & n20632 ;
  assign n20634 = n20633 ^ n14603 ^ 1'b0 ;
  assign n20635 = n9080 & ~n16581 ;
  assign n20636 = n16037 & n20635 ;
  assign n20638 = n5994 & ~n17958 ;
  assign n20637 = n19569 ^ n7131 ^ 1'b0 ;
  assign n20639 = n20638 ^ n20637 ^ 1'b0 ;
  assign n20640 = n1231 | n10201 ;
  assign n20641 = n5497 & ~n20640 ;
  assign n20642 = n2764 & n11285 ;
  assign n20643 = ( n5659 & n10684 ) | ( n5659 & ~n10904 ) | ( n10684 & ~n10904 ) ;
  assign n20644 = n4965 ^ n1233 ^ 1'b0 ;
  assign n20645 = n20643 | n20644 ;
  assign n20646 = n12386 ^ n4356 ^ 1'b0 ;
  assign n20647 = ( ~n1957 & n6740 ) | ( ~n1957 & n8839 ) | ( n6740 & n8839 ) ;
  assign n20648 = n10242 ^ n10072 ^ 1'b0 ;
  assign n20649 = n16968 ^ n3026 ^ 1'b0 ;
  assign n20650 = n4316 | n15153 ;
  assign n20651 = n3753 & ~n20650 ;
  assign n20652 = n3806 | n6456 ;
  assign n20653 = n20651 & ~n20652 ;
  assign n20654 = ~n1246 & n8625 ;
  assign n20655 = ~n1447 & n20654 ;
  assign n20656 = n7892 & ~n14477 ;
  assign n20657 = n4183 & n20656 ;
  assign n20658 = ( n5219 & n8234 ) | ( n5219 & ~n11097 ) | ( n8234 & ~n11097 ) ;
  assign n20659 = n20658 ^ n2170 ^ n307 ;
  assign n20660 = ~x180 & n20659 ;
  assign n20661 = ( n20655 & ~n20657 ) | ( n20655 & n20660 ) | ( ~n20657 & n20660 ) ;
  assign n20662 = ~n4890 & n7028 ;
  assign n20663 = n3765 & n20662 ;
  assign n20664 = n20663 ^ n19708 ^ n8964 ;
  assign n20665 = n20664 ^ n14959 ^ n3736 ;
  assign n20666 = n855 & n3940 ;
  assign n20667 = n9145 ^ n8370 ^ 1'b0 ;
  assign n20668 = n20666 & ~n20667 ;
  assign n20669 = ~n10466 & n11381 ;
  assign n20670 = n17934 & n20669 ;
  assign n20671 = n20670 ^ n14008 ^ 1'b0 ;
  assign n20672 = ~n15378 & n20671 ;
  assign n20673 = n11451 ^ n2716 ^ 1'b0 ;
  assign n20674 = n20673 ^ n1558 ^ 1'b0 ;
  assign n20675 = n19779 & ~n20674 ;
  assign n20676 = n2585 & n4224 ;
  assign n20677 = n20676 ^ n4341 ^ 1'b0 ;
  assign n20678 = ~n2982 & n13643 ;
  assign n20679 = n2498 & n20678 ;
  assign n20680 = ( n1723 & n20677 ) | ( n1723 & n20679 ) | ( n20677 & n20679 ) ;
  assign n20681 = n20668 ^ n9434 ^ 1'b0 ;
  assign n20682 = n4579 & ~n20681 ;
  assign n20683 = n17556 ^ n4860 ^ n4017 ;
  assign n20684 = n20683 ^ n7225 ^ n6397 ;
  assign n20685 = ~n4680 & n8049 ;
  assign n20686 = n20685 ^ n7754 ^ n3472 ;
  assign n20687 = ( ~n11589 & n14689 ) | ( ~n11589 & n20686 ) | ( n14689 & n20686 ) ;
  assign n20688 = n13461 ^ n1233 ^ 1'b0 ;
  assign n20689 = ( ~n8658 & n11411 ) | ( ~n8658 & n11482 ) | ( n11411 & n11482 ) ;
  assign n20690 = n20688 & n20689 ;
  assign n20691 = ( n1451 & ~n2836 ) | ( n1451 & n3874 ) | ( ~n2836 & n3874 ) ;
  assign n20692 = n20563 & ~n20691 ;
  assign n20693 = n914 & n20692 ;
  assign n20694 = n17682 ^ n12941 ^ 1'b0 ;
  assign n20695 = ( ~n1330 & n3727 ) | ( ~n1330 & n5532 ) | ( n3727 & n5532 ) ;
  assign n20696 = ( n1077 & ~n15749 ) | ( n1077 & n20695 ) | ( ~n15749 & n20695 ) ;
  assign n20697 = n7980 & n14769 ;
  assign n20698 = ~n8435 & n20697 ;
  assign n20699 = n1380 & n11990 ;
  assign n20700 = n20699 ^ n5085 ^ 1'b0 ;
  assign n20701 = n18707 ^ n14644 ^ 1'b0 ;
  assign n20702 = n1812 & n14016 ;
  assign n20703 = n20702 ^ n11332 ^ 1'b0 ;
  assign n20704 = n4966 & ~n7055 ;
  assign n20705 = n20704 ^ n11077 ^ 1'b0 ;
  assign n20706 = ~n648 & n20705 ;
  assign n20707 = n20706 ^ n17937 ^ n3548 ;
  assign n20708 = n20707 ^ n20178 ^ 1'b0 ;
  assign n20709 = n20708 ^ n3619 ^ n1594 ;
  assign n20710 = n6114 ^ n1378 ^ n1377 ;
  assign n20711 = ~n6264 & n20710 ;
  assign n20712 = n16150 & n20711 ;
  assign n20713 = n20712 ^ n6346 ^ 1'b0 ;
  assign n20714 = ~n10419 & n20713 ;
  assign n20715 = n4890 & n20714 ;
  assign n20716 = ( n8800 & ~n17076 ) | ( n8800 & n18319 ) | ( ~n17076 & n18319 ) ;
  assign n20717 = n6886 | n10396 ;
  assign n20718 = n12649 & ~n20717 ;
  assign n20719 = ( ~n11294 & n13382 ) | ( ~n11294 & n20718 ) | ( n13382 & n20718 ) ;
  assign n20720 = n8970 | n17618 ;
  assign n20721 = n16115 & ~n20720 ;
  assign n20722 = n12658 | n20721 ;
  assign n20723 = n12738 | n20722 ;
  assign n20724 = n17026 ^ n13571 ^ n9970 ;
  assign n20725 = n8336 & ~n12917 ;
  assign n20726 = ~n16484 & n20725 ;
  assign n20727 = n20724 & n20726 ;
  assign n20728 = n8206 | n10732 ;
  assign n20729 = n20583 | n20728 ;
  assign n20730 = n20727 & ~n20729 ;
  assign n20731 = ~n1941 & n8739 ;
  assign n20732 = n19633 ^ n7869 ^ 1'b0 ;
  assign n20733 = n20731 & n20732 ;
  assign n20734 = n20733 ^ n13538 ^ n8408 ;
  assign n20735 = ( n4919 & ~n7518 ) | ( n4919 & n15482 ) | ( ~n7518 & n15482 ) ;
  assign n20736 = n20735 ^ n8331 ^ n446 ;
  assign n20737 = ~n7917 & n20736 ;
  assign n20738 = n1597 | n1748 ;
  assign n20739 = ( n2560 & ~n20194 ) | ( n2560 & n20738 ) | ( ~n20194 & n20738 ) ;
  assign n20740 = n20739 ^ n12826 ^ 1'b0 ;
  assign n20741 = ( n3630 & n6120 ) | ( n3630 & n7521 ) | ( n6120 & n7521 ) ;
  assign n20742 = n2925 | n20741 ;
  assign n20743 = n20742 ^ n6173 ^ 1'b0 ;
  assign n20744 = n7740 | n8244 ;
  assign n20745 = n3844 & ~n20744 ;
  assign n20746 = ( n293 & ~n6098 ) | ( n293 & n20745 ) | ( ~n6098 & n20745 ) ;
  assign n20747 = ( n1916 & n6344 ) | ( n1916 & n8062 ) | ( n6344 & n8062 ) ;
  assign n20748 = ( ~n4695 & n20177 ) | ( ~n4695 & n20747 ) | ( n20177 & n20747 ) ;
  assign n20749 = n8976 ^ n4560 ^ n1393 ;
  assign n20750 = ~n7039 & n20749 ;
  assign n20751 = n20750 ^ n12503 ^ 1'b0 ;
  assign n20752 = n6785 ^ n855 ^ 1'b0 ;
  assign n20753 = n7819 ^ n6358 ^ 1'b0 ;
  assign n20754 = n4470 | n20753 ;
  assign n20755 = n19077 | n20754 ;
  assign n20756 = n20752 & ~n20755 ;
  assign n20757 = n11604 & ~n17859 ;
  assign n20758 = n20757 ^ n3008 ^ 1'b0 ;
  assign n20759 = ( ~n3830 & n18666 ) | ( ~n3830 & n19282 ) | ( n18666 & n19282 ) ;
  assign n20760 = n6463 & n11263 ;
  assign n20761 = n20760 ^ n13776 ^ 1'b0 ;
  assign n20762 = n12356 ^ n7165 ^ 1'b0 ;
  assign n20763 = n5201 & ~n20762 ;
  assign n20764 = n20763 ^ n299 ^ 1'b0 ;
  assign n20765 = n12474 & ~n20764 ;
  assign n20766 = n14739 ^ n8699 ^ n6149 ;
  assign n20767 = ( n1111 & n16616 ) | ( n1111 & ~n20766 ) | ( n16616 & ~n20766 ) ;
  assign n20768 = n20765 & n20767 ;
  assign n20771 = n3126 & ~n7003 ;
  assign n20772 = n20771 ^ n10681 ^ 1'b0 ;
  assign n20769 = n10557 ^ n4306 ^ n4254 ;
  assign n20770 = ( n7564 & n17553 ) | ( n7564 & ~n20769 ) | ( n17553 & ~n20769 ) ;
  assign n20773 = n20772 ^ n20770 ^ n8658 ;
  assign n20774 = n12740 ^ n1028 ^ 1'b0 ;
  assign n20775 = n4234 & ~n20774 ;
  assign n20776 = n2977 & n7427 ;
  assign n20777 = n20776 ^ n3496 ^ 1'b0 ;
  assign n20778 = n20777 ^ n17571 ^ 1'b0 ;
  assign n20779 = n1867 & ~n3056 ;
  assign n20780 = n20779 ^ n12140 ^ 1'b0 ;
  assign n20781 = n2475 & n17561 ;
  assign n20782 = n5604 | n20781 ;
  assign n20783 = ~n12150 & n20782 ;
  assign n20784 = ~n20780 & n20783 ;
  assign n20785 = n13785 & ~n20784 ;
  assign n20786 = n20785 ^ n19867 ^ 1'b0 ;
  assign n20787 = ( n799 & n1558 ) | ( n799 & ~n4055 ) | ( n1558 & ~n4055 ) ;
  assign n20788 = n8754 & ~n20787 ;
  assign n20789 = n20788 ^ n10610 ^ 1'b0 ;
  assign n20790 = n3868 & n4291 ;
  assign n20791 = n352 & n20790 ;
  assign n20792 = n3197 | n20791 ;
  assign n20793 = n20789 & ~n20792 ;
  assign n20794 = n11359 & ~n20793 ;
  assign n20795 = n20794 ^ n17509 ^ n5460 ;
  assign n20798 = n7317 ^ n2840 ^ n1211 ;
  assign n20796 = n12288 | n19994 ;
  assign n20797 = n20796 ^ n9944 ^ 1'b0 ;
  assign n20799 = n20798 ^ n20797 ^ 1'b0 ;
  assign n20800 = n17035 & ~n20799 ;
  assign n20801 = n7837 & n12088 ;
  assign n20802 = n20801 ^ n9472 ^ 1'b0 ;
  assign n20803 = n7191 & ~n12116 ;
  assign n20804 = n20803 ^ n8518 ^ 1'b0 ;
  assign n20805 = n20804 ^ n7024 ^ 1'b0 ;
  assign n20806 = n5655 | n20805 ;
  assign n20807 = n20806 ^ x87 ^ 1'b0 ;
  assign n20808 = n11086 & n16827 ;
  assign n20809 = ~n20807 & n20808 ;
  assign n20810 = ( n14313 & ~n20802 ) | ( n14313 & n20809 ) | ( ~n20802 & n20809 ) ;
  assign n20811 = n7574 ^ n5125 ^ 1'b0 ;
  assign n20812 = ~n18922 & n20811 ;
  assign n20813 = n6607 ^ x59 ^ 1'b0 ;
  assign n20814 = n3613 | n20813 ;
  assign n20815 = ~n1513 & n20814 ;
  assign n20816 = n3795 & n7884 ;
  assign n20817 = n20315 ^ n14758 ^ n7218 ;
  assign n20818 = ( ~n5751 & n6566 ) | ( ~n5751 & n8580 ) | ( n6566 & n8580 ) ;
  assign n20819 = ~n13092 & n20818 ;
  assign n20820 = ~n3543 & n20819 ;
  assign n20821 = ( n15523 & n20817 ) | ( n15523 & n20820 ) | ( n20817 & n20820 ) ;
  assign n20822 = ( ~n10478 & n14571 ) | ( ~n10478 & n20821 ) | ( n14571 & n20821 ) ;
  assign n20823 = n20822 ^ n583 ^ 1'b0 ;
  assign n20824 = n13571 ^ n12014 ^ n3347 ;
  assign n20825 = n8566 | n20824 ;
  assign n20826 = n5499 & ~n20825 ;
  assign n20827 = n20826 ^ n14097 ^ 1'b0 ;
  assign n20828 = x176 & ~n20827 ;
  assign n20829 = n20828 ^ n757 ^ 1'b0 ;
  assign n20830 = n3230 | n3856 ;
  assign n20831 = n20830 ^ n7031 ^ n5107 ;
  assign n20832 = n2567 ^ n1763 ^ 1'b0 ;
  assign n20833 = ~n2523 & n20832 ;
  assign n20834 = n20833 ^ n608 ^ 1'b0 ;
  assign n20835 = ~n20831 & n20834 ;
  assign n20836 = ( n4042 & ~n4089 ) | ( n4042 & n5755 ) | ( ~n4089 & n5755 ) ;
  assign n20837 = n20836 ^ n1907 ^ n1192 ;
  assign n20838 = n11428 ^ n11118 ^ 1'b0 ;
  assign n20839 = ~n8630 & n20838 ;
  assign n20840 = ( n936 & n8655 ) | ( n936 & n8828 ) | ( n8655 & n8828 ) ;
  assign n20841 = n20840 ^ n2704 ^ 1'b0 ;
  assign n20842 = n8068 & ~n18538 ;
  assign n20843 = n13201 | n20842 ;
  assign n20844 = n20843 ^ n15603 ^ 1'b0 ;
  assign n20845 = n6384 & n11704 ;
  assign n20846 = n7713 ^ n2336 ^ 1'b0 ;
  assign n20847 = ~n6891 & n20846 ;
  assign n20848 = n20847 ^ n18495 ^ n734 ;
  assign n20849 = n3604 | n14782 ;
  assign n20850 = n20848 & ~n20849 ;
  assign n20851 = ( n3030 & n16268 ) | ( n3030 & ~n20850 ) | ( n16268 & ~n20850 ) ;
  assign n20852 = ~n20845 & n20851 ;
  assign n20853 = ~n12946 & n20852 ;
  assign n20854 = ~n11294 & n11572 ;
  assign n20855 = n6495 ^ n2693 ^ n656 ;
  assign n20856 = ( ~n3507 & n7140 ) | ( ~n3507 & n20855 ) | ( n7140 & n20855 ) ;
  assign n20857 = n11956 ^ n6168 ^ 1'b0 ;
  assign n20858 = n1093 & ~n20857 ;
  assign n20859 = ( n8235 & n10612 ) | ( n8235 & ~n20858 ) | ( n10612 & ~n20858 ) ;
  assign n20860 = ( n5889 & n20856 ) | ( n5889 & n20859 ) | ( n20856 & n20859 ) ;
  assign n20861 = n20860 ^ n1191 ^ 1'b0 ;
  assign n20862 = ( x221 & ~n818 ) | ( x221 & n849 ) | ( ~n818 & n849 ) ;
  assign n20863 = ~n8076 & n13223 ;
  assign n20864 = n20863 ^ n4540 ^ 1'b0 ;
  assign n20865 = n4419 | n20864 ;
  assign n20866 = n20865 ^ x26 ^ 1'b0 ;
  assign n20867 = n20866 ^ n19053 ^ x208 ;
  assign n20868 = ( ~n4204 & n20862 ) | ( ~n4204 & n20867 ) | ( n20862 & n20867 ) ;
  assign n20874 = ( n3902 & n4666 ) | ( n3902 & n11480 ) | ( n4666 & n11480 ) ;
  assign n20875 = ~n2509 & n8447 ;
  assign n20876 = n20875 ^ n6555 ^ 1'b0 ;
  assign n20877 = n5607 ^ n4016 ^ 1'b0 ;
  assign n20878 = ~n5239 & n20877 ;
  assign n20879 = n20878 ^ x103 ^ 1'b0 ;
  assign n20880 = n18670 & n20879 ;
  assign n20881 = ( n20874 & n20876 ) | ( n20874 & ~n20880 ) | ( n20876 & ~n20880 ) ;
  assign n20869 = n14090 ^ n10531 ^ n8204 ;
  assign n20870 = n20869 ^ n9764 ^ n4641 ;
  assign n20871 = n20870 ^ n15994 ^ n6832 ;
  assign n20872 = n20871 ^ n17687 ^ 1'b0 ;
  assign n20873 = n15556 | n20872 ;
  assign n20882 = n20881 ^ n20873 ^ 1'b0 ;
  assign n20885 = ( n4830 & n7135 ) | ( n4830 & ~n11122 ) | ( n7135 & ~n11122 ) ;
  assign n20883 = n282 & n3026 ;
  assign n20884 = n8975 & n20883 ;
  assign n20886 = n20885 ^ n20884 ^ n7089 ;
  assign n20887 = ( ~n4966 & n5840 ) | ( ~n4966 & n7439 ) | ( n5840 & n7439 ) ;
  assign n20888 = ( n1873 & n6406 ) | ( n1873 & ~n19609 ) | ( n6406 & ~n19609 ) ;
  assign n20889 = n20887 & ~n20888 ;
  assign n20890 = ~n11680 & n20889 ;
  assign n20891 = n20886 & n20890 ;
  assign n20892 = n11165 | n13738 ;
  assign n20893 = n11044 ^ n8677 ^ 1'b0 ;
  assign n20894 = n20893 ^ n13758 ^ n5559 ;
  assign n20895 = n12312 ^ n4414 ^ 1'b0 ;
  assign n20896 = n1363 | n20895 ;
  assign n20897 = ~n11093 & n12883 ;
  assign n20898 = n2119 & n20897 ;
  assign n20899 = ~n1037 & n20898 ;
  assign n20900 = ( ~n20894 & n20896 ) | ( ~n20894 & n20899 ) | ( n20896 & n20899 ) ;
  assign n20901 = ~n9473 & n18206 ;
  assign n20902 = ~n12111 & n20901 ;
  assign n20903 = n14522 ^ n8658 ^ 1'b0 ;
  assign n20904 = ( n579 & ~n4507 ) | ( n579 & n14697 ) | ( ~n4507 & n14697 ) ;
  assign n20905 = ~n20128 & n20904 ;
  assign n20906 = n9398 & n14671 ;
  assign n20907 = ~n2011 & n20906 ;
  assign n20908 = n20907 ^ x90 ^ 1'b0 ;
  assign n20909 = n20905 | n20908 ;
  assign n20910 = ( n4498 & n4937 ) | ( n4498 & n8461 ) | ( n4937 & n8461 ) ;
  assign n20911 = ( ~n816 & n3967 ) | ( ~n816 & n14671 ) | ( n3967 & n14671 ) ;
  assign n20912 = ( n2947 & n9341 ) | ( n2947 & ~n20911 ) | ( n9341 & ~n20911 ) ;
  assign n20913 = n20912 ^ n17329 ^ 1'b0 ;
  assign n20914 = n20910 | n20913 ;
  assign n20915 = ~n5926 & n12634 ;
  assign n20916 = ~n8469 & n20915 ;
  assign n20917 = n20916 ^ n12109 ^ 1'b0 ;
  assign n20918 = x181 & n17113 ;
  assign n20919 = n20918 ^ n3801 ^ 1'b0 ;
  assign n20920 = n20919 ^ n11855 ^ n9929 ;
  assign n20922 = n10581 ^ n4028 ^ 1'b0 ;
  assign n20923 = n3196 | n20922 ;
  assign n20921 = n3125 ^ n2682 ^ n2499 ;
  assign n20924 = n20923 ^ n20921 ^ n18989 ;
  assign n20925 = ~n12615 & n19327 ;
  assign n20926 = n20925 ^ n3411 ^ 1'b0 ;
  assign n20927 = n12383 & ~n17828 ;
  assign n20928 = n20524 & n20927 ;
  assign n20929 = ( ~n3697 & n7151 ) | ( ~n3697 & n20351 ) | ( n7151 & n20351 ) ;
  assign n20930 = n5126 & ~n6891 ;
  assign n20931 = ~n10077 & n20930 ;
  assign n20932 = n9457 | n10107 ;
  assign n20933 = n9479 | n20932 ;
  assign n20934 = n5436 & n20933 ;
  assign n20935 = ( n4340 & n20931 ) | ( n4340 & n20934 ) | ( n20931 & n20934 ) ;
  assign n20939 = ~n2317 & n15357 ;
  assign n20940 = n20939 ^ n9633 ^ 1'b0 ;
  assign n20941 = n14776 | n20940 ;
  assign n20936 = n2709 & ~n6136 ;
  assign n20937 = n20936 ^ n13628 ^ n5749 ;
  assign n20938 = n7692 | n20937 ;
  assign n20942 = n20941 ^ n20938 ^ 1'b0 ;
  assign n20943 = n5508 & n20942 ;
  assign n20944 = n3332 & ~n20816 ;
  assign n20945 = n20943 & n20944 ;
  assign n20946 = ~n5571 & n14364 ;
  assign n20947 = ( n4163 & n10163 ) | ( n4163 & ~n12293 ) | ( n10163 & ~n12293 ) ;
  assign n20948 = n6100 & n20947 ;
  assign n20949 = n20948 ^ n16058 ^ n10789 ;
  assign n20950 = n9337 ^ n5793 ^ 1'b0 ;
  assign n20951 = n578 & n20950 ;
  assign n20952 = ( n5316 & n13419 ) | ( n5316 & n20951 ) | ( n13419 & n20951 ) ;
  assign n20953 = n11029 & n20855 ;
  assign n20954 = ~n20952 & n20953 ;
  assign n20955 = n6515 ^ n2638 ^ 1'b0 ;
  assign n20956 = n552 | n20955 ;
  assign n20957 = n20956 ^ n16711 ^ n5441 ;
  assign n20958 = n3258 | n4153 ;
  assign n20959 = n9302 & ~n20958 ;
  assign n20962 = ( n499 & n5272 ) | ( n499 & ~n18382 ) | ( n5272 & ~n18382 ) ;
  assign n20963 = n6598 & n12635 ;
  assign n20964 = ~n10928 & n20963 ;
  assign n20965 = ~n20962 & n20964 ;
  assign n20960 = n11937 | n17522 ;
  assign n20961 = n20960 ^ n12304 ^ 1'b0 ;
  assign n20966 = n20965 ^ n20961 ^ 1'b0 ;
  assign n20967 = n20670 ^ n11156 ^ 1'b0 ;
  assign n20968 = ~n3830 & n20967 ;
  assign n20969 = n9113 & n11057 ;
  assign n20970 = ~x184 & n20969 ;
  assign n20971 = n9145 & ~n20970 ;
  assign n20972 = ~n8105 & n20971 ;
  assign n20973 = ( ~n16512 & n20968 ) | ( ~n16512 & n20972 ) | ( n20968 & n20972 ) ;
  assign n20974 = ( x173 & ~n595 ) | ( x173 & n12991 ) | ( ~n595 & n12991 ) ;
  assign n20975 = n20974 ^ n3159 ^ 1'b0 ;
  assign n20976 = n12073 & n20975 ;
  assign n20977 = ( n4594 & n7523 ) | ( n4594 & n19404 ) | ( n7523 & n19404 ) ;
  assign n20978 = n19319 ^ n3713 ^ 1'b0 ;
  assign n20979 = n14708 | n20978 ;
  assign n20980 = n20979 ^ n10024 ^ 1'b0 ;
  assign n20981 = ~n20977 & n20980 ;
  assign n20982 = ( n2484 & ~n6697 ) | ( n2484 & n10163 ) | ( ~n6697 & n10163 ) ;
  assign n20983 = n7913 | n20982 ;
  assign n20984 = n20983 ^ n6238 ^ 1'b0 ;
  assign n20985 = n1932 | n3133 ;
  assign n20986 = n20985 ^ n6586 ^ 1'b0 ;
  assign n20987 = ~n17971 & n20986 ;
  assign n20988 = n1406 & n20987 ;
  assign n20989 = n20988 ^ n14379 ^ n6560 ;
  assign n20990 = n4238 & n6615 ;
  assign n20991 = n20990 ^ n5143 ^ 1'b0 ;
  assign n20992 = ~n10869 & n20991 ;
  assign n20993 = n4137 ^ n1759 ^ 1'b0 ;
  assign n20994 = x246 & ~n12459 ;
  assign n20995 = n7759 ^ n5524 ^ n1950 ;
  assign n20996 = ~n15727 & n20995 ;
  assign n20998 = n4067 & n8297 ;
  assign n20999 = ~n1812 & n20998 ;
  assign n21000 = n19708 & n20999 ;
  assign n20997 = n523 & ~n8659 ;
  assign n21001 = n21000 ^ n20997 ^ 1'b0 ;
  assign n21002 = n19960 ^ n17952 ^ n5816 ;
  assign n21009 = n17239 ^ n5662 ^ 1'b0 ;
  assign n21010 = ~n18402 & n21009 ;
  assign n21011 = ( n8881 & n13624 ) | ( n8881 & n21010 ) | ( n13624 & n21010 ) ;
  assign n21012 = n21011 ^ n7201 ^ n1277 ;
  assign n21013 = ~n2246 & n5635 ;
  assign n21014 = n21013 ^ n5474 ^ 1'b0 ;
  assign n21015 = n21014 ^ n2486 ^ 1'b0 ;
  assign n21016 = n8631 | n21015 ;
  assign n21017 = ~n9743 & n19120 ;
  assign n21018 = n21016 & n21017 ;
  assign n21019 = n21012 | n21018 ;
  assign n21020 = n626 | n21019 ;
  assign n21003 = ~n8803 & n9754 ;
  assign n21004 = n13528 & n21003 ;
  assign n21005 = n6526 & ~n21004 ;
  assign n21006 = n21005 ^ n2322 ^ 1'b0 ;
  assign n21007 = n21006 ^ n4864 ^ 1'b0 ;
  assign n21008 = ~n9598 & n21007 ;
  assign n21021 = n21020 ^ n21008 ^ 1'b0 ;
  assign n21022 = x42 & ~n1401 ;
  assign n21023 = n16153 ^ n12776 ^ 1'b0 ;
  assign n21024 = x248 & ~n21023 ;
  assign n21025 = n21024 ^ n10968 ^ 1'b0 ;
  assign n21026 = ( n13950 & ~n21022 ) | ( n13950 & n21025 ) | ( ~n21022 & n21025 ) ;
  assign n21027 = n21026 ^ n9394 ^ 1'b0 ;
  assign n21028 = n21027 ^ n923 ^ 1'b0 ;
  assign n21029 = n14401 ^ n6046 ^ 1'b0 ;
  assign n21030 = n19940 & ~n21029 ;
  assign n21031 = n11591 ^ n11111 ^ n1214 ;
  assign n21032 = ( n1570 & n12421 ) | ( n1570 & n21031 ) | ( n12421 & n21031 ) ;
  assign n21034 = n2286 & ~n9531 ;
  assign n21033 = x238 & ~n20338 ;
  assign n21035 = n21034 ^ n21033 ^ 1'b0 ;
  assign n21036 = ~n4557 & n4653 ;
  assign n21037 = n6390 & ~n21036 ;
  assign n21038 = n21037 ^ n17345 ^ 1'b0 ;
  assign n21039 = ~n10763 & n14791 ;
  assign n21040 = n2890 & n8733 ;
  assign n21041 = ~n6666 & n21040 ;
  assign n21043 = n9618 ^ n1640 ^ n343 ;
  assign n21042 = n20192 ^ n10852 ^ n3921 ;
  assign n21044 = n21043 ^ n21042 ^ n2616 ;
  assign n21048 = n2047 ^ n988 ^ 1'b0 ;
  assign n21045 = n1501 | n2924 ;
  assign n21046 = n21045 ^ n6606 ^ 1'b0 ;
  assign n21047 = n5107 & ~n21046 ;
  assign n21049 = n21048 ^ n21047 ^ 1'b0 ;
  assign n21050 = n21049 ^ n9131 ^ 1'b0 ;
  assign n21051 = n5850 | n21050 ;
  assign n21052 = n21051 ^ n8688 ^ 1'b0 ;
  assign n21053 = n21052 ^ n14963 ^ n6163 ;
  assign n21054 = n3940 ^ n2793 ^ 1'b0 ;
  assign n21055 = ~n7727 & n21054 ;
  assign n21056 = n19656 & n21055 ;
  assign n21057 = ~n8285 & n21056 ;
  assign n21058 = ( ~n7762 & n15587 ) | ( ~n7762 & n18256 ) | ( n15587 & n18256 ) ;
  assign n21059 = n10626 ^ n9603 ^ n3754 ;
  assign n21060 = n21059 ^ n9365 ^ 1'b0 ;
  assign n21061 = n13945 & n21060 ;
  assign n21062 = x89 & ~n7738 ;
  assign n21063 = n21062 ^ n16544 ^ 1'b0 ;
  assign n21064 = n884 | n21063 ;
  assign n21065 = ( n1489 & n7192 ) | ( n1489 & ~n7706 ) | ( n7192 & ~n7706 ) ;
  assign n21066 = n15348 & ~n21065 ;
  assign n21067 = n21066 ^ n10104 ^ 1'b0 ;
  assign n21068 = ( ~n4180 & n4557 ) | ( ~n4180 & n21067 ) | ( n4557 & n21067 ) ;
  assign n21069 = ( n6683 & ~n15835 ) | ( n6683 & n18233 ) | ( ~n15835 & n18233 ) ;
  assign n21070 = n21069 ^ n15855 ^ 1'b0 ;
  assign n21071 = n13456 ^ n4794 ^ 1'b0 ;
  assign n21072 = n17498 ^ n15373 ^ 1'b0 ;
  assign n21073 = n21071 | n21072 ;
  assign n21075 = ( n8163 & n8751 ) | ( n8163 & n19579 ) | ( n8751 & n19579 ) ;
  assign n21074 = n8717 ^ n5743 ^ 1'b0 ;
  assign n21076 = n21075 ^ n21074 ^ 1'b0 ;
  assign n21077 = n13321 | n21076 ;
  assign n21078 = ( n6064 & n14082 ) | ( n6064 & n21077 ) | ( n14082 & n21077 ) ;
  assign n21079 = ( n6708 & n11300 ) | ( n6708 & ~n21078 ) | ( n11300 & ~n21078 ) ;
  assign n21080 = n18457 ^ n10193 ^ 1'b0 ;
  assign n21081 = ~n7367 & n21080 ;
  assign n21082 = n21081 ^ n20739 ^ n12826 ;
  assign n21083 = ( n3368 & n11718 ) | ( n3368 & ~n18370 ) | ( n11718 & ~n18370 ) ;
  assign n21084 = n11367 ^ n5797 ^ 1'b0 ;
  assign n21085 = n8468 | n21084 ;
  assign n21086 = n19308 & ~n21085 ;
  assign n21087 = ~n21083 & n21086 ;
  assign n21088 = n8854 ^ x242 ^ 1'b0 ;
  assign n21089 = n21087 | n21088 ;
  assign n21090 = n11251 ^ x236 ^ 1'b0 ;
  assign n21091 = ( n7401 & ~n16924 ) | ( n7401 & n21090 ) | ( ~n16924 & n21090 ) ;
  assign n21092 = n8462 | n21091 ;
  assign n21093 = n15543 | n21092 ;
  assign n21094 = n4077 ^ n2434 ^ n2389 ;
  assign n21095 = n4476 | n10372 ;
  assign n21096 = n21094 | n21095 ;
  assign n21097 = n21096 ^ n16894 ^ n9633 ;
  assign n21098 = n12249 & n21097 ;
  assign n21099 = ~n20780 & n21098 ;
  assign n21100 = n21099 ^ n10104 ^ n1268 ;
  assign n21101 = n5276 & ~n11165 ;
  assign n21104 = ~n1012 & n2530 ;
  assign n21105 = n19924 & n21104 ;
  assign n21102 = n2066 & ~n14824 ;
  assign n21103 = n13976 & n21102 ;
  assign n21106 = n21105 ^ n21103 ^ 1'b0 ;
  assign n21107 = ( ~n4629 & n10404 ) | ( ~n4629 & n15525 ) | ( n10404 & n15525 ) ;
  assign n21108 = n5678 & n21107 ;
  assign n21109 = n7612 ^ n7246 ^ 1'b0 ;
  assign n21110 = ~n21108 & n21109 ;
  assign n21111 = n17926 ^ n14818 ^ n7083 ;
  assign n21112 = n3010 ^ x230 ^ 1'b0 ;
  assign n21115 = ( ~n7223 & n8937 ) | ( ~n7223 & n16255 ) | ( n8937 & n16255 ) ;
  assign n21113 = n18734 ^ n13764 ^ n3648 ;
  assign n21114 = ( n8786 & n12194 ) | ( n8786 & n21113 ) | ( n12194 & n21113 ) ;
  assign n21116 = n21115 ^ n21114 ^ n6216 ;
  assign n21117 = n1028 | n6458 ;
  assign n21118 = n4984 | n21117 ;
  assign n21119 = n21118 ^ n7697 ^ 1'b0 ;
  assign n21120 = n21119 ^ n10673 ^ 1'b0 ;
  assign n21121 = n13326 & ~n21120 ;
  assign n21122 = ( n7748 & n11161 ) | ( n7748 & n15230 ) | ( n11161 & n15230 ) ;
  assign n21123 = n503 | n1919 ;
  assign n21124 = n4930 & ~n8558 ;
  assign n21125 = n8754 & n21124 ;
  assign n21126 = n21125 ^ n12244 ^ n2068 ;
  assign n21127 = n320 | n6607 ;
  assign n21128 = n8554 ^ n8413 ^ n6207 ;
  assign n21129 = n21127 | n21128 ;
  assign n21130 = n15364 ^ n6736 ^ 1'b0 ;
  assign n21131 = ~n7929 & n15927 ;
  assign n21132 = n12335 & n18132 ;
  assign n21133 = ~n21131 & n21132 ;
  assign n21134 = n21133 ^ n19098 ^ n2270 ;
  assign n21135 = n21134 ^ n6021 ^ 1'b0 ;
  assign n21136 = n4956 | n5193 ;
  assign n21137 = n21136 ^ n12322 ^ 1'b0 ;
  assign n21138 = n16917 ^ n11953 ^ n5510 ;
  assign n21139 = n6209 & ~n21138 ;
  assign n21140 = n21139 ^ n14838 ^ 1'b0 ;
  assign n21141 = n18218 ^ n7152 ^ n2566 ;
  assign n21142 = n18683 & ~n21141 ;
  assign n21143 = n21142 ^ n14955 ^ 1'b0 ;
  assign n21144 = n5975 ^ n3037 ^ 1'b0 ;
  assign n21145 = n16248 | n21144 ;
  assign n21146 = n21145 ^ n19709 ^ n5238 ;
  assign n21147 = n12622 & ~n15200 ;
  assign n21148 = n15041 ^ n14894 ^ 1'b0 ;
  assign n21149 = ( ~n15511 & n19852 ) | ( ~n15511 & n21148 ) | ( n19852 & n21148 ) ;
  assign n21150 = n11439 ^ n3655 ^ 1'b0 ;
  assign n21151 = n14377 ^ n10095 ^ 1'b0 ;
  assign n21152 = n8564 & ~n21151 ;
  assign n21153 = ~n19127 & n21152 ;
  assign n21154 = n10800 & n17911 ;
  assign n21155 = n17422 & ~n21154 ;
  assign n21156 = ~n21153 & n21155 ;
  assign n21157 = ~n2819 & n5608 ;
  assign n21158 = ( ~n3927 & n8530 ) | ( ~n3927 & n21157 ) | ( n8530 & n21157 ) ;
  assign n21159 = n18897 ^ n7428 ^ 1'b0 ;
  assign n21160 = n5820 ^ n2711 ^ 1'b0 ;
  assign n21161 = n4717 ^ n741 ^ 1'b0 ;
  assign n21162 = ~n5709 & n21161 ;
  assign n21163 = n21160 & n21162 ;
  assign n21164 = n21159 & n21163 ;
  assign n21165 = n11460 ^ n9249 ^ n1164 ;
  assign n21166 = n21165 ^ n10379 ^ 1'b0 ;
  assign n21167 = ( n5597 & n10559 ) | ( n5597 & n17117 ) | ( n10559 & n17117 ) ;
  assign n21168 = ( n8896 & n11044 ) | ( n8896 & ~n14170 ) | ( n11044 & ~n14170 ) ;
  assign n21169 = n6013 & n21168 ;
  assign n21170 = n11140 & ~n21169 ;
  assign n21171 = n1062 & n13844 ;
  assign n21172 = n14689 ^ n6296 ^ 1'b0 ;
  assign n21173 = ~n14807 & n18424 ;
  assign n21174 = n8448 & n8923 ;
  assign n21175 = n4476 & n21174 ;
  assign n21176 = n1091 & n1580 ;
  assign n21177 = n21176 ^ n15956 ^ 1'b0 ;
  assign n21178 = n18097 ^ n6199 ^ 1'b0 ;
  assign n21179 = n21178 ^ n10209 ^ n6553 ;
  assign n21180 = ( n16054 & ~n21177 ) | ( n16054 & n21179 ) | ( ~n21177 & n21179 ) ;
  assign n21181 = ~n8044 & n19695 ;
  assign n21182 = n18151 ^ n7490 ^ n1277 ;
  assign n21184 = n8775 ^ n3055 ^ 1'b0 ;
  assign n21185 = n10570 & n21184 ;
  assign n21186 = n12789 | n21185 ;
  assign n21183 = n660 | n7701 ;
  assign n21187 = n21186 ^ n21183 ^ n13092 ;
  assign n21188 = n9622 & n21187 ;
  assign n21189 = n21188 ^ n9056 ^ 1'b0 ;
  assign n21190 = ~n21182 & n21189 ;
  assign n21191 = n11683 & n18315 ;
  assign n21192 = n21191 ^ n8159 ^ 1'b0 ;
  assign n21193 = n21081 ^ x193 ^ 1'b0 ;
  assign n21194 = ( n7215 & n8369 ) | ( n7215 & n15247 ) | ( n8369 & n15247 ) ;
  assign n21195 = n20731 & n21194 ;
  assign n21196 = n4394 & n8811 ;
  assign n21197 = ~n10921 & n21196 ;
  assign n21198 = n908 & ~n12251 ;
  assign n21199 = x248 | n8496 ;
  assign n21200 = n21198 | n21199 ;
  assign n21201 = n6942 & n7170 ;
  assign n21202 = n21201 ^ n16191 ^ 1'b0 ;
  assign n21203 = n15827 | n16605 ;
  assign n21204 = n21202 | n21203 ;
  assign n21205 = n17484 ^ n13371 ^ n5706 ;
  assign n21206 = ( x184 & n2956 ) | ( x184 & n13718 ) | ( n2956 & n13718 ) ;
  assign n21207 = n4675 & n21206 ;
  assign n21208 = n21207 ^ n16001 ^ 1'b0 ;
  assign n21209 = n13317 & n21208 ;
  assign n21210 = n15041 ^ n8163 ^ n8029 ;
  assign n21211 = n479 & n6568 ;
  assign n21212 = ~n21210 & n21211 ;
  assign n21213 = ( ~x169 & n21209 ) | ( ~x169 & n21212 ) | ( n21209 & n21212 ) ;
  assign n21214 = n7270 ^ n4307 ^ 1'b0 ;
  assign n21215 = n14321 ^ n11159 ^ 1'b0 ;
  assign n21216 = n4970 & ~n21215 ;
  assign n21217 = ~n14095 & n21216 ;
  assign n21218 = n1159 & n21217 ;
  assign n21219 = n14731 ^ n11616 ^ 1'b0 ;
  assign n21220 = n9275 ^ n428 ^ x111 ;
  assign n21221 = n10659 & n21220 ;
  assign n21222 = ~n21219 & n21221 ;
  assign n21223 = n5078 ^ n2369 ^ 1'b0 ;
  assign n21224 = n19961 & ~n21223 ;
  assign n21225 = n2704 & n21224 ;
  assign n21226 = n21225 ^ n1355 ^ 1'b0 ;
  assign n21227 = n14443 & n21226 ;
  assign n21228 = n12414 ^ n9717 ^ 1'b0 ;
  assign n21229 = n21228 ^ n11093 ^ 1'b0 ;
  assign n21230 = n5076 & ~n16628 ;
  assign n21231 = ~n17911 & n21230 ;
  assign n21232 = ( n607 & n3665 ) | ( n607 & ~n4011 ) | ( n3665 & ~n4011 ) ;
  assign n21233 = n21232 ^ n1451 ^ 1'b0 ;
  assign n21234 = n21233 ^ n3336 ^ 1'b0 ;
  assign n21235 = n834 & n11912 ;
  assign n21236 = n9276 ^ n2628 ^ 1'b0 ;
  assign n21237 = n21236 ^ n9568 ^ n3453 ;
  assign n21238 = ( ~n3324 & n21235 ) | ( ~n3324 & n21237 ) | ( n21235 & n21237 ) ;
  assign n21239 = n11464 & n17960 ;
  assign n21244 = n10727 & n17362 ;
  assign n21243 = n3418 ^ n353 ^ 1'b0 ;
  assign n21245 = n21244 ^ n21243 ^ 1'b0 ;
  assign n21241 = n1764 & ~n16737 ;
  assign n21240 = n1617 | n9420 ;
  assign n21242 = n21241 ^ n21240 ^ 1'b0 ;
  assign n21246 = n21245 ^ n21242 ^ n4450 ;
  assign n21248 = n4934 ^ n4066 ^ 1'b0 ;
  assign n21247 = ( n15680 & ~n15973 ) | ( n15680 & n18668 ) | ( ~n15973 & n18668 ) ;
  assign n21249 = n21248 ^ n21247 ^ 1'b0 ;
  assign n21250 = ~n2573 & n21249 ;
  assign n21251 = n2359 | n8137 ;
  assign n21254 = n1995 | n9964 ;
  assign n21252 = n4760 ^ n726 ^ 1'b0 ;
  assign n21253 = n21252 ^ n9754 ^ 1'b0 ;
  assign n21255 = n21254 ^ n21253 ^ 1'b0 ;
  assign n21256 = n21251 | n21255 ;
  assign n21257 = n3479 | n20974 ;
  assign n21258 = n21257 ^ n21224 ^ 1'b0 ;
  assign n21259 = n2335 | n17000 ;
  assign n21260 = n7682 & ~n21259 ;
  assign n21261 = n17407 & ~n21260 ;
  assign n21262 = n16608 | n21261 ;
  assign n21263 = n21262 ^ n2836 ^ 1'b0 ;
  assign n21264 = n3376 ^ n3302 ^ 1'b0 ;
  assign n21265 = ~n3099 & n4238 ;
  assign n21266 = n21265 ^ n9911 ^ n4118 ;
  assign n21267 = ~n1217 & n5188 ;
  assign n21268 = n21267 ^ n16641 ^ 1'b0 ;
  assign n21269 = n21268 ^ n12098 ^ 1'b0 ;
  assign n21270 = n1390 & n8512 ;
  assign n21271 = n21270 ^ n4499 ^ 1'b0 ;
  assign n21272 = x127 & ~n989 ;
  assign n21273 = ~n17901 & n21272 ;
  assign n21274 = n291 & ~n16488 ;
  assign n21275 = n21274 ^ n9914 ^ n6353 ;
  assign n21276 = n21275 ^ n3967 ^ n3809 ;
  assign n21277 = ~n6128 & n8406 ;
  assign n21278 = n21277 ^ n4062 ^ 1'b0 ;
  assign n21279 = n4918 & ~n21278 ;
  assign n21280 = ( ~n21273 & n21276 ) | ( ~n21273 & n21279 ) | ( n21276 & n21279 ) ;
  assign n21281 = n8165 ^ n7510 ^ n6441 ;
  assign n21282 = n15820 ^ n5384 ^ 1'b0 ;
  assign n21283 = n2544 | n21282 ;
  assign n21284 = n21281 | n21283 ;
  assign n21285 = n21284 ^ n16822 ^ n2273 ;
  assign n21286 = n21285 ^ n15407 ^ n5317 ;
  assign n21287 = n3792 & ~n3960 ;
  assign n21288 = ~n21286 & n21287 ;
  assign n21289 = n6440 | n8405 ;
  assign n21290 = n19834 ^ n2562 ^ n1363 ;
  assign n21291 = ( ~n435 & n7743 ) | ( ~n435 & n21290 ) | ( n7743 & n21290 ) ;
  assign n21292 = ( n1197 & n2740 ) | ( n1197 & ~n9118 ) | ( n2740 & ~n9118 ) ;
  assign n21293 = n19830 ^ n18106 ^ n17126 ;
  assign n21294 = n12465 ^ n7405 ^ 1'b0 ;
  assign n21295 = n8805 | n21294 ;
  assign n21296 = n6279 | n21295 ;
  assign n21297 = n21296 ^ n7011 ^ 1'b0 ;
  assign n21298 = n10756 ^ n5261 ^ 1'b0 ;
  assign n21299 = n13424 | n21298 ;
  assign n21300 = ( n5799 & n21297 ) | ( n5799 & ~n21299 ) | ( n21297 & ~n21299 ) ;
  assign n21301 = ( n16844 & ~n18710 ) | ( n16844 & n21300 ) | ( ~n18710 & n21300 ) ;
  assign n21302 = n1568 ^ n607 ^ 1'b0 ;
  assign n21303 = n1949 & ~n21302 ;
  assign n21304 = n3583 & n21303 ;
  assign n21305 = ~n5539 & n21304 ;
  assign n21306 = n21305 ^ n430 ^ 1'b0 ;
  assign n21307 = ~n17762 & n21306 ;
  assign n21308 = ~n20553 & n21307 ;
  assign n21309 = n2699 | n17713 ;
  assign n21310 = n11181 ^ n10337 ^ 1'b0 ;
  assign n21311 = n21309 & n21310 ;
  assign n21314 = n9890 ^ n6021 ^ 1'b0 ;
  assign n21312 = n5272 & n6666 ;
  assign n21313 = ~n5026 & n21312 ;
  assign n21315 = n21314 ^ n21313 ^ 1'b0 ;
  assign n21316 = n9015 & ~n21315 ;
  assign n21317 = ( n6184 & n12576 ) | ( n6184 & ~n17366 ) | ( n12576 & ~n17366 ) ;
  assign n21318 = n21317 ^ n7178 ^ n3604 ;
  assign n21321 = n6108 ^ n3485 ^ 1'b0 ;
  assign n21319 = n5680 ^ n2634 ^ n997 ;
  assign n21320 = n9532 | n21319 ;
  assign n21322 = n21321 ^ n21320 ^ n2654 ;
  assign n21323 = ( n864 & ~n8819 ) | ( n864 & n21322 ) | ( ~n8819 & n21322 ) ;
  assign n21324 = n8515 & n21323 ;
  assign n21325 = ( n5937 & n12123 ) | ( n5937 & n13145 ) | ( n12123 & n13145 ) ;
  assign n21326 = n6928 ^ n4954 ^ 1'b0 ;
  assign n21327 = ( n10964 & n13034 ) | ( n10964 & n21326 ) | ( n13034 & n21326 ) ;
  assign n21328 = ~n2146 & n11548 ;
  assign n21329 = ~n7494 & n21328 ;
  assign n21330 = n21327 | n21329 ;
  assign n21331 = n2617 & ~n21330 ;
  assign n21332 = n16108 | n21331 ;
  assign n21333 = n15133 | n21332 ;
  assign n21334 = n3761 & ~n15063 ;
  assign n21335 = n7617 & n21334 ;
  assign n21336 = n20856 & ~n21335 ;
  assign n21337 = n19858 & n21336 ;
  assign n21338 = n4378 | n14588 ;
  assign n21339 = n18691 & ~n21338 ;
  assign n21340 = n10150 ^ n8517 ^ 1'b0 ;
  assign n21341 = ~n9732 & n14883 ;
  assign n21342 = n21340 & ~n21341 ;
  assign n21343 = n17651 ^ n10945 ^ 1'b0 ;
  assign n21344 = n3650 | n21343 ;
  assign n21345 = n2367 | n10919 ;
  assign n21346 = n21344 & ~n21345 ;
  assign n21347 = n2017 & n9504 ;
  assign n21348 = n21347 ^ n1776 ^ n1585 ;
  assign n21349 = n21348 ^ n473 ^ 1'b0 ;
  assign n21350 = n11549 & n21349 ;
  assign n21351 = n4818 | n21350 ;
  assign n21362 = n15044 ^ n14221 ^ 1'b0 ;
  assign n21359 = ~n1607 & n13303 ;
  assign n21360 = n21359 ^ n5723 ^ 1'b0 ;
  assign n21361 = ~n2635 & n21360 ;
  assign n21355 = n3229 & ~n18665 ;
  assign n21356 = n21355 ^ n14516 ^ n7329 ;
  assign n21353 = ( n6852 & n13857 ) | ( n6852 & ~n20923 ) | ( n13857 & ~n20923 ) ;
  assign n21354 = n21353 ^ n19614 ^ 1'b0 ;
  assign n21352 = ~n15682 & n19649 ;
  assign n21357 = n21356 ^ n21354 ^ n21352 ;
  assign n21358 = n21357 ^ n9304 ^ n6475 ;
  assign n21363 = n21362 ^ n21361 ^ n21358 ;
  assign n21364 = n2423 ^ n2073 ^ x190 ;
  assign n21365 = n11049 & ~n16112 ;
  assign n21366 = n21365 ^ n8942 ^ 1'b0 ;
  assign n21367 = n6266 & n21366 ;
  assign n21368 = ( n4187 & n6156 ) | ( n4187 & n21367 ) | ( n6156 & n21367 ) ;
  assign n21369 = n20473 ^ n12207 ^ 1'b0 ;
  assign n21370 = n21166 & n21369 ;
  assign n21372 = ~n2293 & n5490 ;
  assign n21373 = n1425 & n21372 ;
  assign n21371 = n1634 | n11356 ;
  assign n21374 = n21373 ^ n21371 ^ n19857 ;
  assign n21375 = n7050 ^ n4592 ^ n1206 ;
  assign n21376 = n1973 & ~n21375 ;
  assign n21377 = ~n3645 & n21376 ;
  assign n21379 = n13419 & ~n18531 ;
  assign n21378 = ( n804 & n868 ) | ( n804 & n18042 ) | ( n868 & n18042 ) ;
  assign n21380 = n21379 ^ n21378 ^ 1'b0 ;
  assign n21381 = ~n1853 & n9228 ;
  assign n21382 = n21381 ^ n3846 ^ 1'b0 ;
  assign n21383 = n21382 ^ n20598 ^ 1'b0 ;
  assign n21384 = n9287 & n21383 ;
  assign n21385 = n21384 ^ n13418 ^ 1'b0 ;
  assign n21386 = ( n10085 & ~n11592 ) | ( n10085 & n21385 ) | ( ~n11592 & n21385 ) ;
  assign n21387 = n13499 & ~n21386 ;
  assign n21388 = n15428 & n20358 ;
  assign n21389 = n7926 ^ n2460 ^ 1'b0 ;
  assign n21390 = n21389 ^ x197 ^ 1'b0 ;
  assign n21391 = n11766 & n21390 ;
  assign n21392 = n11001 ^ n1393 ^ 1'b0 ;
  assign n21393 = n7349 | n21392 ;
  assign n21394 = n21393 ^ n19526 ^ 1'b0 ;
  assign n21395 = ~n5176 & n21394 ;
  assign n21396 = n21395 ^ n9877 ^ 1'b0 ;
  assign n21397 = n8756 & ~n17640 ;
  assign n21401 = ( n1146 & n1934 ) | ( n1146 & n6531 ) | ( n1934 & n6531 ) ;
  assign n21402 = n7762 & ~n21401 ;
  assign n21403 = n5250 & n21402 ;
  assign n21398 = n17958 ^ n679 ^ 1'b0 ;
  assign n21399 = n13061 & n21398 ;
  assign n21400 = n6046 & n21399 ;
  assign n21404 = n21403 ^ n21400 ^ 1'b0 ;
  assign n21405 = n19347 ^ n7379 ^ n2388 ;
  assign n21406 = n16005 ^ n12726 ^ 1'b0 ;
  assign n21407 = ( n21404 & n21405 ) | ( n21404 & ~n21406 ) | ( n21405 & ~n21406 ) ;
  assign n21408 = ~n17617 & n19420 ;
  assign n21409 = n21408 ^ n19091 ^ n12666 ;
  assign n21410 = ( n2502 & ~n6701 ) | ( n2502 & n11349 ) | ( ~n6701 & n11349 ) ;
  assign n21411 = n21409 & n21410 ;
  assign n21412 = n8231 ^ n7852 ^ n6777 ;
  assign n21413 = ( n2160 & n4310 ) | ( n2160 & ~n21412 ) | ( n4310 & ~n21412 ) ;
  assign n21414 = n21413 ^ n2740 ^ 1'b0 ;
  assign n21415 = n21414 ^ n11150 ^ n8396 ;
  assign n21416 = n9605 ^ n7840 ^ 1'b0 ;
  assign n21417 = n21416 ^ n4728 ^ 1'b0 ;
  assign n21418 = x246 & n10559 ;
  assign n21419 = n6235 & n21418 ;
  assign n21420 = n7288 ^ n4638 ^ 1'b0 ;
  assign n21421 = n21419 & n21420 ;
  assign n21422 = n3982 & n14166 ;
  assign n21423 = n21422 ^ n1075 ^ 1'b0 ;
  assign n21424 = ~n20951 & n21423 ;
  assign n21425 = ( n424 & n7136 ) | ( n424 & n21424 ) | ( n7136 & n21424 ) ;
  assign n21431 = n6056 ^ n5523 ^ 1'b0 ;
  assign n21430 = ~n10851 & n15113 ;
  assign n21427 = ~n8548 & n21011 ;
  assign n21428 = ~n7854 & n21427 ;
  assign n21429 = ( n3782 & n5082 ) | ( n3782 & n21428 ) | ( n5082 & n21428 ) ;
  assign n21432 = n21431 ^ n21430 ^ n21429 ;
  assign n21426 = n8940 | n13272 ;
  assign n21433 = n21432 ^ n21426 ^ 1'b0 ;
  assign n21434 = n8429 ^ n6719 ^ 1'b0 ;
  assign n21435 = ~n3016 & n21434 ;
  assign n21436 = n9394 & n12230 ;
  assign n21437 = ~n6693 & n21436 ;
  assign n21438 = ( n2967 & n21435 ) | ( n2967 & n21437 ) | ( n21435 & n21437 ) ;
  assign n21439 = n11619 & ~n21438 ;
  assign n21440 = n6527 | n21125 ;
  assign n21441 = n16514 & ~n21440 ;
  assign n21442 = n19038 & n21441 ;
  assign n21443 = n19257 ^ n6204 ^ n1192 ;
  assign n21444 = n2399 & ~n18614 ;
  assign n21445 = ~n9015 & n21444 ;
  assign n21446 = n21445 ^ n16918 ^ 1'b0 ;
  assign n21447 = n4247 & ~n21446 ;
  assign n21453 = n2613 | n7943 ;
  assign n21454 = ( n14186 & n15183 ) | ( n14186 & ~n20763 ) | ( n15183 & ~n20763 ) ;
  assign n21455 = n13351 ^ n10003 ^ n4187 ;
  assign n21456 = ( n21453 & n21454 ) | ( n21453 & n21455 ) | ( n21454 & n21455 ) ;
  assign n21457 = ( n2081 & n4057 ) | ( n2081 & ~n21456 ) | ( n4057 & ~n21456 ) ;
  assign n21449 = n10563 ^ n9053 ^ n2151 ;
  assign n21448 = n12489 ^ n9343 ^ n7395 ;
  assign n21450 = n21449 ^ n21448 ^ 1'b0 ;
  assign n21451 = ~n11157 & n21450 ;
  assign n21452 = ~n7991 & n21451 ;
  assign n21458 = n21457 ^ n21452 ^ 1'b0 ;
  assign n21475 = ( x65 & n1345 ) | ( x65 & ~n12670 ) | ( n1345 & ~n12670 ) ;
  assign n21474 = n2858 & ~n11111 ;
  assign n21476 = n21475 ^ n21474 ^ 1'b0 ;
  assign n21462 = n11735 & ~n16141 ;
  assign n21463 = n3481 & n21462 ;
  assign n21464 = n21463 ^ n5987 ^ 1'b0 ;
  assign n21461 = n6488 & ~n18764 ;
  assign n21465 = n21464 ^ n21461 ^ 1'b0 ;
  assign n21459 = n8006 & n18063 ;
  assign n21460 = n21459 ^ n3416 ^ n2754 ;
  assign n21466 = n21465 ^ n21460 ^ 1'b0 ;
  assign n21469 = n4219 | n4528 ;
  assign n21470 = n10297 & ~n21469 ;
  assign n21471 = n1258 | n21470 ;
  assign n21467 = n5474 & n13976 ;
  assign n21468 = n21467 ^ n20711 ^ 1'b0 ;
  assign n21472 = n21471 ^ n21468 ^ 1'b0 ;
  assign n21473 = ~n21466 & n21472 ;
  assign n21477 = n21476 ^ n21473 ^ 1'b0 ;
  assign n21478 = n8836 ^ n3672 ^ 1'b0 ;
  assign n21479 = ~n4073 & n21478 ;
  assign n21480 = n8887 | n21479 ;
  assign n21481 = n541 | n6763 ;
  assign n21482 = n3322 | n21481 ;
  assign n21483 = n8073 | n18763 ;
  assign n21484 = n21482 | n21483 ;
  assign n21485 = n8230 ^ n2353 ^ x161 ;
  assign n21486 = x55 & n17823 ;
  assign n21487 = n21486 ^ n21118 ^ 1'b0 ;
  assign n21488 = n21319 ^ n14086 ^ n7834 ;
  assign n21489 = ( ~n11103 & n16170 ) | ( ~n11103 & n21488 ) | ( n16170 & n21488 ) ;
  assign n21490 = n21487 & ~n21489 ;
  assign n21491 = ( n8813 & ~n16656 ) | ( n8813 & n21490 ) | ( ~n16656 & n21490 ) ;
  assign n21492 = n7370 | n9546 ;
  assign n21493 = n10797 & ~n21492 ;
  assign n21494 = ~n5509 & n19462 ;
  assign n21495 = ( ~n2905 & n6156 ) | ( ~n2905 & n21494 ) | ( n6156 & n21494 ) ;
  assign n21496 = n3144 & ~n6787 ;
  assign n21510 = n11518 ^ n9095 ^ 1'b0 ;
  assign n21497 = ( ~x156 & n3428 ) | ( ~x156 & n15446 ) | ( n3428 & n15446 ) ;
  assign n21502 = n16112 ^ n2606 ^ 1'b0 ;
  assign n21498 = n5629 ^ x13 ^ 1'b0 ;
  assign n21499 = ~n537 & n21498 ;
  assign n21500 = n21499 ^ n7257 ^ 1'b0 ;
  assign n21501 = ( n2122 & n4550 ) | ( n2122 & ~n21500 ) | ( n4550 & ~n21500 ) ;
  assign n21503 = n21502 ^ n21501 ^ n11601 ;
  assign n21506 = n7383 ^ n2412 ^ 1'b0 ;
  assign n21504 = n15302 ^ n4369 ^ n1296 ;
  assign n21505 = ( ~n3483 & n7669 ) | ( ~n3483 & n21504 ) | ( n7669 & n21504 ) ;
  assign n21507 = n21506 ^ n21505 ^ 1'b0 ;
  assign n21508 = n21503 | n21507 ;
  assign n21509 = ( ~n15556 & n21497 ) | ( ~n15556 & n21508 ) | ( n21497 & n21508 ) ;
  assign n21511 = n21510 ^ n21509 ^ 1'b0 ;
  assign n21512 = n21496 & ~n21511 ;
  assign n21513 = ( n6666 & ~n16502 ) | ( n6666 & n19956 ) | ( ~n16502 & n19956 ) ;
  assign n21514 = n18839 ^ n11124 ^ n6081 ;
  assign n21515 = n11257 ^ n7464 ^ n5504 ;
  assign n21516 = n21515 ^ n20266 ^ 1'b0 ;
  assign n21517 = n18264 & n21516 ;
  assign n21518 = n1730 ^ n1496 ^ 1'b0 ;
  assign n21519 = n14910 & ~n21518 ;
  assign n21520 = n2699 & n3641 ;
  assign n21521 = ( n7402 & n16268 ) | ( n7402 & n21520 ) | ( n16268 & n21520 ) ;
  assign n21522 = n13183 ^ n3557 ^ 1'b0 ;
  assign n21523 = n21522 ^ n6197 ^ n3068 ;
  assign n21524 = n4779 | n21523 ;
  assign n21525 = n3764 & ~n21524 ;
  assign n21527 = n7403 ^ n2077 ^ 1'b0 ;
  assign n21526 = n4443 | n21014 ;
  assign n21528 = n21527 ^ n21526 ^ 1'b0 ;
  assign n21529 = n1099 & n11285 ;
  assign n21530 = n13996 & ~n18876 ;
  assign n21531 = n17708 & n21530 ;
  assign n21532 = ~n4097 & n7790 ;
  assign n21533 = ( n1469 & ~n8132 ) | ( n1469 & n21532 ) | ( ~n8132 & n21532 ) ;
  assign n21534 = n21533 ^ n20362 ^ n16280 ;
  assign n21535 = ~n6940 & n19317 ;
  assign n21536 = ( n13223 & ~n14007 ) | ( n13223 & n16271 ) | ( ~n14007 & n16271 ) ;
  assign n21537 = n10527 ^ n4958 ^ n3359 ;
  assign n21538 = n21537 ^ n13398 ^ 1'b0 ;
  assign n21539 = n21536 | n21538 ;
  assign n21540 = n21539 ^ n963 ^ 1'b0 ;
  assign n21541 = ~n639 & n5086 ;
  assign n21542 = n21541 ^ n8297 ^ 1'b0 ;
  assign n21543 = ( ~n5418 & n14030 ) | ( ~n5418 & n21542 ) | ( n14030 & n21542 ) ;
  assign n21544 = n21543 ^ n1469 ^ 1'b0 ;
  assign n21545 = n12457 | n20502 ;
  assign n21546 = n21545 ^ n13317 ^ 1'b0 ;
  assign n21547 = n10202 ^ n9671 ^ n6941 ;
  assign n21548 = ( n1264 & n2021 ) | ( n1264 & ~n5022 ) | ( n2021 & ~n5022 ) ;
  assign n21549 = n3637 ^ n1743 ^ 1'b0 ;
  assign n21550 = n14349 & ~n21549 ;
  assign n21551 = ~n8292 & n21550 ;
  assign n21552 = n21551 ^ n14617 ^ n5441 ;
  assign n21553 = n21552 ^ n16761 ^ 1'b0 ;
  assign n21554 = n15550 ^ n4443 ^ 1'b0 ;
  assign n21555 = n21554 ^ n9168 ^ n3297 ;
  assign n21556 = n21555 ^ n19721 ^ 1'b0 ;
  assign n21557 = n14151 & n21556 ;
  assign n21558 = ~n14157 & n14166 ;
  assign n21559 = n21558 ^ n13317 ^ 1'b0 ;
  assign n21560 = n13204 ^ n4360 ^ 1'b0 ;
  assign n21561 = ( n2893 & ~n7510 ) | ( n2893 & n21560 ) | ( ~n7510 & n21560 ) ;
  assign n21562 = ( n1485 & n10445 ) | ( n1485 & ~n21561 ) | ( n10445 & ~n21561 ) ;
  assign n21563 = ( ~n8413 & n16236 ) | ( ~n8413 & n21562 ) | ( n16236 & n21562 ) ;
  assign n21564 = n8946 ^ n2423 ^ n1510 ;
  assign n21565 = n3776 & ~n4410 ;
  assign n21566 = n21565 ^ n21236 ^ 1'b0 ;
  assign n21567 = ~n19893 & n21566 ;
  assign n21568 = ( ~n3819 & n9524 ) | ( ~n3819 & n18402 ) | ( n9524 & n18402 ) ;
  assign n21569 = n21568 ^ n9199 ^ n2815 ;
  assign n21570 = ( n14533 & ~n14816 ) | ( n14533 & n21569 ) | ( ~n14816 & n21569 ) ;
  assign n21571 = n6472 & ~n14945 ;
  assign n21572 = n11212 ^ n8410 ^ n7046 ;
  assign n21573 = ( n378 & n11794 ) | ( n378 & ~n19499 ) | ( n11794 & ~n19499 ) ;
  assign n21574 = n21573 ^ n17474 ^ n11738 ;
  assign n21575 = n9827 ^ n2032 ^ 1'b0 ;
  assign n21576 = x1 & n21575 ;
  assign n21577 = n10479 & ~n21576 ;
  assign n21578 = ( n345 & n4503 ) | ( n345 & n11348 ) | ( n4503 & n11348 ) ;
  assign n21579 = ( n16175 & ~n21577 ) | ( n16175 & n21578 ) | ( ~n21577 & n21578 ) ;
  assign n21580 = n3862 ^ n397 ^ n311 ;
  assign n21581 = n21580 ^ n13943 ^ n8691 ;
  assign n21582 = ( n1292 & ~n2052 ) | ( n1292 & n3112 ) | ( ~n2052 & n3112 ) ;
  assign n21583 = n21582 ^ n11263 ^ 1'b0 ;
  assign n21584 = ~n21581 & n21583 ;
  assign n21585 = n443 & ~n3905 ;
  assign n21586 = n21585 ^ n13721 ^ 1'b0 ;
  assign n21587 = ~n7900 & n13698 ;
  assign n21588 = ~n1270 & n3771 ;
  assign n21589 = n21588 ^ n3316 ^ 1'b0 ;
  assign n21590 = n21589 ^ n15969 ^ n10474 ;
  assign n21591 = n2199 & ~n4982 ;
  assign n21592 = n5389 & n21591 ;
  assign n21593 = ~n6423 & n6470 ;
  assign n21594 = ~n13905 & n21593 ;
  assign n21595 = n12311 ^ n915 ^ 1'b0 ;
  assign n21596 = n10699 ^ n2839 ^ 1'b0 ;
  assign n21597 = ~n2061 & n21596 ;
  assign n21598 = n21597 ^ n19607 ^ 1'b0 ;
  assign n21599 = ( ~n1806 & n16483 ) | ( ~n1806 & n16978 ) | ( n16483 & n16978 ) ;
  assign n21600 = ~n7882 & n13236 ;
  assign n21601 = ~n10045 & n21600 ;
  assign n21602 = n1447 & ~n13969 ;
  assign n21603 = n8413 & n21602 ;
  assign n21604 = n12470 & ~n20136 ;
  assign n21605 = ~n14848 & n21604 ;
  assign n21606 = ( n4871 & n6458 ) | ( n4871 & ~n18420 ) | ( n6458 & ~n18420 ) ;
  assign n21607 = n4774 ^ n779 ^ 1'b0 ;
  assign n21608 = x3 & ~n21607 ;
  assign n21609 = ( n20015 & n21606 ) | ( n20015 & n21608 ) | ( n21606 & n21608 ) ;
  assign n21610 = n13915 ^ n8447 ^ 1'b0 ;
  assign n21611 = n3083 & ~n14398 ;
  assign n21612 = x50 & n21611 ;
  assign n21613 = ~n12080 & n19686 ;
  assign n21614 = n17438 & n21613 ;
  assign n21615 = ( n8593 & n15529 ) | ( n8593 & n17025 ) | ( n15529 & n17025 ) ;
  assign n21616 = x99 & ~n12239 ;
  assign n21617 = n2793 & n21616 ;
  assign n21618 = n21617 ^ n10087 ^ n8097 ;
  assign n21619 = n11632 ^ n5474 ^ 1'b0 ;
  assign n21620 = n15750 ^ n4970 ^ 1'b0 ;
  assign n21621 = n7925 | n19511 ;
  assign n21622 = n1285 & n7741 ;
  assign n21623 = n13506 ^ n3380 ^ n3330 ;
  assign n21624 = ( n2469 & n21622 ) | ( n2469 & n21623 ) | ( n21622 & n21623 ) ;
  assign n21625 = ( n16650 & n21621 ) | ( n16650 & n21624 ) | ( n21621 & n21624 ) ;
  assign n21626 = n21625 ^ n14123 ^ n2280 ;
  assign n21627 = n8644 ^ x63 ^ 1'b0 ;
  assign n21628 = n17384 ^ n2389 ^ 1'b0 ;
  assign n21629 = n21628 ^ n7241 ^ n7239 ;
  assign n21630 = n5376 | n9089 ;
  assign n21631 = n21629 | n21630 ;
  assign n21633 = ( n1816 & n4231 ) | ( n1816 & ~n4928 ) | ( n4231 & ~n4928 ) ;
  assign n21634 = n21633 ^ n19927 ^ n10731 ;
  assign n21635 = n21634 ^ n18048 ^ n16552 ;
  assign n21632 = ~n12593 & n14740 ;
  assign n21636 = n21635 ^ n21632 ^ 1'b0 ;
  assign n21639 = n7354 | n20604 ;
  assign n21637 = n10335 ^ n4438 ^ n3446 ;
  assign n21638 = n21637 ^ n5874 ^ 1'b0 ;
  assign n21640 = n21639 ^ n21638 ^ x126 ;
  assign n21641 = n17049 ^ n5323 ^ 1'b0 ;
  assign n21642 = n9936 ^ n6641 ^ 1'b0 ;
  assign n21643 = n2321 & n9120 ;
  assign n21644 = n21643 ^ n2646 ^ 1'b0 ;
  assign n21645 = n2195 & n21644 ;
  assign n21646 = ~n12101 & n21645 ;
  assign n21647 = n21646 ^ n3887 ^ x175 ;
  assign n21648 = n21647 ^ n1406 ^ 1'b0 ;
  assign n21649 = ~n5311 & n21648 ;
  assign n21650 = n21642 | n21649 ;
  assign n21651 = n17297 ^ n5481 ^ x107 ;
  assign n21652 = ~n4053 & n16662 ;
  assign n21653 = n8230 & n21652 ;
  assign n21654 = n21653 ^ n11148 ^ n9044 ;
  assign n21655 = ~n5179 & n20249 ;
  assign n21656 = n21655 ^ n9217 ^ 1'b0 ;
  assign n21657 = n10354 ^ n2685 ^ 1'b0 ;
  assign n21658 = ~n10671 & n15322 ;
  assign n21659 = n21658 ^ n7375 ^ 1'b0 ;
  assign n21663 = n1826 | n19084 ;
  assign n21664 = n21663 ^ n7542 ^ 1'b0 ;
  assign n21660 = ( ~n2965 & n8198 ) | ( ~n2965 & n14139 ) | ( n8198 & n14139 ) ;
  assign n21661 = ~n7406 & n21660 ;
  assign n21662 = n1328 & n21661 ;
  assign n21665 = n21664 ^ n21662 ^ 1'b0 ;
  assign n21666 = n15967 ^ n7605 ^ 1'b0 ;
  assign n21667 = n21666 ^ n18171 ^ n3665 ;
  assign n21668 = n2730 & ~n20456 ;
  assign n21669 = ( n2255 & n4064 ) | ( n2255 & ~n9087 ) | ( n4064 & ~n9087 ) ;
  assign n21670 = ~n2075 & n21669 ;
  assign n21671 = ~n9015 & n21670 ;
  assign n21672 = n14054 & ~n21671 ;
  assign n21673 = n2721 & n21672 ;
  assign n21674 = n2811 & ~n5791 ;
  assign n21675 = n21674 ^ n14034 ^ 1'b0 ;
  assign n21676 = n12373 ^ n9997 ^ 1'b0 ;
  assign n21677 = n4237 | n8835 ;
  assign n21683 = n2386 & n8293 ;
  assign n21678 = n10265 ^ n8094 ^ n4438 ;
  assign n21679 = x101 & n13169 ;
  assign n21680 = n21678 & n21679 ;
  assign n21681 = n21680 ^ n13043 ^ n7442 ;
  assign n21682 = n17218 | n21681 ;
  assign n21684 = n21683 ^ n21682 ^ 1'b0 ;
  assign n21685 = n6384 | n15152 ;
  assign n21686 = n4924 | n21685 ;
  assign n21687 = ( n2252 & ~n6312 ) | ( n2252 & n21686 ) | ( ~n6312 & n21686 ) ;
  assign n21688 = n21687 ^ n11061 ^ 1'b0 ;
  assign n21690 = n1199 & n14829 ;
  assign n21689 = n2363 | n5905 ;
  assign n21691 = n21690 ^ n21689 ^ 1'b0 ;
  assign n21692 = ( n1598 & ~n8097 ) | ( n1598 & n11476 ) | ( ~n8097 & n11476 ) ;
  assign n21693 = ~n8414 & n21692 ;
  assign n21694 = n7081 & n21693 ;
  assign n21695 = n16720 ^ n3661 ^ 1'b0 ;
  assign n21696 = n19724 & ~n21695 ;
  assign n21697 = n8816 ^ n6809 ^ n6018 ;
  assign n21698 = ( n6847 & ~n11131 ) | ( n6847 & n21697 ) | ( ~n11131 & n21697 ) ;
  assign n21699 = n17431 ^ n1231 ^ 1'b0 ;
  assign n21700 = ~n20974 & n21699 ;
  assign n21701 = n21700 ^ n6594 ^ 1'b0 ;
  assign n21702 = n21698 & n21701 ;
  assign n21703 = ( n633 & n7130 ) | ( n633 & ~n9113 ) | ( n7130 & ~n9113 ) ;
  assign n21704 = n8114 | n13642 ;
  assign n21705 = n21704 ^ n1672 ^ 1'b0 ;
  assign n21706 = n9257 & n21705 ;
  assign n21707 = n21706 ^ n15926 ^ n8926 ;
  assign n21708 = ( ~n5100 & n11476 ) | ( ~n5100 & n21707 ) | ( n11476 & n21707 ) ;
  assign n21709 = ( x247 & n7248 ) | ( x247 & ~n7537 ) | ( n7248 & ~n7537 ) ;
  assign n21710 = n2092 & ~n21709 ;
  assign n21711 = n21710 ^ n19810 ^ 1'b0 ;
  assign n21712 = n11313 & ~n21711 ;
  assign n21713 = x53 & ~n7998 ;
  assign n21714 = ~n2943 & n21713 ;
  assign n21715 = ( n6103 & n21712 ) | ( n6103 & ~n21714 ) | ( n21712 & ~n21714 ) ;
  assign n21716 = ~n13285 & n15147 ;
  assign n21717 = n21716 ^ n3687 ^ 1'b0 ;
  assign n21718 = n18603 ^ n554 ^ 1'b0 ;
  assign n21719 = ~n4690 & n21718 ;
  assign n21720 = n20888 ^ n19419 ^ n8539 ;
  assign n21721 = ( n13581 & ~n21680 ) | ( n13581 & n21720 ) | ( ~n21680 & n21720 ) ;
  assign n21722 = ( n2745 & n8933 ) | ( n2745 & ~n10523 ) | ( n8933 & ~n10523 ) ;
  assign n21723 = n18237 & ~n21722 ;
  assign n21724 = ~n21721 & n21723 ;
  assign n21725 = n13699 & n15807 ;
  assign n21726 = ~n7910 & n21725 ;
  assign n21727 = n21726 ^ n8783 ^ n1352 ;
  assign n21729 = ( n1276 & n2666 ) | ( n1276 & ~n16003 ) | ( n2666 & ~n16003 ) ;
  assign n21728 = ( ~n6575 & n11112 ) | ( ~n6575 & n19478 ) | ( n11112 & n19478 ) ;
  assign n21730 = n21729 ^ n21728 ^ 1'b0 ;
  assign n21731 = n21730 ^ n257 ^ 1'b0 ;
  assign n21732 = n21727 & ~n21731 ;
  assign n21733 = n14813 & n21732 ;
  assign n21734 = ~n829 & n21733 ;
  assign n21735 = n19917 ^ n4307 ^ 1'b0 ;
  assign n21736 = n20046 ^ n10170 ^ 1'b0 ;
  assign n21737 = n2597 & n6804 ;
  assign n21738 = n21736 & n21737 ;
  assign n21739 = n7071 & n21738 ;
  assign n21744 = n17037 ^ n1383 ^ 1'b0 ;
  assign n21745 = n21744 ^ n3169 ^ n1133 ;
  assign n21740 = ~n2613 & n8047 ;
  assign n21741 = ~n1913 & n21740 ;
  assign n21742 = n21741 ^ n10993 ^ n8191 ;
  assign n21743 = n11350 & n21742 ;
  assign n21746 = n21745 ^ n21743 ^ 1'b0 ;
  assign n21747 = ~n21739 & n21746 ;
  assign n21748 = n3495 & ~n6634 ;
  assign n21749 = n15763 & n21748 ;
  assign n21750 = n12092 ^ n3476 ^ 1'b0 ;
  assign n21751 = ~n18756 & n21750 ;
  assign n21753 = ( n967 & n2796 ) | ( n967 & ~n12705 ) | ( n2796 & ~n12705 ) ;
  assign n21752 = ( ~n4341 & n9061 ) | ( ~n4341 & n15181 ) | ( n9061 & n15181 ) ;
  assign n21754 = n21753 ^ n21752 ^ n19875 ;
  assign n21755 = n11151 ^ n8243 ^ n838 ;
  assign n21756 = n21755 ^ n9856 ^ 1'b0 ;
  assign n21757 = n21754 & n21756 ;
  assign n21758 = ( n8162 & ~n21751 ) | ( n8162 & n21757 ) | ( ~n21751 & n21757 ) ;
  assign n21764 = n706 | n8710 ;
  assign n21765 = n4989 & ~n21764 ;
  assign n21766 = n12088 | n21765 ;
  assign n21767 = ~n14259 & n14972 ;
  assign n21768 = n21766 & n21767 ;
  assign n21769 = n16800 | n21768 ;
  assign n21770 = ( n16973 & n17739 ) | ( n16973 & ~n21769 ) | ( n17739 & ~n21769 ) ;
  assign n21759 = n3105 & ~n15845 ;
  assign n21760 = ~n1652 & n21759 ;
  assign n21761 = n9662 & n21760 ;
  assign n21762 = n2676 | n10573 ;
  assign n21763 = n21761 & ~n21762 ;
  assign n21771 = n21770 ^ n21763 ^ 1'b0 ;
  assign n21772 = n16780 & n21771 ;
  assign n21773 = n1365 & ~n21108 ;
  assign n21774 = n21773 ^ n5457 ^ 1'b0 ;
  assign n21775 = n21125 ^ n15809 ^ n4528 ;
  assign n21776 = ( n2197 & n3678 ) | ( n2197 & ~n21775 ) | ( n3678 & ~n21775 ) ;
  assign n21777 = ~n14210 & n21776 ;
  assign n21778 = ( ~n1186 & n2423 ) | ( ~n1186 & n13780 ) | ( n2423 & n13780 ) ;
  assign n21779 = n21778 ^ n11689 ^ 1'b0 ;
  assign n21780 = ( ~n436 & n6872 ) | ( ~n436 & n20194 ) | ( n6872 & n20194 ) ;
  assign n21781 = n21780 ^ n2096 ^ 1'b0 ;
  assign n21782 = n21779 & ~n21781 ;
  assign n21784 = n1289 & ~n20754 ;
  assign n21783 = ( n404 & n16989 ) | ( n404 & ~n18359 ) | ( n16989 & ~n18359 ) ;
  assign n21785 = n21784 ^ n21783 ^ n1673 ;
  assign n21786 = n8854 ^ n3450 ^ 1'b0 ;
  assign n21787 = n11597 ^ n3121 ^ 1'b0 ;
  assign n21788 = n21787 ^ n11661 ^ n5063 ;
  assign n21789 = n936 & ~n5701 ;
  assign n21790 = n967 & n21789 ;
  assign n21791 = ( n381 & ~n12672 ) | ( n381 & n21790 ) | ( ~n12672 & n21790 ) ;
  assign n21792 = n21791 ^ n5681 ^ x187 ;
  assign n21793 = ( n7745 & n12355 ) | ( n7745 & ~n21792 ) | ( n12355 & ~n21792 ) ;
  assign n21794 = n11704 & ~n12726 ;
  assign n21795 = n7000 & n21794 ;
  assign n21796 = n21795 ^ n3120 ^ n2955 ;
  assign n21797 = n3243 | n13497 ;
  assign n21799 = n11719 ^ n4315 ^ 1'b0 ;
  assign n21800 = n7930 | n21799 ;
  assign n21798 = n8422 ^ n7377 ^ n6593 ;
  assign n21801 = n21800 ^ n21798 ^ 1'b0 ;
  assign n21802 = n21797 | n21801 ;
  assign n21803 = n13969 ^ n2179 ^ n1331 ;
  assign n21804 = n21803 ^ n2689 ^ 1'b0 ;
  assign n21805 = n11257 | n21804 ;
  assign n21806 = n9237 ^ n4759 ^ 1'b0 ;
  assign n21807 = n16167 ^ n8760 ^ n8733 ;
  assign n21808 = ( n2329 & ~n5860 ) | ( n2329 & n21807 ) | ( ~n5860 & n21807 ) ;
  assign n21809 = ( n6764 & n8517 ) | ( n6764 & ~n21808 ) | ( n8517 & ~n21808 ) ;
  assign n21810 = ( n2377 & ~n6883 ) | ( n2377 & n13778 ) | ( ~n6883 & n13778 ) ;
  assign n21811 = n21810 ^ n3347 ^ 1'b0 ;
  assign n21812 = n18928 | n21811 ;
  assign n21813 = n7453 | n10023 ;
  assign n21814 = n8055 | n21813 ;
  assign n21815 = n21471 ^ n18588 ^ 1'b0 ;
  assign n21816 = ~n10307 & n21815 ;
  assign n21817 = n18790 ^ n2532 ^ 1'b0 ;
  assign n21818 = n5565 & ~n21817 ;
  assign n21819 = n16098 ^ n10038 ^ 1'b0 ;
  assign n21820 = n21818 & ~n21819 ;
  assign n21821 = n18814 ^ n11279 ^ n9727 ;
  assign n21822 = n8658 ^ n5919 ^ 1'b0 ;
  assign n21823 = ~n7223 & n21822 ;
  assign n21824 = n21823 ^ n19397 ^ 1'b0 ;
  assign n21825 = n3515 & n10388 ;
  assign n21826 = ( n4688 & ~n5480 ) | ( n4688 & n21825 ) | ( ~n5480 & n21825 ) ;
  assign n21827 = n21826 ^ n20262 ^ n16271 ;
  assign n21828 = n619 & ~n8027 ;
  assign n21829 = n21828 ^ n5965 ^ 1'b0 ;
  assign n21830 = n8702 ^ n2958 ^ n1444 ;
  assign n21831 = n21830 ^ n2215 ^ n322 ;
  assign n21832 = n12226 ^ n3138 ^ 1'b0 ;
  assign n21833 = ~n6111 & n21832 ;
  assign n21834 = n9949 & ~n21833 ;
  assign n21835 = n7978 ^ n2946 ^ 1'b0 ;
  assign n21836 = n9473 ^ n413 ^ 1'b0 ;
  assign n21837 = ~n21835 & n21836 ;
  assign n21838 = ( n21831 & n21834 ) | ( n21831 & ~n21837 ) | ( n21834 & ~n21837 ) ;
  assign n21839 = n966 & ~n21838 ;
  assign n21840 = n1866 & ~n10911 ;
  assign n21841 = n21840 ^ n2119 ^ 1'b0 ;
  assign n21842 = n2623 & n15555 ;
  assign n21850 = ( ~n2441 & n3141 ) | ( ~n2441 & n6503 ) | ( n3141 & n6503 ) ;
  assign n21843 = n2363 & ~n15365 ;
  assign n21844 = n20063 ^ n8297 ^ 1'b0 ;
  assign n21845 = ( ~n3023 & n21843 ) | ( ~n3023 & n21844 ) | ( n21843 & n21844 ) ;
  assign n21846 = n9726 ^ n7688 ^ n5397 ;
  assign n21847 = ~n10617 & n21846 ;
  assign n21848 = ~n21845 & n21847 ;
  assign n21849 = ~n12690 & n21848 ;
  assign n21851 = n21850 ^ n21849 ^ 1'b0 ;
  assign n21852 = ( n1337 & n11059 ) | ( n1337 & n11515 ) | ( n11059 & n11515 ) ;
  assign n21853 = n7040 | n21852 ;
  assign n21854 = n17132 ^ n14601 ^ 1'b0 ;
  assign n21864 = n3100 | n15066 ;
  assign n21865 = n3476 & ~n21864 ;
  assign n21861 = n3568 & ~n11021 ;
  assign n21862 = n5453 & n21861 ;
  assign n21863 = n18582 | n21862 ;
  assign n21866 = n21865 ^ n21863 ^ n8780 ;
  assign n21855 = ( n7708 & n12410 ) | ( n7708 & n14476 ) | ( n12410 & n14476 ) ;
  assign n21858 = n14266 ^ n3455 ^ n2947 ;
  assign n21856 = ~n1555 & n2208 ;
  assign n21857 = n16906 | n21856 ;
  assign n21859 = n21858 ^ n21857 ^ 1'b0 ;
  assign n21860 = n21855 | n21859 ;
  assign n21867 = n21866 ^ n21860 ^ 1'b0 ;
  assign n21872 = n13154 ^ n8937 ^ n1630 ;
  assign n21873 = n21872 ^ n16797 ^ n11594 ;
  assign n21868 = ~n2445 & n9843 ;
  assign n21869 = n21868 ^ n19993 ^ 1'b0 ;
  assign n21870 = ( n15105 & n15614 ) | ( n15105 & n21869 ) | ( n15614 & n21869 ) ;
  assign n21871 = ( n8484 & n17301 ) | ( n8484 & ~n21870 ) | ( n17301 & ~n21870 ) ;
  assign n21874 = n21873 ^ n21871 ^ n20563 ;
  assign n21875 = n4177 ^ n857 ^ x225 ;
  assign n21876 = n18761 ^ n12372 ^ n3857 ;
  assign n21877 = n1075 | n21876 ;
  assign n21878 = n17141 | n21877 ;
  assign n21879 = ~n13894 & n21878 ;
  assign n21880 = ( n4911 & n21875 ) | ( n4911 & ~n21879 ) | ( n21875 & ~n21879 ) ;
  assign n21881 = n21880 ^ n21506 ^ n13028 ;
  assign n21882 = n1028 | n3117 ;
  assign n21883 = ( n4837 & n9540 ) | ( n4837 & ~n15712 ) | ( n9540 & ~n15712 ) ;
  assign n21884 = ( n711 & n12841 ) | ( n711 & n21883 ) | ( n12841 & n21883 ) ;
  assign n21885 = n9788 ^ n9366 ^ 1'b0 ;
  assign n21886 = n3650 | n13125 ;
  assign n21887 = n21886 ^ n12705 ^ 1'b0 ;
  assign n21888 = n14924 ^ n12053 ^ n4457 ;
  assign n21893 = n5765 & ~n7840 ;
  assign n21894 = ( ~n12391 & n17170 ) | ( ~n12391 & n21893 ) | ( n17170 & n21893 ) ;
  assign n21889 = n5918 & ~n6964 ;
  assign n21890 = n3048 & n21889 ;
  assign n21891 = n21890 ^ n9322 ^ 1'b0 ;
  assign n21892 = ~n9018 & n21891 ;
  assign n21895 = n21894 ^ n21892 ^ 1'b0 ;
  assign n21896 = n21888 & ~n21895 ;
  assign n21897 = n14849 ^ n11560 ^ 1'b0 ;
  assign n21898 = n7753 & ~n21897 ;
  assign n21899 = ( n7505 & ~n16385 ) | ( n7505 & n19192 ) | ( ~n16385 & n19192 ) ;
  assign n21900 = ( n365 & n10316 ) | ( n365 & n20076 ) | ( n10316 & n20076 ) ;
  assign n21901 = n2679 & n21900 ;
  assign n21902 = ( n12237 & ~n20498 ) | ( n12237 & n21871 ) | ( ~n20498 & n21871 ) ;
  assign n21903 = n17744 ^ n1192 ^ n663 ;
  assign n21904 = n12403 ^ n3433 ^ n394 ;
  assign n21905 = n15011 & n21904 ;
  assign n21906 = n11124 ^ n9658 ^ n6267 ;
  assign n21907 = ~n10781 & n21906 ;
  assign n21908 = n7974 ^ n5062 ^ 1'b0 ;
  assign n21909 = ( x188 & n1934 ) | ( x188 & n21908 ) | ( n1934 & n21908 ) ;
  assign n21910 = ( n9103 & ~n21907 ) | ( n9103 & n21909 ) | ( ~n21907 & n21909 ) ;
  assign n21911 = n17095 ^ n16555 ^ 1'b0 ;
  assign n21912 = n21911 ^ n10956 ^ 1'b0 ;
  assign n21913 = n3190 & ~n4794 ;
  assign n21914 = n7823 ^ n3776 ^ 1'b0 ;
  assign n21915 = ( n18899 & n21913 ) | ( n18899 & ~n21914 ) | ( n21913 & ~n21914 ) ;
  assign n21916 = n940 & n10233 ;
  assign n21917 = n21916 ^ n19496 ^ n9072 ;
  assign n21918 = n21917 ^ n15291 ^ 1'b0 ;
  assign n21919 = n17689 & ~n21918 ;
  assign n21920 = ~n1464 & n21919 ;
  assign n21921 = n8377 ^ n1026 ^ x4 ;
  assign n21922 = ( n8103 & ~n9066 ) | ( n8103 & n21921 ) | ( ~n9066 & n21921 ) ;
  assign n21923 = n11498 & n21922 ;
  assign n21924 = n21870 ^ n10921 ^ 1'b0 ;
  assign n21925 = n21923 & ~n21924 ;
  assign n21926 = n5032 | n5311 ;
  assign n21927 = n11727 & ~n21926 ;
  assign n21928 = x18 & ~n21927 ;
  assign n21929 = n21928 ^ n12255 ^ 1'b0 ;
  assign n21930 = ( ~n10867 & n18806 ) | ( ~n10867 & n21929 ) | ( n18806 & n21929 ) ;
  assign n21931 = n10633 | n12263 ;
  assign n21932 = n21931 ^ n18615 ^ 1'b0 ;
  assign n21933 = n15666 & ~n21932 ;
  assign n21934 = n21933 ^ n19539 ^ 1'b0 ;
  assign n21935 = n20763 ^ n5318 ^ n4455 ;
  assign n21936 = n21935 ^ n18121 ^ n6988 ;
  assign n21937 = n21936 ^ n15631 ^ 1'b0 ;
  assign n21938 = ( n4897 & n17092 ) | ( n4897 & n18493 ) | ( n17092 & n18493 ) ;
  assign n21939 = x189 & ~n21625 ;
  assign n21940 = n13692 & ~n14880 ;
  assign n21941 = ~n7689 & n10843 ;
  assign n21942 = n5480 | n17136 ;
  assign n21943 = n2982 & ~n21942 ;
  assign n21944 = n4860 ^ n1746 ^ 1'b0 ;
  assign n21945 = ~n4648 & n5929 ;
  assign n21946 = n21944 & ~n21945 ;
  assign n21947 = n21943 & n21946 ;
  assign n21948 = ( ~n6512 & n21941 ) | ( ~n6512 & n21947 ) | ( n21941 & n21947 ) ;
  assign n21949 = n7783 ^ n7085 ^ n4443 ;
  assign n21950 = n1175 & ~n21949 ;
  assign n21951 = n15883 ^ n2406 ^ 1'b0 ;
  assign n21952 = n21951 ^ n15666 ^ x11 ;
  assign n21953 = ( n2179 & ~n21950 ) | ( n2179 & n21952 ) | ( ~n21950 & n21952 ) ;
  assign n21954 = n11027 | n14389 ;
  assign n21955 = n14915 | n21954 ;
  assign n21956 = n4626 | n14095 ;
  assign n21957 = n6823 & ~n21956 ;
  assign n21958 = n11433 ^ n9777 ^ 1'b0 ;
  assign n21959 = n5676 | n21958 ;
  assign n21960 = n21959 ^ n1317 ^ 1'b0 ;
  assign n21961 = ~n883 & n5486 ;
  assign n21962 = n793 & n21961 ;
  assign n21963 = ( n8810 & ~n19759 ) | ( n8810 & n21962 ) | ( ~n19759 & n21962 ) ;
  assign n21964 = n17147 ^ n9969 ^ 1'b0 ;
  assign n21965 = n10638 & n21964 ;
  assign n21966 = ~n7941 & n21965 ;
  assign n21967 = n21966 ^ n2980 ^ 1'b0 ;
  assign n21968 = ( n11157 & ~n21139 ) | ( n11157 & n21967 ) | ( ~n21139 & n21967 ) ;
  assign n21969 = n3780 | n12304 ;
  assign n21970 = n3388 | n21969 ;
  assign n21971 = ( n2017 & n8766 ) | ( n2017 & n9327 ) | ( n8766 & n9327 ) ;
  assign n21972 = n18216 ^ n11909 ^ 1'b0 ;
  assign n21973 = n21971 & ~n21972 ;
  assign n21974 = n21970 & ~n21973 ;
  assign n21975 = n6211 | n21974 ;
  assign n21976 = n21968 | n21975 ;
  assign n21977 = n21976 ^ n1311 ^ 1'b0 ;
  assign n21978 = n7689 | n18737 ;
  assign n21979 = n21978 ^ n13490 ^ 1'b0 ;
  assign n21980 = n3671 & n15426 ;
  assign n21981 = n21980 ^ n8337 ^ 1'b0 ;
  assign n21982 = n7812 | n21981 ;
  assign n21983 = ( x93 & ~n6043 ) | ( x93 & n21982 ) | ( ~n6043 & n21982 ) ;
  assign n21984 = ~n6423 & n8458 ;
  assign n21985 = n3652 & n3945 ;
  assign n21986 = n21985 ^ n4794 ^ 1'b0 ;
  assign n21987 = ~n4813 & n21986 ;
  assign n21988 = ( ~n21983 & n21984 ) | ( ~n21983 & n21987 ) | ( n21984 & n21987 ) ;
  assign n21990 = ( n4900 & n5402 ) | ( n4900 & n11751 ) | ( n5402 & n11751 ) ;
  assign n21989 = n9992 & ~n12789 ;
  assign n21991 = n21990 ^ n21989 ^ 1'b0 ;
  assign n21992 = n17014 ^ n4779 ^ 1'b0 ;
  assign n21993 = n10890 & n21992 ;
  assign n21994 = n18841 & n21993 ;
  assign n21995 = n21991 | n21994 ;
  assign n21996 = n15003 ^ n6306 ^ 1'b0 ;
  assign n21997 = ( n8727 & n11747 ) | ( n8727 & ~n14901 ) | ( n11747 & ~n14901 ) ;
  assign n21998 = n3061 & n13544 ;
  assign n21999 = n11618 & n21998 ;
  assign n22000 = n21999 ^ n2880 ^ 1'b0 ;
  assign n22001 = n11463 ^ n4060 ^ 1'b0 ;
  assign n22002 = n3967 ^ n3807 ^ 1'b0 ;
  assign n22003 = ~n22001 & n22002 ;
  assign n22004 = n22003 ^ n20270 ^ 1'b0 ;
  assign n22005 = n22004 ^ n2559 ^ 1'b0 ;
  assign n22007 = n5189 ^ n4536 ^ 1'b0 ;
  assign n22008 = x237 & ~n22007 ;
  assign n22006 = n8070 ^ n6286 ^ 1'b0 ;
  assign n22009 = n22008 ^ n22006 ^ 1'b0 ;
  assign n22010 = n13976 & ~n22009 ;
  assign n22011 = n16807 ^ n11796 ^ 1'b0 ;
  assign n22012 = n5554 | n11504 ;
  assign n22013 = ( n5607 & ~n13326 ) | ( n5607 & n22012 ) | ( ~n13326 & n22012 ) ;
  assign n22014 = n22013 ^ n16117 ^ n8187 ;
  assign n22015 = n13317 & n22014 ;
  assign n22016 = n22015 ^ n18521 ^ 1'b0 ;
  assign n22017 = n22016 ^ n19824 ^ 1'b0 ;
  assign n22020 = n13713 ^ n5070 ^ 1'b0 ;
  assign n22021 = n15098 & n22020 ;
  assign n22022 = n22021 ^ n4666 ^ 1'b0 ;
  assign n22018 = n9019 ^ n7586 ^ 1'b0 ;
  assign n22019 = ( n1123 & ~n10995 ) | ( n1123 & n22018 ) | ( ~n10995 & n22018 ) ;
  assign n22023 = n22022 ^ n22019 ^ n4072 ;
  assign n22024 = ( ~n2170 & n12103 ) | ( ~n2170 & n13086 ) | ( n12103 & n13086 ) ;
  assign n22025 = n22024 ^ n6415 ^ 1'b0 ;
  assign n22026 = n3839 | n11627 ;
  assign n22027 = ( n4150 & n22025 ) | ( n4150 & ~n22026 ) | ( n22025 & ~n22026 ) ;
  assign n22028 = n9205 ^ n1183 ^ 1'b0 ;
  assign n22029 = n22028 ^ n9485 ^ 1'b0 ;
  assign n22030 = n17351 & n22029 ;
  assign n22034 = n19324 ^ n8200 ^ n4393 ;
  assign n22035 = ~n10740 & n22034 ;
  assign n22031 = n20283 ^ n1483 ^ 1'b0 ;
  assign n22032 = n22031 ^ n4566 ^ 1'b0 ;
  assign n22033 = ( n3863 & ~n17132 ) | ( n3863 & n22032 ) | ( ~n17132 & n22032 ) ;
  assign n22036 = n22035 ^ n22033 ^ n5966 ;
  assign n22041 = n14685 ^ n3415 ^ 1'b0 ;
  assign n22042 = n6974 | n22041 ;
  assign n22043 = ( n10206 & ~n13313 ) | ( n10206 & n22042 ) | ( ~n13313 & n22042 ) ;
  assign n22037 = n20235 ^ n12428 ^ n2515 ;
  assign n22038 = n5504 | n9793 ;
  assign n22039 = n16740 & ~n22038 ;
  assign n22040 = n22037 & ~n22039 ;
  assign n22044 = n22043 ^ n22040 ^ 1'b0 ;
  assign n22045 = ~n1660 & n5276 ;
  assign n22046 = n2194 & ~n9370 ;
  assign n22047 = ~n10939 & n22046 ;
  assign n22048 = n3280 | n5979 ;
  assign n22049 = n22048 ^ n4280 ^ 1'b0 ;
  assign n22050 = ( ~n9671 & n12344 ) | ( ~n9671 & n22049 ) | ( n12344 & n22049 ) ;
  assign n22051 = ( n15572 & n22047 ) | ( n15572 & ~n22050 ) | ( n22047 & ~n22050 ) ;
  assign n22052 = n2423 & ~n12755 ;
  assign n22053 = ( n750 & ~n12729 ) | ( n750 & n19874 ) | ( ~n12729 & n19874 ) ;
  assign n22054 = n22053 ^ n20588 ^ n1780 ;
  assign n22055 = ( n2716 & ~n7742 ) | ( n2716 & n8603 ) | ( ~n7742 & n8603 ) ;
  assign n22056 = ~n12947 & n21365 ;
  assign n22057 = n15405 & n22056 ;
  assign n22058 = ~n4501 & n15552 ;
  assign n22059 = n6070 & ~n10835 ;
  assign n22060 = n22059 ^ n7453 ^ 1'b0 ;
  assign n22061 = ( ~n11984 & n22058 ) | ( ~n11984 & n22060 ) | ( n22058 & n22060 ) ;
  assign n22062 = n22061 ^ n6056 ^ 1'b0 ;
  assign n22063 = ~n8548 & n22062 ;
  assign n22064 = n4670 & n22063 ;
  assign n22065 = n22064 ^ n2639 ^ 1'b0 ;
  assign n22066 = ( n22055 & n22057 ) | ( n22055 & ~n22065 ) | ( n22057 & ~n22065 ) ;
  assign n22067 = n3381 & ~n12701 ;
  assign n22068 = ~n10757 & n22067 ;
  assign n22069 = ( x105 & ~x201 ) | ( x105 & n22068 ) | ( ~x201 & n22068 ) ;
  assign n22070 = ~n5770 & n22069 ;
  assign n22071 = ( ~x10 & n4240 ) | ( ~x10 & n20791 ) | ( n4240 & n20791 ) ;
  assign n22072 = ( ~n6246 & n6978 ) | ( ~n6246 & n22071 ) | ( n6978 & n22071 ) ;
  assign n22073 = n20433 ^ n17284 ^ n9749 ;
  assign n22074 = ( n12526 & n13467 ) | ( n12526 & ~n17009 ) | ( n13467 & ~n17009 ) ;
  assign n22075 = ( n4070 & ~n5061 ) | ( n4070 & n6235 ) | ( ~n5061 & n6235 ) ;
  assign n22076 = n19238 ^ n6367 ^ 1'b0 ;
  assign n22077 = n22075 | n22076 ;
  assign n22078 = n22077 ^ n10794 ^ n1175 ;
  assign n22079 = n20350 ^ n15731 ^ n12200 ;
  assign n22080 = ~n871 & n22079 ;
  assign n22081 = n2146 ^ n713 ^ 1'b0 ;
  assign n22082 = ( n1226 & n6856 ) | ( n1226 & n10418 ) | ( n6856 & n10418 ) ;
  assign n22083 = n22081 | n22082 ;
  assign n22084 = ( n15719 & n20229 ) | ( n15719 & ~n22083 ) | ( n20229 & ~n22083 ) ;
  assign n22085 = n15510 | n21154 ;
  assign n22086 = n6030 & ~n22085 ;
  assign n22087 = n5456 & ~n11226 ;
  assign n22088 = n22087 ^ n2544 ^ 1'b0 ;
  assign n22089 = ( n2006 & n5376 ) | ( n2006 & ~n5508 ) | ( n5376 & ~n5508 ) ;
  assign n22090 = n22089 ^ n3042 ^ 1'b0 ;
  assign n22091 = n13985 ^ n355 ^ 1'b0 ;
  assign n22092 = ~n22090 & n22091 ;
  assign n22093 = n2816 & n22092 ;
  assign n22094 = ~n22088 & n22093 ;
  assign n22099 = ~x106 & n5526 ;
  assign n22100 = ~n4664 & n22099 ;
  assign n22098 = n14129 ^ n13011 ^ n4756 ;
  assign n22101 = n22100 ^ n22098 ^ n2559 ;
  assign n22095 = n11843 ^ n7363 ^ n4226 ;
  assign n22096 = ~n12524 & n22095 ;
  assign n22097 = n10826 | n22096 ;
  assign n22102 = n22101 ^ n22097 ^ 1'b0 ;
  assign n22103 = n12759 & n20532 ;
  assign n22110 = x232 & ~n3728 ;
  assign n22111 = n4481 & n22110 ;
  assign n22104 = n3346 | n22057 ;
  assign n22105 = n22104 ^ n15360 ^ 1'b0 ;
  assign n22106 = n17618 ^ n17493 ^ 1'b0 ;
  assign n22107 = n22106 ^ n15921 ^ n6181 ;
  assign n22108 = n22107 ^ n2595 ^ 1'b0 ;
  assign n22109 = ~n22105 & n22108 ;
  assign n22112 = n22111 ^ n22109 ^ n5463 ;
  assign n22113 = n9820 ^ n6044 ^ x86 ;
  assign n22114 = ~n4974 & n22113 ;
  assign n22115 = n6064 & n22114 ;
  assign n22118 = n10358 ^ n7185 ^ n1743 ;
  assign n22119 = n10628 ^ n1388 ^ 1'b0 ;
  assign n22120 = ~n22118 & n22119 ;
  assign n22121 = n1930 | n22120 ;
  assign n22116 = n9084 ^ n2498 ^ n276 ;
  assign n22117 = ( ~n10351 & n20601 ) | ( ~n10351 & n22116 ) | ( n20601 & n22116 ) ;
  assign n22122 = n22121 ^ n22117 ^ n6705 ;
  assign n22123 = n2965 & ~n20621 ;
  assign n22124 = n6384 & n8878 ;
  assign n22125 = n19928 ^ n9297 ^ n619 ;
  assign n22126 = n22125 ^ n11269 ^ n10077 ;
  assign n22127 = n22126 ^ n12037 ^ 1'b0 ;
  assign n22128 = ( n16864 & n22124 ) | ( n16864 & ~n22127 ) | ( n22124 & ~n22127 ) ;
  assign n22132 = n910 & ~n1446 ;
  assign n22133 = n2240 & n22132 ;
  assign n22134 = ( n552 & ~n7542 ) | ( n552 & n22133 ) | ( ~n7542 & n22133 ) ;
  assign n22131 = n14365 ^ n10620 ^ n6359 ;
  assign n22135 = n22134 ^ n22131 ^ n10731 ;
  assign n22129 = n14731 ^ n3209 ^ n294 ;
  assign n22130 = n7274 & n22129 ;
  assign n22136 = n22135 ^ n22130 ^ n19065 ;
  assign n22137 = n22136 ^ n20772 ^ n900 ;
  assign n22138 = n1485 | n3035 ;
  assign n22139 = n22138 ^ n10804 ^ 1'b0 ;
  assign n22140 = ~n6681 & n22139 ;
  assign n22141 = n13141 ^ n9084 ^ n3328 ;
  assign n22142 = ( n2450 & n6548 ) | ( n2450 & ~n22141 ) | ( n6548 & ~n22141 ) ;
  assign n22143 = ~n21354 & n22142 ;
  assign n22144 = n22143 ^ n19152 ^ 1'b0 ;
  assign n22145 = n12360 ^ n2642 ^ 1'b0 ;
  assign n22146 = n19009 & ~n22145 ;
  assign n22147 = n20940 ^ n2540 ^ 1'b0 ;
  assign n22148 = n22147 ^ n18493 ^ n16481 ;
  assign n22149 = n3496 | n4473 ;
  assign n22150 = n22149 ^ n9855 ^ n6173 ;
  assign n22151 = n3915 & ~n22150 ;
  assign n22152 = n22151 ^ n7216 ^ 1'b0 ;
  assign n22153 = n17114 & n22152 ;
  assign n22154 = n5455 & n11104 ;
  assign n22155 = ( n7220 & ~n22153 ) | ( n7220 & n22154 ) | ( ~n22153 & n22154 ) ;
  assign n22156 = n7174 & n22155 ;
  assign n22157 = n21788 ^ n18873 ^ 1'b0 ;
  assign n22161 = n12718 ^ n8359 ^ 1'b0 ;
  assign n22158 = n5563 ^ n1461 ^ 1'b0 ;
  assign n22159 = ~n4364 & n22158 ;
  assign n22160 = n22159 ^ n2820 ^ n2649 ;
  assign n22162 = n22161 ^ n22160 ^ n1889 ;
  assign n22163 = n5068 & n16077 ;
  assign n22164 = n22163 ^ n16378 ^ 1'b0 ;
  assign n22165 = n22164 ^ n3089 ^ 1'b0 ;
  assign n22166 = n22162 & n22165 ;
  assign n22167 = n6624 ^ n3530 ^ n870 ;
  assign n22168 = ( n5674 & ~n15019 ) | ( n5674 & n22167 ) | ( ~n15019 & n22167 ) ;
  assign n22169 = n22168 ^ n14634 ^ n1330 ;
  assign n22170 = ( ~n800 & n5349 ) | ( ~n800 & n6045 ) | ( n5349 & n6045 ) ;
  assign n22172 = n17164 ^ n13351 ^ n2709 ;
  assign n22173 = n22172 ^ n3536 ^ x186 ;
  assign n22171 = ( n5809 & n12225 ) | ( n5809 & ~n17109 ) | ( n12225 & ~n17109 ) ;
  assign n22174 = n22173 ^ n22171 ^ n15407 ;
  assign n22175 = ( n6349 & n22170 ) | ( n6349 & n22174 ) | ( n22170 & n22174 ) ;
  assign n22176 = n18801 ^ n16266 ^ n14446 ;
  assign n22177 = n3928 | n21261 ;
  assign n22181 = n8520 & ~n8593 ;
  assign n22182 = n14406 & ~n22181 ;
  assign n22179 = n1854 & ~n15809 ;
  assign n22180 = n22179 ^ n17707 ^ 1'b0 ;
  assign n22178 = ( x82 & n7503 ) | ( x82 & ~n11193 ) | ( n7503 & ~n11193 ) ;
  assign n22183 = n22182 ^ n22180 ^ n22178 ;
  assign n22184 = n15587 & n21471 ;
  assign n22185 = ~n15024 & n22184 ;
  assign n22186 = ~n7345 & n22185 ;
  assign n22188 = n19098 ^ n13909 ^ n703 ;
  assign n22187 = n7511 & ~n15221 ;
  assign n22189 = n22188 ^ n22187 ^ n11412 ;
  assign n22194 = n5458 ^ n5097 ^ 1'b0 ;
  assign n22195 = n8047 & n22194 ;
  assign n22190 = n4800 & n6103 ;
  assign n22191 = n756 | n15011 ;
  assign n22192 = n22191 ^ n14803 ^ 1'b0 ;
  assign n22193 = n22190 & ~n22192 ;
  assign n22196 = n22195 ^ n22193 ^ n15573 ;
  assign n22197 = n19587 ^ n4143 ^ n1102 ;
  assign n22198 = n21603 ^ n21464 ^ 1'b0 ;
  assign n22199 = n10183 ^ n2955 ^ 1'b0 ;
  assign n22200 = n1387 & ~n22199 ;
  assign n22202 = n2606 & ~n10584 ;
  assign n22203 = ( ~n13152 & n13326 ) | ( ~n13152 & n22202 ) | ( n13326 & n22202 ) ;
  assign n22201 = ~n11487 & n15166 ;
  assign n22204 = n22203 ^ n22201 ^ 1'b0 ;
  assign n22205 = ~n7115 & n12020 ;
  assign n22207 = n20609 ^ n6411 ^ 1'b0 ;
  assign n22208 = n12899 & ~n22207 ;
  assign n22206 = n4982 & ~n8947 ;
  assign n22209 = n22208 ^ n22206 ^ n745 ;
  assign n22210 = ( n7994 & ~n14644 ) | ( n7994 & n19910 ) | ( ~n14644 & n19910 ) ;
  assign n22211 = n2823 ^ n1050 ^ 1'b0 ;
  assign n22212 = n6432 | n22211 ;
  assign n22213 = n7017 ^ n4524 ^ 1'b0 ;
  assign n22214 = n7353 | n22213 ;
  assign n22215 = n22212 | n22214 ;
  assign n22216 = n22215 ^ n14815 ^ 1'b0 ;
  assign n22217 = n22216 ^ n20014 ^ 1'b0 ;
  assign n22218 = ~n22210 & n22217 ;
  assign n22220 = ( n5544 & n7320 ) | ( n5544 & ~n10102 ) | ( n7320 & ~n10102 ) ;
  assign n22219 = n7892 & ~n11037 ;
  assign n22221 = n22220 ^ n22219 ^ 1'b0 ;
  assign n22222 = n16638 ^ n1184 ^ 1'b0 ;
  assign n22223 = n22221 & n22222 ;
  assign n22224 = n22223 ^ n2746 ^ n488 ;
  assign n22225 = n16904 ^ n13487 ^ 1'b0 ;
  assign n22226 = n22225 ^ n10254 ^ n1383 ;
  assign n22227 = ( n320 & n19806 ) | ( n320 & n21950 ) | ( n19806 & n21950 ) ;
  assign n22228 = ( n10499 & ~n22226 ) | ( n10499 & n22227 ) | ( ~n22226 & n22227 ) ;
  assign n22229 = ~n4540 & n13675 ;
  assign n22230 = n22229 ^ n19716 ^ 1'b0 ;
  assign n22231 = ~n8080 & n22230 ;
  assign n22232 = ( ~n14991 & n21051 ) | ( ~n14991 & n22231 ) | ( n21051 & n22231 ) ;
  assign n22233 = n7467 | n10633 ;
  assign n22234 = n22233 ^ n16272 ^ 1'b0 ;
  assign n22235 = n22234 ^ n11136 ^ n2361 ;
  assign n22236 = n22235 ^ n15631 ^ n7854 ;
  assign n22237 = n1752 | n2388 ;
  assign n22238 = n22237 ^ n14123 ^ 1'b0 ;
  assign n22239 = n22024 ^ n2553 ^ 1'b0 ;
  assign n22240 = n18431 | n22239 ;
  assign n22241 = n22238 | n22240 ;
  assign n22242 = n22241 ^ n17779 ^ 1'b0 ;
  assign n22243 = n1342 ^ n280 ^ 1'b0 ;
  assign n22244 = n19834 ^ n6699 ^ 1'b0 ;
  assign n22246 = ( ~n9178 & n11476 ) | ( ~n9178 & n11493 ) | ( n11476 & n11493 ) ;
  assign n22245 = n11026 | n12009 ;
  assign n22247 = n22246 ^ n22245 ^ 1'b0 ;
  assign n22248 = n306 & n17956 ;
  assign n22251 = ~n470 & n6015 ;
  assign n22252 = n470 & n22251 ;
  assign n22253 = n22252 ^ n1348 ^ 1'b0 ;
  assign n22249 = n5114 | n11503 ;
  assign n22250 = n11503 & ~n22249 ;
  assign n22254 = n22253 ^ n22250 ^ 1'b0 ;
  assign n22255 = n7252 & n16951 ;
  assign n22256 = n8515 & ~n12142 ;
  assign n22257 = n3583 & ~n22256 ;
  assign n22258 = ( n1046 & ~n9240 ) | ( n1046 & n10461 ) | ( ~n9240 & n10461 ) ;
  assign n22259 = ( n6393 & n22257 ) | ( n6393 & n22258 ) | ( n22257 & n22258 ) ;
  assign n22260 = n5722 & ~n22259 ;
  assign n22261 = n22260 ^ n16794 ^ 1'b0 ;
  assign n22262 = n2277 & n2892 ;
  assign n22263 = n22262 ^ n17737 ^ 1'b0 ;
  assign n22264 = ( n2131 & ~n12867 ) | ( n2131 & n15976 ) | ( ~n12867 & n15976 ) ;
  assign n22265 = n22264 ^ n20349 ^ 1'b0 ;
  assign n22266 = ~n536 & n1303 ;
  assign n22267 = ( n17367 & n18341 ) | ( n17367 & n22266 ) | ( n18341 & n22266 ) ;
  assign n22268 = n9300 ^ n4934 ^ 1'b0 ;
  assign n22269 = ( n436 & n3312 ) | ( n436 & n4910 ) | ( n3312 & n4910 ) ;
  assign n22270 = n22269 ^ n5196 ^ 1'b0 ;
  assign n22271 = ~n350 & n7373 ;
  assign n22272 = n22271 ^ n14462 ^ 1'b0 ;
  assign n22273 = n22272 ^ n12016 ^ 1'b0 ;
  assign n22274 = n10259 & ~n22273 ;
  assign n22275 = n2085 & n22274 ;
  assign n22276 = n22275 ^ n9755 ^ 1'b0 ;
  assign n22277 = ( n7004 & n9446 ) | ( n7004 & n20951 ) | ( n9446 & n20951 ) ;
  assign n22278 = n22277 ^ n21389 ^ 1'b0 ;
  assign n22279 = n18862 & n22278 ;
  assign n22280 = n2169 | n7991 ;
  assign n22281 = n15157 | n22280 ;
  assign n22282 = n4398 ^ n1876 ^ n1149 ;
  assign n22283 = x236 & ~n6077 ;
  assign n22284 = n8707 & n22283 ;
  assign n22285 = n22284 ^ n20685 ^ n7414 ;
  assign n22286 = n22285 ^ n11853 ^ n9522 ;
  assign n22287 = ( n9147 & n22282 ) | ( n9147 & n22286 ) | ( n22282 & n22286 ) ;
  assign n22288 = n9122 & ~n22287 ;
  assign n22289 = ~n22281 & n22288 ;
  assign n22290 = n2417 ^ n420 ^ 1'b0 ;
  assign n22291 = n813 & n22290 ;
  assign n22292 = n15826 ^ n10359 ^ n6523 ;
  assign n22293 = n22291 | n22292 ;
  assign n22294 = n22293 ^ n8595 ^ 1'b0 ;
  assign n22295 = n13554 | n22294 ;
  assign n22296 = ( ~n3823 & n9114 ) | ( ~n3823 & n16259 ) | ( n9114 & n16259 ) ;
  assign n22297 = n12107 ^ n11872 ^ n3225 ;
  assign n22298 = n22297 ^ n15290 ^ n9477 ;
  assign n22299 = ~n16007 & n22298 ;
  assign n22300 = x148 & ~n1337 ;
  assign n22301 = n22300 ^ n5294 ^ 1'b0 ;
  assign n22302 = n3873 ^ n637 ^ 1'b0 ;
  assign n22303 = n22302 ^ n2704 ^ 1'b0 ;
  assign n22304 = n22301 & n22303 ;
  assign n22305 = n22304 ^ n12443 ^ 1'b0 ;
  assign n22306 = n22305 ^ n21000 ^ 1'b0 ;
  assign n22307 = n22299 & ~n22306 ;
  assign n22314 = n17145 ^ n5085 ^ 1'b0 ;
  assign n22308 = ( n954 & n2527 ) | ( n954 & n3413 ) | ( n2527 & n3413 ) ;
  assign n22309 = x51 & n22308 ;
  assign n22310 = ~n3870 & n22309 ;
  assign n22311 = n17179 | n22310 ;
  assign n22312 = n13239 & ~n22311 ;
  assign n22313 = n22312 ^ n5407 ^ n2692 ;
  assign n22315 = n22314 ^ n22313 ^ n9075 ;
  assign n22316 = n17671 ^ n2523 ^ 1'b0 ;
  assign n22317 = n629 & ~n22316 ;
  assign n22318 = n2427 & ~n22001 ;
  assign n22319 = n17329 & n22318 ;
  assign n22320 = x48 & n3157 ;
  assign n22321 = n1868 & n22320 ;
  assign n22322 = n22321 ^ n16047 ^ n11863 ;
  assign n22323 = n9878 ^ n733 ^ 1'b0 ;
  assign n22324 = n12905 & ~n22323 ;
  assign n22325 = n1052 & ~n3324 ;
  assign n22326 = n1682 & ~n7410 ;
  assign n22327 = ~n14204 & n22326 ;
  assign n22328 = n22325 & n22327 ;
  assign n22329 = n5646 & ~n16034 ;
  assign n22330 = n15860 ^ n6493 ^ x18 ;
  assign n22331 = n2261 | n15562 ;
  assign n22335 = n3491 | n3655 ;
  assign n22336 = x224 | n22335 ;
  assign n22337 = n22336 ^ n2488 ^ 1'b0 ;
  assign n22338 = n9549 | n22337 ;
  assign n22332 = n2966 ^ n2508 ^ 1'b0 ;
  assign n22333 = n22332 ^ n14172 ^ n11241 ;
  assign n22334 = n22333 ^ n2191 ^ n481 ;
  assign n22339 = n22338 ^ n22334 ^ n2274 ;
  assign n22340 = n1649 & n1975 ;
  assign n22341 = n22340 ^ n748 ^ 1'b0 ;
  assign n22342 = ~n1356 & n8675 ;
  assign n22343 = n7461 & n22342 ;
  assign n22344 = n1712 & n9521 ;
  assign n22345 = n899 & n22344 ;
  assign n22346 = n22345 ^ n598 ^ 1'b0 ;
  assign n22347 = n22343 | n22346 ;
  assign n22348 = n12805 ^ n1806 ^ x33 ;
  assign n22349 = n16180 & n22348 ;
  assign n22350 = ( n11703 & n12999 ) | ( n11703 & n13075 ) | ( n12999 & n13075 ) ;
  assign n22351 = n3523 & ~n11669 ;
  assign n22352 = ( ~n7076 & n15234 ) | ( ~n7076 & n22351 ) | ( n15234 & n22351 ) ;
  assign n22353 = ( ~n7783 & n11041 ) | ( ~n7783 & n16156 ) | ( n11041 & n16156 ) ;
  assign n22354 = n13810 & ~n22353 ;
  assign n22355 = n13841 | n22034 ;
  assign n22356 = n11948 ^ n9378 ^ n5913 ;
  assign n22357 = n22356 ^ n18535 ^ n9770 ;
  assign n22358 = n10194 ^ n3813 ^ 1'b0 ;
  assign n22359 = ~n7764 & n22358 ;
  assign n22360 = ( n389 & n7325 ) | ( n389 & n10858 ) | ( n7325 & n10858 ) ;
  assign n22361 = n8212 ^ n7386 ^ 1'b0 ;
  assign n22362 = ~n22360 & n22361 ;
  assign n22363 = n9134 & n22362 ;
  assign n22364 = n22363 ^ n14166 ^ 1'b0 ;
  assign n22365 = n7665 ^ n5242 ^ 1'b0 ;
  assign n22366 = n6395 & ~n22365 ;
  assign n22367 = n2220 & n22366 ;
  assign n22368 = n18801 & n22367 ;
  assign n22369 = n5557 ^ n5251 ^ n1984 ;
  assign n22370 = n4062 | n22369 ;
  assign n22372 = n7278 | n9034 ;
  assign n22371 = n2262 & ~n8887 ;
  assign n22373 = n22372 ^ n22371 ^ 1'b0 ;
  assign n22374 = n6697 & n17971 ;
  assign n22375 = n22374 ^ n10945 ^ 1'b0 ;
  assign n22376 = ~n2236 & n22375 ;
  assign n22377 = n10250 ^ n5846 ^ 1'b0 ;
  assign n22378 = n14963 | n22377 ;
  assign n22379 = n22378 ^ n13262 ^ 1'b0 ;
  assign n22385 = ( n738 & n7984 ) | ( n738 & n19966 ) | ( n7984 & n19966 ) ;
  assign n22380 = n6335 ^ n4659 ^ 1'b0 ;
  assign n22381 = n15752 | n22380 ;
  assign n22382 = n22381 ^ n18995 ^ 1'b0 ;
  assign n22383 = n22382 ^ n1894 ^ 1'b0 ;
  assign n22384 = ~n8023 & n22383 ;
  assign n22386 = n22385 ^ n22384 ^ n14798 ;
  assign n22387 = n16466 ^ n14913 ^ n7163 ;
  assign n22388 = n22387 ^ x154 ^ 1'b0 ;
  assign n22389 = n18965 ^ n11837 ^ n10433 ;
  assign n22390 = n13740 & ~n22389 ;
  assign n22391 = n979 & ~n22390 ;
  assign n22392 = n2740 & ~n20136 ;
  assign n22393 = n22392 ^ n6642 ^ 1'b0 ;
  assign n22394 = n5650 ^ n861 ^ 1'b0 ;
  assign n22395 = n22394 ^ n17201 ^ n445 ;
  assign n22396 = n1359 | n22395 ;
  assign n22397 = n2243 & ~n10606 ;
  assign n22398 = x205 & n22397 ;
  assign n22399 = n5862 & n22398 ;
  assign n22400 = n8306 & n22399 ;
  assign n22401 = n9328 ^ n7713 ^ 1'b0 ;
  assign n22402 = n22401 ^ n8490 ^ 1'b0 ;
  assign n22403 = n16427 ^ n10557 ^ 1'b0 ;
  assign n22404 = ~n3878 & n13496 ;
  assign n22405 = ~n3783 & n22404 ;
  assign n22406 = ( n2724 & n5288 ) | ( n2724 & ~n14091 ) | ( n5288 & ~n14091 ) ;
  assign n22407 = n12319 & ~n14836 ;
  assign n22408 = ( n851 & n22406 ) | ( n851 & ~n22407 ) | ( n22406 & ~n22407 ) ;
  assign n22409 = n15150 ^ n9380 ^ 1'b0 ;
  assign n22410 = n20844 & ~n22409 ;
  assign n22411 = n12733 ^ n11544 ^ 1'b0 ;
  assign n22412 = n6025 & n22411 ;
  assign n22413 = ( n3117 & ~n9814 ) | ( n3117 & n16959 ) | ( ~n9814 & n16959 ) ;
  assign n22414 = ~n607 & n14579 ;
  assign n22415 = n9299 & n22414 ;
  assign n22416 = ( n5425 & ~n22413 ) | ( n5425 & n22415 ) | ( ~n22413 & n22415 ) ;
  assign n22417 = n6009 & ~n22416 ;
  assign n22418 = ( n3323 & n9882 ) | ( n3323 & n10160 ) | ( n9882 & n10160 ) ;
  assign n22419 = ~n12869 & n17928 ;
  assign n22420 = ~n1010 & n22419 ;
  assign n22421 = ~n22418 & n22420 ;
  assign n22422 = n22111 ^ n8789 ^ n3897 ;
  assign n22423 = n22422 ^ n17586 ^ n16863 ;
  assign n22424 = n17014 ^ n11245 ^ n464 ;
  assign n22425 = ( n9351 & n18803 ) | ( n9351 & n22424 ) | ( n18803 & n22424 ) ;
  assign n22426 = ~n8343 & n10037 ;
  assign n22427 = ~n2685 & n22426 ;
  assign n22428 = n13776 ^ n12750 ^ n4212 ;
  assign n22429 = ( n573 & n916 ) | ( n573 & ~n16456 ) | ( n916 & ~n16456 ) ;
  assign n22430 = n21990 ^ n8175 ^ 1'b0 ;
  assign n22431 = n14029 ^ n3366 ^ 1'b0 ;
  assign n22432 = n8148 & ~n22431 ;
  assign n22433 = n2497 | n7064 ;
  assign n22434 = n22433 ^ n10976 ^ n1503 ;
  assign n22435 = n15663 | n22434 ;
  assign n22437 = n7673 ^ n2565 ^ 1'b0 ;
  assign n22438 = n2815 & n22437 ;
  assign n22439 = n2576 & ~n22438 ;
  assign n22436 = ~n3730 & n17140 ;
  assign n22440 = n22439 ^ n22436 ^ n675 ;
  assign n22441 = x105 | n495 ;
  assign n22442 = ( n16587 & n21720 ) | ( n16587 & ~n22441 ) | ( n21720 & ~n22441 ) ;
  assign n22443 = ( n6791 & n12071 ) | ( n6791 & ~n14975 ) | ( n12071 & ~n14975 ) ;
  assign n22444 = n16486 ^ n15068 ^ 1'b0 ;
  assign n22445 = n22443 | n22444 ;
  assign n22447 = n1687 | n16529 ;
  assign n22448 = n22447 ^ n14578 ^ 1'b0 ;
  assign n22446 = n5492 | n10492 ;
  assign n22449 = n22448 ^ n22446 ^ 1'b0 ;
  assign n22450 = n7577 ^ x60 ^ 1'b0 ;
  assign n22451 = n9193 & ~n22450 ;
  assign n22452 = ( n12558 & n12745 ) | ( n12558 & ~n22451 ) | ( n12745 & ~n22451 ) ;
  assign n22453 = n6023 & ~n22452 ;
  assign n22454 = n22449 & ~n22453 ;
  assign n22455 = ~n18281 & n22454 ;
  assign n22456 = n10299 ^ n6008 ^ 1'b0 ;
  assign n22457 = n22456 ^ n12622 ^ 1'b0 ;
  assign n22458 = n20026 | n21938 ;
  assign n22459 = n22457 | n22458 ;
  assign n22460 = ~n10714 & n19060 ;
  assign n22461 = ( ~n9798 & n13496 ) | ( ~n9798 & n22460 ) | ( n13496 & n22460 ) ;
  assign n22462 = n1173 & ~n17651 ;
  assign n22463 = n22462 ^ n4346 ^ 1'b0 ;
  assign n22464 = n22463 ^ n18258 ^ 1'b0 ;
  assign n22465 = ~n17509 & n22464 ;
  assign n22466 = n22465 ^ n1701 ^ n600 ;
  assign n22468 = ( n414 & ~n8301 ) | ( n414 & n21800 ) | ( ~n8301 & n21800 ) ;
  assign n22469 = ~n13459 & n22468 ;
  assign n22470 = n22469 ^ n12862 ^ 1'b0 ;
  assign n22471 = n17323 & ~n22470 ;
  assign n22472 = ( n9300 & ~n9907 ) | ( n9300 & n11527 ) | ( ~n9907 & n11527 ) ;
  assign n22473 = n22472 ^ n7528 ^ n6493 ;
  assign n22474 = ~n17803 & n22473 ;
  assign n22475 = n22471 & n22474 ;
  assign n22467 = ( n434 & n9098 ) | ( n434 & n15558 ) | ( n9098 & n15558 ) ;
  assign n22476 = n22475 ^ n22467 ^ n13546 ;
  assign n22477 = ~n9420 & n12798 ;
  assign n22478 = n12861 & n22477 ;
  assign n22479 = ( n5961 & n12393 ) | ( n5961 & ~n22478 ) | ( n12393 & ~n22478 ) ;
  assign n22480 = n5912 ^ n5682 ^ 1'b0 ;
  assign n22481 = n6066 & n22480 ;
  assign n22482 = n12233 & n16317 ;
  assign n22483 = ~n22481 & n22482 ;
  assign n22484 = n20225 | n21571 ;
  assign n22485 = n22483 & ~n22484 ;
  assign n22486 = n6256 ^ n5284 ^ n4289 ;
  assign n22487 = n3641 ^ n1958 ^ 1'b0 ;
  assign n22488 = n22486 | n22487 ;
  assign n22489 = n22488 ^ n18337 ^ 1'b0 ;
  assign n22490 = ~n713 & n1427 ;
  assign n22491 = n22490 ^ n4265 ^ 1'b0 ;
  assign n22492 = n22491 ^ n5601 ^ n1431 ;
  assign n22493 = n3261 ^ n2944 ^ n322 ;
  assign n22494 = n22493 ^ n16892 ^ 1'b0 ;
  assign n22495 = n15663 | n22494 ;
  assign n22496 = n22495 ^ n1861 ^ n703 ;
  assign n22497 = n22496 ^ n12718 ^ 1'b0 ;
  assign n22498 = ~n15967 & n22497 ;
  assign n22499 = n11809 & n22498 ;
  assign n22500 = n22499 ^ n1037 ^ 1'b0 ;
  assign n22501 = n16555 ^ n16338 ^ 1'b0 ;
  assign n22502 = n6490 & n22501 ;
  assign n22503 = n22343 ^ n17209 ^ n11008 ;
  assign n22504 = n15078 ^ n11990 ^ n9130 ;
  assign n22505 = n22504 ^ n14592 ^ 1'b0 ;
  assign n22506 = n8807 | n22505 ;
  assign n22507 = n6043 | n7160 ;
  assign n22508 = n20750 ^ n2286 ^ 1'b0 ;
  assign n22509 = n8347 & n22508 ;
  assign n22510 = n22509 ^ n7503 ^ 1'b0 ;
  assign n22511 = n22507 | n22510 ;
  assign n22512 = n2740 | n11363 ;
  assign n22513 = ( n7625 & n14233 ) | ( n7625 & ~n22512 ) | ( n14233 & ~n22512 ) ;
  assign n22514 = n22451 ^ n22394 ^ 1'b0 ;
  assign n22515 = n22514 ^ n21465 ^ n6641 ;
  assign n22518 = ( n5012 & n12143 ) | ( n5012 & n17431 ) | ( n12143 & n17431 ) ;
  assign n22516 = n1353 | n12998 ;
  assign n22517 = n10312 & ~n22516 ;
  assign n22519 = n22518 ^ n22517 ^ n13211 ;
  assign n22520 = n22519 ^ n11390 ^ n10728 ;
  assign n22521 = n22520 ^ n19290 ^ n7421 ;
  assign n22522 = ( ~n4573 & n7581 ) | ( ~n4573 & n10988 ) | ( n7581 & n10988 ) ;
  assign n22523 = ( n4845 & n12634 ) | ( n4845 & ~n22522 ) | ( n12634 & ~n22522 ) ;
  assign n22524 = n22523 ^ n17695 ^ n3941 ;
  assign n22525 = n22524 ^ n6843 ^ 1'b0 ;
  assign n22526 = n9427 & ~n22525 ;
  assign n22527 = ( n731 & ~n2788 ) | ( n731 & n9452 ) | ( ~n2788 & n9452 ) ;
  assign n22528 = n887 & n6876 ;
  assign n22529 = n22527 & ~n22528 ;
  assign n22530 = ~n4098 & n22529 ;
  assign n22532 = n20870 ^ n18302 ^ 1'b0 ;
  assign n22533 = n1385 & ~n22532 ;
  assign n22531 = ~n5292 & n16612 ;
  assign n22534 = n22533 ^ n22531 ^ n10699 ;
  assign n22535 = n16434 ^ n16047 ^ 1'b0 ;
  assign n22537 = n12406 ^ n9691 ^ 1'b0 ;
  assign n22536 = n9555 & n18543 ;
  assign n22538 = n22537 ^ n22536 ^ 1'b0 ;
  assign n22539 = ( n21798 & n22535 ) | ( n21798 & ~n22538 ) | ( n22535 & ~n22538 ) ;
  assign n22540 = n1757 | n7342 ;
  assign n22541 = n22540 ^ n1775 ^ 1'b0 ;
  assign n22542 = n5553 ^ n3734 ^ 1'b0 ;
  assign n22543 = n22541 & n22542 ;
  assign n22544 = ~n1269 & n15741 ;
  assign n22545 = n9256 ^ n9003 ^ 1'b0 ;
  assign n22546 = n7014 & ~n22545 ;
  assign n22547 = ( n17476 & n20791 ) | ( n17476 & ~n22546 ) | ( n20791 & ~n22546 ) ;
  assign n22548 = ( ~n1875 & n5000 ) | ( ~n1875 & n12313 ) | ( n5000 & n12313 ) ;
  assign n22549 = ( n3234 & n8008 ) | ( n3234 & ~n22548 ) | ( n8008 & ~n22548 ) ;
  assign n22550 = n7392 | n20851 ;
  assign n22551 = ~n15510 & n22550 ;
  assign n22552 = n22551 ^ n562 ^ 1'b0 ;
  assign n22553 = n10113 & ~n17953 ;
  assign n22554 = n22553 ^ n1421 ^ 1'b0 ;
  assign n22560 = n560 & ~n1997 ;
  assign n22559 = ~n9846 & n13490 ;
  assign n22555 = n1640 & ~n6053 ;
  assign n22556 = n22555 ^ n4123 ^ 1'b0 ;
  assign n22557 = x148 & n22556 ;
  assign n22558 = n22557 ^ n7360 ^ n4970 ;
  assign n22561 = n22560 ^ n22559 ^ n22558 ;
  assign n22562 = ( n14366 & ~n17379 ) | ( n14366 & n22561 ) | ( ~n17379 & n22561 ) ;
  assign n22563 = ( n982 & ~n5880 ) | ( n982 & n13232 ) | ( ~n5880 & n13232 ) ;
  assign n22564 = n2696 | n22563 ;
  assign n22565 = ~n410 & n6935 ;
  assign n22566 = n22565 ^ n12788 ^ 1'b0 ;
  assign n22567 = n22564 & ~n22566 ;
  assign n22568 = n13757 & ~n22567 ;
  assign n22569 = n22568 ^ n21281 ^ 1'b0 ;
  assign n22570 = ( n9013 & n15763 ) | ( n9013 & ~n22569 ) | ( n15763 & ~n22569 ) ;
  assign n22573 = ~n9037 & n15394 ;
  assign n22571 = ( n3409 & n12411 ) | ( n3409 & n14406 ) | ( n12411 & n14406 ) ;
  assign n22572 = ( ~n8848 & n16431 ) | ( ~n8848 & n22571 ) | ( n16431 & n22571 ) ;
  assign n22574 = n22573 ^ n22572 ^ n4490 ;
  assign n22575 = n21505 ^ n16117 ^ 1'b0 ;
  assign n22576 = ( n2194 & n9064 ) | ( n2194 & n22575 ) | ( n9064 & n22575 ) ;
  assign n22577 = n8122 ^ n6793 ^ 1'b0 ;
  assign n22578 = ~n4550 & n22577 ;
  assign n22579 = ~n4129 & n20545 ;
  assign n22580 = ~n22578 & n22579 ;
  assign n22581 = n17999 ^ n7826 ^ 1'b0 ;
  assign n22582 = n22581 ^ n18338 ^ n11488 ;
  assign n22583 = n10935 ^ n915 ^ 1'b0 ;
  assign n22584 = n4554 | n22583 ;
  assign n22585 = n11574 ^ n2110 ^ 1'b0 ;
  assign n22586 = ~n5457 & n12053 ;
  assign n22587 = n22585 & n22586 ;
  assign n22588 = n19928 ^ n19299 ^ 1'b0 ;
  assign n22589 = n7947 & ~n12843 ;
  assign n22590 = n4871 & n22589 ;
  assign n22591 = n22590 ^ n9217 ^ 1'b0 ;
  assign n22592 = ( n4152 & ~n8781 ) | ( n4152 & n9399 ) | ( ~n8781 & n9399 ) ;
  assign n22593 = n21168 ^ n7231 ^ 1'b0 ;
  assign n22594 = ( n4556 & n13227 ) | ( n4556 & ~n22593 ) | ( n13227 & ~n22593 ) ;
  assign n22595 = ~n706 & n12750 ;
  assign n22596 = ~n22594 & n22595 ;
  assign n22597 = ~n4816 & n22596 ;
  assign n22598 = ( n20437 & n22592 ) | ( n20437 & n22597 ) | ( n22592 & n22597 ) ;
  assign n22599 = ( n20148 & ~n21890 ) | ( n20148 & n22598 ) | ( ~n21890 & n22598 ) ;
  assign n22600 = x156 & n7235 ;
  assign n22601 = n17971 ^ n9554 ^ 1'b0 ;
  assign n22602 = ~n22600 & n22601 ;
  assign n22603 = ( n2774 & n12740 ) | ( n2774 & ~n22602 ) | ( n12740 & ~n22602 ) ;
  assign n22604 = n3369 & n17837 ;
  assign n22605 = ~n4240 & n22604 ;
  assign n22606 = ~n12466 & n22605 ;
  assign n22607 = x153 & n1277 ;
  assign n22608 = n22607 ^ n19769 ^ n8608 ;
  assign n22609 = n19584 ^ n6245 ^ 1'b0 ;
  assign n22610 = n22608 & n22609 ;
  assign n22611 = n6006 ^ n1412 ^ 1'b0 ;
  assign n22612 = n1401 | n12669 ;
  assign n22613 = n5775 | n22612 ;
  assign n22614 = n14546 ^ n2981 ^ 1'b0 ;
  assign n22615 = n22613 & n22614 ;
  assign n22616 = ( n5122 & ~n19691 ) | ( n5122 & n21585 ) | ( ~n19691 & n21585 ) ;
  assign n22617 = ~n6878 & n22616 ;
  assign n22618 = ~n963 & n7908 ;
  assign n22619 = n284 & n22618 ;
  assign n22620 = n9699 ^ n8399 ^ 1'b0 ;
  assign n22621 = n6809 | n22620 ;
  assign n22622 = n5015 | n22621 ;
  assign n22623 = n20627 & ~n22622 ;
  assign n22624 = n22623 ^ n17875 ^ n2114 ;
  assign n22625 = n9422 | n22624 ;
  assign n22626 = n22619 & ~n22625 ;
  assign n22627 = n13310 ^ n2586 ^ 1'b0 ;
  assign n22628 = ( ~n8431 & n9412 ) | ( ~n8431 & n14390 ) | ( n9412 & n14390 ) ;
  assign n22629 = ( n15391 & ~n18850 ) | ( n15391 & n22628 ) | ( ~n18850 & n22628 ) ;
  assign n22630 = n22629 ^ n8894 ^ 1'b0 ;
  assign n22634 = ( ~n2405 & n6297 ) | ( ~n2405 & n7216 ) | ( n6297 & n7216 ) ;
  assign n22635 = n22634 ^ n13396 ^ 1'b0 ;
  assign n22631 = ( n2260 & ~n10043 ) | ( n2260 & n22034 ) | ( ~n10043 & n22034 ) ;
  assign n22632 = n22631 ^ n3223 ^ 1'b0 ;
  assign n22633 = ~n4080 & n22632 ;
  assign n22636 = n22635 ^ n22633 ^ n21448 ;
  assign n22637 = n4598 & ~n22636 ;
  assign n22638 = ~n5105 & n14114 ;
  assign n22639 = n22638 ^ n2448 ^ 1'b0 ;
  assign n22640 = n384 | n22639 ;
  assign n22641 = n22640 ^ n9304 ^ 1'b0 ;
  assign n22642 = n22641 ^ n10994 ^ 1'b0 ;
  assign n22643 = n3322 | n15022 ;
  assign n22644 = n18351 ^ n1902 ^ 1'b0 ;
  assign n22645 = n908 & n22644 ;
  assign n22646 = n5683 & n22645 ;
  assign n22647 = ~n4093 & n22646 ;
  assign n22648 = n8612 & ~n22647 ;
  assign n22649 = ~n18844 & n22648 ;
  assign n22650 = n22649 ^ n806 ^ 1'b0 ;
  assign n22651 = ~n3012 & n22650 ;
  assign n22652 = ~n16542 & n22651 ;
  assign n22653 = n22652 ^ n3776 ^ 1'b0 ;
  assign n22654 = ~n4051 & n22653 ;
  assign n22655 = n9749 ^ n8754 ^ n4358 ;
  assign n22656 = n12795 & n14415 ;
  assign n22657 = n11542 ^ n4694 ^ 1'b0 ;
  assign n22659 = n2234 & ~n19501 ;
  assign n22660 = ~n10719 & n22659 ;
  assign n22658 = x21 | n608 ;
  assign n22661 = n22660 ^ n22658 ^ n21729 ;
  assign n22662 = n12289 ^ n1249 ^ 1'b0 ;
  assign n22663 = n22662 ^ n11050 ^ n9816 ;
  assign n22664 = n3717 & ~n9776 ;
  assign n22665 = n22664 ^ n20276 ^ 1'b0 ;
  assign n22668 = ( n1475 & n5605 ) | ( n1475 & n18512 ) | ( n5605 & n18512 ) ;
  assign n22669 = ( n8952 & ~n9416 ) | ( n8952 & n22668 ) | ( ~n9416 & n22668 ) ;
  assign n22666 = n12928 ^ n5946 ^ 1'b0 ;
  assign n22667 = n19011 & n22666 ;
  assign n22670 = n22669 ^ n22667 ^ n291 ;
  assign n22671 = ~n13813 & n17526 ;
  assign n22672 = n22671 ^ n20759 ^ 1'b0 ;
  assign n22679 = n21022 ^ n13693 ^ n11996 ;
  assign n22673 = n4267 ^ n4240 ^ 1'b0 ;
  assign n22674 = n8949 & ~n22673 ;
  assign n22675 = ( ~n4932 & n8915 ) | ( ~n4932 & n22021 ) | ( n8915 & n22021 ) ;
  assign n22676 = n22674 & ~n22675 ;
  assign n22677 = n22676 ^ n10382 ^ 1'b0 ;
  assign n22678 = n2252 | n22677 ;
  assign n22680 = n22679 ^ n22678 ^ n16729 ;
  assign n22681 = n22680 ^ n18531 ^ n13272 ;
  assign n22683 = x237 ^ x50 ^ 1'b0 ;
  assign n22682 = n1279 & n15857 ;
  assign n22684 = n22683 ^ n22682 ^ 1'b0 ;
  assign n22685 = n1588 | n7007 ;
  assign n22686 = n8893 ^ n7592 ^ 1'b0 ;
  assign n22687 = ~n1953 & n22686 ;
  assign n22688 = ( n7801 & n22685 ) | ( n7801 & ~n22687 ) | ( n22685 & ~n22687 ) ;
  assign n22689 = n5763 & ~n14393 ;
  assign n22690 = n22689 ^ n3817 ^ 1'b0 ;
  assign n22691 = n22688 | n22690 ;
  assign n22692 = n20767 ^ n8769 ^ 1'b0 ;
  assign n22693 = n5544 & ~n22692 ;
  assign n22694 = n2329 & n22693 ;
  assign n22696 = n9970 ^ n8733 ^ n755 ;
  assign n22695 = n6428 & n12792 ;
  assign n22697 = n22696 ^ n22695 ^ n409 ;
  assign n22698 = n10695 ^ n6108 ^ 1'b0 ;
  assign n22699 = n22698 ^ n20415 ^ 1'b0 ;
  assign n22700 = n1124 ^ n720 ^ x163 ;
  assign n22701 = n14623 & ~n22700 ;
  assign n22702 = n9394 ^ n5034 ^ n4046 ;
  assign n22703 = n7263 & ~n22702 ;
  assign n22704 = ~n9702 & n22703 ;
  assign n22705 = ~n7910 & n22704 ;
  assign n22706 = n3456 | n3946 ;
  assign n22707 = n22706 ^ n11188 ^ 1'b0 ;
  assign n22708 = n11025 | n22707 ;
  assign n22709 = n11025 & ~n22708 ;
  assign n22710 = ~n6423 & n22709 ;
  assign n22711 = n12415 ^ n1461 ^ n1228 ;
  assign n22712 = n22711 ^ n12015 ^ n5683 ;
  assign n22713 = n9739 | n9872 ;
  assign n22714 = n22713 ^ n13972 ^ 1'b0 ;
  assign n22715 = n22712 | n22714 ;
  assign n22716 = ~n4117 & n13456 ;
  assign n22717 = n22716 ^ n5298 ^ 1'b0 ;
  assign n22718 = ~n12728 & n22717 ;
  assign n22719 = n22718 ^ n6871 ^ 1'b0 ;
  assign n22720 = n22719 ^ n15088 ^ n8406 ;
  assign n22721 = n12287 & n22720 ;
  assign n22722 = n14139 ^ n14016 ^ n7148 ;
  assign n22723 = n22722 ^ n2421 ^ n421 ;
  assign n22724 = ( n2551 & n4198 ) | ( n2551 & n4906 ) | ( n4198 & n4906 ) ;
  assign n22725 = n8409 ^ n2509 ^ n1520 ;
  assign n22726 = n22724 & n22725 ;
  assign n22727 = n2602 | n22726 ;
  assign n22728 = n6124 & ~n13170 ;
  assign n22729 = n22728 ^ n20859 ^ 1'b0 ;
  assign n22730 = n15588 ^ x11 ^ 1'b0 ;
  assign n22731 = ( n3937 & n6181 ) | ( n3937 & n11571 ) | ( n6181 & n11571 ) ;
  assign n22732 = n15506 ^ n7264 ^ 1'b0 ;
  assign n22733 = n13668 ^ n11534 ^ 1'b0 ;
  assign n22734 = n22732 | n22733 ;
  assign n22735 = n22734 ^ n14953 ^ n3101 ;
  assign n22736 = n391 & n9863 ;
  assign n22737 = n22736 ^ n21848 ^ 1'b0 ;
  assign n22738 = n11083 ^ n1068 ^ 1'b0 ;
  assign n22739 = n22738 ^ n20182 ^ 1'b0 ;
  assign n22740 = n3679 & ~n22739 ;
  assign n22741 = n11816 ^ n9665 ^ n7913 ;
  assign n22742 = ( n9201 & n16489 ) | ( n9201 & ~n22741 ) | ( n16489 & ~n22741 ) ;
  assign n22743 = n12302 | n22742 ;
  assign n22744 = n14644 | n22743 ;
  assign n22748 = n13575 ^ n5207 ^ n2986 ;
  assign n22745 = ~n586 & n18841 ;
  assign n22746 = n22745 ^ n8557 ^ 1'b0 ;
  assign n22747 = n5406 | n22746 ;
  assign n22749 = n22748 ^ n22747 ^ 1'b0 ;
  assign n22750 = ( ~n3535 & n4281 ) | ( ~n3535 & n10525 ) | ( n4281 & n10525 ) ;
  assign n22751 = n15676 ^ n13474 ^ 1'b0 ;
  assign n22752 = n22750 & ~n22751 ;
  assign n22753 = n8402 ^ n299 ^ 1'b0 ;
  assign n22754 = ~n3492 & n22753 ;
  assign n22755 = ~n22752 & n22754 ;
  assign n22756 = n11348 ^ n10647 ^ 1'b0 ;
  assign n22757 = n22756 ^ n10018 ^ 1'b0 ;
  assign n22758 = n471 | n3196 ;
  assign n22759 = n471 & ~n22758 ;
  assign n22760 = n900 | n13929 ;
  assign n22761 = n22760 ^ n13572 ^ 1'b0 ;
  assign n22762 = ( n1054 & n22759 ) | ( n1054 & ~n22761 ) | ( n22759 & ~n22761 ) ;
  assign n22765 = n9424 & ~n13335 ;
  assign n22763 = n14283 ^ n9782 ^ 1'b0 ;
  assign n22764 = n4080 | n22763 ;
  assign n22766 = n22765 ^ n22764 ^ n3299 ;
  assign n22767 = n1508 & ~n4830 ;
  assign n22768 = ( ~n20112 & n21639 ) | ( ~n20112 & n22767 ) | ( n21639 & n22767 ) ;
  assign n22769 = n19965 ^ n2217 ^ 1'b0 ;
  assign n22770 = ~n14632 & n22769 ;
  assign n22771 = n20940 ^ n18054 ^ n12803 ;
  assign n22772 = ( ~n6139 & n7819 ) | ( ~n6139 & n18841 ) | ( n7819 & n18841 ) ;
  assign n22773 = n19262 ^ n10063 ^ 1'b0 ;
  assign n22774 = ( n13364 & n22772 ) | ( n13364 & ~n22773 ) | ( n22772 & ~n22773 ) ;
  assign n22775 = n22774 ^ n19108 ^ n633 ;
  assign n22776 = n3205 ^ n884 ^ 1'b0 ;
  assign n22777 = n9246 & ~n13417 ;
  assign n22778 = ~n4016 & n22777 ;
  assign n22779 = n1494 & n3796 ;
  assign n22780 = n22779 ^ n11963 ^ n9015 ;
  assign n22781 = n20897 ^ n1059 ^ 1'b0 ;
  assign n22782 = n6428 & ~n12977 ;
  assign n22783 = n18676 ^ n1873 ^ 1'b0 ;
  assign n22784 = ~n10603 & n22783 ;
  assign n22785 = n13364 ^ n10753 ^ 1'b0 ;
  assign n22786 = n22785 ^ n21551 ^ n14120 ;
  assign n22787 = n12740 | n21729 ;
  assign n22788 = n6481 | n10110 ;
  assign n22789 = n10532 | n14892 ;
  assign n22790 = n22789 ^ n20266 ^ 1'b0 ;
  assign n22791 = ( ~n6333 & n22788 ) | ( ~n6333 & n22790 ) | ( n22788 & n22790 ) ;
  assign n22792 = n6064 ^ n4737 ^ 1'b0 ;
  assign n22793 = n22792 ^ n19836 ^ 1'b0 ;
  assign n22794 = n20349 | n22793 ;
  assign n22807 = ( ~n1948 & n2336 ) | ( ~n1948 & n4993 ) | ( n2336 & n4993 ) ;
  assign n22804 = n1327 ^ n749 ^ 1'b0 ;
  assign n22805 = n18349 | n22804 ;
  assign n22806 = n22805 ^ n4952 ^ x254 ;
  assign n22808 = n22807 ^ n22806 ^ n22285 ;
  assign n22796 = n7766 ^ n3775 ^ n1148 ;
  assign n22797 = ~n9666 & n19604 ;
  assign n22798 = ~n10974 & n22797 ;
  assign n22799 = n12020 ^ n4045 ^ 1'b0 ;
  assign n22800 = n12100 ^ n9021 ^ 1'b0 ;
  assign n22801 = n22799 | n22800 ;
  assign n22802 = ( n22796 & n22798 ) | ( n22796 & ~n22801 ) | ( n22798 & ~n22801 ) ;
  assign n22795 = n8063 & ~n15057 ;
  assign n22803 = n22802 ^ n22795 ^ 1'b0 ;
  assign n22809 = n22808 ^ n22803 ^ 1'b0 ;
  assign n22810 = ~n22794 & n22809 ;
  assign n22812 = ( x4 & ~n13717 ) | ( x4 & n14587 ) | ( ~n13717 & n14587 ) ;
  assign n22811 = n6241 | n7487 ;
  assign n22813 = n22812 ^ n22811 ^ 1'b0 ;
  assign n22814 = n12331 ^ n5823 ^ n4516 ;
  assign n22815 = n20428 & ~n22814 ;
  assign n22816 = n10253 ^ n3613 ^ 1'b0 ;
  assign n22817 = n22816 ^ n16047 ^ n11403 ;
  assign n22818 = ~n11620 & n22817 ;
  assign n22819 = n22818 ^ n20467 ^ n2442 ;
  assign n22820 = n6022 | n14938 ;
  assign n22821 = n22820 ^ n13240 ^ n11843 ;
  assign n22822 = n19778 ^ n16448 ^ n13021 ;
  assign n22823 = n22821 | n22822 ;
  assign n22826 = n2268 & n19295 ;
  assign n22827 = n3926 & n15529 ;
  assign n22828 = ~n22826 & n22827 ;
  assign n22829 = n22828 ^ n8729 ^ 1'b0 ;
  assign n22824 = ~n9501 & n9654 ;
  assign n22825 = ~n13563 & n22824 ;
  assign n22830 = n22829 ^ n22825 ^ 1'b0 ;
  assign n22831 = ~n14499 & n21902 ;
  assign n22832 = n22831 ^ n21119 ^ 1'b0 ;
  assign n22833 = n9095 & ~n13039 ;
  assign n22834 = ~n10472 & n22833 ;
  assign n22838 = ~n2051 & n10968 ;
  assign n22835 = ( n1912 & n6066 ) | ( n1912 & n11570 ) | ( n6066 & n11570 ) ;
  assign n22836 = n22835 ^ n19267 ^ n17339 ;
  assign n22837 = n14207 & n22836 ;
  assign n22839 = n22838 ^ n22837 ^ 1'b0 ;
  assign n22840 = x176 & n1595 ;
  assign n22841 = ( n3553 & n8802 ) | ( n3553 & ~n22840 ) | ( n8802 & ~n22840 ) ;
  assign n22842 = n22841 ^ n3496 ^ 1'b0 ;
  assign n22846 = ( n3240 & ~n4526 ) | ( n3240 & n6260 ) | ( ~n4526 & n6260 ) ;
  assign n22847 = ( ~n914 & n6732 ) | ( ~n914 & n22846 ) | ( n6732 & n22846 ) ;
  assign n22848 = ( n15816 & n21081 ) | ( n15816 & n22847 ) | ( n21081 & n22847 ) ;
  assign n22843 = n3247 & ~n6524 ;
  assign n22844 = n22843 ^ n2753 ^ 1'b0 ;
  assign n22845 = n12331 | n22844 ;
  assign n22849 = n22848 ^ n22845 ^ 1'b0 ;
  assign n22850 = n14198 & ~n15656 ;
  assign n22851 = n22850 ^ n11766 ^ 1'b0 ;
  assign n22852 = n5980 ^ n4912 ^ 1'b0 ;
  assign n22853 = ( n2243 & ~n2502 ) | ( n2243 & n5250 ) | ( ~n2502 & n5250 ) ;
  assign n22854 = ( n436 & n2194 ) | ( n436 & n22853 ) | ( n2194 & n22853 ) ;
  assign n22855 = ~n1852 & n22854 ;
  assign n22856 = n7511 ^ n5971 ^ 1'b0 ;
  assign n22857 = n22855 | n22856 ;
  assign n22858 = ( n22851 & ~n22852 ) | ( n22851 & n22857 ) | ( ~n22852 & n22857 ) ;
  assign n22859 = n22820 ^ n22621 ^ 1'b0 ;
  assign n22860 = n22858 | n22859 ;
  assign n22861 = n2970 | n22719 ;
  assign n22862 = ( n6872 & n18318 ) | ( n6872 & n22861 ) | ( n18318 & n22861 ) ;
  assign n22863 = ( ~n1916 & n16959 ) | ( ~n1916 & n22862 ) | ( n16959 & n22862 ) ;
  assign n22864 = ~n1027 & n8442 ;
  assign n22865 = n13177 & ~n18975 ;
  assign n22866 = n22864 & n22865 ;
  assign n22867 = ~n5751 & n22866 ;
  assign n22868 = ( n4409 & ~n16266 ) | ( n4409 & n21591 ) | ( ~n16266 & n21591 ) ;
  assign n22869 = n22867 | n22868 ;
  assign n22870 = n22452 ^ n7252 ^ 1'b0 ;
  assign n22871 = n20104 ^ n5488 ^ n1168 ;
  assign n22872 = n22871 ^ n1184 ^ 1'b0 ;
  assign n22873 = n14653 | n22872 ;
  assign n22874 = ( n16842 & n22870 ) | ( n16842 & n22873 ) | ( n22870 & n22873 ) ;
  assign n22875 = n12819 ^ n5150 ^ 1'b0 ;
  assign n22876 = ~n14742 & n22875 ;
  assign n22877 = n6538 & n12016 ;
  assign n22878 = n22877 ^ n7163 ^ 1'b0 ;
  assign n22879 = n7481 ^ n3299 ^ n594 ;
  assign n22880 = ( n7867 & n11645 ) | ( n7867 & n22879 ) | ( n11645 & n22879 ) ;
  assign n22881 = n15212 & ~n15598 ;
  assign n22882 = ~n4793 & n21971 ;
  assign n22883 = ~n22881 & n22882 ;
  assign n22884 = n17961 ^ n5557 ^ 1'b0 ;
  assign n22885 = n12792 ^ n2515 ^ 1'b0 ;
  assign n22886 = n22885 ^ n17723 ^ n9149 ;
  assign n22887 = ~n5793 & n8055 ;
  assign n22888 = n22887 ^ n5902 ^ 1'b0 ;
  assign n22889 = n22888 ^ n12428 ^ 1'b0 ;
  assign n22890 = ( n4450 & n7009 ) | ( n4450 & ~n12530 ) | ( n7009 & ~n12530 ) ;
  assign n22893 = n10713 ^ n3834 ^ 1'b0 ;
  assign n22894 = ~n9772 & n22893 ;
  assign n22891 = n8484 | n13528 ;
  assign n22892 = n1864 | n22891 ;
  assign n22895 = n22894 ^ n22892 ^ 1'b0 ;
  assign n22896 = n1173 & n13738 ;
  assign n22897 = n22896 ^ n15456 ^ n7173 ;
  assign n22898 = ~n1074 & n1554 ;
  assign n22899 = n22898 ^ x246 ^ 1'b0 ;
  assign n22900 = n22899 ^ n13720 ^ 1'b0 ;
  assign n22901 = ( n5710 & ~n13752 ) | ( n5710 & n18082 ) | ( ~n13752 & n18082 ) ;
  assign n22902 = n11506 ^ n11234 ^ 1'b0 ;
  assign n22903 = ~n5933 & n22902 ;
  assign n22904 = n12737 ^ n5399 ^ 1'b0 ;
  assign n22905 = n22904 ^ n8016 ^ 1'b0 ;
  assign n22906 = n22903 & ~n22905 ;
  assign n22907 = ( x135 & ~n2140 ) | ( x135 & n8262 ) | ( ~n2140 & n8262 ) ;
  assign n22908 = ( ~n452 & n6949 ) | ( ~n452 & n22907 ) | ( n6949 & n22907 ) ;
  assign n22909 = n22908 ^ n9033 ^ n4761 ;
  assign n22910 = n13920 ^ n8508 ^ n2927 ;
  assign n22911 = n11592 ^ n3399 ^ 1'b0 ;
  assign n22912 = n22911 ^ n11702 ^ x153 ;
  assign n22913 = n22912 ^ n5025 ^ 1'b0 ;
  assign n22914 = n21459 & n22913 ;
  assign n22915 = ( n4777 & n5581 ) | ( n4777 & ~n8487 ) | ( n5581 & ~n8487 ) ;
  assign n22916 = ( n1062 & n7138 ) | ( n1062 & n22915 ) | ( n7138 & n22915 ) ;
  assign n22917 = ( n22910 & n22914 ) | ( n22910 & n22916 ) | ( n22914 & n22916 ) ;
  assign n22918 = n2634 | n19640 ;
  assign n22919 = ( n11968 & n12194 ) | ( n11968 & n22918 ) | ( n12194 & n22918 ) ;
  assign n22920 = n22919 ^ n17456 ^ 1'b0 ;
  assign n22922 = n10989 & n14733 ;
  assign n22923 = n22922 ^ n15791 ^ 1'b0 ;
  assign n22921 = ( n1488 & n8531 ) | ( n1488 & n8949 ) | ( n8531 & n8949 ) ;
  assign n22924 = n22923 ^ n22921 ^ 1'b0 ;
  assign n22927 = n13342 ^ n3382 ^ 1'b0 ;
  assign n22928 = n4026 & ~n22927 ;
  assign n22926 = ( n1209 & ~n5097 ) | ( n1209 & n5671 ) | ( ~n5097 & n5671 ) ;
  assign n22929 = n22928 ^ n22926 ^ n5938 ;
  assign n22925 = n8824 ^ n6753 ^ n5222 ;
  assign n22930 = n22929 ^ n22925 ^ n22364 ;
  assign n22931 = n10761 ^ n5646 ^ 1'b0 ;
  assign n22932 = n10504 & n22931 ;
  assign n22933 = n22932 ^ n9953 ^ 1'b0 ;
  assign n22934 = n7347 & n19602 ;
  assign n22935 = n7696 | n22934 ;
  assign n22938 = n1627 | n12483 ;
  assign n22936 = n12837 | n13711 ;
  assign n22937 = n2195 | n22936 ;
  assign n22939 = n22938 ^ n22937 ^ 1'b0 ;
  assign n22940 = n1779 & n22939 ;
  assign n22941 = n2693 ^ n1142 ^ 1'b0 ;
  assign n22942 = n2412 & n22941 ;
  assign n22943 = n6753 ^ n6479 ^ n3999 ;
  assign n22944 = n8328 ^ n6117 ^ n3459 ;
  assign n22945 = n15031 & n22944 ;
  assign n22946 = n22943 & n22945 ;
  assign n22947 = n15132 ^ n1601 ^ 1'b0 ;
  assign n22948 = n21907 | n22947 ;
  assign n22949 = n22948 ^ n5075 ^ n1352 ;
  assign n22950 = n13364 ^ n3068 ^ 1'b0 ;
  assign n22951 = n10335 & n22950 ;
  assign n22952 = n1323 & n6349 ;
  assign n22953 = ~n7650 & n22952 ;
  assign n22954 = n5355 & ~n5688 ;
  assign n22955 = n22934 ^ n3983 ^ 1'b0 ;
  assign n22956 = n17701 & ~n22955 ;
  assign n22957 = ( n6683 & ~n22954 ) | ( n6683 & n22956 ) | ( ~n22954 & n22956 ) ;
  assign n22959 = n21623 ^ n18089 ^ n3562 ;
  assign n22958 = n9777 ^ n8005 ^ n3479 ;
  assign n22960 = n22959 ^ n22958 ^ n10480 ;
  assign n22970 = n4331 | n11556 ;
  assign n22966 = ( n7980 & n14584 ) | ( n7980 & n15708 ) | ( n14584 & n15708 ) ;
  assign n22967 = n22966 ^ n6627 ^ 1'b0 ;
  assign n22968 = n8618 | n22967 ;
  assign n22969 = n7805 & ~n22968 ;
  assign n22971 = n22970 ^ n22969 ^ 1'b0 ;
  assign n22961 = ~n10681 & n11860 ;
  assign n22962 = n648 & ~n4393 ;
  assign n22963 = n22962 ^ n4029 ^ 1'b0 ;
  assign n22964 = n16427 | n22963 ;
  assign n22965 = n22961 | n22964 ;
  assign n22972 = n22971 ^ n22965 ^ n776 ;
  assign n22973 = n353 & ~n8981 ;
  assign n22974 = n7428 & n22973 ;
  assign n22975 = n22974 ^ n14321 ^ 1'b0 ;
  assign n22976 = ( n7555 & ~n9037 ) | ( n7555 & n22975 ) | ( ~n9037 & n22975 ) ;
  assign n22977 = n19220 ^ n17976 ^ n12651 ;
  assign n22978 = n15799 ^ n7616 ^ 1'b0 ;
  assign n22979 = n2403 ^ x45 ^ 1'b0 ;
  assign n22980 = n855 | n22979 ;
  assign n22981 = n11382 ^ n5592 ^ n3737 ;
  assign n22982 = ( n584 & n22980 ) | ( n584 & ~n22981 ) | ( n22980 & ~n22981 ) ;
  assign n22983 = n22982 ^ n14518 ^ n10235 ;
  assign n22984 = ( ~n3085 & n21350 ) | ( ~n3085 & n22983 ) | ( n21350 & n22983 ) ;
  assign n22985 = n22984 ^ n9161 ^ n1093 ;
  assign n22987 = n10479 ^ n3839 ^ 1'b0 ;
  assign n22986 = ~n476 & n22736 ;
  assign n22988 = n22987 ^ n22986 ^ n5944 ;
  assign n22989 = n11482 & ~n22988 ;
  assign n22990 = ~n12106 & n22989 ;
  assign n22991 = n22990 ^ n11486 ^ 1'b0 ;
  assign n22992 = x34 | n2518 ;
  assign n22993 = n22992 ^ n15175 ^ 1'b0 ;
  assign n22994 = ( ~n5197 & n7031 ) | ( ~n5197 & n8317 ) | ( n7031 & n8317 ) ;
  assign n22995 = n18335 | n22649 ;
  assign n22996 = n22995 ^ n7228 ^ 1'b0 ;
  assign n22997 = n22996 ^ n15469 ^ 1'b0 ;
  assign n22998 = n18420 ^ n8110 ^ 1'b0 ;
  assign n22999 = n4270 | n22998 ;
  assign n23000 = n9449 | n14988 ;
  assign n23001 = n8990 ^ n5982 ^ 1'b0 ;
  assign n23002 = n22959 | n23001 ;
  assign n23003 = n4688 & ~n23002 ;
  assign n23004 = n2374 ^ n1446 ^ 1'b0 ;
  assign n23005 = ( ~n5185 & n18756 ) | ( ~n5185 & n23004 ) | ( n18756 & n23004 ) ;
  assign n23006 = n23005 ^ n4364 ^ 1'b0 ;
  assign n23007 = n18262 & n23006 ;
  assign n23008 = ( n14996 & n15464 ) | ( n14996 & n23007 ) | ( n15464 & n23007 ) ;
  assign n23009 = n16256 | n23008 ;
  assign n23010 = n23003 & ~n23009 ;
  assign n23011 = n23010 ^ n1301 ^ 1'b0 ;
  assign n23012 = n20956 & ~n23011 ;
  assign n23013 = ~n3415 & n7579 ;
  assign n23014 = n19928 ^ n11461 ^ 1'b0 ;
  assign n23015 = n479 & ~n23014 ;
  assign n23016 = n9496 ^ n4279 ^ n2913 ;
  assign n23017 = n1557 & ~n23016 ;
  assign n23018 = n23017 ^ n10238 ^ n9148 ;
  assign n23019 = n23018 ^ n20459 ^ n5671 ;
  assign n23020 = n838 & ~n4626 ;
  assign n23021 = n23020 ^ n6379 ^ 1'b0 ;
  assign n23022 = n7988 ^ n6028 ^ 1'b0 ;
  assign n23023 = n17776 & ~n19814 ;
  assign n23024 = n23022 & n23023 ;
  assign n23025 = ( n15975 & ~n23021 ) | ( n15975 & n23024 ) | ( ~n23021 & n23024 ) ;
  assign n23026 = n5338 & n8551 ;
  assign n23027 = n12599 | n14588 ;
  assign n23040 = n14072 ^ n10800 ^ x116 ;
  assign n23041 = n13742 | n23040 ;
  assign n23042 = n17312 & ~n23041 ;
  assign n23033 = n5503 & n6976 ;
  assign n23034 = n23033 ^ n2444 ^ 1'b0 ;
  assign n23035 = n10049 | n23034 ;
  assign n23036 = n17807 & n23035 ;
  assign n23037 = n12748 & ~n23036 ;
  assign n23038 = n18049 & n23037 ;
  assign n23039 = n23038 ^ n4505 ^ 1'b0 ;
  assign n23028 = n12815 ^ n864 ^ 1'b0 ;
  assign n23029 = n17095 & n23028 ;
  assign n23030 = n23029 ^ n4548 ^ n2217 ;
  assign n23031 = n14031 & n23030 ;
  assign n23032 = n23031 ^ n20627 ^ 1'b0 ;
  assign n23043 = n23042 ^ n23039 ^ n23032 ;
  assign n23044 = n1776 & ~n2000 ;
  assign n23045 = n23044 ^ n23017 ^ 1'b0 ;
  assign n23046 = ( n8659 & ~n12215 ) | ( n8659 & n23045 ) | ( ~n12215 & n23045 ) ;
  assign n23047 = ~n3029 & n23046 ;
  assign n23048 = n18169 & n23047 ;
  assign n23051 = n4882 & ~n9066 ;
  assign n23052 = n23051 ^ n276 ^ 1'b0 ;
  assign n23053 = n23052 ^ n5928 ^ 1'b0 ;
  assign n23049 = n1566 & ~n7350 ;
  assign n23050 = n23049 ^ n8828 ^ 1'b0 ;
  assign n23054 = n23053 ^ n23050 ^ n5901 ;
  assign n23055 = ~n3032 & n16090 ;
  assign n23056 = n21534 ^ n17891 ^ 1'b0 ;
  assign n23057 = n23055 | n23056 ;
  assign n23058 = n23054 | n23057 ;
  assign n23059 = n16237 & ~n23058 ;
  assign n23060 = ( n4186 & n12547 ) | ( n4186 & ~n23059 ) | ( n12547 & ~n23059 ) ;
  assign n23061 = n10490 ^ n1409 ^ 1'b0 ;
  assign n23062 = n20832 & n23061 ;
  assign n23063 = ~n2192 & n12578 ;
  assign n23064 = n23063 ^ n14323 ^ 1'b0 ;
  assign n23065 = n2726 & ~n23064 ;
  assign n23066 = n11669 ^ n384 ^ 1'b0 ;
  assign n23067 = n11339 | n23066 ;
  assign n23068 = n16827 & n23067 ;
  assign n23069 = n19476 ^ n12411 ^ 1'b0 ;
  assign n23070 = n8290 ^ n4618 ^ 1'b0 ;
  assign n23071 = n22236 ^ n3995 ^ 1'b0 ;
  assign n23073 = x157 & n7717 ;
  assign n23072 = ~n4316 & n19280 ;
  assign n23074 = n23073 ^ n23072 ^ n7061 ;
  assign n23076 = ( n2336 & ~n2899 ) | ( n2336 & n7595 ) | ( ~n2899 & n7595 ) ;
  assign n23077 = n3424 | n23076 ;
  assign n23075 = n5815 & n22486 ;
  assign n23078 = n23077 ^ n23075 ^ n14818 ;
  assign n23080 = n9766 ^ n7675 ^ 1'b0 ;
  assign n23081 = n8983 | n23080 ;
  assign n23079 = n14284 | n15913 ;
  assign n23082 = n23081 ^ n23079 ^ 1'b0 ;
  assign n23089 = ( x160 & n4208 ) | ( x160 & ~n4704 ) | ( n4208 & ~n4704 ) ;
  assign n23083 = n2178 | n2377 ;
  assign n23084 = n23083 ^ n4838 ^ 1'b0 ;
  assign n23085 = n12773 ^ n1149 ^ 1'b0 ;
  assign n23086 = n12516 & ~n23085 ;
  assign n23087 = ( ~n12491 & n18555 ) | ( ~n12491 & n23086 ) | ( n18555 & n23086 ) ;
  assign n23088 = n23084 | n23087 ;
  assign n23090 = n23089 ^ n23088 ^ 1'b0 ;
  assign n23091 = n9543 & ~n11209 ;
  assign n23092 = n23091 ^ n3569 ^ n3154 ;
  assign n23093 = n17267 | n23092 ;
  assign n23094 = n19296 ^ n6591 ^ n5490 ;
  assign n23095 = n17381 ^ n16036 ^ n13491 ;
  assign n23096 = ( n9642 & ~n19116 ) | ( n9642 & n23095 ) | ( ~n19116 & n23095 ) ;
  assign n23098 = n2514 | n5971 ;
  assign n23099 = n4469 ^ n2376 ^ 1'b0 ;
  assign n23100 = ~n23098 & n23099 ;
  assign n23097 = ~n12329 & n13456 ;
  assign n23101 = n23100 ^ n23097 ^ 1'b0 ;
  assign n23102 = n13291 & n17823 ;
  assign n23103 = n2878 & n23102 ;
  assign n23104 = n23103 ^ n2573 ^ 1'b0 ;
  assign n23106 = n10995 ^ n6037 ^ 1'b0 ;
  assign n23105 = n9740 ^ n3572 ^ 1'b0 ;
  assign n23107 = n23106 ^ n23105 ^ n21292 ;
  assign n23110 = n376 & n12684 ;
  assign n23108 = n5467 | n9424 ;
  assign n23109 = n23108 ^ n4296 ^ 1'b0 ;
  assign n23111 = n23110 ^ n23109 ^ 1'b0 ;
  assign n23112 = n4980 & ~n23111 ;
  assign n23113 = n2341 & n17423 ;
  assign n23114 = n6531 & n23113 ;
  assign n23115 = n23114 ^ n10252 ^ n8280 ;
  assign n23116 = ( ~n12160 & n19689 ) | ( ~n12160 & n22817 ) | ( n19689 & n22817 ) ;
  assign n23117 = ( n1338 & n23115 ) | ( n1338 & n23116 ) | ( n23115 & n23116 ) ;
  assign n23118 = ( n1136 & ~n1558 ) | ( n1136 & n11041 ) | ( ~n1558 & n11041 ) ;
  assign n23119 = n23118 ^ n13244 ^ 1'b0 ;
  assign n23120 = n8339 & n23119 ;
  assign n23121 = n1502 | n11948 ;
  assign n23122 = n6549 | n9024 ;
  assign n23123 = n23122 ^ n18354 ^ 1'b0 ;
  assign n23124 = n7097 | n10631 ;
  assign n23125 = n7301 & ~n23124 ;
  assign n23126 = n6670 | n23125 ;
  assign n23127 = n23123 | n23126 ;
  assign n23128 = n3977 & ~n15455 ;
  assign n23129 = ~n1223 & n23128 ;
  assign n23130 = n23129 ^ n21984 ^ 1'b0 ;
  assign n23131 = n3759 & ~n22910 ;
  assign n23132 = n23131 ^ n16234 ^ 1'b0 ;
  assign n23133 = ~n14320 & n22829 ;
  assign n23134 = ( n5294 & ~n7693 ) | ( n5294 & n11082 ) | ( ~n7693 & n11082 ) ;
  assign n23136 = n1803 | n7707 ;
  assign n23137 = n5036 & ~n23136 ;
  assign n23135 = ( n5062 & ~n15690 ) | ( n5062 & n21157 ) | ( ~n15690 & n21157 ) ;
  assign n23138 = n23137 ^ n23135 ^ n2440 ;
  assign n23139 = n10647 ^ n8446 ^ n1188 ;
  assign n23143 = n12504 ^ n3467 ^ 1'b0 ;
  assign n23144 = ~n1742 & n23143 ;
  assign n23145 = n4787 & ~n23144 ;
  assign n23140 = ( n3689 & n4090 ) | ( n3689 & n8791 ) | ( n4090 & n8791 ) ;
  assign n23141 = n7342 | n23140 ;
  assign n23142 = n23141 ^ n22014 ^ n4566 ;
  assign n23146 = n23145 ^ n23142 ^ n1953 ;
  assign n23147 = x199 | n9299 ;
  assign n23148 = n551 & ~n5585 ;
  assign n23149 = n23148 ^ n5869 ^ 1'b0 ;
  assign n23150 = n23149 ^ n16292 ^ n8199 ;
  assign n23151 = n8540 ^ n335 ^ 1'b0 ;
  assign n23152 = n19580 | n23151 ;
  assign n23153 = n10202 & n14368 ;
  assign n23154 = n23152 & n23153 ;
  assign n23155 = n2507 & n13677 ;
  assign n23156 = n8490 & n23155 ;
  assign n23157 = ( ~n5091 & n13622 ) | ( ~n5091 & n23156 ) | ( n13622 & n23156 ) ;
  assign n23162 = ~n3283 & n3921 ;
  assign n23163 = n23162 ^ n2135 ^ n1957 ;
  assign n23158 = n2647 & n9286 ;
  assign n23159 = ~n8325 & n23158 ;
  assign n23160 = ~n5910 & n22117 ;
  assign n23161 = n23159 & n23160 ;
  assign n23164 = n23163 ^ n23161 ^ n15913 ;
  assign n23165 = n11995 ^ n6330 ^ 1'b0 ;
  assign n23166 = n5828 | n23165 ;
  assign n23167 = n23166 ^ n17667 ^ n7744 ;
  assign n23168 = n6615 & n23167 ;
  assign n23169 = n23168 ^ n2749 ^ 1'b0 ;
  assign n23170 = ~n4230 & n16379 ;
  assign n23171 = n2391 & ~n23170 ;
  assign n23172 = n23171 ^ n2464 ^ 1'b0 ;
  assign n23173 = n6761 ^ n1959 ^ 1'b0 ;
  assign n23174 = n23173 ^ n3297 ^ 1'b0 ;
  assign n23175 = n929 | n12173 ;
  assign n23176 = n23175 ^ n4603 ^ 1'b0 ;
  assign n23179 = n9765 ^ x54 ^ 1'b0 ;
  assign n23177 = n3605 & n12356 ;
  assign n23178 = n23177 ^ n15728 ^ 1'b0 ;
  assign n23180 = n23179 ^ n23178 ^ n5653 ;
  assign n23181 = n3734 & n5249 ;
  assign n23182 = n4343 & ~n23181 ;
  assign n23183 = n19940 ^ n6031 ^ 1'b0 ;
  assign n23184 = ~n22387 & n23183 ;
  assign n23185 = ~n9311 & n9411 ;
  assign n23186 = n13066 & n23185 ;
  assign n23187 = n23186 ^ n12847 ^ 1'b0 ;
  assign n23188 = n6984 ^ n6502 ^ n5516 ;
  assign n23189 = ~n2100 & n16250 ;
  assign n23190 = ( ~n8727 & n11071 ) | ( ~n8727 & n23189 ) | ( n11071 & n23189 ) ;
  assign n23191 = x26 & ~n11778 ;
  assign n23192 = n23191 ^ n6621 ^ 1'b0 ;
  assign n23193 = n23192 ^ n9663 ^ 1'b0 ;
  assign n23194 = n11086 & ~n23193 ;
  assign n23195 = n9729 & n23194 ;
  assign n23196 = ~x190 & n23195 ;
  assign n23197 = n2712 & n9824 ;
  assign n23198 = ~n17209 & n23197 ;
  assign n23199 = n7300 & ~n11058 ;
  assign n23200 = ~n7052 & n23199 ;
  assign n23201 = n23200 ^ n7465 ^ n3951 ;
  assign n23202 = n3176 | n4875 ;
  assign n23203 = n23202 ^ n12955 ^ 1'b0 ;
  assign n23204 = ( n2832 & ~n10756 ) | ( n2832 & n23203 ) | ( ~n10756 & n23203 ) ;
  assign n23205 = n23204 ^ n19171 ^ n16822 ;
  assign n23206 = n2250 & n11498 ;
  assign n23207 = n10204 ^ n1559 ^ n757 ;
  assign n23208 = n12225 | n23207 ;
  assign n23209 = n4748 | n23208 ;
  assign n23210 = n9177 ^ n2985 ^ n966 ;
  assign n23211 = n6245 & ~n23210 ;
  assign n23212 = n23211 ^ n2569 ^ 1'b0 ;
  assign n23213 = n14129 ^ n6008 ^ 1'b0 ;
  assign n23214 = n23212 | n23213 ;
  assign n23215 = n11898 ^ n8327 ^ n681 ;
  assign n23216 = n23215 ^ n18281 ^ n14105 ;
  assign n23217 = n9936 & ~n19127 ;
  assign n23218 = n17379 ^ n7991 ^ 1'b0 ;
  assign n23219 = n8864 & ~n23218 ;
  assign n23220 = ( n10483 & n23217 ) | ( n10483 & ~n23219 ) | ( n23217 & ~n23219 ) ;
  assign n23221 = n10900 | n23220 ;
  assign n23222 = n14836 ^ n7461 ^ n989 ;
  assign n23223 = n23222 ^ n20350 ^ n297 ;
  assign n23224 = ( ~n1945 & n6408 ) | ( ~n1945 & n17607 ) | ( n6408 & n17607 ) ;
  assign n23225 = n2458 & ~n21573 ;
  assign n23226 = n23225 ^ n17560 ^ 1'b0 ;
  assign n23227 = n23226 ^ n4256 ^ 1'b0 ;
  assign n23228 = n1134 & ~n16937 ;
  assign n23229 = n23228 ^ n1303 ^ 1'b0 ;
  assign n23230 = ( n10994 & n19262 ) | ( n10994 & n22841 ) | ( n19262 & n22841 ) ;
  assign n23231 = ~n3632 & n23230 ;
  assign n23232 = n1473 | n15464 ;
  assign n23233 = n23232 ^ n6081 ^ 1'b0 ;
  assign n23234 = n7408 ^ n6265 ^ 1'b0 ;
  assign n23235 = ( n6548 & n13147 ) | ( n6548 & n23234 ) | ( n13147 & n23234 ) ;
  assign n23236 = n23235 ^ n14984 ^ n350 ;
  assign n23247 = n7952 ^ n5264 ^ 1'b0 ;
  assign n23243 = n12895 ^ n12705 ^ 1'b0 ;
  assign n23244 = ( n6408 & ~n7535 ) | ( n6408 & n23243 ) | ( ~n7535 & n23243 ) ;
  assign n23245 = n23244 ^ n2533 ^ 1'b0 ;
  assign n23246 = x44 & n23245 ;
  assign n23248 = n23247 ^ n23246 ^ 1'b0 ;
  assign n23249 = ~n14117 & n23248 ;
  assign n23237 = n12904 ^ n3261 ^ 1'b0 ;
  assign n23238 = n9438 & ~n23237 ;
  assign n23239 = n8625 ^ n2333 ^ 1'b0 ;
  assign n23240 = n4087 & ~n23239 ;
  assign n23241 = ( n20286 & ~n23238 ) | ( n20286 & n23240 ) | ( ~n23238 & n23240 ) ;
  assign n23242 = n23241 ^ n5602 ^ 1'b0 ;
  assign n23250 = n23249 ^ n23242 ^ n3906 ;
  assign n23251 = n3235 ^ n1851 ^ n647 ;
  assign n23252 = n23251 ^ n21055 ^ n2697 ;
  assign n23254 = n16656 ^ n16654 ^ n11309 ;
  assign n23253 = ~n5657 & n13525 ;
  assign n23255 = n23254 ^ n23253 ^ 1'b0 ;
  assign n23256 = ( x109 & n934 ) | ( x109 & n23255 ) | ( n934 & n23255 ) ;
  assign n23257 = ~n2208 & n11685 ;
  assign n23258 = n3475 ^ n1548 ^ 1'b0 ;
  assign n23259 = n1035 | n10157 ;
  assign n23260 = n23258 | n23259 ;
  assign n23261 = n23260 ^ n9857 ^ x85 ;
  assign n23271 = ( ~n4364 & n7759 ) | ( ~n4364 & n7770 ) | ( n7759 & n7770 ) ;
  assign n23262 = n5210 ^ n1476 ^ 1'b0 ;
  assign n23263 = n1682 & n23262 ;
  assign n23264 = n11826 ^ n1810 ^ 1'b0 ;
  assign n23265 = ( ~n11706 & n23263 ) | ( ~n11706 & n23264 ) | ( n23263 & n23264 ) ;
  assign n23266 = n23265 ^ n22717 ^ n2411 ;
  assign n23267 = n18402 ^ n5848 ^ 1'b0 ;
  assign n23268 = n23267 ^ n20607 ^ 1'b0 ;
  assign n23269 = n23266 | n23268 ;
  assign n23270 = n9311 & ~n23269 ;
  assign n23272 = n23271 ^ n23270 ^ n3735 ;
  assign n23273 = n7817 & ~n13309 ;
  assign n23274 = n23273 ^ n15973 ^ 1'b0 ;
  assign n23275 = n23274 ^ n10733 ^ n4266 ;
  assign n23276 = n12976 & n19724 ;
  assign n23277 = n7888 & ~n23276 ;
  assign n23278 = n23277 ^ n15817 ^ n3556 ;
  assign n23279 = n4260 & ~n9620 ;
  assign n23280 = n10738 ^ n1685 ^ 1'b0 ;
  assign n23281 = ~n4215 & n23280 ;
  assign n23282 = n23279 & n23281 ;
  assign n23283 = n13190 ^ n7907 ^ 1'b0 ;
  assign n23284 = n23283 ^ n20606 ^ 1'b0 ;
  assign n23285 = n9109 ^ n6160 ^ n831 ;
  assign n23286 = n23285 ^ n16270 ^ n384 ;
  assign n23287 = n23286 ^ n19592 ^ 1'b0 ;
  assign n23288 = n2436 | n8332 ;
  assign n23289 = n15330 | n23288 ;
  assign n23290 = ( n4432 & n9100 ) | ( n4432 & ~n23289 ) | ( n9100 & ~n23289 ) ;
  assign n23291 = n13989 ^ n2665 ^ 1'b0 ;
  assign n23292 = n23291 ^ n17934 ^ 1'b0 ;
  assign n23293 = ~n6695 & n23292 ;
  assign n23294 = ~n9959 & n19709 ;
  assign n23295 = ~n7476 & n23294 ;
  assign n23296 = n13798 ^ n4989 ^ n4446 ;
  assign n23297 = n23296 ^ n16780 ^ 1'b0 ;
  assign n23298 = ~n647 & n13795 ;
  assign n23299 = n23298 ^ n8709 ^ 1'b0 ;
  assign n23300 = n3903 ^ n1655 ^ 1'b0 ;
  assign n23301 = ~n11916 & n23300 ;
  assign n23302 = n7651 & ~n23301 ;
  assign n23303 = n23302 ^ n22134 ^ n9756 ;
  assign n23304 = n4156 & n18156 ;
  assign n23305 = ~n414 & n23304 ;
  assign n23306 = n23305 ^ n21576 ^ 1'b0 ;
  assign n23307 = n2386 & ~n18481 ;
  assign n23308 = n23307 ^ n11439 ^ 1'b0 ;
  assign n23309 = n1173 & ~n14134 ;
  assign n23310 = ( n4982 & n19402 ) | ( n4982 & n23309 ) | ( n19402 & n23309 ) ;
  assign n23311 = ( ~n3855 & n8504 ) | ( ~n3855 & n18331 ) | ( n8504 & n18331 ) ;
  assign n23312 = n18164 & n23311 ;
  assign n23315 = n21466 ^ n15829 ^ 1'b0 ;
  assign n23316 = n421 | n23315 ;
  assign n23317 = n7173 & ~n23316 ;
  assign n23318 = n23317 ^ n20331 ^ 1'b0 ;
  assign n23319 = ( n5210 & n22765 ) | ( n5210 & n23318 ) | ( n22765 & n23318 ) ;
  assign n23313 = ( n3821 & n19201 ) | ( n3821 & ~n21419 ) | ( n19201 & ~n21419 ) ;
  assign n23314 = ( n15595 & ~n16268 ) | ( n15595 & n23313 ) | ( ~n16268 & n23313 ) ;
  assign n23320 = n23319 ^ n23314 ^ 1'b0 ;
  assign n23321 = n1056 & n14449 ;
  assign n23322 = n10202 & n23321 ;
  assign n23323 = n23322 ^ n3218 ^ 1'b0 ;
  assign n23324 = ~n1730 & n13655 ;
  assign n23325 = n23324 ^ n14491 ^ n10581 ;
  assign n23326 = ~n2241 & n4797 ;
  assign n23327 = n11963 & n23326 ;
  assign n23328 = n23327 ^ n19193 ^ 1'b0 ;
  assign n23329 = n11961 ^ n9517 ^ 1'b0 ;
  assign n23330 = n9886 | n23329 ;
  assign n23331 = x176 & n10527 ;
  assign n23332 = ( n5454 & ~n5576 ) | ( n5454 & n20658 ) | ( ~n5576 & n20658 ) ;
  assign n23333 = n23332 ^ n20528 ^ x163 ;
  assign n23334 = n23331 | n23333 ;
  assign n23335 = n7662 & ~n9642 ;
  assign n23336 = x7 & n4034 ;
  assign n23337 = n3170 & n23336 ;
  assign n23338 = n23335 & n23337 ;
  assign n23339 = n3630 | n14382 ;
  assign n23340 = n23339 ^ n17615 ^ 1'b0 ;
  assign n23341 = ~n20424 & n22515 ;
  assign n23342 = n23341 ^ n9174 ^ 1'b0 ;
  assign n23343 = ~n13743 & n19311 ;
  assign n23344 = n17188 ^ n13792 ^ n9374 ;
  assign n23345 = ~n10985 & n23344 ;
  assign n23346 = n14192 & n23345 ;
  assign n23347 = n23343 | n23346 ;
  assign n23348 = n2369 | n8469 ;
  assign n23349 = ( n4230 & ~n21455 ) | ( n4230 & n21890 ) | ( ~n21455 & n21890 ) ;
  assign n23350 = n3289 & ~n23349 ;
  assign n23351 = ~n23348 & n23350 ;
  assign n23352 = ~n284 & n8727 ;
  assign n23353 = ~n2677 & n5804 ;
  assign n23354 = ~n11924 & n23353 ;
  assign n23355 = ~n23352 & n23354 ;
  assign n23357 = x183 & ~n10334 ;
  assign n23358 = n11132 & n23357 ;
  assign n23359 = n16778 | n23358 ;
  assign n23360 = n4644 | n23359 ;
  assign n23356 = ~n13813 & n20634 ;
  assign n23361 = n23360 ^ n23356 ^ 1'b0 ;
  assign n23362 = n3589 ^ n2773 ^ 1'b0 ;
  assign n23363 = n10754 | n23362 ;
  assign n23364 = n23363 ^ n17578 ^ n11027 ;
  assign n23365 = n20334 ^ n10478 ^ n3077 ;
  assign n23366 = n23365 ^ n3171 ^ 1'b0 ;
  assign n23367 = n8539 ^ n5629 ^ 1'b0 ;
  assign n23368 = n23366 | n23367 ;
  assign n23370 = n4893 | n5448 ;
  assign n23371 = n21177 | n23370 ;
  assign n23372 = ( n939 & n9486 ) | ( n939 & ~n23371 ) | ( n9486 & ~n23371 ) ;
  assign n23369 = n872 & n7925 ;
  assign n23373 = n23372 ^ n23369 ^ 1'b0 ;
  assign n23374 = n3138 & ~n20144 ;
  assign n23375 = n3375 & n10225 ;
  assign n23376 = ( n5040 & n6690 ) | ( n5040 & n23375 ) | ( n6690 & n23375 ) ;
  assign n23377 = ~n5360 & n23376 ;
  assign n23378 = ( ~n3362 & n7051 ) | ( ~n3362 & n15104 ) | ( n7051 & n15104 ) ;
  assign n23379 = n23378 ^ n11041 ^ n4826 ;
  assign n23380 = ~n8860 & n9205 ;
  assign n23381 = n9420 & n23380 ;
  assign n23382 = n4921 | n5675 ;
  assign n23383 = n1037 | n23382 ;
  assign n23384 = n23383 ^ n8226 ^ 1'b0 ;
  assign n23385 = n3798 & n23384 ;
  assign n23386 = n16964 ^ n6646 ^ n4316 ;
  assign n23387 = n23386 ^ n14889 ^ n3425 ;
  assign n23388 = n23387 ^ n290 ^ 1'b0 ;
  assign n23389 = n13293 & ~n19505 ;
  assign n23390 = ~n14298 & n23389 ;
  assign n23391 = n12507 ^ n5724 ^ 1'b0 ;
  assign n23392 = n4776 & n20271 ;
  assign n23393 = n23392 ^ n1225 ^ 1'b0 ;
  assign n23394 = n22873 ^ n4251 ^ 1'b0 ;
  assign n23395 = n19290 ^ n17744 ^ n851 ;
  assign n23403 = ~n939 & n22301 ;
  assign n23400 = n7717 ^ n5238 ^ 1'b0 ;
  assign n23401 = n18838 & ~n23400 ;
  assign n23396 = ~n3658 & n11370 ;
  assign n23397 = n23396 ^ n5688 ^ 1'b0 ;
  assign n23398 = n23397 ^ n14866 ^ n12389 ;
  assign n23399 = ( n4234 & ~n18210 ) | ( n4234 & n23398 ) | ( ~n18210 & n23398 ) ;
  assign n23402 = n23401 ^ n23399 ^ n14281 ;
  assign n23404 = n23403 ^ n23402 ^ 1'b0 ;
  assign n23405 = n22732 ^ n11337 ^ 1'b0 ;
  assign n23406 = n10719 ^ n5573 ^ n2474 ;
  assign n23407 = n3957 & n23406 ;
  assign n23408 = n23407 ^ n1342 ^ 1'b0 ;
  assign n23409 = n11129 ^ n5907 ^ 1'b0 ;
  assign n23410 = n23409 ^ n23397 ^ n12147 ;
  assign n23411 = ( n16803 & ~n23408 ) | ( n16803 & n23410 ) | ( ~n23408 & n23410 ) ;
  assign n23412 = n4355 | n14647 ;
  assign n23413 = n22178 ^ n20817 ^ 1'b0 ;
  assign n23414 = ~n10932 & n19450 ;
  assign n23415 = n8751 ^ n842 ^ 1'b0 ;
  assign n23416 = x167 & ~n23415 ;
  assign n23417 = n15994 ^ n10519 ^ n4504 ;
  assign n23418 = n1263 & ~n5091 ;
  assign n23419 = ~n23417 & n23418 ;
  assign n23420 = n23416 | n23419 ;
  assign n23421 = n15134 ^ n6806 ^ n5642 ;
  assign n23422 = ~n5740 & n23421 ;
  assign n23423 = n18753 ^ n9840 ^ 1'b0 ;
  assign n23424 = n7395 ^ n6330 ^ 1'b0 ;
  assign n23425 = ~n23423 & n23424 ;
  assign n23426 = ( n10521 & ~n12823 ) | ( n10521 & n23425 ) | ( ~n12823 & n23425 ) ;
  assign n23427 = n18770 ^ n6120 ^ 1'b0 ;
  assign n23428 = n23427 ^ n13294 ^ 1'b0 ;
  assign n23429 = n23426 & ~n23428 ;
  assign n23430 = n6639 & n11106 ;
  assign n23431 = n2466 & n3517 ;
  assign n23432 = ~n3123 & n23431 ;
  assign n23433 = n6580 | n23432 ;
  assign n23434 = n23430 | n23433 ;
  assign n23435 = n12607 & n23434 ;
  assign n23436 = n23435 ^ n13223 ^ 1'b0 ;
  assign n23437 = n10712 ^ n9900 ^ n7160 ;
  assign n23438 = ~n14624 & n23437 ;
  assign n23439 = ~n6091 & n23438 ;
  assign n23440 = n23439 ^ n13056 ^ 1'b0 ;
  assign n23441 = n18380 ^ n12459 ^ n1750 ;
  assign n23442 = ~n3858 & n6331 ;
  assign n23443 = n13541 & ~n17590 ;
  assign n23444 = n15677 ^ n12123 ^ 1'b0 ;
  assign n23445 = n23444 ^ x4 ^ 1'b0 ;
  assign n23446 = n1105 & ~n2861 ;
  assign n23447 = ~n10661 & n23446 ;
  assign n23448 = n3049 ^ n1542 ^ x129 ;
  assign n23449 = n10596 | n23448 ;
  assign n23450 = n14675 ^ n4340 ^ 1'b0 ;
  assign n23451 = x70 & ~n23450 ;
  assign n23452 = ~n23449 & n23451 ;
  assign n23453 = n2877 ^ n1796 ^ 1'b0 ;
  assign n23454 = n2654 | n23453 ;
  assign n23455 = n17383 ^ n16314 ^ n2283 ;
  assign n23456 = n1971 | n23455 ;
  assign n23458 = n3589 ^ n2225 ^ n2013 ;
  assign n23457 = ( n9988 & n14792 ) | ( n9988 & ~n15996 ) | ( n14792 & ~n15996 ) ;
  assign n23459 = n23458 ^ n23457 ^ n4744 ;
  assign n23460 = ( n825 & n23456 ) | ( n825 & n23459 ) | ( n23456 & n23459 ) ;
  assign n23461 = n23454 | n23460 ;
  assign n23462 = n23461 ^ n18767 ^ 1'b0 ;
  assign n23463 = n8740 ^ n1064 ^ 1'b0 ;
  assign n23464 = ~n6596 & n10261 ;
  assign n23465 = ~n269 & n23464 ;
  assign n23466 = n2041 & ~n23465 ;
  assign n23468 = n13122 ^ n6914 ^ 1'b0 ;
  assign n23469 = n6388 | n23468 ;
  assign n23470 = n23469 ^ n7012 ^ n3690 ;
  assign n23467 = n17224 ^ n15798 ^ n2156 ;
  assign n23471 = n23470 ^ n23467 ^ n16028 ;
  assign n23472 = n21373 ^ n7183 ^ 1'b0 ;
  assign n23473 = n23472 ^ n21476 ^ 1'b0 ;
  assign n23474 = n4264 & ~n23473 ;
  assign n23475 = n1053 | n2777 ;
  assign n23476 = ( n6552 & n11156 ) | ( n6552 & n23475 ) | ( n11156 & n23475 ) ;
  assign n23477 = n23476 ^ n4286 ^ 1'b0 ;
  assign n23478 = ( n1390 & n17903 ) | ( n1390 & n23477 ) | ( n17903 & n23477 ) ;
  assign n23479 = n13317 & ~n23478 ;
  assign n23480 = ~n23474 & n23479 ;
  assign n23481 = ( ~x249 & n6045 ) | ( ~x249 & n23480 ) | ( n6045 & n23480 ) ;
  assign n23482 = n8429 ^ n2607 ^ n516 ;
  assign n23483 = n11767 ^ n5281 ^ n512 ;
  assign n23484 = n23483 ^ n3110 ^ n2764 ;
  assign n23485 = n23484 ^ n19105 ^ 1'b0 ;
  assign n23486 = n23482 & n23485 ;
  assign n23487 = n23486 ^ n23063 ^ 1'b0 ;
  assign n23488 = ~n3177 & n23487 ;
  assign n23489 = n13675 ^ n12635 ^ n1209 ;
  assign n23490 = n12801 & ~n15351 ;
  assign n23491 = n23489 | n23490 ;
  assign n23492 = n21322 ^ n10707 ^ n4469 ;
  assign n23493 = ( n1766 & ~n2201 ) | ( n1766 & n4809 ) | ( ~n2201 & n4809 ) ;
  assign n23494 = n6030 & ~n9529 ;
  assign n23495 = n12167 | n23494 ;
  assign n23496 = n23495 ^ n16478 ^ 1'b0 ;
  assign n23497 = ( x154 & n23493 ) | ( x154 & n23496 ) | ( n23493 & n23496 ) ;
  assign n23498 = n20326 ^ n5042 ^ n2786 ;
  assign n23499 = n23498 ^ n21951 ^ n16181 ;
  assign n23500 = n21649 & n21775 ;
  assign n23501 = n19476 & n23500 ;
  assign n23502 = n23501 ^ n1462 ^ 1'b0 ;
  assign n23503 = n13459 | n23502 ;
  assign n23504 = n10004 ^ n502 ^ 1'b0 ;
  assign n23505 = n9747 & ~n23504 ;
  assign n23506 = n7505 | n23505 ;
  assign n23507 = ( n684 & ~n7519 ) | ( n684 & n23506 ) | ( ~n7519 & n23506 ) ;
  assign n23508 = n16958 ^ n1877 ^ 1'b0 ;
  assign n23509 = ( n1709 & n9125 ) | ( n1709 & n19976 ) | ( n9125 & n19976 ) ;
  assign n23510 = ( n2325 & n4842 ) | ( n2325 & ~n20182 ) | ( n4842 & ~n20182 ) ;
  assign n23511 = ~n5205 & n21350 ;
  assign n23512 = n23511 ^ n19951 ^ 1'b0 ;
  assign n23513 = ~n23510 & n23512 ;
  assign n23514 = n23513 ^ n6360 ^ 1'b0 ;
  assign n23515 = n6030 & n9904 ;
  assign n23516 = n12455 | n23515 ;
  assign n23517 = n923 & ~n22734 ;
  assign n23518 = n23517 ^ n2642 ^ 1'b0 ;
  assign n23519 = ( ~n732 & n6887 ) | ( ~n732 & n14657 ) | ( n6887 & n14657 ) ;
  assign n23520 = ( n9339 & n23518 ) | ( n9339 & n23519 ) | ( n23518 & n23519 ) ;
  assign n23522 = ( n1488 & n9026 ) | ( n1488 & ~n16429 ) | ( n9026 & ~n16429 ) ;
  assign n23521 = ~n5675 & n7792 ;
  assign n23523 = n23522 ^ n23521 ^ n5418 ;
  assign n23524 = n23523 ^ n18339 ^ n14424 ;
  assign n23525 = ( ~n5945 & n13927 ) | ( ~n5945 & n23524 ) | ( n13927 & n23524 ) ;
  assign n23528 = ( n804 & n6643 ) | ( n804 & ~n15347 ) | ( n6643 & ~n15347 ) ;
  assign n23526 = ( n6488 & n15234 ) | ( n6488 & n17111 ) | ( n15234 & n17111 ) ;
  assign n23527 = n23526 ^ n9484 ^ n8098 ;
  assign n23529 = n23528 ^ n23527 ^ 1'b0 ;
  assign n23530 = n3655 | n23529 ;
  assign n23532 = n6866 ^ n4142 ^ n1585 ;
  assign n23533 = ( n2646 & n3556 ) | ( n2646 & n23532 ) | ( n3556 & n23532 ) ;
  assign n23531 = n1986 & n13479 ;
  assign n23534 = n23533 ^ n23531 ^ 1'b0 ;
  assign n23535 = n1623 & n15409 ;
  assign n23536 = ~n18233 & n23535 ;
  assign n23537 = ( n1216 & ~n1887 ) | ( n1216 & n6136 ) | ( ~n1887 & n6136 ) ;
  assign n23538 = n4601 & ~n23537 ;
  assign n23539 = n23538 ^ n16524 ^ n11974 ;
  assign n23540 = n20651 ^ n18232 ^ 1'b0 ;
  assign n23541 = n3268 & n14653 ;
  assign n23544 = n15682 ^ n9322 ^ n870 ;
  assign n23542 = ~n2657 & n12470 ;
  assign n23543 = n18265 & n23542 ;
  assign n23545 = n23544 ^ n23543 ^ 1'b0 ;
  assign n23546 = n20548 | n23545 ;
  assign n23547 = n19651 ^ n15194 ^ 1'b0 ;
  assign n23548 = ~n262 & n23547 ;
  assign n23549 = n14034 ^ n9567 ^ n8418 ;
  assign n23550 = ( n1643 & n4952 ) | ( n1643 & n10156 ) | ( n4952 & n10156 ) ;
  assign n23551 = ( n6771 & n23549 ) | ( n6771 & n23550 ) | ( n23549 & n23550 ) ;
  assign n23552 = ( n1475 & n16439 ) | ( n1475 & n22560 ) | ( n16439 & n22560 ) ;
  assign n23553 = ( n4898 & n23551 ) | ( n4898 & ~n23552 ) | ( n23551 & ~n23552 ) ;
  assign n23554 = n23270 ^ n12335 ^ n7890 ;
  assign n23555 = ~n1363 & n1915 ;
  assign n23556 = ~n1915 & n23555 ;
  assign n23557 = n21431 ^ n11623 ^ 1'b0 ;
  assign n23558 = n8739 & ~n23557 ;
  assign n23559 = ~n17068 & n23558 ;
  assign n23560 = n23556 & n23559 ;
  assign n23562 = n838 | n12310 ;
  assign n23561 = n17866 ^ n9083 ^ n1261 ;
  assign n23563 = n23562 ^ n23561 ^ n6507 ;
  assign n23564 = n1548 & ~n2662 ;
  assign n23565 = n23564 ^ n9631 ^ 1'b0 ;
  assign n23566 = n23480 & n23565 ;
  assign n23567 = n19927 ^ n6168 ^ 1'b0 ;
  assign n23568 = n6088 | n8861 ;
  assign n23569 = n2754 & ~n23568 ;
  assign n23570 = n15166 & ~n23569 ;
  assign n23571 = n23570 ^ n4364 ^ 1'b0 ;
  assign n23572 = n17466 ^ n12724 ^ n2422 ;
  assign n23575 = ( n4093 & ~n4655 ) | ( n4093 & n16350 ) | ( ~n4655 & n16350 ) ;
  assign n23574 = n8838 ^ n8624 ^ n3250 ;
  assign n23573 = n17631 ^ n15450 ^ n6339 ;
  assign n23576 = n23575 ^ n23574 ^ n23573 ;
  assign n23577 = ( n9518 & ~n17048 ) | ( n9518 & n23576 ) | ( ~n17048 & n23576 ) ;
  assign n23579 = n1252 & n13385 ;
  assign n23580 = n23579 ^ n22034 ^ n13164 ;
  assign n23581 = ( n3415 & ~n5356 ) | ( n3415 & n23580 ) | ( ~n5356 & n23580 ) ;
  assign n23578 = n5035 & n17695 ;
  assign n23582 = n23581 ^ n23578 ^ 1'b0 ;
  assign n23583 = n10523 & ~n23582 ;
  assign n23584 = ( n10926 & n23577 ) | ( n10926 & n23583 ) | ( n23577 & n23583 ) ;
  assign n23585 = n7798 & ~n10146 ;
  assign n23587 = n4388 & n21051 ;
  assign n23586 = x10 | n1226 ;
  assign n23588 = n23587 ^ n23586 ^ 1'b0 ;
  assign n23589 = n19627 ^ n18855 ^ 1'b0 ;
  assign n23592 = ~n262 & n13447 ;
  assign n23590 = n10069 & ~n19810 ;
  assign n23591 = n23590 ^ n17352 ^ n15104 ;
  assign n23593 = n23592 ^ n23591 ^ 1'b0 ;
  assign n23594 = n23589 | n23593 ;
  assign n23595 = n13065 & ~n23594 ;
  assign n23596 = n20321 ^ n4796 ^ 1'b0 ;
  assign n23597 = n9700 ^ n462 ^ 1'b0 ;
  assign n23598 = ~n10283 & n23597 ;
  assign n23599 = x189 & n23598 ;
  assign n23600 = n23596 & n23599 ;
  assign n23601 = n6723 ^ n5353 ^ 1'b0 ;
  assign n23602 = n9835 | n11486 ;
  assign n23603 = n12033 & ~n23602 ;
  assign n23604 = ~n1738 & n14021 ;
  assign n23605 = n10936 & n23604 ;
  assign n23606 = n15372 | n23605 ;
  assign n23607 = n9107 & ~n23606 ;
  assign n23608 = n2649 & ~n8868 ;
  assign n23609 = n15670 & ~n23608 ;
  assign n23610 = n23609 ^ n1919 ^ 1'b0 ;
  assign n23611 = n23610 ^ n20606 ^ 1'b0 ;
  assign n23612 = ( n17776 & n23607 ) | ( n17776 & n23611 ) | ( n23607 & n23611 ) ;
  assign n23613 = n23612 ^ n20332 ^ n7414 ;
  assign n23614 = n6780 ^ n4830 ^ 1'b0 ;
  assign n23615 = ( ~n13741 & n21056 ) | ( ~n13741 & n23614 ) | ( n21056 & n23614 ) ;
  assign n23616 = n15925 & ~n20512 ;
  assign n23617 = n23616 ^ n11088 ^ 1'b0 ;
  assign n23618 = ( ~n1132 & n1159 ) | ( ~n1132 & n2457 ) | ( n1159 & n2457 ) ;
  assign n23619 = n16842 ^ n4875 ^ 1'b0 ;
  assign n23620 = ( x253 & n23618 ) | ( x253 & ~n23619 ) | ( n23618 & ~n23619 ) ;
  assign n23621 = n11899 | n23620 ;
  assign n23622 = n4187 & ~n17522 ;
  assign n23623 = n2389 & n23622 ;
  assign n23624 = n23623 ^ x182 ^ 1'b0 ;
  assign n23625 = ~n5120 & n19107 ;
  assign n23626 = ~n8506 & n23625 ;
  assign n23627 = n23626 ^ n12509 ^ n7596 ;
  assign n23628 = n23627 ^ n10211 ^ 1'b0 ;
  assign n23629 = n6809 | n23628 ;
  assign n23630 = n23629 ^ n2578 ^ 1'b0 ;
  assign n23631 = n4881 & ~n22001 ;
  assign n23632 = n23631 ^ n6692 ^ 1'b0 ;
  assign n23633 = n669 | n3650 ;
  assign n23634 = n23632 | n23633 ;
  assign n23635 = n6402 & n9726 ;
  assign n23636 = n23635 ^ n13967 ^ 1'b0 ;
  assign n23637 = ( x223 & ~n10300 ) | ( x223 & n16198 ) | ( ~n10300 & n16198 ) ;
  assign n23638 = ~n15178 & n23637 ;
  assign n23639 = ~n23636 & n23638 ;
  assign n23642 = ( n276 & n6164 ) | ( n276 & ~n19583 ) | ( n6164 & ~n19583 ) ;
  assign n23640 = n20191 ^ n20141 ^ 1'b0 ;
  assign n23641 = ~n14970 & n23640 ;
  assign n23643 = n23642 ^ n23641 ^ 1'b0 ;
  assign n23645 = n1827 | n6369 ;
  assign n23646 = ( x248 & n15377 ) | ( x248 & ~n23645 ) | ( n15377 & ~n23645 ) ;
  assign n23644 = ~n14483 & n20629 ;
  assign n23647 = n23646 ^ n23644 ^ n19263 ;
  assign n23648 = n22687 ^ n3402 ^ 1'b0 ;
  assign n23649 = ( ~n5657 & n10773 ) | ( ~n5657 & n23648 ) | ( n10773 & n23648 ) ;
  assign n23651 = n8001 & ~n15180 ;
  assign n23652 = n23651 ^ n9518 ^ 1'b0 ;
  assign n23650 = n3126 & ~n22169 ;
  assign n23653 = n23652 ^ n23650 ^ 1'b0 ;
  assign n23654 = ~n5453 & n7323 ;
  assign n23655 = n22160 & n23654 ;
  assign n23656 = ( n6712 & n10301 ) | ( n6712 & n23655 ) | ( n10301 & n23655 ) ;
  assign n23657 = n1934 & n12819 ;
  assign n23659 = n15348 ^ n5057 ^ n4801 ;
  assign n23660 = n23659 ^ n15926 ^ 1'b0 ;
  assign n23658 = x70 & ~n2061 ;
  assign n23661 = n23660 ^ n23658 ^ n17205 ;
  assign n23662 = n5802 | n20112 ;
  assign n23663 = n23662 ^ n5116 ^ 1'b0 ;
  assign n23664 = ( ~n12159 & n16657 ) | ( ~n12159 & n20234 ) | ( n16657 & n20234 ) ;
  assign n23665 = n23664 ^ n5092 ^ n491 ;
  assign n23666 = ~n820 & n2164 ;
  assign n23667 = n18657 & n23666 ;
  assign n23670 = ( n336 & n10714 ) | ( n336 & ~n13740 ) | ( n10714 & ~n13740 ) ;
  assign n23668 = n19308 ^ n16737 ^ n2458 ;
  assign n23669 = n23668 ^ n13471 ^ n8047 ;
  assign n23671 = n23670 ^ n23669 ^ n3138 ;
  assign n23672 = ~n23667 & n23671 ;
  assign n23673 = n5132 & n23672 ;
  assign n23674 = n16640 ^ n6296 ^ 1'b0 ;
  assign n23675 = ~n15559 & n23674 ;
  assign n23676 = n17651 & n23675 ;
  assign n23677 = n18268 ^ n5500 ^ n3120 ;
  assign n23678 = n1735 & ~n23677 ;
  assign n23679 = ~n22182 & n23678 ;
  assign n23680 = n23676 | n23679 ;
  assign n23681 = n23408 | n23680 ;
  assign n23682 = n11743 ^ n9779 ^ 1'b0 ;
  assign n23683 = n13011 ^ n6615 ^ 1'b0 ;
  assign n23684 = n10393 ^ n9603 ^ n2314 ;
  assign n23687 = ( ~n1725 & n3982 ) | ( ~n1725 & n8091 ) | ( n3982 & n8091 ) ;
  assign n23685 = n4542 ^ n1312 ^ 1'b0 ;
  assign n23686 = n19592 & n23685 ;
  assign n23688 = n23687 ^ n23686 ^ 1'b0 ;
  assign n23689 = n23684 | n23688 ;
  assign n23690 = n20483 & ~n23689 ;
  assign n23691 = ~n15973 & n23690 ;
  assign n23692 = n6160 ^ n5117 ^ 1'b0 ;
  assign n23697 = n1958 & ~n10559 ;
  assign n23694 = ~n7815 & n13628 ;
  assign n23695 = n23694 ^ n9904 ^ 1'b0 ;
  assign n23693 = n1474 | n4338 ;
  assign n23696 = n23695 ^ n23693 ^ 1'b0 ;
  assign n23698 = n23697 ^ n23696 ^ n436 ;
  assign n23701 = n7360 & n10561 ;
  assign n23699 = n5775 & n11659 ;
  assign n23700 = ~n8512 & n23699 ;
  assign n23702 = n23701 ^ n23700 ^ 1'b0 ;
  assign n23703 = n2646 ^ n1127 ^ n1029 ;
  assign n23704 = n7797 & ~n23703 ;
  assign n23705 = n6589 & ~n13328 ;
  assign n23706 = n23704 & n23705 ;
  assign n23709 = n16751 ^ n16363 ^ n10671 ;
  assign n23707 = n9938 | n23590 ;
  assign n23708 = n373 & ~n23707 ;
  assign n23710 = n23709 ^ n23708 ^ 1'b0 ;
  assign n23711 = n21642 ^ n9801 ^ n9239 ;
  assign n23712 = n23711 ^ n20876 ^ n12033 ;
  assign n23713 = n14673 ^ n8494 ^ n7415 ;
  assign n23714 = n7361 & n20235 ;
  assign n23715 = n7522 & n23714 ;
  assign n23716 = n16509 ^ n13007 ^ 1'b0 ;
  assign n23717 = n23716 ^ n11283 ^ n8730 ;
  assign n23718 = n13289 | n18631 ;
  assign n23719 = n22372 | n23718 ;
  assign n23720 = n17720 ^ n12750 ^ n4137 ;
  assign n23721 = n22468 ^ n3257 ^ 1'b0 ;
  assign n23722 = n7215 ^ n3435 ^ x231 ;
  assign n23723 = n15315 | n23722 ;
  assign n23724 = ( ~n3436 & n12952 ) | ( ~n3436 & n14027 ) | ( n12952 & n14027 ) ;
  assign n23725 = n4918 & ~n23724 ;
  assign n23726 = ~n4256 & n23725 ;
  assign n23727 = n14651 & ~n14680 ;
  assign n23728 = ( n5720 & n8278 ) | ( n5720 & n15193 ) | ( n8278 & n15193 ) ;
  assign n23729 = n22847 & n23728 ;
  assign n23730 = n5366 ^ n1632 ^ n506 ;
  assign n23731 = n12472 ^ n4850 ^ 1'b0 ;
  assign n23732 = ( ~n5637 & n13492 ) | ( ~n5637 & n23731 ) | ( n13492 & n23731 ) ;
  assign n23733 = n20017 ^ n12162 ^ 1'b0 ;
  assign n23734 = ( n17913 & n19120 ) | ( n17913 & ~n23733 ) | ( n19120 & ~n23733 ) ;
  assign n23739 = n8537 ^ x89 ^ 1'b0 ;
  assign n23740 = n23739 ^ n17434 ^ n1917 ;
  assign n23735 = n2949 | n7424 ;
  assign n23736 = n23735 ^ n5122 ^ 1'b0 ;
  assign n23737 = n23736 ^ x116 ^ 1'b0 ;
  assign n23738 = ~n10050 & n23737 ;
  assign n23741 = n23740 ^ n23738 ^ 1'b0 ;
  assign n23742 = ( n10785 & n20346 ) | ( n10785 & ~n23741 ) | ( n20346 & ~n23741 ) ;
  assign n23743 = n21512 ^ n5884 ^ 1'b0 ;
  assign n23748 = ~n2388 & n8724 ;
  assign n23749 = n23748 ^ n15078 ^ 1'b0 ;
  assign n23744 = n2919 & ~n20850 ;
  assign n23745 = n6572 & ~n9755 ;
  assign n23746 = n318 | n23745 ;
  assign n23747 = n23744 & ~n23746 ;
  assign n23750 = n23749 ^ n23747 ^ n1713 ;
  assign n23751 = n17666 & ~n23750 ;
  assign n23752 = ~n12719 & n23751 ;
  assign n23753 = ( ~n15326 & n19942 ) | ( ~n15326 & n22035 ) | ( n19942 & n22035 ) ;
  assign n23754 = n6353 ^ n3957 ^ 1'b0 ;
  assign n23755 = n23754 ^ n16412 ^ n4502 ;
  assign n23756 = n1522 & n3679 ;
  assign n23757 = n3384 ^ n2710 ^ 1'b0 ;
  assign n23758 = n21883 ^ n262 ^ 1'b0 ;
  assign n23759 = n17524 ^ n16831 ^ n11597 ;
  assign n23761 = n23448 ^ n2621 ^ n553 ;
  assign n23760 = n4051 ^ n868 ^ 1'b0 ;
  assign n23762 = n23761 ^ n23760 ^ n13718 ;
  assign n23763 = n23759 & ~n23762 ;
  assign n23764 = ~n23758 & n23763 ;
  assign n23765 = n4321 & ~n22514 ;
  assign n23766 = n7115 | n10252 ;
  assign n23767 = n23766 ^ n6331 ^ 1'b0 ;
  assign n23768 = ( ~n2905 & n14007 ) | ( ~n2905 & n23767 ) | ( n14007 & n23767 ) ;
  assign n23769 = n19813 ^ n10371 ^ 1'b0 ;
  assign n23770 = n23769 ^ n16049 ^ n9674 ;
  assign n23771 = ( n680 & ~n2274 ) | ( n680 & n11990 ) | ( ~n2274 & n11990 ) ;
  assign n23772 = n12283 | n23771 ;
  assign n23773 = n23772 ^ n6999 ^ n2530 ;
  assign n23774 = n9997 ^ n3121 ^ 1'b0 ;
  assign n23775 = n23774 ^ n12199 ^ n9180 ;
  assign n23776 = ~n2240 & n9892 ;
  assign n23777 = n23776 ^ n4453 ^ 1'b0 ;
  assign n23778 = n23777 ^ n19884 ^ 1'b0 ;
  assign n23779 = n22063 & ~n23778 ;
  assign n23780 = ~n17358 & n22473 ;
  assign n23781 = n4553 | n6411 ;
  assign n23782 = n8551 | n23781 ;
  assign n23783 = n23782 ^ n7823 ^ n4054 ;
  assign n23784 = n23783 ^ n7388 ^ 1'b0 ;
  assign n23785 = ( ~n23042 & n23780 ) | ( ~n23042 & n23784 ) | ( n23780 & n23784 ) ;
  assign n23786 = n17417 ^ n11490 ^ n1721 ;
  assign n23787 = n15649 ^ n10670 ^ n9804 ;
  assign n23788 = n8663 ^ n5302 ^ 1'b0 ;
  assign n23789 = ~n1857 & n13354 ;
  assign n23790 = n23789 ^ n2050 ^ 1'b0 ;
  assign n23791 = n23790 ^ n379 ^ 1'b0 ;
  assign n23792 = n23788 & ~n23791 ;
  assign n23793 = n14261 | n17312 ;
  assign n23794 = n16480 & ~n23793 ;
  assign n23795 = n10183 ^ n4575 ^ 1'b0 ;
  assign n23796 = n1957 & ~n23795 ;
  assign n23797 = n20951 ^ n13166 ^ n3511 ;
  assign n23798 = ~n9776 & n23797 ;
  assign n23799 = n23798 ^ n17539 ^ 1'b0 ;
  assign n23800 = ~n19965 & n23799 ;
  assign n23801 = ~n15867 & n23800 ;
  assign n23802 = ~n23796 & n23801 ;
  assign n23803 = ( ~n1303 & n4980 ) | ( ~n1303 & n17366 ) | ( n4980 & n17366 ) ;
  assign n23804 = n11832 ^ n5397 ^ 1'b0 ;
  assign n23805 = ~n6671 & n23804 ;
  assign n23806 = n6365 ^ n1281 ^ 1'b0 ;
  assign n23807 = n892 & n23806 ;
  assign n23808 = n23805 & ~n23807 ;
  assign n23809 = ( n11270 & n23803 ) | ( n11270 & ~n23808 ) | ( n23803 & ~n23808 ) ;
  assign n23810 = n23809 ^ n16922 ^ 1'b0 ;
  assign n23811 = n16639 ^ n6251 ^ n4282 ;
  assign n23812 = ( ~n4421 & n9479 ) | ( ~n4421 & n17375 ) | ( n9479 & n17375 ) ;
  assign n23813 = n23812 ^ n23537 ^ 1'b0 ;
  assign n23814 = n4056 & ~n4267 ;
  assign n23815 = ( n3030 & n12042 ) | ( n3030 & ~n23814 ) | ( n12042 & ~n23814 ) ;
  assign n23816 = n11302 | n15520 ;
  assign n23817 = n23815 & ~n23816 ;
  assign n23818 = n12262 & ~n23817 ;
  assign n23819 = n3322 & n23818 ;
  assign n23820 = n3870 & ~n11766 ;
  assign n23821 = ( n4315 & n15304 ) | ( n4315 & ~n23820 ) | ( n15304 & ~n23820 ) ;
  assign n23822 = n305 | n23821 ;
  assign n23823 = n18531 & ~n23822 ;
  assign n23824 = n12794 ^ n7551 ^ 1'b0 ;
  assign n23825 = ~n8860 & n23824 ;
  assign n23826 = ~n2179 & n23825 ;
  assign n23827 = n1802 & ~n23826 ;
  assign n23828 = n23823 & n23827 ;
  assign n23829 = n2530 & n13648 ;
  assign n23830 = n23829 ^ n4474 ^ 1'b0 ;
  assign n23831 = n23830 ^ n6967 ^ n6331 ;
  assign n23832 = n3958 ^ n1299 ^ 1'b0 ;
  assign n23833 = n2943 & ~n23832 ;
  assign n23834 = n23833 ^ n22308 ^ n11042 ;
  assign n23836 = n782 & n3666 ;
  assign n23837 = n11461 & ~n23836 ;
  assign n23835 = n16492 ^ n8484 ^ n487 ;
  assign n23838 = n23837 ^ n23835 ^ 1'b0 ;
  assign n23839 = n966 & ~n1098 ;
  assign n23840 = ~n23838 & n23839 ;
  assign n23841 = n4607 ^ n4053 ^ 1'b0 ;
  assign n23842 = n23841 ^ n23313 ^ 1'b0 ;
  assign n23843 = ~n2914 & n23842 ;
  assign n23844 = n8671 ^ n7196 ^ 1'b0 ;
  assign n23845 = ( n554 & ~n2357 ) | ( n554 & n3502 ) | ( ~n2357 & n3502 ) ;
  assign n23846 = n10398 | n23845 ;
  assign n23847 = n23844 | n23846 ;
  assign n23848 = ~n3012 & n12180 ;
  assign n23849 = n23848 ^ n9790 ^ 1'b0 ;
  assign n23850 = ~n5935 & n23849 ;
  assign n23851 = n8936 & n23850 ;
  assign n23852 = ~n14041 & n16043 ;
  assign n23853 = n14047 | n23852 ;
  assign n23854 = n23853 ^ n3927 ^ 1'b0 ;
  assign n23855 = ~n23851 & n23854 ;
  assign n23856 = n4710 & n23855 ;
  assign n23857 = n947 & ~n13091 ;
  assign n23858 = n977 | n23857 ;
  assign n23859 = n18634 & ~n23858 ;
  assign n23860 = n23859 ^ n16721 ^ 1'b0 ;
  assign n23861 = n12830 | n23860 ;
  assign n23865 = n13147 ^ n3614 ^ 1'b0 ;
  assign n23866 = ~n18456 & n23865 ;
  assign n23867 = n13077 & n23866 ;
  assign n23863 = n7269 ^ n1906 ^ 1'b0 ;
  assign n23864 = n21244 & n23863 ;
  assign n23862 = n13999 ^ n8977 ^ 1'b0 ;
  assign n23868 = n23867 ^ n23864 ^ n23862 ;
  assign n23869 = n6125 | n23868 ;
  assign n23870 = n10970 | n23869 ;
  assign n23871 = n5371 & ~n6091 ;
  assign n23872 = ~n5622 & n23871 ;
  assign n23873 = n16278 ^ n9771 ^ n3305 ;
  assign n23874 = n23873 ^ n7060 ^ 1'b0 ;
  assign n23875 = n1489 & n23874 ;
  assign n23876 = n23875 ^ n9089 ^ n4520 ;
  assign n23877 = ( n3468 & ~n6928 ) | ( n3468 & n17840 ) | ( ~n6928 & n17840 ) ;
  assign n23878 = ~n5296 & n7927 ;
  assign n23879 = n1823 ^ n1591 ^ 1'b0 ;
  assign n23880 = ( n9904 & n14858 ) | ( n9904 & ~n23879 ) | ( n14858 & ~n23879 ) ;
  assign n23882 = n4355 | n4583 ;
  assign n23881 = ~n21599 & n22408 ;
  assign n23883 = n23882 ^ n23881 ^ 1'b0 ;
  assign n23884 = n9077 ^ n5781 ^ 1'b0 ;
  assign n23885 = n18901 ^ n2223 ^ 1'b0 ;
  assign n23886 = n18789 | n23885 ;
  assign n23887 = ( n19299 & n20145 ) | ( n19299 & ~n23886 ) | ( n20145 & ~n23886 ) ;
  assign n23888 = ( n7481 & ~n7581 ) | ( n7481 & n14900 ) | ( ~n7581 & n14900 ) ;
  assign n23889 = n18907 ^ n10017 ^ 1'b0 ;
  assign n23890 = n21807 | n23889 ;
  assign n23891 = n23890 ^ n7719 ^ 1'b0 ;
  assign n23892 = ~n7962 & n23891 ;
  assign n23893 = ( ~n4438 & n10320 ) | ( ~n4438 & n13831 ) | ( n10320 & n13831 ) ;
  assign n23894 = n15799 ^ n12813 ^ n8312 ;
  assign n23895 = n18615 ^ n15841 ^ 1'b0 ;
  assign n23896 = n23894 & n23895 ;
  assign n23897 = n23896 ^ n16459 ^ n8311 ;
  assign n23898 = ( n363 & n10481 ) | ( n363 & ~n19436 ) | ( n10481 & ~n19436 ) ;
  assign n23899 = ( n2553 & n12310 ) | ( n2553 & n23898 ) | ( n12310 & n23898 ) ;
  assign n23900 = ( n770 & ~n2186 ) | ( n770 & n13717 ) | ( ~n2186 & n13717 ) ;
  assign n23901 = n2260 & ~n13460 ;
  assign n23902 = n23900 | n23901 ;
  assign n23903 = x209 & n4506 ;
  assign n23904 = ~n9814 & n23903 ;
  assign n23905 = n1436 & ~n23904 ;
  assign n23906 = n16851 & n23905 ;
  assign n23907 = n8337 ^ n6705 ^ 1'b0 ;
  assign n23908 = ~n23906 & n23907 ;
  assign n23909 = ( n10149 & n14315 ) | ( n10149 & n16282 ) | ( n14315 & n16282 ) ;
  assign n23910 = ~n952 & n6373 ;
  assign n23911 = n23910 ^ n12515 ^ 1'b0 ;
  assign n23912 = n9714 ^ x112 ^ 1'b0 ;
  assign n23913 = n11464 & ~n23912 ;
  assign n23914 = ~n14551 & n23913 ;
  assign n23915 = n4765 & ~n19606 ;
  assign n23916 = n21342 ^ n12922 ^ 1'b0 ;
  assign n23917 = n10063 ^ n8179 ^ 1'b0 ;
  assign n23918 = ( n2103 & n5902 ) | ( n2103 & n20503 ) | ( n5902 & n20503 ) ;
  assign n23919 = n15507 ^ n4219 ^ 1'b0 ;
  assign n23920 = n6662 & ~n7388 ;
  assign n23921 = n9446 ^ n8091 ^ n1785 ;
  assign n23922 = n5581 & ~n23921 ;
  assign n23923 = n23922 ^ n21697 ^ n19810 ;
  assign n23924 = n10770 & n12653 ;
  assign n23925 = n2899 & n23924 ;
  assign n23926 = n23923 | n23925 ;
  assign n23927 = ~n23920 & n23926 ;
  assign n23928 = ( n1099 & ~n2211 ) | ( n1099 & n13317 ) | ( ~n2211 & n13317 ) ;
  assign n23932 = n18615 ^ n7817 ^ n7801 ;
  assign n23930 = n15743 ^ n12805 ^ x236 ;
  assign n23929 = ( n4390 & n19707 ) | ( n4390 & n21809 ) | ( n19707 & n21809 ) ;
  assign n23931 = n23930 ^ n23929 ^ n5585 ;
  assign n23933 = n23932 ^ n23931 ^ 1'b0 ;
  assign n23934 = n23928 & n23933 ;
  assign n23935 = n12460 ^ n2611 ^ 1'b0 ;
  assign n23936 = n12702 | n23935 ;
  assign n23937 = n22535 ^ n8792 ^ 1'b0 ;
  assign n23938 = ( n7413 & n23936 ) | ( n7413 & n23937 ) | ( n23936 & n23937 ) ;
  assign n23939 = n18563 ^ n15446 ^ 1'b0 ;
  assign n23940 = n1158 & n3933 ;
  assign n23941 = ( n1975 & n13529 ) | ( n1975 & n16555 ) | ( n13529 & n16555 ) ;
  assign n23942 = n23941 ^ n23817 ^ 1'b0 ;
  assign n23943 = n23940 & ~n23942 ;
  assign n23946 = ~x226 & n8913 ;
  assign n23947 = n23946 ^ n11281 ^ 1'b0 ;
  assign n23948 = n5068 ^ n860 ^ 1'b0 ;
  assign n23949 = n23947 | n23948 ;
  assign n23944 = n1635 & n2957 ;
  assign n23945 = n23944 ^ n5716 ^ 1'b0 ;
  assign n23950 = n23949 ^ n23945 ^ 1'b0 ;
  assign n23951 = n23950 ^ n18603 ^ n8930 ;
  assign n23953 = n5540 ^ n806 ^ n258 ;
  assign n23952 = ( n4247 & ~n5728 ) | ( n4247 & n23354 ) | ( ~n5728 & n23354 ) ;
  assign n23954 = n23953 ^ n23952 ^ n12116 ;
  assign n23955 = n1838 & ~n4189 ;
  assign n23956 = ~n6815 & n23955 ;
  assign n23957 = n11627 & n16716 ;
  assign n23958 = ~n3655 & n23957 ;
  assign n23959 = n23956 & n23958 ;
  assign n23961 = ~n7482 & n8832 ;
  assign n23960 = ( n3281 & n6153 ) | ( n3281 & ~n11704 ) | ( n6153 & ~n11704 ) ;
  assign n23962 = n23961 ^ n23960 ^ n3371 ;
  assign n23963 = n1868 | n3487 ;
  assign n23964 = n20845 | n23963 ;
  assign n23965 = n19831 ^ n14844 ^ n8563 ;
  assign n23966 = x17 & n8514 ;
  assign n23967 = n23965 & n23966 ;
  assign n23971 = n3080 ^ n668 ^ 1'b0 ;
  assign n23970 = ( n3347 & n4307 ) | ( n3347 & ~n5422 ) | ( n4307 & ~n5422 ) ;
  assign n23972 = n23971 ^ n23970 ^ n15662 ;
  assign n23968 = ( n9109 & ~n14258 ) | ( n9109 & n17489 ) | ( ~n14258 & n17489 ) ;
  assign n23969 = ( n1703 & n11472 ) | ( n1703 & n23968 ) | ( n11472 & n23968 ) ;
  assign n23973 = n23972 ^ n23969 ^ 1'b0 ;
  assign n23974 = n9805 & n11192 ;
  assign n23975 = ( ~n9322 & n10843 ) | ( ~n9322 & n16957 ) | ( n10843 & n16957 ) ;
  assign n23976 = n16811 ^ n11489 ^ n297 ;
  assign n23977 = n2554 ^ n2057 ^ 1'b0 ;
  assign n23978 = n4157 | n23977 ;
  assign n23979 = n23978 ^ n2066 ^ 1'b0 ;
  assign n23980 = ( n404 & n5959 ) | ( n404 & ~n23979 ) | ( n5959 & ~n23979 ) ;
  assign n23981 = n8510 | n23980 ;
  assign n23982 = n10957 & ~n23981 ;
  assign n23983 = n6722 | n23982 ;
  assign n23984 = n23983 ^ n1851 ^ 1'b0 ;
  assign n23985 = n2363 ^ n808 ^ 1'b0 ;
  assign n23986 = n23985 ^ n22493 ^ n4840 ;
  assign n23987 = n23986 ^ n1080 ^ 1'b0 ;
  assign n23988 = ( n3583 & n19806 ) | ( n3583 & n19829 ) | ( n19806 & n19829 ) ;
  assign n23989 = ( n1474 & ~n7659 ) | ( n1474 & n23988 ) | ( ~n7659 & n23988 ) ;
  assign n23990 = n15631 | n23989 ;
  assign n23991 = n4346 & ~n11134 ;
  assign n23992 = n23991 ^ n18277 ^ n4708 ;
  assign n23993 = ( n7562 & n19914 ) | ( n7562 & ~n23992 ) | ( n19914 & ~n23992 ) ;
  assign n23994 = n23953 ^ n9721 ^ 1'b0 ;
  assign n23995 = n11071 | n23994 ;
  assign n23996 = n8941 | n9598 ;
  assign n23997 = n23995 & ~n23996 ;
  assign n23998 = n23997 ^ n5780 ^ 1'b0 ;
  assign n23999 = n21052 ^ n388 ^ 1'b0 ;
  assign n24000 = n2834 & n23999 ;
  assign n24001 = ~n3619 & n5601 ;
  assign n24002 = n24001 ^ n2933 ^ 1'b0 ;
  assign n24003 = x107 & ~n24002 ;
  assign n24004 = n24003 ^ n7701 ^ 1'b0 ;
  assign n24005 = ( ~n7500 & n18279 ) | ( ~n7500 & n24004 ) | ( n18279 & n24004 ) ;
  assign n24006 = ( n10863 & ~n12181 ) | ( n10863 & n22660 ) | ( ~n12181 & n22660 ) ;
  assign n24007 = n24006 ^ n1502 ^ 1'b0 ;
  assign n24008 = n24005 & n24007 ;
  assign n24009 = ( n521 & ~n3177 ) | ( n521 & n5848 ) | ( ~n3177 & n5848 ) ;
  assign n24010 = ( n7315 & ~n14492 ) | ( n7315 & n24009 ) | ( ~n14492 & n24009 ) ;
  assign n24011 = n15319 & n19377 ;
  assign n24012 = n24011 ^ n6517 ^ 1'b0 ;
  assign n24013 = n12550 ^ n3322 ^ 1'b0 ;
  assign n24014 = ( n2154 & ~n5329 ) | ( n2154 & n23526 ) | ( ~n5329 & n23526 ) ;
  assign n24015 = ~n11474 & n24014 ;
  assign n24016 = n2554 & n7052 ;
  assign n24017 = n24016 ^ n3118 ^ 1'b0 ;
  assign n24018 = ~n8301 & n23783 ;
  assign n24019 = n24018 ^ n10757 ^ 1'b0 ;
  assign n24020 = n20276 ^ n8045 ^ 1'b0 ;
  assign n24021 = n652 ^ n334 ^ 1'b0 ;
  assign n24022 = ( ~n5493 & n10233 ) | ( ~n5493 & n24021 ) | ( n10233 & n24021 ) ;
  assign n24023 = n11622 ^ n9769 ^ n5520 ;
  assign n24024 = n24023 ^ n16662 ^ n9494 ;
  assign n24025 = n24024 ^ n16598 ^ n12612 ;
  assign n24027 = n2567 ^ n382 ^ 1'b0 ;
  assign n24028 = n1165 & ~n9568 ;
  assign n24029 = ~n24027 & n24028 ;
  assign n24030 = n12296 | n24029 ;
  assign n24031 = n15813 | n24030 ;
  assign n24026 = ( ~n14685 & n16470 ) | ( ~n14685 & n23576 ) | ( n16470 & n23576 ) ;
  assign n24032 = n24031 ^ n24026 ^ 1'b0 ;
  assign n24033 = n20395 ^ n11459 ^ n1878 ;
  assign n24034 = n24033 ^ n9722 ^ x237 ;
  assign n24035 = n5754 & n5953 ;
  assign n24036 = n15085 ^ n12999 ^ 1'b0 ;
  assign n24037 = n18568 ^ n7801 ^ 1'b0 ;
  assign n24038 = n6744 | n24037 ;
  assign n24039 = n2490 & n2639 ;
  assign n24040 = ~n8962 & n24039 ;
  assign n24041 = n17219 | n24040 ;
  assign n24042 = n24041 ^ n20793 ^ 1'b0 ;
  assign n24043 = n24038 | n24042 ;
  assign n24044 = n24036 | n24043 ;
  assign n24045 = ~n24035 & n24044 ;
  assign n24046 = ~n7421 & n24045 ;
  assign n24047 = n18688 ^ n1532 ^ 1'b0 ;
  assign n24051 = n20937 ^ n17429 ^ n4518 ;
  assign n24056 = ( n1838 & ~n6551 ) | ( n1838 & n8893 ) | ( ~n6551 & n8893 ) ;
  assign n24052 = ( n3647 & ~n4999 ) | ( n3647 & n12726 ) | ( ~n4999 & n12726 ) ;
  assign n24053 = n12125 ^ n3951 ^ 1'b0 ;
  assign n24054 = n24052 | n24053 ;
  assign n24055 = n16568 & ~n24054 ;
  assign n24057 = n24056 ^ n24055 ^ 1'b0 ;
  assign n24058 = ( n14368 & n24051 ) | ( n14368 & ~n24057 ) | ( n24051 & ~n24057 ) ;
  assign n24048 = n2353 | n12532 ;
  assign n24049 = n24048 ^ n14832 ^ n6644 ;
  assign n24050 = n19448 | n24049 ;
  assign n24059 = n24058 ^ n24050 ^ 1'b0 ;
  assign n24060 = n21490 ^ n4106 ^ 1'b0 ;
  assign n24061 = n24059 & n24060 ;
  assign n24062 = n4689 | n21233 ;
  assign n24063 = n24062 ^ n14232 ^ 1'b0 ;
  assign n24064 = x151 & ~n11840 ;
  assign n24066 = n1832 | n19770 ;
  assign n24067 = n24066 ^ n7086 ^ 1'b0 ;
  assign n24065 = ( n5774 & n8377 ) | ( n5774 & ~n17546 ) | ( n8377 & ~n17546 ) ;
  assign n24068 = n24067 ^ n24065 ^ 1'b0 ;
  assign n24069 = ( n24063 & ~n24064 ) | ( n24063 & n24068 ) | ( ~n24064 & n24068 ) ;
  assign n24070 = n19213 ^ n16141 ^ n7356 ;
  assign n24071 = n5744 | n9685 ;
  assign n24072 = n18054 & ~n24071 ;
  assign n24073 = n12547 ^ n10540 ^ 1'b0 ;
  assign n24074 = n23454 ^ n8229 ^ 1'b0 ;
  assign n24075 = n6973 & ~n24074 ;
  assign n24076 = n8435 ^ n5753 ^ 1'b0 ;
  assign n24077 = ( n1403 & ~n16289 ) | ( n1403 & n24076 ) | ( ~n16289 & n24076 ) ;
  assign n24078 = n16488 ^ n11487 ^ 1'b0 ;
  assign n24079 = n15899 | n24078 ;
  assign n24080 = ( n2315 & n21162 ) | ( n2315 & ~n24079 ) | ( n21162 & ~n24079 ) ;
  assign n24081 = n15953 & n24080 ;
  assign n24082 = n19073 ^ n17987 ^ n7987 ;
  assign n24083 = n5853 & n10359 ;
  assign n24084 = n24083 ^ n19940 ^ n3787 ;
  assign n24085 = n4398 | n10641 ;
  assign n24086 = ( n20479 & n23050 ) | ( n20479 & ~n24085 ) | ( n23050 & ~n24085 ) ;
  assign n24087 = n17881 ^ n7929 ^ n4261 ;
  assign n24088 = n21634 ^ n17132 ^ 1'b0 ;
  assign n24089 = ( ~n10976 & n24087 ) | ( ~n10976 & n24088 ) | ( n24087 & n24088 ) ;
  assign n24090 = ( x79 & n24086 ) | ( x79 & ~n24089 ) | ( n24086 & ~n24089 ) ;
  assign n24091 = ( n7325 & ~n7593 ) | ( n7325 & n14470 ) | ( ~n7593 & n14470 ) ;
  assign n24092 = n24091 ^ n20316 ^ 1'b0 ;
  assign n24093 = n14401 & ~n24092 ;
  assign n24094 = ~n12350 & n22685 ;
  assign n24095 = n18348 ^ n13694 ^ n3275 ;
  assign n24096 = ~n3450 & n14041 ;
  assign n24097 = ~n675 & n24096 ;
  assign n24098 = ( n15616 & ~n24095 ) | ( n15616 & n24097 ) | ( ~n24095 & n24097 ) ;
  assign n24099 = ( ~n396 & n20923 ) | ( ~n396 & n24098 ) | ( n20923 & n24098 ) ;
  assign n24100 = n24099 ^ x238 ^ 1'b0 ;
  assign n24101 = n24094 & n24100 ;
  assign n24102 = n2105 | n7771 ;
  assign n24103 = n15264 | n24102 ;
  assign n24104 = ~n11853 & n24103 ;
  assign n24105 = n21314 ^ n12000 ^ 1'b0 ;
  assign n24106 = n5966 & n9611 ;
  assign n24107 = n24106 ^ n7943 ^ 1'b0 ;
  assign n24108 = n10086 | n18955 ;
  assign n24109 = n9131 & ~n24108 ;
  assign n24110 = n15662 & ~n24109 ;
  assign n24111 = ~n15662 & n24110 ;
  assign n24112 = n20065 & ~n24111 ;
  assign n24113 = ~n17678 & n24112 ;
  assign n24114 = n12881 ^ n8905 ^ 1'b0 ;
  assign n24115 = ~n11084 & n24114 ;
  assign n24116 = n24115 ^ n23639 ^ n7420 ;
  assign n24118 = ( x42 & ~n3141 ) | ( x42 & n8117 ) | ( ~n3141 & n8117 ) ;
  assign n24117 = n22385 ^ n10934 ^ n7682 ;
  assign n24119 = n24118 ^ n24117 ^ n11719 ;
  assign n24120 = n15254 ^ n14395 ^ n8910 ;
  assign n24121 = n13358 ^ n9907 ^ 1'b0 ;
  assign n24122 = n24120 & ~n24121 ;
  assign n24123 = n20300 & n24122 ;
  assign n24124 = n1475 | n9197 ;
  assign n24125 = n24124 ^ n6802 ^ 1'b0 ;
  assign n24126 = n24125 ^ n13488 ^ n4259 ;
  assign n24127 = n24126 ^ n13593 ^ 1'b0 ;
  assign n24128 = ( n7453 & n9505 ) | ( n7453 & n12561 ) | ( n9505 & n12561 ) ;
  assign n24129 = n20907 ^ n16559 ^ n6361 ;
  assign n24130 = n282 & ~n7049 ;
  assign n24131 = n24130 ^ n3515 ^ 1'b0 ;
  assign n24132 = ~n11543 & n24131 ;
  assign n24133 = n24129 & n24132 ;
  assign n24134 = n4882 & n5303 ;
  assign n24135 = n14278 & ~n14620 ;
  assign n24136 = ( n8262 & n24134 ) | ( n8262 & ~n24135 ) | ( n24134 & ~n24135 ) ;
  assign n24137 = n12059 ^ n5209 ^ 1'b0 ;
  assign n24138 = n5682 & n24137 ;
  assign n24139 = n24138 ^ n5464 ^ 1'b0 ;
  assign n24140 = n10533 & ~n24139 ;
  assign n24141 = n24140 ^ n532 ^ 1'b0 ;
  assign n24142 = n8477 ^ n1738 ^ 1'b0 ;
  assign n24143 = n5876 | n24142 ;
  assign n24144 = ~n1020 & n5945 ;
  assign n24145 = n731 & n24144 ;
  assign n24146 = n24145 ^ n2252 ^ n886 ;
  assign n24147 = ( ~n4439 & n11175 ) | ( ~n4439 & n24146 ) | ( n11175 & n24146 ) ;
  assign n24148 = ( n12532 & ~n23716 ) | ( n12532 & n24147 ) | ( ~n23716 & n24147 ) ;
  assign n24149 = n7050 ^ n4568 ^ 1'b0 ;
  assign n24150 = n6694 | n24149 ;
  assign n24151 = ( n17866 & n20609 ) | ( n17866 & ~n24150 ) | ( n20609 & ~n24150 ) ;
  assign n24152 = n19167 ^ n8409 ^ 1'b0 ;
  assign n24154 = ( n1667 & n2469 ) | ( n1667 & ~n3891 ) | ( n2469 & ~n3891 ) ;
  assign n24155 = ( n3803 & ~n6218 ) | ( n3803 & n24154 ) | ( ~n6218 & n24154 ) ;
  assign n24156 = n24155 ^ n1879 ^ 1'b0 ;
  assign n24157 = n24156 ^ n11725 ^ n9858 ;
  assign n24158 = n24157 ^ n13483 ^ n9929 ;
  assign n24153 = n10551 | n13804 ;
  assign n24159 = n24158 ^ n24153 ^ 1'b0 ;
  assign n24160 = n5425 & ~n9274 ;
  assign n24161 = ( ~n5694 & n11231 ) | ( ~n5694 & n12107 ) | ( n11231 & n12107 ) ;
  assign n24162 = ~n7584 & n12535 ;
  assign n24163 = n11300 & ~n21671 ;
  assign n24164 = ~n24162 & n24163 ;
  assign n24165 = ~n14945 & n24164 ;
  assign n24166 = n9170 & ~n24165 ;
  assign n24167 = n24161 & n24166 ;
  assign n24168 = n15142 ^ n12640 ^ n10958 ;
  assign n24169 = n24168 ^ n20533 ^ n1470 ;
  assign n24170 = ~n11244 & n24169 ;
  assign n24171 = ~n23039 & n24170 ;
  assign n24172 = n632 & ~n3409 ;
  assign n24173 = n24172 ^ n5741 ^ 1'b0 ;
  assign n24174 = n1608 & n2807 ;
  assign n24175 = n18939 ^ n4041 ^ n1264 ;
  assign n24176 = n24175 ^ n10379 ^ n4596 ;
  assign n24177 = x242 & n4206 ;
  assign n24178 = n24177 ^ n20860 ^ 1'b0 ;
  assign n24179 = n22848 & ~n24178 ;
  assign n24180 = n24179 ^ n13580 ^ 1'b0 ;
  assign n24181 = n15345 & ~n24180 ;
  assign n24182 = ~n410 & n13294 ;
  assign n24185 = n11790 ^ n11340 ^ 1'b0 ;
  assign n24183 = n1719 ^ n709 ^ 1'b0 ;
  assign n24184 = n9322 | n24183 ;
  assign n24186 = n24185 ^ n24184 ^ n4471 ;
  assign n24197 = ( n6645 & n17096 ) | ( n6645 & n18700 ) | ( n17096 & n18700 ) ;
  assign n24190 = n12317 ^ n6213 ^ n2995 ;
  assign n24191 = x23 & n24190 ;
  assign n24192 = ~n5366 & n24191 ;
  assign n24193 = ~n5411 & n8882 ;
  assign n24194 = n24192 & n24193 ;
  assign n24195 = n4086 & n24194 ;
  assign n24196 = n7437 & ~n24195 ;
  assign n24198 = n24197 ^ n24196 ^ 1'b0 ;
  assign n24187 = n18900 ^ x133 ^ 1'b0 ;
  assign n24188 = ~n8566 & n24187 ;
  assign n24189 = n24188 ^ n3100 ^ 1'b0 ;
  assign n24199 = n24198 ^ n24189 ^ n21056 ;
  assign n24201 = n16772 & ~n17069 ;
  assign n24200 = n10903 ^ n10485 ^ n6549 ;
  assign n24202 = n24201 ^ n24200 ^ 1'b0 ;
  assign n24203 = n2683 & ~n15870 ;
  assign n24205 = n1344 ^ n943 ^ 1'b0 ;
  assign n24206 = x82 & n24205 ;
  assign n24204 = n10679 | n22910 ;
  assign n24207 = n24206 ^ n24204 ^ 1'b0 ;
  assign n24208 = n18463 & n24207 ;
  assign n24209 = n12624 & n24208 ;
  assign n24210 = n24209 ^ n23413 ^ 1'b0 ;
  assign n24211 = n18643 ^ n1398 ^ 1'b0 ;
  assign n24212 = n17208 ^ n11112 ^ n11032 ;
  assign n24213 = n24212 ^ n9522 ^ n7874 ;
  assign n24214 = n14739 ^ n3557 ^ 1'b0 ;
  assign n24215 = n16283 ^ n12790 ^ 1'b0 ;
  assign n24216 = n24214 & n24215 ;
  assign n24217 = ( n19189 & n24213 ) | ( n19189 & ~n24216 ) | ( n24213 & ~n24216 ) ;
  assign n24218 = n4011 | n16315 ;
  assign n24219 = n24218 ^ n7060 ^ n2127 ;
  assign n24220 = n2282 & ~n10095 ;
  assign n24221 = ~n17470 & n24220 ;
  assign n24222 = n24221 ^ n8424 ^ 1'b0 ;
  assign n24223 = n6762 & ~n24222 ;
  assign n24224 = n2107 & ~n21297 ;
  assign n24225 = n5682 & n9803 ;
  assign n24226 = n24225 ^ n1221 ^ 1'b0 ;
  assign n24227 = ~n15153 & n24226 ;
  assign n24228 = n16746 | n24227 ;
  assign n24229 = n24224 & n24228 ;
  assign n24230 = n24229 ^ x164 ^ 1'b0 ;
  assign n24231 = ( ~n6921 & n7544 ) | ( ~n6921 & n12542 ) | ( n7544 & n12542 ) ;
  assign n24232 = n24231 ^ n22522 ^ n12579 ;
  assign n24233 = ( n1975 & ~n4579 ) | ( n1975 & n6586 ) | ( ~n4579 & n6586 ) ;
  assign n24234 = n13328 | n16161 ;
  assign n24235 = n24233 | n24234 ;
  assign n24236 = ~n15783 & n24235 ;
  assign n24237 = n4379 | n4805 ;
  assign n24238 = n4962 & ~n24237 ;
  assign n24239 = ~n9248 & n14247 ;
  assign n24240 = n24239 ^ n4253 ^ 1'b0 ;
  assign n24241 = n24240 ^ n18836 ^ 1'b0 ;
  assign n24242 = n22703 ^ n4845 ^ 1'b0 ;
  assign n24243 = n483 ^ n428 ^ 1'b0 ;
  assign n24244 = n9986 & ~n24243 ;
  assign n24245 = ( n8234 & ~n10631 ) | ( n8234 & n24244 ) | ( ~n10631 & n24244 ) ;
  assign n24246 = n14506 ^ n7373 ^ n3579 ;
  assign n24247 = n7787 ^ n3465 ^ 1'b0 ;
  assign n24248 = ( n21494 & n24246 ) | ( n21494 & ~n24247 ) | ( n24246 & ~n24247 ) ;
  assign n24249 = ~n3406 & n3509 ;
  assign n24250 = ~n24248 & n24249 ;
  assign n24251 = n17275 ^ n11669 ^ 1'b0 ;
  assign n24252 = ~n1241 & n12393 ;
  assign n24253 = ~n15021 & n24252 ;
  assign n24254 = n22491 | n24253 ;
  assign n24255 = n21660 ^ n13223 ^ n1915 ;
  assign n24256 = n24255 ^ n17044 ^ n5362 ;
  assign n24257 = n13571 ^ n2836 ^ n2534 ;
  assign n24258 = n2886 & n14256 ;
  assign n24259 = ~n4376 & n13423 ;
  assign n24260 = n5026 & n24259 ;
  assign n24261 = n24260 ^ n16483 ^ 1'b0 ;
  assign n24262 = n24261 ^ n14710 ^ n1358 ;
  assign n24263 = n21220 ^ n17677 ^ n6740 ;
  assign n24264 = ( x75 & ~n9397 ) | ( x75 & n12222 ) | ( ~n9397 & n12222 ) ;
  assign n24273 = n1229 & n19602 ;
  assign n24274 = n24273 ^ n5491 ^ 1'b0 ;
  assign n24275 = ( n4266 & ~n11325 ) | ( n4266 & n24274 ) | ( ~n11325 & n24274 ) ;
  assign n24268 = n12884 | n13496 ;
  assign n24269 = ~n10289 & n14197 ;
  assign n24270 = ~n1806 & n24269 ;
  assign n24271 = n7949 & ~n24270 ;
  assign n24272 = ~n24268 & n24271 ;
  assign n24265 = ~n4921 & n22433 ;
  assign n24266 = n24265 ^ n10769 ^ 1'b0 ;
  assign n24267 = ~n9446 & n24266 ;
  assign n24276 = n24275 ^ n24272 ^ n24267 ;
  assign n24277 = n10734 & n19196 ;
  assign n24278 = n24277 ^ n17883 ^ 1'b0 ;
  assign n24279 = n8882 & n18550 ;
  assign n24280 = n24279 ^ n3666 ^ 1'b0 ;
  assign n24281 = ~n1353 & n13104 ;
  assign n24282 = n24280 & n24281 ;
  assign n24283 = n11719 ^ n5706 ^ n1377 ;
  assign n24287 = n17517 ^ n7785 ^ n6807 ;
  assign n24288 = n2788 & ~n8635 ;
  assign n24289 = n24288 ^ n11031 ^ 1'b0 ;
  assign n24290 = n24287 & n24289 ;
  assign n24291 = ( n16282 & n17255 ) | ( n16282 & n24290 ) | ( n17255 & n24290 ) ;
  assign n24285 = ~n8996 & n12111 ;
  assign n24286 = n24285 ^ n3548 ^ 1'b0 ;
  assign n24284 = n19483 ^ n14692 ^ 1'b0 ;
  assign n24292 = n24291 ^ n24286 ^ n24284 ;
  assign n24293 = n20271 ^ n10102 ^ n2638 ;
  assign n24294 = n14846 ^ n7902 ^ 1'b0 ;
  assign n24295 = n11138 | n24294 ;
  assign n24296 = n18878 ^ n6490 ^ 1'b0 ;
  assign n24297 = n24296 ^ n10312 ^ 1'b0 ;
  assign n24298 = n1056 ^ x200 ^ 1'b0 ;
  assign n24299 = n21775 & ~n24298 ;
  assign n24300 = ~n24065 & n24299 ;
  assign n24301 = n24300 ^ n14381 ^ 1'b0 ;
  assign n24303 = ~n4235 & n20423 ;
  assign n24302 = n18324 & n21965 ;
  assign n24304 = n24303 ^ n24302 ^ 1'b0 ;
  assign n24306 = n8374 & n19973 ;
  assign n24307 = n3571 & n24306 ;
  assign n24305 = n8441 & n8956 ;
  assign n24308 = n24307 ^ n24305 ^ 1'b0 ;
  assign n24309 = n4604 ^ n2939 ^ 1'b0 ;
  assign n24310 = n8675 ^ n1274 ^ 1'b0 ;
  assign n24311 = ~n1429 & n24310 ;
  assign n24312 = n24311 ^ n5882 ^ 1'b0 ;
  assign n24313 = ( n22472 & ~n24309 ) | ( n22472 & n24312 ) | ( ~n24309 & n24312 ) ;
  assign n24314 = n10518 ^ n2492 ^ 1'b0 ;
  assign n24315 = n24313 | n24314 ;
  assign n24316 = ~n3038 & n3205 ;
  assign n24317 = n9695 ^ n6380 ^ 1'b0 ;
  assign n24318 = ( n2187 & ~n8023 ) | ( n2187 & n19496 ) | ( ~n8023 & n19496 ) ;
  assign n24319 = ( n7844 & ~n10852 ) | ( n7844 & n24318 ) | ( ~n10852 & n24318 ) ;
  assign n24320 = ( n12461 & n13385 ) | ( n12461 & ~n20999 ) | ( n13385 & ~n20999 ) ;
  assign n24321 = n23523 ^ n21935 ^ n3881 ;
  assign n24322 = n4582 & ~n12759 ;
  assign n24323 = ( ~n4707 & n5205 ) | ( ~n4707 & n17498 ) | ( n5205 & n17498 ) ;
  assign n24327 = n5929 & ~n21890 ;
  assign n24328 = n24327 ^ n18828 ^ 1'b0 ;
  assign n24324 = ~n7026 & n8834 ;
  assign n24325 = n24324 ^ n5303 ^ n5088 ;
  assign n24326 = ~n23200 & n24325 ;
  assign n24329 = n24328 ^ n24326 ^ 1'b0 ;
  assign n24330 = n10436 ^ n9708 ^ 1'b0 ;
  assign n24331 = n11881 | n11997 ;
  assign n24332 = n24330 & ~n24331 ;
  assign n24333 = n18467 & ~n18763 ;
  assign n24335 = n11035 ^ n1783 ^ 1'b0 ;
  assign n24336 = n315 | n23605 ;
  assign n24337 = n24336 ^ n15965 ^ 1'b0 ;
  assign n24338 = n24337 ^ n14671 ^ n7019 ;
  assign n24339 = ( n2770 & n24335 ) | ( n2770 & n24338 ) | ( n24335 & n24338 ) ;
  assign n24334 = ~n4116 & n5308 ;
  assign n24340 = n24339 ^ n24334 ^ 1'b0 ;
  assign n24341 = n12780 & ~n13283 ;
  assign n24342 = ( ~x242 & n2045 ) | ( ~x242 & n4989 ) | ( n2045 & n4989 ) ;
  assign n24343 = n24342 ^ n12400 ^ n2192 ;
  assign n24344 = n24343 ^ n14739 ^ 1'b0 ;
  assign n24345 = ( ~n6815 & n14829 ) | ( ~n6815 & n16449 ) | ( n14829 & n16449 ) ;
  assign n24346 = n24344 & ~n24345 ;
  assign n24347 = x14 & n18978 ;
  assign n24348 = n24347 ^ n2113 ^ 1'b0 ;
  assign n24349 = ~n24346 & n24348 ;
  assign n24350 = n1667 & n14555 ;
  assign n24351 = n24350 ^ n14557 ^ 1'b0 ;
  assign n24352 = n6051 & ~n11181 ;
  assign n24353 = ~n3541 & n24352 ;
  assign n24354 = n7678 ^ n5264 ^ n4259 ;
  assign n24355 = n279 & ~n24354 ;
  assign n24356 = n22851 ^ n14912 ^ 1'b0 ;
  assign n24357 = n7431 ^ n1017 ^ 1'b0 ;
  assign n24358 = n24356 & ~n24357 ;
  assign n24359 = ~n9706 & n24358 ;
  assign n24360 = n24359 ^ n4119 ^ 1'b0 ;
  assign n24361 = n24360 ^ n2639 ^ 1'b0 ;
  assign n24362 = n24355 & ~n24361 ;
  assign n24363 = n24362 ^ n22122 ^ 1'b0 ;
  assign n24364 = ~n24353 & n24363 ;
  assign n24365 = n15194 ^ n14894 ^ n12114 ;
  assign n24366 = n15676 ^ n12829 ^ 1'b0 ;
  assign n24367 = ( n13886 & n17852 ) | ( n13886 & n24366 ) | ( n17852 & n24366 ) ;
  assign n24370 = n3563 & n9780 ;
  assign n24368 = n13720 ^ n7166 ^ n2295 ;
  assign n24369 = ~n5457 & n24368 ;
  assign n24371 = n24370 ^ n24369 ^ 1'b0 ;
  assign n24372 = n24371 ^ n6001 ^ 1'b0 ;
  assign n24373 = n12094 & n24372 ;
  assign n24374 = n7500 | n7843 ;
  assign n24375 = n24374 ^ n10661 ^ 1'b0 ;
  assign n24376 = n340 | n632 ;
  assign n24377 = n24376 ^ x152 ^ 1'b0 ;
  assign n24378 = n19224 & n24377 ;
  assign n24379 = ~n15975 & n24378 ;
  assign n24380 = n11303 | n14206 ;
  assign n24381 = ~n977 & n24380 ;
  assign n24382 = ( n14922 & ~n24379 ) | ( n14922 & n24381 ) | ( ~n24379 & n24381 ) ;
  assign n24383 = n16336 ^ n9801 ^ n2234 ;
  assign n24384 = n24383 ^ n4374 ^ n1108 ;
  assign n24385 = n11350 & n14178 ;
  assign n24386 = x114 & n17321 ;
  assign n24387 = n12329 & n24386 ;
  assign n24388 = n24387 ^ n21790 ^ 1'b0 ;
  assign n24389 = ~n3919 & n24388 ;
  assign n24390 = n24389 ^ n7840 ^ 1'b0 ;
  assign n24391 = n14049 ^ n9827 ^ n5660 ;
  assign n24392 = ~n2050 & n24391 ;
  assign n24393 = n24390 & n24392 ;
  assign n24394 = n9857 ^ x87 ^ 1'b0 ;
  assign n24396 = n3599 ^ n1795 ^ 1'b0 ;
  assign n24395 = n22563 ^ n18002 ^ 1'b0 ;
  assign n24397 = n24396 ^ n24395 ^ 1'b0 ;
  assign n24398 = n12311 ^ n12003 ^ 1'b0 ;
  assign n24399 = n4821 ^ n709 ^ 1'b0 ;
  assign n24400 = ~n1764 & n24399 ;
  assign n24401 = n24398 & n24400 ;
  assign n24402 = n23120 | n24401 ;
  assign n24403 = n24397 | n24402 ;
  assign n24404 = n16848 ^ n16421 ^ n1146 ;
  assign n24405 = ( n3492 & ~n4871 ) | ( n3492 & n19309 ) | ( ~n4871 & n19309 ) ;
  assign n24406 = ~n3967 & n24405 ;
  assign n24407 = n1317 | n10647 ;
  assign n24408 = n8484 ^ n5729 ^ 1'b0 ;
  assign n24409 = n18482 ^ n9729 ^ n1072 ;
  assign n24410 = n3960 | n16296 ;
  assign n24411 = n24410 ^ n1531 ^ 1'b0 ;
  assign n24412 = n6545 & ~n24411 ;
  assign n24413 = n10062 ^ n8024 ^ 1'b0 ;
  assign n24414 = n7110 ^ n6690 ^ 1'b0 ;
  assign n24415 = ( n11408 & n12424 ) | ( n11408 & n24414 ) | ( n12424 & n24414 ) ;
  assign n24416 = ( ~n3301 & n4212 ) | ( ~n3301 & n17707 ) | ( n4212 & n17707 ) ;
  assign n24417 = ( x189 & ~n16402 ) | ( x189 & n19134 ) | ( ~n16402 & n19134 ) ;
  assign n24418 = ~n24416 & n24417 ;
  assign n24419 = n21855 & n24418 ;
  assign n24420 = ~n1166 & n13457 ;
  assign n24421 = ( ~n7481 & n9309 ) | ( ~n7481 & n24420 ) | ( n9309 & n24420 ) ;
  assign n24422 = n24421 ^ n23416 ^ n11376 ;
  assign n24423 = n20325 | n24422 ;
  assign n24424 = n24423 ^ n16929 ^ 1'b0 ;
  assign n24425 = n22563 ^ n14532 ^ 1'b0 ;
  assign n24426 = n24425 ^ n17011 ^ 1'b0 ;
  assign n24427 = ~n8999 & n24426 ;
  assign n24428 = n24427 ^ n16837 ^ 1'b0 ;
  assign n24429 = n13907 ^ n11447 ^ 1'b0 ;
  assign n24435 = ~n1297 & n7479 ;
  assign n24436 = n24435 ^ n21982 ^ 1'b0 ;
  assign n24434 = ~n10448 & n24044 ;
  assign n24430 = n14905 ^ n9433 ^ n7538 ;
  assign n24431 = n24430 ^ n12798 ^ n11584 ;
  assign n24432 = ~n22988 & n23270 ;
  assign n24433 = ( n11216 & n24431 ) | ( n11216 & ~n24432 ) | ( n24431 & ~n24432 ) ;
  assign n24437 = n24436 ^ n24434 ^ n24433 ;
  assign n24438 = n2027 & n3874 ;
  assign n24439 = n5444 & ~n12718 ;
  assign n24440 = n24439 ^ n4777 ^ 1'b0 ;
  assign n24441 = n16310 ^ n1721 ^ 1'b0 ;
  assign n24442 = ( n4575 & n13744 ) | ( n4575 & ~n20698 ) | ( n13744 & ~n20698 ) ;
  assign n24443 = n9620 ^ n4540 ^ n1921 ;
  assign n24444 = n24443 ^ n4346 ^ n1428 ;
  assign n24447 = ( n13232 & n19569 ) | ( n13232 & n23807 ) | ( n19569 & n23807 ) ;
  assign n24445 = ( ~n1934 & n3734 ) | ( ~n1934 & n9220 ) | ( n3734 & n9220 ) ;
  assign n24446 = n24445 ^ n4745 ^ x199 ;
  assign n24448 = n24447 ^ n24446 ^ n23590 ;
  assign n24449 = n23116 | n24448 ;
  assign n24450 = ( n7564 & n7994 ) | ( n7564 & ~n9073 ) | ( n7994 & ~n9073 ) ;
  assign n24451 = n24450 ^ n17467 ^ 1'b0 ;
  assign n24452 = n24451 ^ n5154 ^ 1'b0 ;
  assign n24453 = n9247 | n21465 ;
  assign n24454 = n19056 & n23296 ;
  assign n24455 = n24454 ^ n10283 ^ 1'b0 ;
  assign n24456 = n5958 | n10881 ;
  assign n24457 = n23833 | n24456 ;
  assign n24458 = n24457 ^ n17509 ^ 1'b0 ;
  assign n24459 = n8935 | n24458 ;
  assign n24460 = n4470 ^ n1939 ^ 1'b0 ;
  assign n24461 = n9374 & ~n24460 ;
  assign n24462 = ( n329 & n4674 ) | ( n329 & n21741 ) | ( n4674 & n21741 ) ;
  assign n24463 = n24462 ^ n8005 ^ 1'b0 ;
  assign n24464 = n24463 ^ n5613 ^ 1'b0 ;
  assign n24465 = n21399 & ~n24464 ;
  assign n24466 = ~n6998 & n12946 ;
  assign n24467 = ( n3042 & ~n22079 ) | ( n3042 & n24466 ) | ( ~n22079 & n24466 ) ;
  assign n24468 = n3763 & n11140 ;
  assign n24469 = n24468 ^ n15260 ^ 1'b0 ;
  assign n24470 = ~n7531 & n24469 ;
  assign n24471 = ~n13104 & n24470 ;
  assign n24472 = n5456 & n17137 ;
  assign n24473 = n24471 & ~n24472 ;
  assign n24474 = ( n13483 & ~n21219 ) | ( n13483 & n24473 ) | ( ~n21219 & n24473 ) ;
  assign n24475 = ~n2903 & n12977 ;
  assign n24476 = ~n13690 & n24475 ;
  assign n24477 = ( n10896 & n21503 ) | ( n10896 & n22590 ) | ( n21503 & n22590 ) ;
  assign n24478 = n24477 ^ n24182 ^ 1'b0 ;
  assign n24479 = n15078 ^ n6369 ^ n5706 ;
  assign n24480 = n24479 ^ n524 ^ 1'b0 ;
  assign n24481 = ( x99 & n2112 ) | ( x99 & ~n15263 ) | ( n2112 & ~n15263 ) ;
  assign n24482 = n24481 ^ n18369 ^ 1'b0 ;
  assign n24483 = ~n17778 & n24482 ;
  assign n24484 = n24483 ^ n365 ^ 1'b0 ;
  assign n24487 = ( ~n2890 & n4774 ) | ( ~n2890 & n5029 ) | ( n4774 & n5029 ) ;
  assign n24488 = ( n10207 & n13915 ) | ( n10207 & ~n24487 ) | ( n13915 & ~n24487 ) ;
  assign n24486 = n7718 & ~n11047 ;
  assign n24489 = n24488 ^ n24486 ^ 1'b0 ;
  assign n24485 = n15137 | n16252 ;
  assign n24490 = n24489 ^ n24485 ^ 1'b0 ;
  assign n24491 = ~n4194 & n24490 ;
  assign n24492 = ~n8346 & n24491 ;
  assign n24493 = n14306 & n22372 ;
  assign n24494 = n10337 & n24493 ;
  assign n24495 = ( ~n3167 & n7703 ) | ( ~n3167 & n21202 ) | ( n7703 & n21202 ) ;
  assign n24496 = n18883 ^ n2533 ^ 1'b0 ;
  assign n24501 = ~n734 & n12635 ;
  assign n24502 = n24501 ^ n19647 ^ 1'b0 ;
  assign n24497 = n12266 ^ n6528 ^ n2705 ;
  assign n24498 = n14868 ^ n7500 ^ n7181 ;
  assign n24499 = n24498 ^ n22799 ^ n3173 ;
  assign n24500 = ( n18419 & n24497 ) | ( n18419 & ~n24499 ) | ( n24497 & ~n24499 ) ;
  assign n24503 = n24502 ^ n24500 ^ n22722 ;
  assign n24504 = n8410 & ~n21646 ;
  assign n24507 = ~n3144 & n8614 ;
  assign n24505 = n1563 & ~n6648 ;
  assign n24506 = ~n6219 & n24505 ;
  assign n24508 = n24507 ^ n24506 ^ 1'b0 ;
  assign n24509 = n24508 ^ n10026 ^ 1'b0 ;
  assign n24510 = n24504 & n24509 ;
  assign n24511 = n9849 ^ n4441 ^ 1'b0 ;
  assign n24512 = n22256 & ~n24511 ;
  assign n24513 = n6216 & n21034 ;
  assign n24514 = n22584 ^ n18481 ^ 1'b0 ;
  assign n24515 = n24513 & ~n24514 ;
  assign n24516 = n24337 ^ n9057 ^ 1'b0 ;
  assign n24517 = n16152 & ~n24516 ;
  assign n24518 = n8908 | n10924 ;
  assign n24519 = n12110 & n14487 ;
  assign n24520 = ( n15861 & n23639 ) | ( n15861 & ~n24519 ) | ( n23639 & ~n24519 ) ;
  assign n24521 = ( ~n20187 & n24518 ) | ( ~n20187 & n24520 ) | ( n24518 & n24520 ) ;
  assign n24522 = n19464 ^ n8385 ^ n1903 ;
  assign n24523 = n10438 & ~n20341 ;
  assign n24524 = n21244 ^ n8455 ^ 1'b0 ;
  assign n24525 = ~n1896 & n6347 ;
  assign n24526 = ~n24524 & n24525 ;
  assign n24527 = n18351 ^ n8140 ^ 1'b0 ;
  assign n24528 = n17413 ^ n1569 ^ 1'b0 ;
  assign n24529 = n24527 & n24528 ;
  assign n24530 = ( ~n3062 & n6176 ) | ( ~n3062 & n24529 ) | ( n6176 & n24529 ) ;
  assign n24531 = ( n5944 & n24526 ) | ( n5944 & ~n24530 ) | ( n24526 & ~n24530 ) ;
  assign n24532 = ( n5488 & n9052 ) | ( n5488 & n16794 ) | ( n9052 & n16794 ) ;
  assign n24533 = n22835 ^ n7169 ^ 1'b0 ;
  assign n24534 = ~n24532 & n24533 ;
  assign n24535 = n12515 | n13581 ;
  assign n24536 = n24535 ^ n12222 ^ n3474 ;
  assign n24537 = n13929 ^ n11629 ^ 1'b0 ;
  assign n24538 = n13173 & n24537 ;
  assign n24539 = n24538 ^ n7206 ^ n1839 ;
  assign n24541 = n8043 ^ n3765 ^ 1'b0 ;
  assign n24542 = ~n17010 & n17141 ;
  assign n24543 = ~n24541 & n24542 ;
  assign n24540 = n21910 ^ n19704 ^ 1'b0 ;
  assign n24544 = n24543 ^ n24540 ^ n11006 ;
  assign n24545 = ( ~n1311 & n9048 ) | ( ~n1311 & n19655 ) | ( n9048 & n19655 ) ;
  assign n24546 = n8059 ^ n327 ^ 1'b0 ;
  assign n24547 = n3337 & n24546 ;
  assign n24548 = ( n11474 & ~n17840 ) | ( n11474 & n24547 ) | ( ~n17840 & n24547 ) ;
  assign n24549 = ( n10273 & ~n13743 ) | ( n10273 & n20651 ) | ( ~n13743 & n20651 ) ;
  assign n24550 = n2108 ^ n1822 ^ 1'b0 ;
  assign n24551 = n24549 & ~n24550 ;
  assign n24552 = ~n12751 & n24551 ;
  assign n24553 = n7542 & ~n10589 ;
  assign n24554 = ~n11993 & n24553 ;
  assign n24555 = n6153 ^ n5953 ^ x48 ;
  assign n24556 = ( ~n2908 & n5295 ) | ( ~n2908 & n24555 ) | ( n5295 & n24555 ) ;
  assign n24559 = n8423 ^ n5951 ^ 1'b0 ;
  assign n24560 = n8577 & ~n24559 ;
  assign n24557 = n1698 & n13720 ;
  assign n24558 = ~n21379 & n24557 ;
  assign n24561 = n24560 ^ n24558 ^ n8413 ;
  assign n24563 = ( n18909 & n20410 ) | ( n18909 & ~n23207 ) | ( n20410 & ~n23207 ) ;
  assign n24562 = ( n5840 & ~n14873 ) | ( n5840 & n21927 ) | ( ~n14873 & n21927 ) ;
  assign n24564 = n24563 ^ n24562 ^ n12594 ;
  assign n24565 = n5809 & n11747 ;
  assign n24566 = ~n4416 & n24565 ;
  assign n24567 = ~n12521 & n24566 ;
  assign n24568 = n24567 ^ n23702 ^ n12415 ;
  assign n24569 = n7711 & ~n7827 ;
  assign n24570 = ( ~n9174 & n17225 ) | ( ~n9174 & n19274 ) | ( n17225 & n19274 ) ;
  assign n24571 = n24569 & n24570 ;
  assign n24572 = ( n17635 & n23455 ) | ( n17635 & ~n24338 ) | ( n23455 & ~n24338 ) ;
  assign n24573 = ~n13875 & n24572 ;
  assign n24574 = n3160 & n15590 ;
  assign n24575 = n10631 ^ n9570 ^ n6430 ;
  assign n24576 = ~n4879 & n24575 ;
  assign n24577 = n24576 ^ n17337 ^ 1'b0 ;
  assign n24578 = ( ~n3314 & n6825 ) | ( ~n3314 & n8222 ) | ( n6825 & n8222 ) ;
  assign n24579 = n14273 | n24578 ;
  assign n24580 = n14273 & ~n24579 ;
  assign n24581 = n4332 & ~n24580 ;
  assign n24583 = ~n4117 & n4733 ;
  assign n24584 = ~n4733 & n24583 ;
  assign n24582 = n10757 & n14093 ;
  assign n24585 = n24584 ^ n24582 ^ 1'b0 ;
  assign n24586 = ( ~n3997 & n24581 ) | ( ~n3997 & n24585 ) | ( n24581 & n24585 ) ;
  assign n24587 = n11215 | n12503 ;
  assign n24588 = n24586 | n24587 ;
  assign n24589 = n6910 ^ n1654 ^ 1'b0 ;
  assign n24590 = n15912 | n20459 ;
  assign n24591 = n24589 | n24590 ;
  assign n24592 = n13903 ^ n6321 ^ n4187 ;
  assign n24593 = n24592 ^ n7526 ^ 1'b0 ;
  assign n24594 = ~n12796 & n24593 ;
  assign n24595 = n4840 ^ n2040 ^ 1'b0 ;
  assign n24596 = n24595 ^ n3807 ^ 1'b0 ;
  assign n24597 = n11120 & n24596 ;
  assign n24598 = n24597 ^ n17980 ^ n2682 ;
  assign n24599 = n4311 ^ n3568 ^ 1'b0 ;
  assign n24600 = ( ~n832 & n5070 ) | ( ~n832 & n6370 ) | ( n5070 & n6370 ) ;
  assign n24601 = ~n24599 & n24600 ;
  assign n24602 = n8929 ^ n5205 ^ 1'b0 ;
  assign n24603 = n3174 & n24602 ;
  assign n24604 = n24603 ^ n4860 ^ 1'b0 ;
  assign n24605 = ~n8947 & n14072 ;
  assign n24606 = n9450 & n24605 ;
  assign n24607 = n24606 ^ n5026 ^ 1'b0 ;
  assign n24608 = n7802 & ~n24607 ;
  assign n24609 = n4543 & n13499 ;
  assign n24611 = n11820 ^ n5363 ^ n3629 ;
  assign n24610 = ~n5399 & n8437 ;
  assign n24612 = n24611 ^ n24610 ^ 1'b0 ;
  assign n24613 = n16555 & ~n24612 ;
  assign n24614 = n24613 ^ n19091 ^ x39 ;
  assign n24615 = ( n3033 & ~n24609 ) | ( n3033 & n24614 ) | ( ~n24609 & n24614 ) ;
  assign n24616 = x170 & ~n3633 ;
  assign n24617 = ( n321 & ~n2574 ) | ( n321 & n21275 ) | ( ~n2574 & n21275 ) ;
  assign n24618 = n8512 & ~n9997 ;
  assign n24619 = ~n11291 & n24618 ;
  assign n24620 = n24619 ^ n20797 ^ 1'b0 ;
  assign n24621 = n15806 ^ n12565 ^ 1'b0 ;
  assign n24622 = n24244 | n24621 ;
  assign n24623 = n14102 ^ n12999 ^ n11498 ;
  assign n24624 = n14436 ^ n6458 ^ n4240 ;
  assign n24625 = n24624 ^ n3754 ^ n1202 ;
  assign n24626 = n7625 | n10478 ;
  assign n24627 = n24626 ^ n2143 ^ 1'b0 ;
  assign n24628 = n24627 ^ n14336 ^ n7439 ;
  assign n24629 = n4461 & n24628 ;
  assign n24630 = n1045 | n7599 ;
  assign n24631 = n3257 | n24630 ;
  assign n24632 = ( n1857 & n24629 ) | ( n1857 & ~n24631 ) | ( n24629 & ~n24631 ) ;
  assign n24633 = n10889 ^ n1020 ^ 1'b0 ;
  assign n24634 = n24633 ^ n977 ^ x147 ;
  assign n24635 = n24634 ^ n7007 ^ 1'b0 ;
  assign n24636 = n17334 | n24635 ;
  assign n24637 = n12946 | n24636 ;
  assign n24638 = n3301 & n20858 ;
  assign n24639 = n20063 & n24638 ;
  assign n24640 = n24639 ^ n1327 ^ 1'b0 ;
  assign n24641 = ~n9646 & n24640 ;
  assign n24642 = ~n12968 & n15786 ;
  assign n24643 = n24642 ^ n8219 ^ 1'b0 ;
  assign n24644 = n24643 ^ n23605 ^ 1'b0 ;
  assign n24645 = ~n21071 & n24644 ;
  assign n24646 = ( n2160 & n5054 ) | ( n2160 & n9012 ) | ( n5054 & n9012 ) ;
  assign n24647 = n24646 ^ x230 ^ 1'b0 ;
  assign n24648 = n7369 | n22867 ;
  assign n24649 = n15962 & ~n24648 ;
  assign n24650 = ~n10284 & n24649 ;
  assign n24651 = ( ~n1537 & n3196 ) | ( ~n1537 & n16772 ) | ( n3196 & n16772 ) ;
  assign n24652 = ~n19950 & n24651 ;
  assign n24653 = n24652 ^ n2039 ^ 1'b0 ;
  assign n24654 = n24198 ^ n16915 ^ n2949 ;
  assign n24655 = n2948 | n24654 ;
  assign n24656 = n3623 | n5937 ;
  assign n24657 = n10423 | n24656 ;
  assign n24658 = ~n820 & n24657 ;
  assign n24659 = n24658 ^ n722 ^ 1'b0 ;
  assign n24660 = ~n19381 & n24659 ;
  assign n24661 = ~n3623 & n4093 ;
  assign n24662 = n5658 & n24661 ;
  assign n24663 = n24662 ^ n4499 ^ 1'b0 ;
  assign n24664 = ( n9225 & n12344 ) | ( n9225 & n24663 ) | ( n12344 & n24663 ) ;
  assign n24665 = n24664 ^ n10899 ^ n9389 ;
  assign n24666 = n8588 ^ n7403 ^ 1'b0 ;
  assign n24667 = n305 & ~n24666 ;
  assign n24668 = n6249 & ~n9298 ;
  assign n24669 = ~n5309 & n24668 ;
  assign n24670 = n19845 ^ n14041 ^ n1229 ;
  assign n24671 = n19642 ^ n6686 ^ x170 ;
  assign n24672 = n24671 ^ n16148 ^ 1'b0 ;
  assign n24673 = n12126 & n24672 ;
  assign n24674 = ( n8008 & n9188 ) | ( n8008 & n24673 ) | ( n9188 & n24673 ) ;
  assign n24675 = n21075 ^ n8735 ^ n2093 ;
  assign n24676 = n15816 ^ n13327 ^ 1'b0 ;
  assign n24677 = n5357 & n24676 ;
  assign n24678 = n290 & ~n7998 ;
  assign n24679 = ~n3200 & n4977 ;
  assign n24680 = n24679 ^ n4911 ^ 1'b0 ;
  assign n24681 = n2412 | n20754 ;
  assign n24682 = n24681 ^ n18184 ^ n7370 ;
  assign n24683 = n5259 | n7461 ;
  assign n24684 = n16937 & ~n24683 ;
  assign n24685 = ( ~n3966 & n16826 ) | ( ~n3966 & n24684 ) | ( n16826 & n24684 ) ;
  assign n24686 = n14844 ^ n13056 ^ n3245 ;
  assign n24687 = ( n18399 & n24685 ) | ( n18399 & n24686 ) | ( n24685 & n24686 ) ;
  assign n24688 = n2557 | n16594 ;
  assign n24689 = n24564 & ~n24688 ;
  assign n24690 = n2880 & ~n20591 ;
  assign n24691 = n8159 & n9146 ;
  assign n24692 = n24690 & n24691 ;
  assign n24693 = ~n11146 & n13970 ;
  assign n24694 = n24693 ^ n8861 ^ 1'b0 ;
  assign n24695 = ( n6808 & n8969 ) | ( n6808 & n9264 ) | ( n8969 & n9264 ) ;
  assign n24696 = n24694 & ~n24695 ;
  assign n24697 = n2914 | n24696 ;
  assign n24698 = n7445 | n15596 ;
  assign n24699 = ( n1542 & ~n15704 ) | ( n1542 & n24698 ) | ( ~n15704 & n24698 ) ;
  assign n24700 = n18101 ^ n5762 ^ x196 ;
  assign n24701 = n8139 ^ n361 ^ 1'b0 ;
  assign n24702 = n24700 | n24701 ;
  assign n24703 = ( ~n18231 & n21333 ) | ( ~n18231 & n24702 ) | ( n21333 & n24702 ) ;
  assign n24705 = n7959 & ~n8184 ;
  assign n24706 = ~n5070 & n24705 ;
  assign n24704 = ~n9835 & n10004 ;
  assign n24707 = n24706 ^ n24704 ^ 1'b0 ;
  assign n24708 = n24707 ^ n17719 ^ n6153 ;
  assign n24709 = n23477 | n24708 ;
  assign n24710 = n20461 ^ n11300 ^ n4732 ;
  assign n24711 = n753 | n12826 ;
  assign n24712 = n24711 ^ n5196 ^ 1'b0 ;
  assign n24713 = n5389 | n6664 ;
  assign n24714 = n24713 ^ n3605 ^ 1'b0 ;
  assign n24715 = ~n7086 & n24714 ;
  assign n24716 = n24715 ^ n8593 ^ 1'b0 ;
  assign n24717 = n24716 ^ n19813 ^ n2524 ;
  assign n24718 = n19270 & n24717 ;
  assign n24719 = n24718 ^ n2558 ^ 1'b0 ;
  assign n24720 = n5272 & ~n17762 ;
  assign n24721 = ~n24436 & n24720 ;
  assign n24722 = n10996 & n11169 ;
  assign n24725 = n15300 ^ n428 ^ x157 ;
  assign n24723 = ~n2028 & n12121 ;
  assign n24724 = ~n10561 & n24723 ;
  assign n24726 = n24725 ^ n24724 ^ n19917 ;
  assign n24729 = n3790 & n19165 ;
  assign n24727 = n12166 | n24221 ;
  assign n24728 = n24727 ^ n4091 ^ 1'b0 ;
  assign n24730 = n24729 ^ n24728 ^ 1'b0 ;
  assign n24731 = ~n18663 & n24730 ;
  assign n24732 = ~n2393 & n2685 ;
  assign n24733 = n19653 & n24732 ;
  assign n24734 = n6554 ^ n4879 ^ n1406 ;
  assign n24735 = n24734 ^ n20866 ^ n8070 ;
  assign n24739 = n9411 ^ n6523 ^ 1'b0 ;
  assign n24740 = n2263 & ~n24739 ;
  assign n24741 = n7476 ^ n4910 ^ 1'b0 ;
  assign n24742 = n24740 & ~n24741 ;
  assign n24738 = n4421 | n5528 ;
  assign n24743 = n24742 ^ n24738 ^ 1'b0 ;
  assign n24736 = n14844 ^ n13776 ^ 1'b0 ;
  assign n24737 = n20012 & n24736 ;
  assign n24744 = n24743 ^ n24737 ^ n22470 ;
  assign n24747 = n889 & n1405 ;
  assign n24748 = n24747 ^ n9067 ^ 1'b0 ;
  assign n24749 = n6876 | n24748 ;
  assign n24745 = ( n2630 & n4564 ) | ( n2630 & ~n11874 ) | ( n4564 & ~n11874 ) ;
  assign n24746 = n7565 & ~n24745 ;
  assign n24750 = n24749 ^ n24746 ^ 1'b0 ;
  assign n24751 = n24750 ^ n9543 ^ n9101 ;
  assign n24752 = n14854 & n24751 ;
  assign n24753 = n6425 ^ n3581 ^ 1'b0 ;
  assign n24754 = n24752 | n24753 ;
  assign n24755 = n14122 | n20663 ;
  assign n24756 = n3235 | n8364 ;
  assign n24757 = n4038 | n24756 ;
  assign n24758 = n24757 ^ n14715 ^ 1'b0 ;
  assign n24759 = n12491 & ~n24758 ;
  assign n24760 = n23343 ^ n2725 ^ 1'b0 ;
  assign n24761 = ( n14207 & ~n24759 ) | ( n14207 & n24760 ) | ( ~n24759 & n24760 ) ;
  assign n24762 = n2564 & ~n22879 ;
  assign n24763 = ( ~n9394 & n15670 ) | ( ~n9394 & n24762 ) | ( n15670 & n24762 ) ;
  assign n24764 = n24763 ^ n14700 ^ n8446 ;
  assign n24765 = n4006 ^ n3501 ^ 1'b0 ;
  assign n24766 = n19270 & ~n24765 ;
  assign n24769 = ( n8347 & n18441 ) | ( n8347 & n19256 ) | ( n18441 & n19256 ) ;
  assign n24767 = n14959 | n18304 ;
  assign n24768 = n24767 ^ n10415 ^ 1'b0 ;
  assign n24770 = n24769 ^ n24768 ^ 1'b0 ;
  assign n24771 = ( ~n17561 & n20809 ) | ( ~n17561 & n23004 ) | ( n20809 & n23004 ) ;
  assign n24772 = ( ~n9559 & n15469 ) | ( ~n9559 & n24771 ) | ( n15469 & n24771 ) ;
  assign n24773 = n4240 | n7101 ;
  assign n24774 = n17316 & n24773 ;
  assign n24775 = n2928 | n14804 ;
  assign n24776 = n24775 ^ n20789 ^ 1'b0 ;
  assign n24777 = n15996 & ~n24776 ;
  assign n24778 = ( ~n1047 & n2232 ) | ( ~n1047 & n3315 ) | ( n2232 & n3315 ) ;
  assign n24779 = ( n5751 & n19770 ) | ( n5751 & ~n24778 ) | ( n19770 & ~n24778 ) ;
  assign n24780 = n6018 | n20766 ;
  assign n24781 = n11330 & ~n24780 ;
  assign n24785 = ( n5315 & ~n10702 ) | ( n5315 & n15631 ) | ( ~n10702 & n15631 ) ;
  assign n24786 = n10794 ^ n1132 ^ 1'b0 ;
  assign n24787 = ~n24785 & n24786 ;
  assign n24788 = ~n19117 & n24787 ;
  assign n24789 = n22441 & n24788 ;
  assign n24783 = n5834 | n11956 ;
  assign n24784 = n7729 & ~n24783 ;
  assign n24782 = ( n15915 & ~n18634 ) | ( n15915 & n21642 ) | ( ~n18634 & n21642 ) ;
  assign n24790 = n24789 ^ n24784 ^ n24782 ;
  assign n24791 = ~n24781 & n24790 ;
  assign n24792 = n10128 ^ n8397 ^ 1'b0 ;
  assign n24793 = ( x104 & n4959 ) | ( x104 & n6556 ) | ( n4959 & n6556 ) ;
  assign n24794 = ( n23242 & ~n24792 ) | ( n23242 & n24793 ) | ( ~n24792 & n24793 ) ;
  assign n24795 = n13792 & n14883 ;
  assign n24796 = ( ~n18085 & n19851 ) | ( ~n18085 & n24795 ) | ( n19851 & n24795 ) ;
  assign n24797 = n12999 ^ n4266 ^ 1'b0 ;
  assign n24798 = ( ~n12873 & n13546 ) | ( ~n12873 & n24797 ) | ( n13546 & n24797 ) ;
  assign n24799 = n11609 | n13945 ;
  assign n24800 = n18385 & ~n24799 ;
  assign n24801 = n4526 ^ n3569 ^ 1'b0 ;
  assign n24802 = n17427 | n24801 ;
  assign n24803 = n4469 & ~n24802 ;
  assign n24804 = n10480 & n10509 ;
  assign n24805 = n24804 ^ n1484 ^ 1'b0 ;
  assign n24806 = n20794 & ~n24805 ;
  assign n24807 = n1687 & n2402 ;
  assign n24808 = n5048 & ~n19660 ;
  assign n24809 = ~n2764 & n24808 ;
  assign n24810 = ( n6629 & n24807 ) | ( n6629 & n24809 ) | ( n24807 & n24809 ) ;
  assign n24811 = n15334 ^ n14486 ^ n13423 ;
  assign n24812 = ~n11921 & n16375 ;
  assign n24813 = ~n10177 & n24812 ;
  assign n24814 = n2363 ^ n1309 ^ 1'b0 ;
  assign n24815 = n9903 | n24814 ;
  assign n24816 = n16760 & ~n24815 ;
  assign n24817 = n983 ^ n636 ^ 1'b0 ;
  assign n24818 = n1574 & ~n24817 ;
  assign n24819 = n24818 ^ n11999 ^ 1'b0 ;
  assign n24820 = n17226 | n24819 ;
  assign n24821 = n24816 & ~n24820 ;
  assign n24822 = n1667 & ~n17375 ;
  assign n24823 = ~n19708 & n24822 ;
  assign n24824 = n24823 ^ n17589 ^ n9317 ;
  assign n24825 = ( n1047 & ~n5982 ) | ( n1047 & n7510 ) | ( ~n5982 & n7510 ) ;
  assign n24826 = n16978 | n24825 ;
  assign n24827 = n23626 ^ n16906 ^ 1'b0 ;
  assign n24828 = n24826 & ~n24827 ;
  assign n24829 = n24828 ^ x171 ^ 1'b0 ;
  assign n24830 = n10562 ^ n4530 ^ n1159 ;
  assign n24831 = n22460 ^ n3016 ^ 1'b0 ;
  assign n24832 = n12278 ^ n2211 ^ n2128 ;
  assign n24833 = n24832 ^ n23988 ^ n9451 ;
  assign n24834 = n24833 ^ n12124 ^ 1'b0 ;
  assign n24835 = n4794 | n24834 ;
  assign n24836 = n1704 | n11811 ;
  assign n24837 = n24836 ^ n17049 ^ 1'b0 ;
  assign n24838 = n7935 ^ n5635 ^ 1'b0 ;
  assign n24839 = n24837 & n24838 ;
  assign n24840 = n24839 ^ n1924 ^ 1'b0 ;
  assign n24841 = n10777 ^ n1649 ^ 1'b0 ;
  assign n24842 = n4124 & n20855 ;
  assign n24843 = n4067 & ~n12924 ;
  assign n24844 = n12155 & n24843 ;
  assign n24845 = n17455 & ~n24844 ;
  assign n24846 = n24845 ^ n14639 ^ 1'b0 ;
  assign n24847 = ( n24841 & n24842 ) | ( n24841 & n24846 ) | ( n24842 & n24846 ) ;
  assign n24848 = n4935 | n9430 ;
  assign n24849 = n24848 ^ n6851 ^ n776 ;
  assign n24850 = n14052 ^ n6911 ^ 1'b0 ;
  assign n24851 = n24850 ^ n7280 ^ 1'b0 ;
  assign n24852 = n24851 ^ n16453 ^ 1'b0 ;
  assign n24853 = n4588 ^ n1588 ^ 1'b0 ;
  assign n24854 = n21476 | n24853 ;
  assign n24855 = n24852 | n24854 ;
  assign n24856 = n4237 | n10808 ;
  assign n24857 = n1813 | n24856 ;
  assign n24858 = n3038 & n24857 ;
  assign n24859 = ~n11860 & n24858 ;
  assign n24860 = n22395 & ~n24859 ;
  assign n24861 = n3696 & ~n16673 ;
  assign n24862 = n12886 | n24861 ;
  assign n24863 = ( n2509 & ~n13585 ) | ( n2509 & n19604 ) | ( ~n13585 & n19604 ) ;
  assign n24864 = n11134 | n13616 ;
  assign n24865 = n24864 ^ n18466 ^ 1'b0 ;
  assign n24866 = n12551 & n24865 ;
  assign n24867 = n14701 & n24866 ;
  assign n24868 = n4208 ^ n3048 ^ 1'b0 ;
  assign n24869 = n24868 ^ n310 ^ 1'b0 ;
  assign n24870 = ~n820 & n24869 ;
  assign n24871 = n20355 ^ n13020 ^ n10862 ;
  assign n24872 = n23194 ^ n15975 ^ n11298 ;
  assign n24873 = n13970 ^ n1496 ^ 1'b0 ;
  assign n24874 = n21908 | n24873 ;
  assign n24879 = n5877 | n13506 ;
  assign n24880 = n24466 & ~n24879 ;
  assign n24881 = n24880 ^ n16997 ^ n10799 ;
  assign n24875 = ~n6432 & n7243 ;
  assign n24876 = n24875 ^ n11339 ^ 1'b0 ;
  assign n24877 = n24876 ^ n5100 ^ 1'b0 ;
  assign n24878 = n12032 & ~n24877 ;
  assign n24882 = n24881 ^ n24878 ^ 1'b0 ;
  assign n24883 = n21500 ^ n15451 ^ n6428 ;
  assign n24884 = ( n10549 & n19436 ) | ( n10549 & n24883 ) | ( n19436 & n24883 ) ;
  assign n24885 = ( ~n617 & n6705 ) | ( ~n617 & n24884 ) | ( n6705 & n24884 ) ;
  assign n24886 = n7452 ^ n284 ^ 1'b0 ;
  assign n24887 = ~n19530 & n24886 ;
  assign n24889 = n21984 ^ n9690 ^ n5931 ;
  assign n24888 = n15456 | n16654 ;
  assign n24890 = n24889 ^ n24888 ^ 1'b0 ;
  assign n24891 = ( n1484 & n24887 ) | ( n1484 & n24890 ) | ( n24887 & n24890 ) ;
  assign n24892 = n5081 | n15985 ;
  assign n24893 = n24892 ^ n7211 ^ 1'b0 ;
  assign n24894 = n15838 ^ n7213 ^ n6076 ;
  assign n24895 = ( x167 & ~n15860 ) | ( x167 & n24894 ) | ( ~n15860 & n24894 ) ;
  assign n24896 = ~n19814 & n24895 ;
  assign n24897 = ~n24893 & n24896 ;
  assign n24898 = n4550 | n24897 ;
  assign n24899 = n19483 | n24898 ;
  assign n24900 = n2039 | n4555 ;
  assign n24901 = n24900 ^ n23573 ^ n17505 ;
  assign n24902 = n19947 ^ n941 ^ 1'b0 ;
  assign n24905 = n12121 & n15292 ;
  assign n24906 = ~n11287 & n24905 ;
  assign n24903 = ( x187 & n9794 ) | ( x187 & n15353 ) | ( n9794 & n15353 ) ;
  assign n24904 = n24425 & ~n24903 ;
  assign n24907 = n24906 ^ n24904 ^ 1'b0 ;
  assign n24908 = n10953 | n24907 ;
  assign n24909 = n4601 | n24908 ;
  assign n24910 = n11044 & ~n16156 ;
  assign n24911 = n24909 & n24910 ;
  assign n24912 = n1950 & n21633 ;
  assign n24913 = n6176 & n24912 ;
  assign n24914 = n24913 ^ n18622 ^ n7028 ;
  assign n24915 = n14833 ^ n8243 ^ n8110 ;
  assign n24916 = ( n3214 & n22519 ) | ( n3214 & ~n22742 ) | ( n22519 & ~n22742 ) ;
  assign n24917 = ( n10939 & n21029 ) | ( n10939 & n24916 ) | ( n21029 & n24916 ) ;
  assign n24918 = n24915 & n24917 ;
  assign n24921 = n6091 ^ n482 ^ 1'b0 ;
  assign n24922 = n21644 & ~n24921 ;
  assign n24923 = n8704 & n24922 ;
  assign n24924 = n24923 ^ n8518 ^ 1'b0 ;
  assign n24919 = n10513 & ~n13308 ;
  assign n24920 = n16161 | n24919 ;
  assign n24925 = n24924 ^ n24920 ^ 1'b0 ;
  assign n24926 = n6520 | n10961 ;
  assign n24927 = ~n10000 & n21265 ;
  assign n24929 = n7988 | n19973 ;
  assign n24930 = n24929 ^ n11272 ^ 1'b0 ;
  assign n24931 = n17325 & ~n24930 ;
  assign n24928 = ( n758 & n15017 ) | ( n758 & n18734 ) | ( n15017 & n18734 ) ;
  assign n24932 = n24931 ^ n24928 ^ 1'b0 ;
  assign n24933 = ~n24927 & n24932 ;
  assign n24934 = n1067 | n6868 ;
  assign n24935 = n24934 ^ n13569 ^ 1'b0 ;
  assign n24936 = n2231 & n15843 ;
  assign n24937 = ~n14240 & n24936 ;
  assign n24938 = n24937 ^ n13925 ^ n9845 ;
  assign n24939 = ( ~n8029 & n14489 ) | ( ~n8029 & n24938 ) | ( n14489 & n24938 ) ;
  assign n24940 = n1585 & n14467 ;
  assign n24941 = n2666 & n4304 ;
  assign n24942 = n24941 ^ n1442 ^ 1'b0 ;
  assign n24943 = ~n7920 & n24942 ;
  assign n24944 = n5531 ^ n1985 ^ 1'b0 ;
  assign n24945 = n318 | n24944 ;
  assign n24946 = ( ~n14008 & n14916 ) | ( ~n14008 & n17761 ) | ( n14916 & n17761 ) ;
  assign n24947 = ( ~n954 & n13857 ) | ( ~n954 & n15455 ) | ( n13857 & n15455 ) ;
  assign n24949 = ~n3032 & n13316 ;
  assign n24950 = ( ~n4724 & n18143 ) | ( ~n4724 & n24949 ) | ( n18143 & n24949 ) ;
  assign n24948 = n11580 ^ n4906 ^ n3106 ;
  assign n24951 = n24950 ^ n24948 ^ n12411 ;
  assign n24952 = n18291 ^ n14395 ^ 1'b0 ;
  assign n24953 = ~n10710 & n17768 ;
  assign n24954 = ~n24952 & n24953 ;
  assign n24955 = ~n3279 & n5372 ;
  assign n24959 = ( ~x7 & n894 ) | ( ~x7 & n7655 ) | ( n894 & n7655 ) ;
  assign n24960 = n4325 | n9872 ;
  assign n24961 = n10967 | n24960 ;
  assign n24962 = ( n10566 & ~n24959 ) | ( n10566 & n24961 ) | ( ~n24959 & n24961 ) ;
  assign n24956 = n14298 ^ n12295 ^ 1'b0 ;
  assign n24957 = ~n24785 & n24956 ;
  assign n24958 = n24957 ^ n3498 ^ 1'b0 ;
  assign n24963 = n24962 ^ n24958 ^ n18338 ;
  assign n24964 = n14141 & ~n24963 ;
  assign n24965 = n24955 & n24964 ;
  assign n24966 = ( n1787 & ~n9710 ) | ( n1787 & n16114 ) | ( ~n9710 & n16114 ) ;
  assign n24967 = ( n7633 & n15333 ) | ( n7633 & n21594 ) | ( n15333 & n21594 ) ;
  assign n24968 = n8390 ^ n3857 ^ n1739 ;
  assign n24969 = n24968 ^ n3161 ^ 1'b0 ;
  assign n24970 = x187 & n20448 ;
  assign n24971 = ~n1374 & n6466 ;
  assign n24972 = n24971 ^ n22495 ^ 1'b0 ;
  assign n24973 = n22293 & n24972 ;
  assign n24974 = n24973 ^ n24924 ^ n12220 ;
  assign n24975 = ( n681 & n11683 ) | ( n681 & n14602 ) | ( n11683 & n14602 ) ;
  assign n24976 = n10727 & ~n24975 ;
  assign n24978 = n2567 | n4430 ;
  assign n24979 = n668 | n24978 ;
  assign n24980 = n24979 ^ n5399 ^ n3042 ;
  assign n24977 = n1098 | n8525 ;
  assign n24981 = n24980 ^ n24977 ^ 1'b0 ;
  assign n24982 = n1938 ^ n1891 ^ 1'b0 ;
  assign n24986 = ~n987 & n10786 ;
  assign n24983 = n1480 & n4286 ;
  assign n24984 = n18841 & ~n24983 ;
  assign n24985 = n24984 ^ n4101 ^ 1'b0 ;
  assign n24987 = n24986 ^ n24985 ^ 1'b0 ;
  assign n24988 = n24982 | n24987 ;
  assign n24990 = ( ~n1331 & n11307 ) | ( ~n1331 & n13749 ) | ( n11307 & n13749 ) ;
  assign n24991 = n1475 & n24990 ;
  assign n24992 = n24991 ^ n12984 ^ 1'b0 ;
  assign n24993 = n24992 ^ n7944 ^ 1'b0 ;
  assign n24989 = n2682 ^ n2457 ^ n397 ;
  assign n24994 = n24993 ^ n24989 ^ n20822 ;
  assign n24995 = n4060 ^ n1930 ^ 1'b0 ;
  assign n24996 = ( n2280 & n16314 ) | ( n2280 & n24995 ) | ( n16314 & n24995 ) ;
  assign n25002 = n17058 ^ n2796 ^ 1'b0 ;
  assign n25000 = ( ~n496 & n7084 ) | ( ~n496 & n10669 ) | ( n7084 & n10669 ) ;
  assign n24997 = n20123 ^ n2613 ^ 1'b0 ;
  assign n24998 = n24997 ^ n13539 ^ 1'b0 ;
  assign n24999 = n4942 | n24998 ;
  assign n25001 = n25000 ^ n24999 ^ n2321 ;
  assign n25003 = n25002 ^ n25001 ^ n3184 ;
  assign n25004 = n25003 ^ n9151 ^ n7877 ;
  assign n25005 = n3571 | n18990 ;
  assign n25006 = n25005 ^ n4788 ^ 1'b0 ;
  assign n25007 = n9002 & ~n25006 ;
  assign n25008 = ~n7515 & n25007 ;
  assign n25009 = n7913 ^ n756 ^ 1'b0 ;
  assign n25010 = ( n642 & ~n8442 ) | ( n642 & n11501 ) | ( ~n8442 & n11501 ) ;
  assign n25011 = n25010 ^ n12607 ^ 1'b0 ;
  assign n25012 = n25011 ^ n7458 ^ 1'b0 ;
  assign n25013 = n6959 & n25012 ;
  assign n25014 = n13830 ^ n4813 ^ 1'b0 ;
  assign n25015 = ~n20115 & n25014 ;
  assign n25018 = n10351 & n10973 ;
  assign n25019 = n5141 | n25018 ;
  assign n25020 = n25019 ^ n8068 ^ 1'b0 ;
  assign n25016 = n16720 ^ n8975 ^ 1'b0 ;
  assign n25017 = n18429 & ~n25016 ;
  assign n25021 = n25020 ^ n25017 ^ 1'b0 ;
  assign n25022 = ~n12729 & n22340 ;
  assign n25023 = ~n25021 & n25022 ;
  assign n25024 = ~n11849 & n11898 ;
  assign n25025 = n25024 ^ n18434 ^ 1'b0 ;
  assign n25026 = n1268 | n3003 ;
  assign n25027 = n25025 | n25026 ;
  assign n25028 = n24185 | n25027 ;
  assign n25029 = n9276 | n17336 ;
  assign n25033 = n1173 ^ n1164 ^ n895 ;
  assign n25030 = n13535 ^ n7818 ^ n734 ;
  assign n25031 = n6979 ^ n5805 ^ 1'b0 ;
  assign n25032 = n25030 & n25031 ;
  assign n25034 = n25033 ^ n25032 ^ n8743 ;
  assign n25035 = ~n9469 & n25034 ;
  assign n25036 = n25035 ^ n17924 ^ 1'b0 ;
  assign n25037 = n614 & n17381 ;
  assign n25038 = n25037 ^ n24288 ^ 1'b0 ;
  assign n25039 = n2231 & ~n3699 ;
  assign n25040 = n749 & ~n4838 ;
  assign n25041 = n21233 & n25040 ;
  assign n25044 = n14790 ^ n10714 ^ n1589 ;
  assign n25045 = ~n12673 & n25044 ;
  assign n25042 = n2444 ^ n1374 ^ 1'b0 ;
  assign n25043 = n7177 & ~n25042 ;
  assign n25046 = n25045 ^ n25043 ^ n10706 ;
  assign n25047 = n24414 ^ n21932 ^ n7350 ;
  assign n25049 = ~n2293 & n24657 ;
  assign n25050 = n25049 ^ n1363 ^ 1'b0 ;
  assign n25048 = ~n11930 & n15634 ;
  assign n25051 = n25050 ^ n25048 ^ 1'b0 ;
  assign n25052 = n22259 ^ n19773 ^ n10189 ;
  assign n25053 = ( n732 & n5160 ) | ( n732 & n5840 ) | ( n5160 & n5840 ) ;
  assign n25054 = n2368 & n3725 ;
  assign n25055 = n12525 ^ n3805 ^ 1'b0 ;
  assign n25056 = n22388 ^ n15187 ^ 1'b0 ;
  assign n25057 = n9628 ^ n8142 ^ n3476 ;
  assign n25058 = ~n1150 & n1928 ;
  assign n25059 = n4278 & ~n6523 ;
  assign n25060 = n19476 & n25059 ;
  assign n25061 = ( ~n5620 & n25058 ) | ( ~n5620 & n25060 ) | ( n25058 & n25060 ) ;
  assign n25062 = n25057 | n25061 ;
  assign n25065 = ~n6476 & n22692 ;
  assign n25063 = n7916 ^ n1511 ^ 1'b0 ;
  assign n25064 = n25063 ^ n7123 ^ 1'b0 ;
  assign n25066 = n25065 ^ n25064 ^ n8008 ;
  assign n25067 = n22765 ^ n17297 ^ n2066 ;
  assign n25068 = n7213 & ~n7900 ;
  assign n25069 = ~n24206 & n25068 ;
  assign n25072 = n2113 & ~n11849 ;
  assign n25073 = n25072 ^ n6847 ^ 1'b0 ;
  assign n25070 = n14906 ^ n9451 ^ n2026 ;
  assign n25071 = ( n14297 & n16527 ) | ( n14297 & n25070 ) | ( n16527 & n25070 ) ;
  assign n25074 = n25073 ^ n25071 ^ 1'b0 ;
  assign n25075 = n25074 ^ n24603 ^ n12348 ;
  assign n25076 = n25075 ^ n11061 ^ 1'b0 ;
  assign n25077 = n25069 | n25076 ;
  assign n25078 = n4620 & ~n11197 ;
  assign n25079 = ( ~n5141 & n7325 ) | ( ~n5141 & n25078 ) | ( n7325 & n25078 ) ;
  assign n25080 = n15786 & n25079 ;
  assign n25081 = n25080 ^ n8854 ^ 1'b0 ;
  assign n25082 = n1279 | n9024 ;
  assign n25083 = x126 & ~n1369 ;
  assign n25084 = ~n1907 & n25083 ;
  assign n25085 = n10090 | n25084 ;
  assign n25086 = ~n9594 & n10137 ;
  assign n25087 = n18537 ^ n11212 ^ 1'b0 ;
  assign n25088 = ( n4017 & n6793 ) | ( n4017 & n9769 ) | ( n6793 & n9769 ) ;
  assign n25089 = n11946 & ~n16914 ;
  assign n25090 = ( n7061 & n19000 ) | ( n7061 & ~n25089 ) | ( n19000 & ~n25089 ) ;
  assign n25091 = ~n20977 & n22075 ;
  assign n25092 = n12626 | n25091 ;
  assign n25093 = ~n25090 & n25092 ;
  assign n25094 = n11013 ^ n7085 ^ n4629 ;
  assign n25095 = ~n12387 & n25094 ;
  assign n25096 = n4434 & n23040 ;
  assign n25097 = n23451 ^ n18829 ^ 1'b0 ;
  assign n25098 = n25096 & ~n25097 ;
  assign n25099 = n25098 ^ n18523 ^ 1'b0 ;
  assign n25100 = n12480 ^ n5470 ^ n1212 ;
  assign n25103 = ~n1591 & n5439 ;
  assign n25104 = n25103 ^ n7892 ^ 1'b0 ;
  assign n25102 = n9113 ^ n8203 ^ n5781 ;
  assign n25105 = n25104 ^ n25102 ^ n5701 ;
  assign n25101 = n9341 & ~n20482 ;
  assign n25106 = n25105 ^ n25101 ^ 1'b0 ;
  assign n25107 = n24044 ^ n23607 ^ 1'b0 ;
  assign n25108 = n3611 | n10608 ;
  assign n25109 = n25108 ^ n19893 ^ 1'b0 ;
  assign n25110 = n11414 & n25109 ;
  assign n25111 = n1478 & ~n2406 ;
  assign n25112 = n25111 ^ n3377 ^ 1'b0 ;
  assign n25113 = ( n2430 & n3389 ) | ( n2430 & ~n9693 ) | ( n3389 & ~n9693 ) ;
  assign n25114 = ( n350 & n875 ) | ( n350 & n25113 ) | ( n875 & n25113 ) ;
  assign n25115 = n25112 | n25114 ;
  assign n25116 = n20169 | n25115 ;
  assign n25117 = n25116 ^ n6901 ^ 1'b0 ;
  assign n25118 = ( ~n4016 & n17181 ) | ( ~n4016 & n19478 ) | ( n17181 & n19478 ) ;
  assign n25119 = n1527 & n8194 ;
  assign n25120 = ~n16195 & n19773 ;
  assign n25121 = ( n8447 & n12988 ) | ( n8447 & n14415 ) | ( n12988 & n14415 ) ;
  assign n25122 = n25121 ^ n9690 ^ 1'b0 ;
  assign n25123 = n25120 | n25122 ;
  assign n25124 = ~n19076 & n23906 ;
  assign n25125 = ( n6545 & n22202 ) | ( n6545 & n23841 ) | ( n22202 & n23841 ) ;
  assign n25126 = n25125 ^ n24819 ^ n4429 ;
  assign n25127 = n18282 ^ n10907 ^ n3794 ;
  assign n25128 = n23575 ^ n10186 ^ 1'b0 ;
  assign n25129 = n25127 & n25128 ;
  assign n25130 = n25129 ^ n20888 ^ n8375 ;
  assign n25131 = n10819 | n25130 ;
  assign n25132 = n2725 | n25131 ;
  assign n25137 = n8851 | n9907 ;
  assign n25138 = n4026 | n25137 ;
  assign n25133 = n2343 & n13534 ;
  assign n25134 = n7490 & n25133 ;
  assign n25135 = n25134 ^ n2892 ^ n1448 ;
  assign n25136 = n25135 ^ n21766 ^ n10477 ;
  assign n25139 = n25138 ^ n25136 ^ n16755 ;
  assign n25140 = n10105 ^ n4027 ^ 1'b0 ;
  assign n25141 = n25139 | n25140 ;
  assign n25148 = n10546 ^ n939 ^ 1'b0 ;
  assign n25147 = ( n6859 & n8387 ) | ( n6859 & n16466 ) | ( n8387 & n16466 ) ;
  assign n25143 = n21074 ^ n12611 ^ n8068 ;
  assign n25142 = n18812 & ~n21642 ;
  assign n25144 = n25143 ^ n25142 ^ 1'b0 ;
  assign n25145 = n25144 ^ n18666 ^ 1'b0 ;
  assign n25146 = ~n14694 & n25145 ;
  assign n25149 = n25148 ^ n25147 ^ n25146 ;
  assign n25150 = n2843 | n4801 ;
  assign n25151 = n18287 & ~n25150 ;
  assign n25152 = n25151 ^ n24235 ^ 1'b0 ;
  assign n25153 = n10659 | n11100 ;
  assign n25163 = n7067 ^ n1864 ^ 1'b0 ;
  assign n25154 = n378 & n2231 ;
  assign n25155 = n25154 ^ n6893 ^ 1'b0 ;
  assign n25156 = ~n7148 & n25155 ;
  assign n25157 = n25156 ^ n5376 ^ 1'b0 ;
  assign n25158 = n17565 & ~n25157 ;
  assign n25159 = n7131 & n14012 ;
  assign n25160 = ~n2865 & n25159 ;
  assign n25161 = n25158 & ~n25160 ;
  assign n25162 = n3598 & n25161 ;
  assign n25164 = n25163 ^ n25162 ^ 1'b0 ;
  assign n25165 = n17573 ^ n14290 ^ 1'b0 ;
  assign n25166 = n25165 ^ n8236 ^ 1'b0 ;
  assign n25167 = ~n3854 & n25166 ;
  assign n25168 = n25167 ^ n18394 ^ n7500 ;
  assign n25177 = ~n1192 & n4506 ;
  assign n25178 = n25177 ^ n2532 ^ 1'b0 ;
  assign n25179 = n25178 ^ n13851 ^ 1'b0 ;
  assign n25180 = ~n3656 & n25179 ;
  assign n25181 = n8122 & ~n25180 ;
  assign n25169 = n2151 & n3175 ;
  assign n25170 = n25169 ^ n4954 ^ n1906 ;
  assign n25174 = n9264 ^ n7751 ^ n3716 ;
  assign n25171 = n20376 ^ n7867 ^ 1'b0 ;
  assign n25172 = n6587 & ~n25171 ;
  assign n25173 = n25172 ^ n6625 ^ 1'b0 ;
  assign n25175 = n25174 ^ n25173 ^ n18289 ;
  assign n25176 = ( n11157 & n25170 ) | ( n11157 & n25175 ) | ( n25170 & n25175 ) ;
  assign n25182 = n25181 ^ n25176 ^ n2763 ;
  assign n25184 = n9644 & ~n24611 ;
  assign n25183 = n10426 ^ n3409 ^ n1360 ;
  assign n25185 = n25184 ^ n25183 ^ n23268 ;
  assign n25186 = ( ~n6362 & n12234 ) | ( ~n6362 & n25185 ) | ( n12234 & n25185 ) ;
  assign n25187 = n4384 & ~n8234 ;
  assign n25188 = n5530 ^ n5516 ^ n932 ;
  assign n25189 = n25188 ^ n24138 ^ n277 ;
  assign n25190 = x170 | n10682 ;
  assign n25191 = n25190 ^ n20759 ^ n4153 ;
  assign n25192 = ~n11883 & n18127 ;
  assign n25193 = ~n16903 & n25192 ;
  assign n25194 = n1608 | n24377 ;
  assign n25195 = n11762 ^ n10110 ^ n1097 ;
  assign n25196 = n25195 ^ n9110 ^ 1'b0 ;
  assign n25197 = n3030 & ~n13657 ;
  assign n25198 = n22182 ^ n17921 ^ n9881 ;
  assign n25204 = n7194 ^ n1042 ^ 1'b0 ;
  assign n25205 = ( n12824 & n14064 ) | ( n12824 & n25204 ) | ( n14064 & n25204 ) ;
  assign n25199 = n25184 ^ n9540 ^ 1'b0 ;
  assign n25200 = ~n7306 & n25199 ;
  assign n25201 = n779 & n25200 ;
  assign n25202 = n25201 ^ n14708 ^ 1'b0 ;
  assign n25203 = n13994 & n25202 ;
  assign n25206 = n25205 ^ n25203 ^ n4363 ;
  assign n25207 = ( n3553 & n14789 ) | ( n3553 & n23417 ) | ( n14789 & n23417 ) ;
  assign n25208 = n8997 & n25207 ;
  assign n25209 = n4003 & n25208 ;
  assign n25210 = n25209 ^ n16720 ^ 1'b0 ;
  assign n25211 = n8394 & ~n8539 ;
  assign n25212 = n25211 ^ n10994 ^ 1'b0 ;
  assign n25213 = n16647 ^ n11534 ^ n4328 ;
  assign n25214 = n11872 ^ n6809 ^ 1'b0 ;
  assign n25215 = n15526 & n25214 ;
  assign n25216 = n25215 ^ n20270 ^ n8296 ;
  assign n25217 = n7547 ^ n5542 ^ n3021 ;
  assign n25218 = n22959 ^ n9501 ^ n7139 ;
  assign n25219 = ~n5826 & n25218 ;
  assign n25220 = ( n316 & n3910 ) | ( n316 & ~n20312 ) | ( n3910 & ~n20312 ) ;
  assign n25221 = n9771 & ~n15763 ;
  assign n25222 = ( ~n4323 & n8836 ) | ( ~n4323 & n10477 ) | ( n8836 & n10477 ) ;
  assign n25223 = n25222 ^ n6333 ^ 1'b0 ;
  assign n25224 = ( n10248 & ~n12070 ) | ( n10248 & n19473 ) | ( ~n12070 & n19473 ) ;
  assign n25227 = n21728 ^ n12651 ^ 1'b0 ;
  assign n25228 = n8497 & n25227 ;
  assign n25225 = ~n5155 & n8519 ;
  assign n25226 = n25225 ^ n18901 ^ n11978 ;
  assign n25229 = n25228 ^ n25226 ^ 1'b0 ;
  assign n25230 = n25229 ^ x248 ^ 1'b0 ;
  assign n25231 = n12739 & n25230 ;
  assign n25232 = n1363 | n13317 ;
  assign n25234 = ~n5638 & n20951 ;
  assign n25235 = n1943 & n25234 ;
  assign n25236 = n25235 ^ n12326 ^ 1'b0 ;
  assign n25233 = n20814 | n22328 ;
  assign n25237 = n25236 ^ n25233 ^ 1'b0 ;
  assign n25238 = n18550 ^ n2710 ^ 1'b0 ;
  assign n25239 = n11370 & n25238 ;
  assign n25240 = n25239 ^ n20719 ^ 1'b0 ;
  assign n25241 = n5624 ^ n5574 ^ 1'b0 ;
  assign n25242 = n17118 ^ n4876 ^ 1'b0 ;
  assign n25243 = n25242 ^ n10753 ^ 1'b0 ;
  assign n25244 = n25243 ^ n7551 ^ n4316 ;
  assign n25245 = n8345 & n17423 ;
  assign n25246 = ~n6071 & n25245 ;
  assign n25247 = ~n4132 & n12687 ;
  assign n25248 = n22767 | n25247 ;
  assign n25249 = ( n3803 & ~n9009 ) | ( n3803 & n9193 ) | ( ~n9009 & n9193 ) ;
  assign n25250 = n14007 ^ n9668 ^ 1'b0 ;
  assign n25251 = n3336 & n25250 ;
  assign n25252 = ( n8644 & ~n25249 ) | ( n8644 & n25251 ) | ( ~n25249 & n25251 ) ;
  assign n25253 = n15036 & n25252 ;
  assign n25254 = n18082 & n25253 ;
  assign n25255 = n1108 | n22792 ;
  assign n25256 = ( n1827 & n5343 ) | ( n1827 & ~n7164 ) | ( n5343 & ~n7164 ) ;
  assign n25257 = n25256 ^ n4390 ^ 1'b0 ;
  assign n25258 = ( n8869 & ~n9119 ) | ( n8869 & n13731 ) | ( ~n9119 & n13731 ) ;
  assign n25259 = n25258 ^ n268 ^ 1'b0 ;
  assign n25260 = ( n8398 & n25257 ) | ( n8398 & n25259 ) | ( n25257 & n25259 ) ;
  assign n25261 = x8 & n393 ;
  assign n25262 = n4706 ^ n2692 ^ 1'b0 ;
  assign n25263 = n25261 | n25262 ;
  assign n25264 = ~n5724 & n5851 ;
  assign n25265 = ~n5851 & n25264 ;
  assign n25266 = n5250 & ~n25265 ;
  assign n25267 = n23430 ^ n2518 ^ 1'b0 ;
  assign n25268 = x164 & ~n25267 ;
  assign n25269 = ~n3583 & n25268 ;
  assign n25270 = n25269 ^ n21273 ^ 1'b0 ;
  assign n25271 = ~n25266 & n25270 ;
  assign n25272 = n25271 ^ n24398 ^ 1'b0 ;
  assign n25273 = n4343 | n14267 ;
  assign n25274 = n3980 | n25273 ;
  assign n25275 = n25274 ^ n4177 ^ n340 ;
  assign n25276 = n23711 ^ n22867 ^ n9499 ;
  assign n25277 = n21042 & n25276 ;
  assign n25278 = n25277 ^ n20911 ^ 1'b0 ;
  assign n25279 = ( n5597 & n25275 ) | ( n5597 & ~n25278 ) | ( n25275 & ~n25278 ) ;
  assign n25280 = n22053 ^ n17084 ^ n16548 ;
  assign n25281 = ~n580 & n8162 ;
  assign n25282 = n24295 & ~n25281 ;
  assign n25283 = n10141 | n16085 ;
  assign n25284 = n21096 | n25283 ;
  assign n25285 = n25284 ^ n17810 ^ 1'b0 ;
  assign n25286 = n14132 | n25285 ;
  assign n25287 = n19911 ^ n4040 ^ 1'b0 ;
  assign n25288 = ( n3016 & ~n5321 ) | ( n3016 & n25287 ) | ( ~n5321 & n25287 ) ;
  assign n25289 = ( ~n6697 & n12207 ) | ( ~n6697 & n14973 ) | ( n12207 & n14973 ) ;
  assign n25290 = n17287 | n22051 ;
  assign n25291 = n7883 & ~n25290 ;
  assign n25292 = ~n13049 & n18649 ;
  assign n25294 = n12993 ^ n9268 ^ 1'b0 ;
  assign n25295 = n1179 & n25294 ;
  assign n25293 = ( ~n3875 & n17077 ) | ( ~n3875 & n18793 ) | ( n17077 & n18793 ) ;
  assign n25296 = n25295 ^ n25293 ^ 1'b0 ;
  assign n25297 = ( n8695 & ~n11104 ) | ( n8695 & n25296 ) | ( ~n11104 & n25296 ) ;
  assign n25298 = n9700 & n23462 ;
  assign n25299 = n5293 & ~n8600 ;
  assign n25300 = n16031 & n25299 ;
  assign n25301 = n5271 & ~n11230 ;
  assign n25302 = ( ~n3520 & n25300 ) | ( ~n3520 & n25301 ) | ( n25300 & n25301 ) ;
  assign n25303 = n25302 ^ n10621 ^ 1'b0 ;
  assign n25304 = ~n1889 & n8614 ;
  assign n25305 = n12685 | n25304 ;
  assign n25306 = ~n6862 & n25305 ;
  assign n25307 = n10873 ^ n5484 ^ n591 ;
  assign n25308 = n15821 | n25307 ;
  assign n25309 = n25308 ^ n6055 ^ 1'b0 ;
  assign n25310 = ~n3775 & n23073 ;
  assign n25311 = n10797 & n25310 ;
  assign n25312 = ( ~n404 & n7375 ) | ( ~n404 & n7903 ) | ( n7375 & n7903 ) ;
  assign n25313 = ~n3115 & n13080 ;
  assign n25314 = ( n2502 & n13981 ) | ( n2502 & n25313 ) | ( n13981 & n25313 ) ;
  assign n25315 = n3170 ^ n1409 ^ 1'b0 ;
  assign n25316 = n7980 & n25315 ;
  assign n25317 = n25316 ^ n1277 ^ 1'b0 ;
  assign n25318 = ~n22796 & n25317 ;
  assign n25319 = ( ~n10456 & n25314 ) | ( ~n10456 & n25318 ) | ( n25314 & n25318 ) ;
  assign n25320 = ~n350 & n4708 ;
  assign n25321 = n2359 & ~n25320 ;
  assign n25322 = n25321 ^ n6555 ^ n3891 ;
  assign n25323 = ( ~n495 & n8337 ) | ( ~n495 & n12901 ) | ( n8337 & n12901 ) ;
  assign n25324 = n24421 ^ n12070 ^ 1'b0 ;
  assign n25325 = n25323 & n25324 ;
  assign n25326 = ( ~n7291 & n17783 ) | ( ~n7291 & n25325 ) | ( n17783 & n25325 ) ;
  assign n25327 = ~n15305 & n16433 ;
  assign n25328 = n25327 ^ n17601 ^ 1'b0 ;
  assign n25329 = n16333 ^ n4750 ^ 1'b0 ;
  assign n25330 = n25328 & ~n25329 ;
  assign n25331 = ~n3625 & n18827 ;
  assign n25332 = n25331 ^ n15945 ^ 1'b0 ;
  assign n25333 = n1634 | n7165 ;
  assign n25334 = n25333 ^ n18288 ^ 1'b0 ;
  assign n25335 = n5674 & n10128 ;
  assign n25336 = n1040 & n25335 ;
  assign n25337 = n6182 | n13824 ;
  assign n25338 = n25337 ^ n16981 ^ 1'b0 ;
  assign n25339 = n20032 ^ n1333 ^ 1'b0 ;
  assign n25340 = ( n9637 & n25338 ) | ( n9637 & ~n25339 ) | ( n25338 & ~n25339 ) ;
  assign n25341 = n25340 ^ n16124 ^ n14957 ;
  assign n25342 = ( n8824 & n11009 ) | ( n8824 & n14052 ) | ( n11009 & n14052 ) ;
  assign n25343 = n25342 ^ n19966 ^ 1'b0 ;
  assign n25344 = n17823 & ~n25343 ;
  assign n25345 = n1385 & n15221 ;
  assign n25346 = n4796 ^ n2289 ^ 1'b0 ;
  assign n25347 = ( n7241 & n19086 ) | ( n7241 & ~n25346 ) | ( n19086 & ~n25346 ) ;
  assign n25348 = ( n9234 & ~n19198 ) | ( n9234 & n25347 ) | ( ~n19198 & n25347 ) ;
  assign n25349 = n19106 ^ n738 ^ 1'b0 ;
  assign n25350 = ~n13114 & n25349 ;
  assign n25351 = n15869 & n25350 ;
  assign n25352 = ( n6143 & ~n9503 ) | ( n6143 & n10511 ) | ( ~n9503 & n10511 ) ;
  assign n25353 = ~n687 & n25352 ;
  assign n25354 = ~n19099 & n25353 ;
  assign n25355 = n9209 & n19258 ;
  assign n25356 = n11116 | n25355 ;
  assign n25357 = n4733 & ~n10916 ;
  assign n25358 = n9966 & n25357 ;
  assign n25359 = n25358 ^ n12076 ^ 1'b0 ;
  assign n25360 = ( ~n774 & n18631 ) | ( ~n774 & n25359 ) | ( n18631 & n25359 ) ;
  assign n25361 = n6162 ^ n1438 ^ n992 ;
  assign n25362 = n11816 | n25361 ;
  assign n25363 = n13034 ^ n1517 ^ 1'b0 ;
  assign n25364 = n1622 & ~n25363 ;
  assign n25365 = n2220 & ~n25364 ;
  assign n25375 = n277 & ~n6782 ;
  assign n25376 = n25375 ^ n8278 ^ 1'b0 ;
  assign n25372 = n1381 & n6311 ;
  assign n25373 = n9042 & n25372 ;
  assign n25374 = n25373 ^ n21059 ^ n13376 ;
  assign n25366 = n10760 ^ n1047 ^ 1'b0 ;
  assign n25367 = n5363 & n25366 ;
  assign n25368 = n4937 & n10570 ;
  assign n25369 = n25368 ^ n6331 ^ 1'b0 ;
  assign n25370 = ~n2641 & n25369 ;
  assign n25371 = ~n25367 & n25370 ;
  assign n25377 = n25376 ^ n25374 ^ n25371 ;
  assign n25378 = n13205 ^ n5551 ^ n5162 ;
  assign n25379 = n25378 ^ n14471 ^ n12483 ;
  assign n25380 = ( ~n8743 & n15594 ) | ( ~n8743 & n21871 ) | ( n15594 & n21871 ) ;
  assign n25381 = n5653 & n9093 ;
  assign n25382 = ~n12726 & n25381 ;
  assign n25383 = ( n13655 & ~n22980 ) | ( n13655 & n25382 ) | ( ~n22980 & n25382 ) ;
  assign n25384 = n2256 ^ n1266 ^ 1'b0 ;
  assign n25385 = x70 & n25384 ;
  assign n25386 = ( n16281 & n18075 ) | ( n16281 & n25385 ) | ( n18075 & n25385 ) ;
  assign n25387 = n25383 & ~n25386 ;
  assign n25388 = ( n10016 & ~n12580 ) | ( n10016 & n17896 ) | ( ~n12580 & n17896 ) ;
  assign n25389 = n9654 | n25388 ;
  assign n25390 = n16590 | n25292 ;
  assign n25391 = n10984 & ~n25390 ;
  assign n25392 = n11363 ^ n4875 ^ 1'b0 ;
  assign n25393 = n9285 | n25392 ;
  assign n25394 = n3752 | n25393 ;
  assign n25395 = ~n7488 & n11704 ;
  assign n25396 = ( n4975 & n13430 ) | ( n4975 & n25395 ) | ( n13430 & n25395 ) ;
  assign n25397 = n19756 ^ n6707 ^ 1'b0 ;
  assign n25398 = n10360 ^ n2122 ^ 1'b0 ;
  assign n25399 = n3799 | n25398 ;
  assign n25400 = n25397 & ~n25399 ;
  assign n25401 = n5921 & n25400 ;
  assign n25402 = n10759 & ~n18081 ;
  assign n25403 = ( n12560 & n25401 ) | ( n12560 & ~n25402 ) | ( n25401 & ~n25402 ) ;
  assign n25404 = n1298 ^ n814 ^ 1'b0 ;
  assign n25405 = n14896 & n25404 ;
  assign n25406 = n25405 ^ n13875 ^ 1'b0 ;
  assign n25407 = n5308 & n9740 ;
  assign n25408 = n25407 ^ n2812 ^ 1'b0 ;
  assign n25409 = ( n3796 & n11272 ) | ( n3796 & n18201 ) | ( n11272 & n18201 ) ;
  assign n25410 = n25408 & n25409 ;
  assign n25411 = ~n14582 & n25410 ;
  assign n25412 = ~n6011 & n9868 ;
  assign n25413 = n14022 ^ n8442 ^ 1'b0 ;
  assign n25414 = ( n8333 & n14658 ) | ( n8333 & ~n25413 ) | ( n14658 & ~n25413 ) ;
  assign n25415 = ( n11153 & ~n12247 ) | ( n11153 & n25414 ) | ( ~n12247 & n25414 ) ;
  assign n25416 = n9225 | n13818 ;
  assign n25417 = n25416 ^ n9339 ^ 1'b0 ;
  assign n25418 = n4730 ^ n756 ^ 1'b0 ;
  assign n25419 = n3393 | n25418 ;
  assign n25420 = ~n25417 & n25419 ;
  assign n25421 = ~n9288 & n13150 ;
  assign n25422 = n25421 ^ n6474 ^ 1'b0 ;
  assign n25423 = n25422 ^ n19887 ^ 1'b0 ;
  assign n25424 = n8671 ^ n6659 ^ 1'b0 ;
  assign n25425 = ( n7853 & ~n14448 ) | ( n7853 & n21707 ) | ( ~n14448 & n21707 ) ;
  assign n25426 = n21004 ^ n20017 ^ n3101 ;
  assign n25427 = n1467 & ~n2876 ;
  assign n25428 = n21275 ^ n8318 ^ 1'b0 ;
  assign n25433 = n25373 ^ n18390 ^ n7480 ;
  assign n25434 = n22724 & n25433 ;
  assign n25435 = n17494 & n25434 ;
  assign n25429 = n4848 ^ n4005 ^ 1'b0 ;
  assign n25430 = n17164 ^ n13831 ^ 1'b0 ;
  assign n25431 = n25429 & n25430 ;
  assign n25432 = n17314 & ~n25431 ;
  assign n25436 = n25435 ^ n25432 ^ n19266 ;
  assign n25437 = ~n13331 & n24685 ;
  assign n25438 = n25437 ^ n11607 ^ 1'b0 ;
  assign n25439 = n12424 & n24307 ;
  assign n25440 = ( ~n6334 & n21478 ) | ( ~n6334 & n22153 ) | ( n21478 & n22153 ) ;
  assign n25441 = n25440 ^ n8828 ^ n5300 ;
  assign n25443 = n7198 & n7994 ;
  assign n25444 = n25443 ^ n2112 ^ 1'b0 ;
  assign n25445 = n25444 ^ n7719 ^ n4359 ;
  assign n25442 = ( n2121 & n4307 ) | ( n2121 & ~n23360 ) | ( n4307 & ~n23360 ) ;
  assign n25446 = n25445 ^ n25442 ^ n24950 ;
  assign n25447 = ( ~n13285 & n14587 ) | ( ~n13285 & n17168 ) | ( n14587 & n17168 ) ;
  assign n25448 = n25447 ^ n19924 ^ 1'b0 ;
  assign n25449 = n4182 & ~n25448 ;
  assign n25450 = n13616 | n22925 ;
  assign n25451 = n25450 ^ n19462 ^ 1'b0 ;
  assign n25452 = n5026 ^ n615 ^ 1'b0 ;
  assign n25453 = n25452 ^ n2684 ^ 1'b0 ;
  assign n25454 = ( n1056 & n6205 ) | ( n1056 & ~n15323 ) | ( n6205 & ~n15323 ) ;
  assign n25455 = n25454 ^ n3401 ^ 1'b0 ;
  assign n25456 = ~n1725 & n25455 ;
  assign n25457 = ( n22178 & n25453 ) | ( n22178 & n25456 ) | ( n25453 & n25456 ) ;
  assign n25458 = n657 | n1864 ;
  assign n25459 = n2450 | n25458 ;
  assign n25460 = n20888 ^ n17224 ^ n13569 ;
  assign n25461 = n16840 & n25460 ;
  assign n25462 = n25459 & ~n25461 ;
  assign n25463 = n25462 ^ n1391 ^ 1'b0 ;
  assign n25464 = n2747 & ~n14836 ;
  assign n25465 = n25464 ^ n16222 ^ 1'b0 ;
  assign n25466 = n25465 ^ n12086 ^ 1'b0 ;
  assign n25467 = ~n7657 & n25466 ;
  assign n25468 = n6083 & n8298 ;
  assign n25469 = n25468 ^ n3231 ^ 1'b0 ;
  assign n25470 = n6074 | n6758 ;
  assign n25471 = ( n4638 & ~n13599 ) | ( n4638 & n25470 ) | ( ~n13599 & n25470 ) ;
  assign n25474 = n14829 ^ n1720 ^ 1'b0 ;
  assign n25475 = ( n13324 & ~n14168 ) | ( n13324 & n25474 ) | ( ~n14168 & n25474 ) ;
  assign n25472 = ~n4900 & n15750 ;
  assign n25473 = ~n5341 & n25472 ;
  assign n25476 = n25475 ^ n25473 ^ n24749 ;
  assign n25477 = ( ~n25469 & n25471 ) | ( ~n25469 & n25476 ) | ( n25471 & n25476 ) ;
  assign n25478 = ( n1808 & n14311 ) | ( n1808 & ~n20067 ) | ( n14311 & ~n20067 ) ;
  assign n25479 = n16348 ^ n15550 ^ 1'b0 ;
  assign n25480 = n5530 & n25479 ;
  assign n25481 = ( n12607 & n19446 ) | ( n12607 & ~n25480 ) | ( n19446 & ~n25480 ) ;
  assign n25482 = ~n3693 & n5038 ;
  assign n25483 = n25482 ^ n25422 ^ 1'b0 ;
  assign n25484 = ~n6637 & n25483 ;
  assign n25489 = n22170 ^ n4544 ^ 1'b0 ;
  assign n25490 = ~n2876 & n25489 ;
  assign n25491 = ~n24447 & n25490 ;
  assign n25492 = ~n6852 & n25491 ;
  assign n25485 = n18460 ^ n4364 ^ n2525 ;
  assign n25486 = n20359 ^ n16451 ^ n10167 ;
  assign n25487 = ( n10835 & n22557 ) | ( n10835 & n25486 ) | ( n22557 & n25486 ) ;
  assign n25488 = ( n15532 & ~n25485 ) | ( n15532 & n25487 ) | ( ~n25485 & n25487 ) ;
  assign n25493 = n25492 ^ n25488 ^ n17212 ;
  assign n25494 = n15078 & n25493 ;
  assign n25495 = n21752 ^ n14358 ^ 1'b0 ;
  assign n25496 = n8119 & n11832 ;
  assign n25498 = ~n1934 & n15012 ;
  assign n25497 = x179 & n8125 ;
  assign n25499 = n25498 ^ n25497 ^ 1'b0 ;
  assign n25503 = n12080 ^ n3459 ^ 1'b0 ;
  assign n25504 = ~n2267 & n25503 ;
  assign n25500 = n688 | n18048 ;
  assign n25501 = n25500 ^ n12113 ^ 1'b0 ;
  assign n25502 = ~n6754 & n25501 ;
  assign n25505 = n25504 ^ n25502 ^ 1'b0 ;
  assign n25506 = n20141 ^ n14275 ^ 1'b0 ;
  assign n25507 = ~n25505 & n25506 ;
  assign n25509 = n9217 ^ n7026 ^ 1'b0 ;
  assign n25510 = ~n19289 & n25509 ;
  assign n25508 = n9470 & n12322 ;
  assign n25511 = n25510 ^ n25508 ^ 1'b0 ;
  assign n25513 = n1539 & n4684 ;
  assign n25514 = n25513 ^ n24527 ^ 1'b0 ;
  assign n25515 = n13748 ^ n10968 ^ 1'b0 ;
  assign n25516 = ~n25514 & n25515 ;
  assign n25517 = n17428 ^ n6156 ^ n4849 ;
  assign n25518 = n492 & n25517 ;
  assign n25519 = n25518 ^ n7358 ^ 1'b0 ;
  assign n25520 = n25519 ^ n19207 ^ n750 ;
  assign n25521 = ( n5042 & n25516 ) | ( n5042 & ~n25520 ) | ( n25516 & ~n25520 ) ;
  assign n25512 = n24504 ^ n1202 ^ 1'b0 ;
  assign n25522 = n25521 ^ n25512 ^ n1630 ;
  assign n25525 = n9500 & n12381 ;
  assign n25523 = n8068 ^ x216 ^ 1'b0 ;
  assign n25524 = n25523 ^ n9648 ^ n4325 ;
  assign n25526 = n25525 ^ n25524 ^ n9591 ;
  assign n25527 = n25526 ^ n3166 ^ 1'b0 ;
  assign n25528 = n25522 & ~n25527 ;
  assign n25529 = n25528 ^ n22678 ^ n9970 ;
  assign n25530 = ~n12472 & n13127 ;
  assign n25531 = n18699 ^ n8760 ^ n4588 ;
  assign n25534 = n7215 ^ n4835 ^ 1'b0 ;
  assign n25535 = ~n11706 & n25534 ;
  assign n25533 = n19369 ^ n9273 ^ 1'b0 ;
  assign n25536 = n25535 ^ n25533 ^ n8594 ;
  assign n25532 = ( n5388 & n9640 ) | ( n5388 & ~n23575 ) | ( n9640 & ~n23575 ) ;
  assign n25537 = n25536 ^ n25532 ^ 1'b0 ;
  assign n25538 = ~n25531 & n25537 ;
  assign n25539 = n25530 | n25538 ;
  assign n25540 = n6994 & ~n17976 ;
  assign n25541 = n7108 ^ n5491 ^ n668 ;
  assign n25542 = ~n18216 & n25541 ;
  assign n25543 = n17154 & n25542 ;
  assign n25544 = n2506 & n4350 ;
  assign n25545 = n25544 ^ n826 ^ 1'b0 ;
  assign n25546 = ( n8116 & n10325 ) | ( n8116 & ~n25545 ) | ( n10325 & ~n25545 ) ;
  assign n25547 = ~n2146 & n25546 ;
  assign n25548 = n25543 & n25547 ;
  assign n25549 = n13452 ^ n2450 ^ 1'b0 ;
  assign n25550 = n22798 ^ n19879 ^ 1'b0 ;
  assign n25551 = n25550 ^ n22660 ^ 1'b0 ;
  assign n25552 = ~n25549 & n25551 ;
  assign n25553 = n25552 ^ n2394 ^ 1'b0 ;
  assign n25554 = n9687 & ~n25553 ;
  assign n25555 = n590 | n11197 ;
  assign n25556 = n25555 ^ n13046 ^ 1'b0 ;
  assign n25557 = ~n20793 & n25556 ;
  assign n25558 = n18944 | n25557 ;
  assign n25559 = n8848 ^ n5984 ^ 1'b0 ;
  assign n25560 = n25559 ^ n23684 ^ n1532 ;
  assign n25564 = n8538 | n14689 ;
  assign n25561 = ( n2236 & n2621 ) | ( n2236 & ~n24303 ) | ( n2621 & ~n24303 ) ;
  assign n25562 = n25561 ^ n3535 ^ 1'b0 ;
  assign n25563 = ~n3913 & n25562 ;
  assign n25565 = n25564 ^ n25563 ^ n2117 ;
  assign n25566 = n2417 & n18230 ;
  assign n25567 = n24401 ^ n14192 ^ n3683 ;
  assign n25568 = ( ~n10472 & n25566 ) | ( ~n10472 & n25567 ) | ( n25566 & n25567 ) ;
  assign n25569 = n8484 & ~n11412 ;
  assign n25570 = n24529 ^ n8754 ^ 1'b0 ;
  assign n25571 = ~n25569 & n25570 ;
  assign n25572 = n21354 ^ n5799 ^ 1'b0 ;
  assign n25573 = n616 ^ x67 ^ 1'b0 ;
  assign n25574 = n6079 & n25573 ;
  assign n25575 = n20586 & n25574 ;
  assign n25579 = ~n5403 & n12437 ;
  assign n25580 = ( ~n2234 & n25367 ) | ( ~n2234 & n25579 ) | ( n25367 & n25579 ) ;
  assign n25576 = ( ~n1634 & n8244 ) | ( ~n1634 & n9746 ) | ( n8244 & n9746 ) ;
  assign n25577 = n8612 | n25576 ;
  assign n25578 = ~n12565 & n25577 ;
  assign n25581 = n25580 ^ n25578 ^ 1'b0 ;
  assign n25582 = n7421 & ~n11972 ;
  assign n25583 = ~n2894 & n25582 ;
  assign n25589 = n10997 ^ n591 ^ n579 ;
  assign n25586 = n9503 & ~n15234 ;
  assign n25587 = n25586 ^ n17892 ^ 1'b0 ;
  assign n25588 = n10524 & n25587 ;
  assign n25590 = n25589 ^ n25588 ^ 1'b0 ;
  assign n25584 = n24186 ^ n16348 ^ 1'b0 ;
  assign n25585 = n14858 | n25584 ;
  assign n25591 = n25590 ^ n25585 ^ 1'b0 ;
  assign n25592 = ( n2987 & ~n17875 ) | ( n2987 & n19049 ) | ( ~n17875 & n19049 ) ;
  assign n25593 = ( n4282 & ~n18608 ) | ( n4282 & n25592 ) | ( ~n18608 & n25592 ) ;
  assign n25594 = ( n14207 & ~n21692 ) | ( n14207 & n25593 ) | ( ~n21692 & n25593 ) ;
  assign n25595 = n11091 & n17420 ;
  assign n25596 = ~n11853 & n25595 ;
  assign n25597 = n22687 ^ n9293 ^ 1'b0 ;
  assign n25598 = n25597 ^ n18530 ^ n12193 ;
  assign n25599 = n18323 ^ n12957 ^ n10150 ;
  assign n25600 = n8622 ^ n7852 ^ 1'b0 ;
  assign n25601 = ~n25599 & n25600 ;
  assign n25602 = n12573 & ~n18335 ;
  assign n25603 = ~n22340 & n25602 ;
  assign n25604 = n18661 ^ n14974 ^ n8506 ;
  assign n25605 = n25604 ^ n20096 ^ n14602 ;
  assign n25606 = n2699 & n22202 ;
  assign n25607 = n16826 & n25606 ;
  assign n25608 = n25607 ^ n23823 ^ 1'b0 ;
  assign n25609 = ( n9384 & ~n23118 ) | ( n9384 & n24036 ) | ( ~n23118 & n24036 ) ;
  assign n25610 = n25609 ^ n17713 ^ n16732 ;
  assign n25611 = n9494 ^ n3964 ^ 1'b0 ;
  assign n25612 = ~n23645 & n25611 ;
  assign n25613 = ( n2332 & n9625 ) | ( n2332 & n16136 ) | ( n9625 & n16136 ) ;
  assign n25614 = n25613 ^ n23592 ^ 1'b0 ;
  assign n25615 = n20742 & ~n25614 ;
  assign n25616 = n3358 | n7240 ;
  assign n25617 = n15513 | n25616 ;
  assign n25618 = ( n1036 & n12362 ) | ( n1036 & n25617 ) | ( n12362 & n25617 ) ;
  assign n25619 = n19708 & n25618 ;
  assign n25620 = n6247 | n16466 ;
  assign n25621 = n25619 & ~n25620 ;
  assign n25622 = n23799 ^ n6237 ^ 1'b0 ;
  assign n25623 = n10759 ^ n4760 ^ 1'b0 ;
  assign n25624 = n13449 ^ n10755 ^ n6797 ;
  assign n25625 = ~n12941 & n25624 ;
  assign n25626 = n2035 & ~n3389 ;
  assign n25627 = n25626 ^ n4090 ^ 1'b0 ;
  assign n25628 = ( n4870 & n9040 ) | ( n4870 & ~n25627 ) | ( n9040 & ~n25627 ) ;
  assign n25629 = ( n1911 & n15684 ) | ( n1911 & ~n25628 ) | ( n15684 & ~n25628 ) ;
  assign n25630 = n16662 ^ n7422 ^ n6132 ;
  assign n25631 = n25630 ^ n5910 ^ n1640 ;
  assign n25633 = n4732 | n5840 ;
  assign n25634 = n25079 ^ n1449 ^ 1'b0 ;
  assign n25635 = n25633 & n25634 ;
  assign n25632 = n883 | n14973 ;
  assign n25636 = n25635 ^ n25632 ^ 1'b0 ;
  assign n25637 = n8780 | n20805 ;
  assign n25638 = n8523 ^ n6562 ^ 1'b0 ;
  assign n25639 = n25637 & n25638 ;
  assign n25640 = ~n4527 & n25639 ;
  assign n25641 = n25640 ^ n11295 ^ 1'b0 ;
  assign n25642 = n9163 ^ n2561 ^ 1'b0 ;
  assign n25643 = n9740 & n18659 ;
  assign n25644 = ~n25642 & n25643 ;
  assign n25645 = n5956 | n14803 ;
  assign n25646 = ( n10418 & ~n10750 ) | ( n10418 & n25645 ) | ( ~n10750 & n25645 ) ;
  assign n25647 = n4568 | n17643 ;
  assign n25648 = n12319 | n25647 ;
  assign n25649 = n25648 ^ n9827 ^ n7146 ;
  assign n25650 = n25649 ^ n5962 ^ n4046 ;
  assign n25651 = n6279 | n22387 ;
  assign n25652 = n24769 | n25651 ;
  assign n25653 = n21617 | n25652 ;
  assign n25654 = n1787 | n6887 ;
  assign n25655 = n1673 & ~n25654 ;
  assign n25656 = n21792 | n21995 ;
  assign n25657 = n20805 ^ n19258 ^ n8120 ;
  assign n25658 = ( n3319 & ~n9665 ) | ( n3319 & n19525 ) | ( ~n9665 & n19525 ) ;
  assign n25659 = n25658 ^ n19241 ^ n10022 ;
  assign n25660 = ( n1763 & n5094 ) | ( n1763 & ~n8857 ) | ( n5094 & ~n8857 ) ;
  assign n25661 = n25660 ^ n10844 ^ 1'b0 ;
  assign n25662 = n25661 ^ n18512 ^ 1'b0 ;
  assign n25663 = n25662 ^ n17643 ^ n11193 ;
  assign n25664 = n2824 & n25663 ;
  assign n25665 = ~x254 & n25664 ;
  assign n25668 = n9246 | n16276 ;
  assign n25669 = n9251 & ~n25668 ;
  assign n25670 = ~n12386 & n25669 ;
  assign n25666 = ( n8249 & n13354 ) | ( n8249 & n18282 ) | ( n13354 & n18282 ) ;
  assign n25667 = ~n2388 & n25666 ;
  assign n25671 = n25670 ^ n25667 ^ 1'b0 ;
  assign n25675 = n4575 ^ n1352 ^ x235 ;
  assign n25676 = n2362 & n25675 ;
  assign n25677 = n14243 & n25676 ;
  assign n25672 = n337 & n3719 ;
  assign n25673 = ~n12210 & n25672 ;
  assign n25674 = n4675 & ~n25673 ;
  assign n25678 = n25677 ^ n25674 ^ 1'b0 ;
  assign n25679 = ( n3921 & ~n10114 ) | ( n3921 & n15502 ) | ( ~n10114 & n15502 ) ;
  assign n25680 = ~n3075 & n25679 ;
  assign n25681 = ~n13303 & n25680 ;
  assign n25691 = n14686 & ~n16479 ;
  assign n25692 = n25691 ^ n4714 ^ 1'b0 ;
  assign n25690 = n5737 & ~n15128 ;
  assign n25683 = n3541 ^ n2849 ^ 1'b0 ;
  assign n25684 = x223 & n25683 ;
  assign n25685 = n15413 & n25684 ;
  assign n25682 = n11079 | n13824 ;
  assign n25686 = n25685 ^ n25682 ^ 1'b0 ;
  assign n25687 = ( n7548 & n8995 ) | ( n7548 & ~n24131 ) | ( n8995 & ~n24131 ) ;
  assign n25688 = n6228 | n25687 ;
  assign n25689 = n25686 & ~n25688 ;
  assign n25693 = n25692 ^ n25690 ^ n25689 ;
  assign n25694 = n17362 ^ n1400 ^ 1'b0 ;
  assign n25695 = ~n25576 & n25694 ;
  assign n25696 = ~n24002 & n25695 ;
  assign n25697 = n7226 & n25696 ;
  assign n25698 = n6725 & n21599 ;
  assign n25699 = n7965 ^ n2340 ^ 1'b0 ;
  assign n25700 = n15041 | n25699 ;
  assign n25701 = n11332 | n25700 ;
  assign n25702 = n20839 & n25701 ;
  assign n25703 = ~n345 & n25702 ;
  assign n25704 = n373 & n1198 ;
  assign n25705 = n7784 & n25704 ;
  assign n25706 = n15653 & ~n25705 ;
  assign n25707 = n20028 & ~n24221 ;
  assign n25708 = n25707 ^ n13954 ^ 1'b0 ;
  assign n25709 = ~n12861 & n25708 ;
  assign n25710 = n15085 & n25709 ;
  assign n25711 = n25710 ^ n20274 ^ 1'b0 ;
  assign n25712 = n11316 ^ n258 ^ 1'b0 ;
  assign n25713 = n8015 & ~n25712 ;
  assign n25714 = ~n6580 & n25713 ;
  assign n25715 = n262 & n25714 ;
  assign n25716 = n11871 | n25715 ;
  assign n25717 = n9992 | n25716 ;
  assign n25718 = ( ~n675 & n3091 ) | ( ~n675 & n10167 ) | ( n3091 & n10167 ) ;
  assign n25719 = ( n15843 & ~n25717 ) | ( n15843 & n25718 ) | ( ~n25717 & n25718 ) ;
  assign n25720 = n5086 | n6977 ;
  assign n25721 = ( ~n10119 & n13589 ) | ( ~n10119 & n14664 ) | ( n13589 & n14664 ) ;
  assign n25723 = n7806 & n13752 ;
  assign n25724 = n25723 ^ n6495 ^ 1'b0 ;
  assign n25725 = ~n3016 & n25724 ;
  assign n25726 = n11804 ^ n8533 ^ 1'b0 ;
  assign n25727 = n20951 & ~n25726 ;
  assign n25728 = n25727 ^ n2613 ^ 1'b0 ;
  assign n25729 = n3496 | n25728 ;
  assign n25730 = n25725 | n25729 ;
  assign n25722 = n1964 & n10477 ;
  assign n25731 = n25730 ^ n25722 ^ 1'b0 ;
  assign n25732 = n8915 & ~n16329 ;
  assign n25733 = n12811 | n19584 ;
  assign n25734 = n8397 | n25733 ;
  assign n25735 = n25636 ^ n6476 ^ 1'b0 ;
  assign n25736 = ~n327 & n15125 ;
  assign n25737 = n25736 ^ n17971 ^ n5481 ;
  assign n25738 = n25737 ^ n16855 ^ x19 ;
  assign n25739 = n10121 & n25738 ;
  assign n25740 = n3805 ^ n3272 ^ n435 ;
  assign n25741 = n19375 & n25740 ;
  assign n25742 = ~n11689 & n25741 ;
  assign n25743 = ~n11289 & n14163 ;
  assign n25744 = n25743 ^ n16945 ^ n1838 ;
  assign n25745 = n25744 ^ n20227 ^ n8383 ;
  assign n25746 = n9949 ^ n2808 ^ n287 ;
  assign n25747 = n25746 ^ n14834 ^ 1'b0 ;
  assign n25748 = n25745 & n25747 ;
  assign n25749 = ~n23005 & n25748 ;
  assign n25753 = ~n6843 & n24893 ;
  assign n25750 = n19146 ^ n16338 ^ 1'b0 ;
  assign n25751 = ~n20633 & n25750 ;
  assign n25752 = n19547 & n25751 ;
  assign n25754 = n25753 ^ n25752 ^ 1'b0 ;
  assign n25755 = n4173 | n11585 ;
  assign n25756 = n21682 | n25755 ;
  assign n25757 = ~n15041 & n18641 ;
  assign n25758 = n1497 & n4501 ;
  assign n25759 = n25758 ^ n2504 ^ 1'b0 ;
  assign n25760 = n25759 ^ n8122 ^ n1643 ;
  assign n25761 = ( n8461 & n8754 ) | ( n8461 & ~n25589 ) | ( n8754 & ~n25589 ) ;
  assign n25762 = n11365 ^ x34 ^ 1'b0 ;
  assign n25763 = n10645 & n25762 ;
  assign n25764 = n15942 ^ n2333 ^ 1'b0 ;
  assign n25765 = ( ~x4 & n25763 ) | ( ~x4 & n25764 ) | ( n25763 & n25764 ) ;
  assign n25766 = n15251 & ~n25765 ;
  assign n25767 = n14854 & n25766 ;
  assign n25768 = n25767 ^ n9008 ^ 1'b0 ;
  assign n25769 = x103 | n4641 ;
  assign n25770 = n25769 ^ n4779 ^ 1'b0 ;
  assign n25771 = n16737 | n25770 ;
  assign n25772 = ( ~n3273 & n5009 ) | ( ~n3273 & n6310 ) | ( n5009 & n6310 ) ;
  assign n25773 = n25772 ^ n1281 ^ 1'b0 ;
  assign n25774 = ( n13367 & n25771 ) | ( n13367 & n25773 ) | ( n25771 & n25773 ) ;
  assign n25775 = n25774 ^ n20696 ^ 1'b0 ;
  assign n25776 = n1541 | n25775 ;
  assign n25777 = n10461 | n19278 ;
  assign n25778 = n25777 ^ n22084 ^ 1'b0 ;
  assign n25779 = n789 | n25778 ;
  assign n25780 = n7116 ^ n637 ^ 1'b0 ;
  assign n25781 = n25780 ^ n9589 ^ 1'b0 ;
  assign n25782 = n25781 ^ n17132 ^ n10259 ;
  assign n25783 = ( n4165 & n10487 ) | ( n4165 & ~n19445 ) | ( n10487 & ~n19445 ) ;
  assign n25784 = n25783 ^ n6085 ^ 1'b0 ;
  assign n25785 = n25784 ^ n6205 ^ 1'b0 ;
  assign n25786 = n5530 & n9315 ;
  assign n25787 = n25786 ^ n14290 ^ 1'b0 ;
  assign n25788 = n25787 ^ n3608 ^ 1'b0 ;
  assign n25789 = n19293 ^ n2354 ^ 1'b0 ;
  assign n25790 = ~n25788 & n25789 ;
  assign n25791 = n2036 & n12411 ;
  assign n25792 = n23496 | n25791 ;
  assign n25793 = ( ~n3785 & n8370 ) | ( ~n3785 & n17589 ) | ( n8370 & n17589 ) ;
  assign n25794 = n25793 ^ n16021 ^ n8500 ;
  assign n25795 = n25794 ^ n22340 ^ n14583 ;
  assign n25796 = n9211 | n20137 ;
  assign n25797 = n17607 ^ n10107 ^ 1'b0 ;
  assign n25798 = n1971 | n25797 ;
  assign n25799 = n6962 ^ n4590 ^ n4356 ;
  assign n25800 = n9702 ^ n3832 ^ 1'b0 ;
  assign n25801 = n2630 | n25800 ;
  assign n25802 = n25801 ^ n22191 ^ n15044 ;
  assign n25803 = n10597 ^ n322 ^ 1'b0 ;
  assign n25804 = n2402 & n3222 ;
  assign n25805 = n25804 ^ n4163 ^ 1'b0 ;
  assign n25806 = n25805 ^ n4089 ^ 1'b0 ;
  assign n25807 = n17383 | n25806 ;
  assign n25808 = n25807 ^ n3767 ^ 1'b0 ;
  assign n25809 = n13603 | n25808 ;
  assign n25810 = n5541 & n14107 ;
  assign n25811 = n4346 | n14268 ;
  assign n25812 = n25810 & ~n25811 ;
  assign n25813 = n18317 & n24023 ;
  assign n25815 = n10798 & ~n11542 ;
  assign n25816 = n9989 ^ n1557 ^ 1'b0 ;
  assign n25817 = ~n25815 & n25816 ;
  assign n25814 = n4895 & ~n17847 ;
  assign n25818 = n25817 ^ n25814 ^ n20397 ;
  assign n25819 = n19047 ^ n13071 ^ 1'b0 ;
  assign n25820 = n2097 ^ n579 ^ 1'b0 ;
  assign n25821 = ( n455 & n2822 ) | ( n455 & ~n3120 ) | ( n2822 & ~n3120 ) ;
  assign n25822 = n2283 & n25821 ;
  assign n25823 = ~n7646 & n25822 ;
  assign n25824 = n2216 & n25823 ;
  assign n25825 = n11031 ^ n8882 ^ 1'b0 ;
  assign n25826 = n25139 | n25825 ;
  assign n25831 = n21868 ^ n18116 ^ 1'b0 ;
  assign n25827 = n7595 | n8080 ;
  assign n25828 = n17098 | n25827 ;
  assign n25829 = n25828 ^ n5462 ^ 1'b0 ;
  assign n25830 = ( n4688 & n20794 ) | ( n4688 & n25829 ) | ( n20794 & n25829 ) ;
  assign n25832 = n25831 ^ n25830 ^ n10278 ;
  assign n25833 = ( n3581 & n7143 ) | ( n3581 & n11866 ) | ( n7143 & n11866 ) ;
  assign n25834 = ~n15696 & n25833 ;
  assign n25835 = n15455 & n25834 ;
  assign n25836 = n25835 ^ n24863 ^ 1'b0 ;
  assign n25837 = n17332 & n25836 ;
  assign n25840 = n1868 ^ n468 ^ 1'b0 ;
  assign n25838 = n6332 & ~n9010 ;
  assign n25839 = n9867 & n25838 ;
  assign n25841 = n25840 ^ n25839 ^ n22082 ;
  assign n25842 = n25841 ^ n19049 ^ 1'b0 ;
  assign n25843 = n6529 ^ n1922 ^ 1'b0 ;
  assign n25844 = n17718 & n25843 ;
  assign n25845 = n9093 & n9745 ;
  assign n25846 = ~n25844 & n25845 ;
  assign n25847 = n20909 ^ n18046 ^ n8251 ;
  assign n25848 = ( n5901 & n25846 ) | ( n5901 & n25847 ) | ( n25846 & n25847 ) ;
  assign n25849 = n5362 & n25848 ;
  assign n25850 = n2492 ^ n2103 ^ 1'b0 ;
  assign n25851 = n11106 & ~n22274 ;
  assign n25852 = ( n7075 & ~n22567 ) | ( n7075 & n25576 ) | ( ~n22567 & n25576 ) ;
  assign n25853 = ~n7127 & n10443 ;
  assign n25854 = ~n25852 & n25853 ;
  assign n25855 = n17029 & n25854 ;
  assign n25858 = ~n7128 & n7256 ;
  assign n25859 = n25858 ^ n626 ^ 1'b0 ;
  assign n25860 = ~n17014 & n25859 ;
  assign n25861 = n25860 ^ n14836 ^ 1'b0 ;
  assign n25862 = n25861 ^ n12946 ^ n7214 ;
  assign n25856 = ( n8273 & n14669 ) | ( n8273 & n21751 ) | ( n14669 & n21751 ) ;
  assign n25857 = n3583 & ~n25856 ;
  assign n25863 = n25862 ^ n25857 ^ 1'b0 ;
  assign n25864 = ~n14259 & n25320 ;
  assign n25865 = n25864 ^ n2408 ^ 1'b0 ;
  assign n25866 = n25863 & ~n25865 ;
  assign n25867 = n22911 ^ n22135 ^ n6846 ;
  assign n25868 = n25867 ^ n17649 ^ 1'b0 ;
  assign n25869 = ~n279 & n11560 ;
  assign n25870 = n25869 ^ n5268 ^ 1'b0 ;
  assign n25874 = n6357 ^ n4741 ^ 1'b0 ;
  assign n25871 = n13935 ^ n9936 ^ 1'b0 ;
  assign n25872 = n24611 & ~n25871 ;
  assign n25873 = n2201 & n25872 ;
  assign n25875 = n25874 ^ n25873 ^ 1'b0 ;
  assign n25876 = ~n3767 & n13623 ;
  assign n25877 = n25876 ^ n16176 ^ 1'b0 ;
  assign n25878 = ~n10308 & n12850 ;
  assign n25879 = n25877 & n25878 ;
  assign n25880 = n2227 & n25879 ;
  assign n25881 = n10792 ^ n2000 ^ 1'b0 ;
  assign n25882 = ~n13211 & n16740 ;
  assign n25883 = n9427 ^ n1688 ^ x230 ;
  assign n25884 = n25883 ^ n5364 ^ 1'b0 ;
  assign n25885 = ( n25881 & ~n25882 ) | ( n25881 & n25884 ) | ( ~n25882 & n25884 ) ;
  assign n25886 = n25885 ^ n18730 ^ 1'b0 ;
  assign n25887 = ( n867 & n19161 ) | ( n867 & n25886 ) | ( n19161 & n25886 ) ;
  assign n25895 = n3330 | n9337 ;
  assign n25896 = n25895 ^ n1537 ^ 1'b0 ;
  assign n25892 = n9288 ^ n6061 ^ 1'b0 ;
  assign n25893 = n18265 | n25892 ;
  assign n25890 = n400 & ~n2016 ;
  assign n25891 = n25890 ^ n14232 ^ 1'b0 ;
  assign n25894 = n25893 ^ n25891 ^ n2475 ;
  assign n25888 = n21808 ^ n1948 ^ 1'b0 ;
  assign n25889 = n813 & ~n25888 ;
  assign n25897 = n25896 ^ n25894 ^ n25889 ;
  assign n25898 = n9278 & ~n10955 ;
  assign n25899 = ( n13743 & ~n14849 ) | ( n13743 & n16654 ) | ( ~n14849 & n16654 ) ;
  assign n25900 = ~n1276 & n19347 ;
  assign n25901 = n10988 & ~n14963 ;
  assign n25902 = n25900 & n25901 ;
  assign n25903 = n25902 ^ n5030 ^ 1'b0 ;
  assign n25904 = ~n25899 & n25903 ;
  assign n25905 = ( n1121 & n25898 ) | ( n1121 & ~n25904 ) | ( n25898 & ~n25904 ) ;
  assign n25906 = n15433 ^ n8614 ^ n3360 ;
  assign n25907 = n16302 & n25906 ;
  assign n25908 = n9837 & n25907 ;
  assign n25909 = ( n9148 & n9675 ) | ( n9148 & n24095 ) | ( n9675 & n24095 ) ;
  assign n25910 = n25909 ^ n17049 ^ 1'b0 ;
  assign n25911 = n25910 ^ n9322 ^ 1'b0 ;
  assign n25912 = n25908 | n25911 ;
  assign n25913 = n2071 & ~n4974 ;
  assign n25914 = ( ~n7138 & n14136 ) | ( ~n7138 & n25913 ) | ( n14136 & n25913 ) ;
  assign n25915 = n25914 ^ n19164 ^ n3363 ;
  assign n25916 = ~n20996 & n25915 ;
  assign n25917 = n25916 ^ x140 ^ 1'b0 ;
  assign n25918 = ~n21006 & n25917 ;
  assign n25919 = ( n19464 & ~n22184 ) | ( n19464 & n25918 ) | ( ~n22184 & n25918 ) ;
  assign n25920 = ~n1111 & n21846 ;
  assign n25921 = n25920 ^ n19797 ^ 1'b0 ;
  assign n25922 = n540 | n25921 ;
  assign n25923 = n25922 ^ n12140 ^ 1'b0 ;
  assign n25924 = n20225 & ~n22720 ;
  assign n25925 = ( ~n1146 & n11966 ) | ( ~n1146 & n22202 ) | ( n11966 & n22202 ) ;
  assign n25926 = x144 & n25925 ;
  assign n25927 = n9605 ^ n5775 ^ n2697 ;
  assign n25928 = n3954 & ~n25927 ;
  assign n25929 = ~n3805 & n25928 ;
  assign n25930 = n25929 ^ n18900 ^ 1'b0 ;
  assign n25931 = n12646 | n21355 ;
  assign n25932 = ( n12899 & n25930 ) | ( n12899 & n25931 ) | ( n25930 & n25931 ) ;
  assign n25933 = ( n6196 & ~n24349 ) | ( n6196 & n24476 ) | ( ~n24349 & n24476 ) ;
  assign n25934 = n21403 & ~n25060 ;
  assign n25935 = n8651 & n25934 ;
  assign n25936 = n3949 | n5758 ;
  assign n25937 = n25538 ^ n20959 ^ n5181 ;
  assign n25939 = n13075 ^ n8206 ^ n1462 ;
  assign n25938 = n4049 & n17401 ;
  assign n25940 = n25939 ^ n25938 ^ 1'b0 ;
  assign n25941 = n12963 ^ n7630 ^ n1323 ;
  assign n25942 = n25941 ^ n11365 ^ 1'b0 ;
  assign n25943 = n3872 | n25942 ;
  assign n25944 = ( ~n7815 & n8800 ) | ( ~n7815 & n14839 ) | ( n8800 & n14839 ) ;
  assign n25945 = n25944 ^ n552 ^ 1'b0 ;
  assign n25946 = n14441 & ~n17639 ;
  assign n25947 = n25946 ^ n15678 ^ 1'b0 ;
  assign n25948 = ( n14707 & n25945 ) | ( n14707 & n25947 ) | ( n25945 & n25947 ) ;
  assign n25949 = ( n3826 & n7314 ) | ( n3826 & n25295 ) | ( n7314 & n25295 ) ;
  assign n25950 = ( ~n7349 & n25810 ) | ( ~n7349 & n25949 ) | ( n25810 & n25949 ) ;
  assign n25951 = n22799 ^ n19478 ^ 1'b0 ;
  assign n25952 = n25951 ^ n13587 ^ n1435 ;
  assign n25953 = ( ~n19616 & n25950 ) | ( ~n19616 & n25952 ) | ( n25950 & n25952 ) ;
  assign n25954 = n3297 | n18002 ;
  assign n25955 = n6727 & ~n25954 ;
  assign n25956 = n15627 | n25955 ;
  assign n25957 = n8783 | n25956 ;
  assign n25958 = n10581 & ~n12596 ;
  assign n25959 = ~n25957 & n25958 ;
  assign n25960 = ( n5078 & n18467 ) | ( n5078 & ~n24307 ) | ( n18467 & ~n24307 ) ;
  assign n25961 = n10183 ^ n892 ^ 1'b0 ;
  assign n25962 = n338 & ~n25961 ;
  assign n25963 = n25962 ^ n668 ^ 1'b0 ;
  assign n25964 = n6710 ^ n5445 ^ 1'b0 ;
  assign n25965 = n11798 & ~n25964 ;
  assign n25968 = n24662 ^ n13423 ^ 1'b0 ;
  assign n25967 = n13358 & ~n20272 ;
  assign n25966 = ~n15767 & n17596 ;
  assign n25969 = n25968 ^ n25967 ^ n25966 ;
  assign n25970 = n24505 ^ n2834 ^ 1'b0 ;
  assign n25971 = n1137 & ~n3966 ;
  assign n25972 = n25971 ^ n16089 ^ n1152 ;
  assign n25973 = n18623 | n18863 ;
  assign n25974 = n20664 & n25973 ;
  assign n25975 = ~n19918 & n25598 ;
  assign n25976 = n24477 ^ n16365 ^ n1078 ;
  assign n25977 = n13766 | n19005 ;
  assign n25978 = n25977 ^ n13039 ^ 1'b0 ;
  assign n25979 = n8008 & ~n22387 ;
  assign n25980 = n4444 & ~n6771 ;
  assign n25981 = n6019 & n25980 ;
  assign n25982 = n25981 ^ x90 ^ 1'b0 ;
  assign n25983 = n13332 | n25982 ;
  assign n25984 = n625 | n13831 ;
  assign n25985 = n25984 ^ n7424 ^ 1'b0 ;
  assign n25987 = n1573 ^ x135 ^ 1'b0 ;
  assign n25986 = ( ~n2187 & n5409 ) | ( ~n2187 & n16769 ) | ( n5409 & n16769 ) ;
  assign n25988 = n25987 ^ n25986 ^ 1'b0 ;
  assign n25989 = n25985 | n25988 ;
  assign n25990 = ( n12146 & ~n14826 ) | ( n12146 & n25989 ) | ( ~n14826 & n25989 ) ;
  assign n25991 = n25918 ^ n14502 ^ 1'b0 ;
  assign n25992 = n4967 & ~n9954 ;
  assign n25993 = n25992 ^ n15920 ^ n15838 ;
  assign n25996 = n14396 ^ n715 ^ 1'b0 ;
  assign n25997 = n25996 ^ n13646 ^ 1'b0 ;
  assign n25994 = n365 | n807 ;
  assign n25995 = n9001 & ~n25994 ;
  assign n25998 = n25997 ^ n25995 ^ n1513 ;
  assign n25999 = n18447 ^ n488 ^ 1'b0 ;
  assign n26000 = n25459 ^ n10663 ^ 1'b0 ;
  assign n26001 = ( n8506 & ~n25999 ) | ( n8506 & n26000 ) | ( ~n25999 & n26000 ) ;
  assign n26002 = ~n23378 & n23636 ;
  assign n26003 = n26002 ^ n14832 ^ n8657 ;
  assign n26004 = n26003 ^ n12524 ^ n2265 ;
  assign n26005 = n9542 & ~n13927 ;
  assign n26006 = n5536 & ~n6634 ;
  assign n26007 = ~n1585 & n26006 ;
  assign n26008 = n10534 ^ n6623 ^ 1'b0 ;
  assign n26009 = n18997 | n26008 ;
  assign n26010 = n26009 ^ n1331 ^ 1'b0 ;
  assign n26011 = n26007 & ~n26010 ;
  assign n26012 = n18121 ^ n940 ^ 1'b0 ;
  assign n26013 = n7642 ^ n1537 ^ 1'b0 ;
  assign n26014 = n6641 & n26013 ;
  assign n26015 = ~n26012 & n26014 ;
  assign n26016 = n14898 | n23196 ;
  assign n26017 = n21519 & n25405 ;
  assign n26018 = n26017 ^ n11244 ^ 1'b0 ;
  assign n26019 = ( ~n4773 & n6336 ) | ( ~n4773 & n18854 ) | ( n6336 & n18854 ) ;
  assign n26020 = n26019 ^ n16028 ^ n14542 ;
  assign n26021 = n23254 | n24564 ;
  assign n26022 = n26020 | n26021 ;
  assign n26023 = ( n11364 & n26018 ) | ( n11364 & ~n26022 ) | ( n26018 & ~n26022 ) ;
  assign n26024 = n15523 ^ n2314 ^ 1'b0 ;
  assign n26025 = n25877 ^ n19304 ^ n4688 ;
  assign n26026 = n26024 | n26025 ;
  assign n26027 = n26026 ^ n1354 ^ x129 ;
  assign n26028 = ( x140 & n13293 ) | ( x140 & n26027 ) | ( n13293 & n26027 ) ;
  assign n26029 = n1014 & ~n14122 ;
  assign n26030 = n18956 ^ n18285 ^ 1'b0 ;
  assign n26031 = n534 & ~n26030 ;
  assign n26032 = n11164 & ~n18101 ;
  assign n26033 = ~n354 & n1378 ;
  assign n26034 = ~n6269 & n26033 ;
  assign n26035 = ( n5728 & n26032 ) | ( n5728 & ~n26034 ) | ( n26032 & ~n26034 ) ;
  assign n26036 = n1395 ^ n574 ^ 1'b0 ;
  assign n26037 = ~n8642 & n26036 ;
  assign n26038 = ~n21878 & n26037 ;
  assign n26039 = n471 & ~n26038 ;
  assign n26040 = n4566 ^ n1446 ^ 1'b0 ;
  assign n26041 = n26040 ^ n11116 ^ 1'b0 ;
  assign n26042 = n26041 ^ n2189 ^ 1'b0 ;
  assign n26043 = n26042 ^ n11304 ^ n5715 ;
  assign n26044 = ( n1449 & n23244 ) | ( n1449 & n26043 ) | ( n23244 & n26043 ) ;
  assign n26045 = n26044 ^ n23132 ^ 1'b0 ;
  assign n26048 = n18189 & n18781 ;
  assign n26049 = ~n18848 & n26048 ;
  assign n26046 = ( n1902 & n16225 ) | ( n1902 & ~n19530 ) | ( n16225 & ~n19530 ) ;
  assign n26047 = n4575 & n26046 ;
  assign n26050 = n26049 ^ n26047 ^ 1'b0 ;
  assign n26051 = ( n1903 & n2833 ) | ( n1903 & ~n19417 ) | ( n2833 & ~n19417 ) ;
  assign n26052 = n10995 ^ n9793 ^ n2634 ;
  assign n26053 = n13217 | n26052 ;
  assign n26054 = n26051 & ~n26053 ;
  assign n26055 = ~n10446 & n18545 ;
  assign n26056 = ~n11656 & n26055 ;
  assign n26057 = n26056 ^ n14981 ^ 1'b0 ;
  assign n26058 = ~n14532 & n26057 ;
  assign n26059 = ~n17563 & n26058 ;
  assign n26060 = n6823 ^ x44 ^ 1'b0 ;
  assign n26061 = n11301 ^ n7120 ^ n2858 ;
  assign n26062 = n26061 ^ n13536 ^ 1'b0 ;
  assign n26063 = ( ~n25666 & n26060 ) | ( ~n25666 & n26062 ) | ( n26060 & n26062 ) ;
  assign n26064 = ( n8247 & n14081 ) | ( n8247 & ~n26063 ) | ( n14081 & ~n26063 ) ;
  assign n26065 = n10393 ^ n5953 ^ 1'b0 ;
  assign n26066 = n12411 ^ n3050 ^ 1'b0 ;
  assign n26067 = n8790 & n26066 ;
  assign n26068 = ~n18264 & n26067 ;
  assign n26069 = n22590 ^ n15829 ^ n8091 ;
  assign n26070 = n1838 | n26069 ;
  assign n26071 = ~n21690 & n26070 ;
  assign n26072 = n19116 ^ n8069 ^ n4178 ;
  assign n26073 = n21494 ^ n20021 ^ n5231 ;
  assign n26074 = n4982 | n18942 ;
  assign n26075 = n26074 ^ n3717 ^ 1'b0 ;
  assign n26076 = n26075 ^ n10783 ^ n511 ;
  assign n26077 = ~n1345 & n10072 ;
  assign n26078 = n26077 ^ n14373 ^ 1'b0 ;
  assign n26079 = ( n1827 & n19357 ) | ( n1827 & ~n26078 ) | ( n19357 & ~n26078 ) ;
  assign n26080 = n26079 ^ n25034 ^ 1'b0 ;
  assign n26081 = n26076 & ~n26080 ;
  assign n26082 = n14979 | n23605 ;
  assign n26083 = n16663 ^ n4609 ^ n2646 ;
  assign n26084 = n26083 ^ n21759 ^ n13163 ;
  assign n26085 = ~n7943 & n9020 ;
  assign n26086 = ( ~n21706 & n22541 ) | ( ~n21706 & n26085 ) | ( n22541 & n26085 ) ;
  assign n26087 = ( n2564 & n7363 ) | ( n2564 & ~n18443 ) | ( n7363 & ~n18443 ) ;
  assign n26088 = ( x157 & n9112 ) | ( x157 & ~n11627 ) | ( n9112 & ~n11627 ) ;
  assign n26089 = n26088 ^ n20187 ^ 1'b0 ;
  assign n26090 = n25737 & n26089 ;
  assign n26091 = n19541 & n26090 ;
  assign n26092 = n7558 ^ n5347 ^ x125 ;
  assign n26093 = ( n8569 & ~n10806 ) | ( n8569 & n14276 ) | ( ~n10806 & n14276 ) ;
  assign n26096 = ( n1113 & n8268 ) | ( n1113 & n14290 ) | ( n8268 & n14290 ) ;
  assign n26094 = n22008 & n25385 ;
  assign n26095 = ~n7249 & n26094 ;
  assign n26097 = n26096 ^ n26095 ^ n289 ;
  assign n26098 = n3870 & n26097 ;
  assign n26099 = n26098 ^ n7903 ^ n1201 ;
  assign n26100 = n16890 ^ n3030 ^ 1'b0 ;
  assign n26101 = n19864 ^ n6290 ^ 1'b0 ;
  assign n26102 = n18161 & n26101 ;
  assign n26103 = n1400 & ~n2322 ;
  assign n26104 = n26103 ^ n8239 ^ 1'b0 ;
  assign n26105 = ~n13763 & n26104 ;
  assign n26106 = ~n14848 & n26105 ;
  assign n26107 = n14288 ^ n8970 ^ n8927 ;
  assign n26108 = n836 ^ n455 ^ 1'b0 ;
  assign n26109 = ~n26107 & n26108 ;
  assign n26110 = n6376 & n25184 ;
  assign n26111 = n26110 ^ n13201 ^ n5929 ;
  assign n26112 = n9588 ^ n2297 ^ 1'b0 ;
  assign n26113 = n26111 | n26112 ;
  assign n26114 = n9794 ^ n6931 ^ n6442 ;
  assign n26115 = ( x87 & n1280 ) | ( x87 & n5673 ) | ( n1280 & n5673 ) ;
  assign n26116 = n3163 & n26115 ;
  assign n26117 = n26114 | n26116 ;
  assign n26118 = n26117 ^ n16932 ^ 1'b0 ;
  assign n26119 = n7302 & ~n21448 ;
  assign n26120 = x183 & ~n5097 ;
  assign n26121 = ( n8941 & n14995 ) | ( n8941 & n26120 ) | ( n14995 & n26120 ) ;
  assign n26122 = n26121 ^ n2547 ^ 1'b0 ;
  assign n26123 = ( n4232 & n19120 ) | ( n4232 & n25930 ) | ( n19120 & n25930 ) ;
  assign n26124 = n26122 & ~n26123 ;
  assign n26125 = n26124 ^ n12311 ^ 1'b0 ;
  assign n26126 = n26119 | n26125 ;
  assign n26127 = n24818 ^ n2094 ^ 1'b0 ;
  assign n26128 = n26016 & ~n26127 ;
  assign n26129 = ( x10 & n1301 ) | ( x10 & n15631 ) | ( n1301 & n15631 ) ;
  assign n26130 = ( ~n1678 & n1684 ) | ( ~n1678 & n3422 ) | ( n1684 & n3422 ) ;
  assign n26131 = n26130 ^ n24522 ^ n5004 ;
  assign n26132 = n14741 ^ n6364 ^ 1'b0 ;
  assign n26133 = n17973 & ~n26132 ;
  assign n26134 = ( n12401 & n15389 ) | ( n12401 & n26133 ) | ( n15389 & n26133 ) ;
  assign n26135 = ( n15927 & n23207 ) | ( n15927 & ~n26134 ) | ( n23207 & ~n26134 ) ;
  assign n26136 = n24033 ^ n4769 ^ 1'b0 ;
  assign n26137 = n12859 ^ n11764 ^ 1'b0 ;
  assign n26138 = n1153 & ~n26137 ;
  assign n26139 = ( n23291 & n26136 ) | ( n23291 & n26138 ) | ( n26136 & n26138 ) ;
  assign n26140 = ~n21533 & n22703 ;
  assign n26141 = ~n19785 & n26140 ;
  assign n26142 = n14587 ^ n12184 ^ n11138 ;
  assign n26143 = ~n18922 & n26142 ;
  assign n26144 = n10815 ^ x3 ^ 1'b0 ;
  assign n26145 = ~n2871 & n26144 ;
  assign n26146 = n11959 & n26145 ;
  assign n26147 = n26146 ^ n5021 ^ 1'b0 ;
  assign n26148 = n316 | n4059 ;
  assign n26149 = ( ~n26143 & n26147 ) | ( ~n26143 & n26148 ) | ( n26147 & n26148 ) ;
  assign n26150 = ~n5276 & n6816 ;
  assign n26151 = n26150 ^ n6869 ^ 1'b0 ;
  assign n26152 = ( n413 & n3228 ) | ( n413 & ~n5037 ) | ( n3228 & ~n5037 ) ;
  assign n26153 = n5140 & ~n26152 ;
  assign n26154 = ( ~n8702 & n26151 ) | ( ~n8702 & n26153 ) | ( n26151 & n26153 ) ;
  assign n26155 = ( n10519 & n16552 ) | ( n10519 & n26154 ) | ( n16552 & n26154 ) ;
  assign n26156 = ~n12428 & n26155 ;
  assign n26157 = n5381 ^ n4062 ^ 1'b0 ;
  assign n26158 = n26157 ^ n9067 ^ 1'b0 ;
  assign n26159 = n14179 ^ n6260 ^ n725 ;
  assign n26160 = n26159 ^ n25942 ^ n2642 ;
  assign n26161 = ( n3059 & n5019 ) | ( n3059 & n8990 ) | ( n5019 & n8990 ) ;
  assign n26162 = n6077 & ~n26161 ;
  assign n26163 = n26162 ^ n25445 ^ n15078 ;
  assign n26164 = n9020 ^ n2515 ^ 1'b0 ;
  assign n26165 = n3214 | n26164 ;
  assign n26166 = ( n10364 & n18906 ) | ( n10364 & n26165 ) | ( n18906 & n26165 ) ;
  assign n26167 = n4452 ^ n1231 ^ 1'b0 ;
  assign n26168 = n1953 & ~n26167 ;
  assign n26169 = ( x40 & n15953 ) | ( x40 & ~n26168 ) | ( n15953 & ~n26168 ) ;
  assign n26172 = ( ~n749 & n1198 ) | ( ~n749 & n5070 ) | ( n1198 & n5070 ) ;
  assign n26170 = n6693 & ~n19184 ;
  assign n26171 = n26170 ^ n5680 ^ 1'b0 ;
  assign n26173 = n26172 ^ n26171 ^ n4652 ;
  assign n26174 = n1158 & ~n6624 ;
  assign n26175 = n26174 ^ n290 ^ 1'b0 ;
  assign n26176 = n15767 | n26175 ;
  assign n26177 = n26173 | n26176 ;
  assign n26178 = n2607 | n15676 ;
  assign n26179 = n26178 ^ n13480 ^ 1'b0 ;
  assign n26180 = n5035 & ~n23759 ;
  assign n26181 = n7919 ^ n7862 ^ 1'b0 ;
  assign n26182 = ( n925 & ~n4080 ) | ( n925 & n8536 ) | ( ~n4080 & n8536 ) ;
  assign n26183 = n26182 ^ n11458 ^ 1'b0 ;
  assign n26184 = ( n5336 & ~n10820 ) | ( n5336 & n26183 ) | ( ~n10820 & n26183 ) ;
  assign n26185 = n12959 ^ n7878 ^ 1'b0 ;
  assign n26186 = ~n7669 & n26185 ;
  assign n26187 = n26186 ^ n6331 ^ 1'b0 ;
  assign n26188 = ( n5353 & n13223 ) | ( n5353 & n24690 ) | ( n13223 & n24690 ) ;
  assign n26189 = n2606 & ~n26188 ;
  assign n26190 = n3962 & n16626 ;
  assign n26191 = ~x41 & n26190 ;
  assign n26192 = n6803 | n8949 ;
  assign n26193 = ( n584 & n14811 ) | ( n584 & ~n26192 ) | ( n14811 & ~n26192 ) ;
  assign n26194 = ( ~n11248 & n19189 ) | ( ~n11248 & n26193 ) | ( n19189 & n26193 ) ;
  assign n26195 = n3177 | n26194 ;
  assign n26198 = n11294 & n25874 ;
  assign n26199 = n1766 & n20876 ;
  assign n26200 = ~n26198 & n26199 ;
  assign n26201 = n12784 & n26200 ;
  assign n26202 = n25713 ^ n21724 ^ n6906 ;
  assign n26203 = ( n9420 & n26201 ) | ( n9420 & ~n26202 ) | ( n26201 & ~n26202 ) ;
  assign n26196 = n6365 ^ n5355 ^ 1'b0 ;
  assign n26197 = n3887 | n26196 ;
  assign n26204 = n26203 ^ n26197 ^ 1'b0 ;
  assign n26205 = n16291 ^ n4332 ^ 1'b0 ;
  assign n26206 = n3026 ^ n333 ^ 1'b0 ;
  assign n26207 = n2262 & ~n14228 ;
  assign n26208 = n26207 ^ n9363 ^ 1'b0 ;
  assign n26209 = ( ~n3366 & n3891 ) | ( ~n3366 & n4393 ) | ( n3891 & n4393 ) ;
  assign n26210 = n26208 & ~n26209 ;
  assign n26211 = ( n2785 & ~n22191 ) | ( n2785 & n24795 ) | ( ~n22191 & n24795 ) ;
  assign n26212 = ( n15556 & n22713 ) | ( n15556 & n26211 ) | ( n22713 & n26211 ) ;
  assign n26213 = ~n8490 & n26212 ;
  assign n26214 = n26213 ^ n10307 ^ 1'b0 ;
  assign n26216 = n8344 & n24368 ;
  assign n26215 = ~n11590 & n14634 ;
  assign n26217 = n26216 ^ n26215 ^ 1'b0 ;
  assign n26218 = ~n3909 & n22096 ;
  assign n26219 = n2441 & ~n5025 ;
  assign n26220 = n9056 | n26219 ;
  assign n26221 = ( n15564 & n22575 ) | ( n15564 & n26220 ) | ( n22575 & n26220 ) ;
  assign n26222 = n2510 & ~n21291 ;
  assign n26223 = n12030 & n26222 ;
  assign n26224 = n554 | n10566 ;
  assign n26225 = n905 & ~n26224 ;
  assign n26226 = n26225 ^ n16199 ^ 1'b0 ;
  assign n26227 = n11481 & n26226 ;
  assign n26228 = n26227 ^ n1660 ^ 1'b0 ;
  assign n26229 = n22014 ^ n16807 ^ n16417 ;
  assign n26230 = n3117 | n5263 ;
  assign n26231 = ( ~n7315 & n26229 ) | ( ~n7315 & n26230 ) | ( n26229 & n26230 ) ;
  assign n26232 = ~n1873 & n4040 ;
  assign n26233 = ~n4178 & n26232 ;
  assign n26234 = n18803 | n26233 ;
  assign n26235 = n26231 & ~n26234 ;
  assign n26236 = ( n5193 & n13042 ) | ( n5193 & ~n26235 ) | ( n13042 & ~n26235 ) ;
  assign n26237 = n20701 ^ n12470 ^ n2741 ;
  assign n26238 = ~n20501 & n21572 ;
  assign n26239 = n26238 ^ n24955 ^ 1'b0 ;
  assign n26240 = ( n9159 & ~n13679 ) | ( n9159 & n24154 ) | ( ~n13679 & n24154 ) ;
  assign n26241 = n4713 & ~n11693 ;
  assign n26242 = n26241 ^ n25908 ^ n16776 ;
  assign n26243 = n19787 ^ n13923 ^ n1133 ;
  assign n26244 = n11885 & n24851 ;
  assign n26245 = n7709 | n26244 ;
  assign n26246 = n22923 & ~n26245 ;
  assign n26247 = n18795 ^ n15532 ^ n3348 ;
  assign n26248 = ( n18842 & ~n26246 ) | ( n18842 & n26247 ) | ( ~n26246 & n26247 ) ;
  assign n26249 = n14131 | n22756 ;
  assign n26250 = n5074 | n26249 ;
  assign n26251 = ( ~n5307 & n13234 ) | ( ~n5307 & n26250 ) | ( n13234 & n26250 ) ;
  assign n26252 = ( n12053 & n15074 ) | ( n12053 & ~n26251 ) | ( n15074 & ~n26251 ) ;
  assign n26253 = n24895 ^ n13932 ^ n6574 ;
  assign n26254 = n2782 | n8427 ;
  assign n26255 = n4139 | n26254 ;
  assign n26256 = n8603 & n9484 ;
  assign n26257 = n26256 ^ x29 ^ 1'b0 ;
  assign n26258 = n2575 & ~n26257 ;
  assign n26259 = ~n13921 & n26258 ;
  assign n26260 = n4107 | n24762 ;
  assign n26261 = ( n5982 & ~n7221 ) | ( n5982 & n10170 ) | ( ~n7221 & n10170 ) ;
  assign n26262 = n26261 ^ n24488 ^ n17252 ;
  assign n26263 = n26262 ^ n10451 ^ 1'b0 ;
  assign n26264 = ( ~n5229 & n19895 ) | ( ~n5229 & n20630 ) | ( n19895 & n20630 ) ;
  assign n26265 = ( n8090 & n20247 ) | ( n8090 & n26264 ) | ( n20247 & n26264 ) ;
  assign n26273 = n5300 ^ n3831 ^ 1'b0 ;
  assign n26266 = ( n1244 & n14489 ) | ( n1244 & n19366 ) | ( n14489 & n19366 ) ;
  assign n26267 = ~n17203 & n26266 ;
  assign n26268 = n26267 ^ n18723 ^ 1'b0 ;
  assign n26269 = x29 & ~n8235 ;
  assign n26270 = n26269 ^ n16738 ^ 1'b0 ;
  assign n26271 = n16042 & n26270 ;
  assign n26272 = ~n26268 & n26271 ;
  assign n26274 = n26273 ^ n26272 ^ n7071 ;
  assign n26275 = n5894 | n19657 ;
  assign n26276 = n9992 ^ n1428 ^ 1'b0 ;
  assign n26277 = n18209 ^ x18 ^ 1'b0 ;
  assign n26278 = ( ~n15113 & n18854 ) | ( ~n15113 & n26277 ) | ( n18854 & n26277 ) ;
  assign n26279 = ~n26276 & n26278 ;
  assign n26280 = ~n6784 & n26279 ;
  assign n26281 = n17396 ^ n8083 ^ n4740 ;
  assign n26283 = n18457 ^ n11309 ^ 1'b0 ;
  assign n26282 = n18525 ^ n15835 ^ 1'b0 ;
  assign n26284 = n26283 ^ n26282 ^ n19951 ;
  assign n26285 = n21233 ^ n2846 ^ 1'b0 ;
  assign n26286 = ~n7926 & n26285 ;
  assign n26293 = x250 & n3459 ;
  assign n26294 = n23484 ^ n12020 ^ 1'b0 ;
  assign n26295 = n26293 & n26294 ;
  assign n26288 = ( ~n8091 & n8301 ) | ( ~n8091 & n9293 ) | ( n8301 & n9293 ) ;
  assign n26289 = ~n4556 & n13549 ;
  assign n26290 = n15922 | n26289 ;
  assign n26291 = n11048 | n26290 ;
  assign n26292 = n26288 & n26291 ;
  assign n26296 = n26295 ^ n26292 ^ 1'b0 ;
  assign n26287 = x122 & ~n23702 ;
  assign n26297 = n26296 ^ n26287 ^ 1'b0 ;
  assign n26298 = ~n4254 & n12007 ;
  assign n26299 = n26298 ^ n8655 ^ 1'b0 ;
  assign n26300 = n11841 ^ n1775 ^ 1'b0 ;
  assign n26301 = n6228 | n7200 ;
  assign n26302 = n26301 ^ n13200 ^ 1'b0 ;
  assign n26303 = n19112 ^ n9829 ^ n2972 ;
  assign n26304 = n20076 ^ n4748 ^ 1'b0 ;
  assign n26305 = n26303 & n26304 ;
  assign n26306 = n15687 | n19876 ;
  assign n26307 = n26305 | n26306 ;
  assign n26308 = ( n8399 & ~n26302 ) | ( n8399 & n26307 ) | ( ~n26302 & n26307 ) ;
  assign n26309 = ~n2694 & n7401 ;
  assign n26310 = n18226 ^ n615 ^ 1'b0 ;
  assign n26311 = n7324 & n9729 ;
  assign n26312 = n26311 ^ n4291 ^ 1'b0 ;
  assign n26313 = n5954 | n26312 ;
  assign n26314 = n7672 | n26313 ;
  assign n26315 = n11438 | n26314 ;
  assign n26316 = ~n13141 & n26315 ;
  assign n26317 = ( n6681 & n15795 ) | ( n6681 & ~n18443 ) | ( n15795 & ~n18443 ) ;
  assign n26319 = n13039 ^ n9440 ^ 1'b0 ;
  assign n26318 = ~n1004 & n1785 ;
  assign n26320 = n26319 ^ n26318 ^ 1'b0 ;
  assign n26321 = n21893 ^ n13579 ^ n987 ;
  assign n26322 = n3466 & n6380 ;
  assign n26323 = n8496 & n26322 ;
  assign n26324 = ( ~n4785 & n19121 ) | ( ~n4785 & n26323 ) | ( n19121 & n26323 ) ;
  assign n26325 = ( n4830 & n14255 ) | ( n4830 & ~n26324 ) | ( n14255 & ~n26324 ) ;
  assign n26326 = n21460 ^ n16496 ^ 1'b0 ;
  assign n26327 = n409 | n26326 ;
  assign n26328 = ~n3467 & n4061 ;
  assign n26329 = n26328 ^ n295 ^ 1'b0 ;
  assign n26330 = n26329 ^ n22645 ^ 1'b0 ;
  assign n26331 = n1599 & ~n12427 ;
  assign n26332 = n26331 ^ n2007 ^ 1'b0 ;
  assign n26333 = ( n12631 & ~n15199 ) | ( n12631 & n26332 ) | ( ~n15199 & n26332 ) ;
  assign n26337 = ( n8214 & n10404 ) | ( n8214 & ~n10855 ) | ( n10404 & ~n10855 ) ;
  assign n26335 = n11819 | n14892 ;
  assign n26336 = n26335 ^ n3156 ^ n1352 ;
  assign n26334 = n16477 & ~n21831 ;
  assign n26338 = n26337 ^ n26336 ^ n26334 ;
  assign n26339 = n26338 ^ n25349 ^ n6352 ;
  assign n26340 = ~n768 & n14478 ;
  assign n26341 = n13330 ^ n2978 ^ 1'b0 ;
  assign n26342 = n10150 | n26341 ;
  assign n26343 = n26342 ^ n15986 ^ n988 ;
  assign n26344 = ( n1734 & ~n22641 ) | ( n1734 & n26343 ) | ( ~n22641 & n26343 ) ;
  assign n26345 = ( x238 & n5539 ) | ( x238 & n26344 ) | ( n5539 & n26344 ) ;
  assign n26346 = ~n4319 & n12212 ;
  assign n26347 = n26346 ^ n11307 ^ 1'b0 ;
  assign n26348 = ( n722 & n4382 ) | ( n722 & n4827 ) | ( n4382 & n4827 ) ;
  assign n26349 = n26348 ^ n17079 ^ 1'b0 ;
  assign n26350 = ~n6022 & n26349 ;
  assign n26351 = x89 & ~n23207 ;
  assign n26352 = n26351 ^ n915 ^ 1'b0 ;
  assign n26353 = n9073 ^ n5741 ^ 1'b0 ;
  assign n26354 = n6163 | n26353 ;
  assign n26355 = ( x205 & n26352 ) | ( x205 & n26354 ) | ( n26352 & n26354 ) ;
  assign n26356 = n18320 ^ n2732 ^ 1'b0 ;
  assign n26357 = n8423 | n26356 ;
  assign n26358 = n1452 & n26357 ;
  assign n26359 = n26358 ^ n14251 ^ 1'b0 ;
  assign n26360 = ( n4660 & n4881 ) | ( n4660 & ~n13526 ) | ( n4881 & ~n13526 ) ;
  assign n26361 = n7779 & ~n24639 ;
  assign n26362 = ~n2356 & n7578 ;
  assign n26363 = n26362 ^ n2937 ^ 1'b0 ;
  assign n26364 = n26363 ^ n13363 ^ 1'b0 ;
  assign n26365 = ( ~n8558 & n16994 ) | ( ~n8558 & n18283 ) | ( n16994 & n18283 ) ;
  assign n26366 = n12300 | n15768 ;
  assign n26367 = n26365 | n26366 ;
  assign n26368 = n12000 & ~n18266 ;
  assign n26369 = n13580 ^ n8194 ^ 1'b0 ;
  assign n26370 = n1194 & ~n2105 ;
  assign n26371 = n26370 ^ n9423 ^ 1'b0 ;
  assign n26372 = ~n13766 & n26371 ;
  assign n26373 = ~n3022 & n26372 ;
  assign n26374 = ~n26369 & n26373 ;
  assign n26375 = n10181 ^ n4600 ^ n3387 ;
  assign n26376 = ( ~x115 & n17410 ) | ( ~x115 & n26375 ) | ( n17410 & n26375 ) ;
  assign n26377 = n9417 ^ n8810 ^ n320 ;
  assign n26378 = x120 & n26377 ;
  assign n26379 = ( n744 & n14906 ) | ( n744 & n26378 ) | ( n14906 & n26378 ) ;
  assign n26380 = ~n6438 & n26379 ;
  assign n26381 = n16957 & n26380 ;
  assign n26382 = n22584 & ~n26381 ;
  assign n26383 = n26376 & n26382 ;
  assign n26384 = n6854 & n22164 ;
  assign n26385 = n11251 ^ n10318 ^ n8646 ;
  assign n26386 = n26385 ^ n2607 ^ n2097 ;
  assign n26387 = ~n2911 & n21910 ;
  assign n26388 = n26387 ^ n3585 ^ 1'b0 ;
  assign n26389 = ( n4593 & ~n8069 ) | ( n4593 & n26388 ) | ( ~n8069 & n26388 ) ;
  assign n26390 = n26389 ^ n16006 ^ n5008 ;
  assign n26391 = ( n8006 & ~n8881 ) | ( n8006 & n14485 ) | ( ~n8881 & n14485 ) ;
  assign n26392 = n10363 | n25204 ;
  assign n26393 = n1535 & ~n26392 ;
  assign n26394 = n18652 ^ n3506 ^ 1'b0 ;
  assign n26395 = ( n9069 & ~n26393 ) | ( n9069 & n26394 ) | ( ~n26393 & n26394 ) ;
  assign n26396 = ~n10434 & n16374 ;
  assign n26397 = ~n17476 & n26396 ;
  assign n26398 = ~n16890 & n26397 ;
  assign n26399 = n4154 & ~n15030 ;
  assign n26400 = n15177 & n26399 ;
  assign n26401 = n8735 & ~n14051 ;
  assign n26402 = n23633 ^ n16883 ^ 1'b0 ;
  assign n26403 = n11411 & n26402 ;
  assign n26404 = ~n3521 & n23035 ;
  assign n26405 = n1631 & ~n26404 ;
  assign n26406 = n5716 & n24226 ;
  assign n26407 = n26406 ^ n2192 ^ 1'b0 ;
  assign n26408 = n4546 | n26407 ;
  assign n26409 = n13546 & ~n26408 ;
  assign n26410 = n26405 & n26409 ;
  assign n26411 = n14254 ^ n5566 ^ 1'b0 ;
  assign n26412 = ~n11324 & n26411 ;
  assign n26413 = n15621 ^ n4705 ^ 1'b0 ;
  assign n26414 = n12210 & n26413 ;
  assign n26415 = n12315 & n26414 ;
  assign n26416 = ~n26412 & n26415 ;
  assign n26417 = n24448 ^ n13452 ^ n12470 ;
  assign n26418 = n26417 ^ n14821 ^ n7300 ;
  assign n26419 = n22292 ^ n8853 ^ 1'b0 ;
  assign n26420 = n18806 ^ n5040 ^ 1'b0 ;
  assign n26421 = n6701 & n8814 ;
  assign n26422 = n660 & n26421 ;
  assign n26423 = n26422 ^ n2903 ^ 1'b0 ;
  assign n26424 = n26423 ^ n18636 ^ 1'b0 ;
  assign n26425 = n22333 & ~n26424 ;
  assign n26426 = n12046 ^ n5902 ^ 1'b0 ;
  assign n26427 = n16234 ^ n6763 ^ n3268 ;
  assign n26428 = ~n17218 & n25858 ;
  assign n26429 = n11553 ^ n8295 ^ 1'b0 ;
  assign n26430 = n19531 | n26429 ;
  assign n26431 = ( n1629 & n14680 ) | ( n1629 & ~n26430 ) | ( n14680 & ~n26430 ) ;
  assign n26433 = n24040 ^ n2909 ^ 1'b0 ;
  assign n26434 = n9374 & n26433 ;
  assign n26432 = n20789 ^ n18474 ^ n7000 ;
  assign n26435 = n26434 ^ n26432 ^ 1'b0 ;
  assign n26436 = n4432 | n26435 ;
  assign n26437 = n26436 ^ n10922 ^ 1'b0 ;
  assign n26438 = n24611 ^ n8924 ^ n3395 ;
  assign n26439 = n9278 & ~n26438 ;
  assign n26440 = n26439 ^ n8430 ^ 1'b0 ;
  assign n26441 = ( ~n3527 & n7561 ) | ( ~n3527 & n14704 ) | ( n7561 & n14704 ) ;
  assign n26442 = n20942 & n26441 ;
  assign n26444 = ( ~n7617 & n7940 ) | ( ~n7617 & n8916 ) | ( n7940 & n8916 ) ;
  assign n26445 = ( n1775 & n11208 ) | ( n1775 & n26444 ) | ( n11208 & n26444 ) ;
  assign n26443 = ~n8136 & n8159 ;
  assign n26446 = n26445 ^ n26443 ^ n20750 ;
  assign n26447 = n12295 & ~n17840 ;
  assign n26448 = ~n17789 & n26447 ;
  assign n26449 = ( n1438 & n2532 ) | ( n1438 & n26448 ) | ( n2532 & n26448 ) ;
  assign n26450 = n9298 ^ n7833 ^ n363 ;
  assign n26451 = n13961 ^ n2947 ^ 1'b0 ;
  assign n26452 = n19647 ^ n1502 ^ 1'b0 ;
  assign n26453 = n9754 & n26452 ;
  assign n26454 = x49 & ~n12132 ;
  assign n26455 = n26454 ^ n1294 ^ 1'b0 ;
  assign n26456 = n3068 & n26455 ;
  assign n26457 = n24868 & n26456 ;
  assign n26458 = n18642 ^ n11771 ^ 1'b0 ;
  assign n26459 = ~n4590 & n26458 ;
  assign n26460 = ~n17091 & n26459 ;
  assign n26461 = ~n26457 & n26460 ;
  assign n26462 = ~n12488 & n26461 ;
  assign n26463 = x134 & n11941 ;
  assign n26464 = n26463 ^ n1502 ^ 1'b0 ;
  assign n26465 = n26464 ^ n23769 ^ n751 ;
  assign n26466 = n11565 ^ x10 ^ 1'b0 ;
  assign n26467 = n23807 & n26466 ;
  assign n26468 = n26467 ^ n11140 ^ 1'b0 ;
  assign n26469 = n1043 & ~n3682 ;
  assign n26470 = n611 & n26469 ;
  assign n26471 = n26470 ^ n10850 ^ n2939 ;
  assign n26472 = n16333 ^ n8983 ^ n4011 ;
  assign n26473 = n26471 & ~n26472 ;
  assign n26474 = n6852 ^ n4518 ^ 1'b0 ;
  assign n26475 = ~n3496 & n26474 ;
  assign n26476 = n12389 ^ n2924 ^ 1'b0 ;
  assign n26477 = n26475 | n26476 ;
  assign n26478 = n5138 & ~n10212 ;
  assign n26479 = n26478 ^ n16758 ^ x72 ;
  assign n26480 = ( n6520 & ~n6560 ) | ( n6520 & n26479 ) | ( ~n6560 & n26479 ) ;
  assign n26481 = n9615 ^ n7904 ^ 1'b0 ;
  assign n26482 = n24599 ^ n13054 ^ 1'b0 ;
  assign n26483 = ( ~n12484 & n21743 ) | ( ~n12484 & n26482 ) | ( n21743 & n26482 ) ;
  assign n26484 = n24905 ^ n14936 ^ 1'b0 ;
  assign n26485 = n16067 & n26484 ;
  assign n26486 = n26483 & ~n26485 ;
  assign n26487 = n1913 & n3145 ;
  assign n26488 = n2633 & n26487 ;
  assign n26489 = n26488 ^ n11741 ^ 1'b0 ;
  assign n26490 = n26489 ^ n1264 ^ 1'b0 ;
  assign n26491 = ~n3992 & n17105 ;
  assign n26492 = ~n10215 & n26491 ;
  assign n26493 = n25115 | n26492 ;
  assign n26494 = n13957 & ~n26493 ;
  assign n26495 = n15252 | n20556 ;
  assign n26496 = n3186 & ~n26495 ;
  assign n26498 = ~n23626 & n25821 ;
  assign n26497 = n3037 & n11722 ;
  assign n26499 = n26498 ^ n26497 ^ 1'b0 ;
  assign n26500 = n17851 ^ n15989 ^ 1'b0 ;
  assign n26501 = ~n9469 & n26500 ;
  assign n26502 = n26501 ^ n18881 ^ 1'b0 ;
  assign n26503 = n6991 | n17756 ;
  assign n26504 = n26503 ^ n7510 ^ 1'b0 ;
  assign n26505 = n26504 ^ n17494 ^ n10870 ;
  assign n26506 = ( n783 & ~n20727 ) | ( n783 & n26505 ) | ( ~n20727 & n26505 ) ;
  assign n26507 = n4548 ^ n1650 ^ 1'b0 ;
  assign n26508 = ( n1591 & n11168 ) | ( n1591 & ~n26507 ) | ( n11168 & ~n26507 ) ;
  assign n26509 = n841 & n2750 ;
  assign n26510 = n26509 ^ n771 ^ 1'b0 ;
  assign n26511 = ~n16855 & n26510 ;
  assign n26512 = n4045 & ~n20501 ;
  assign n26513 = ( ~n16024 & n26511 ) | ( ~n16024 & n26512 ) | ( n26511 & n26512 ) ;
  assign n26515 = n6132 & n13819 ;
  assign n26516 = n26515 ^ n16075 ^ 1'b0 ;
  assign n26514 = n1552 & n3752 ;
  assign n26517 = n26516 ^ n26514 ^ 1'b0 ;
  assign n26518 = ( n9842 & ~n15943 ) | ( n9842 & n19496 ) | ( ~n15943 & n19496 ) ;
  assign n26519 = n26518 ^ n3424 ^ 1'b0 ;
  assign n26520 = n26519 ^ n19799 ^ 1'b0 ;
  assign n26521 = n2566 | n13330 ;
  assign n26522 = n26521 ^ n3157 ^ 1'b0 ;
  assign n26523 = ~n1834 & n3377 ;
  assign n26524 = ~n15587 & n26523 ;
  assign n26525 = n1511 | n8607 ;
  assign n26526 = n13227 & ~n26525 ;
  assign n26527 = n26526 ^ n13780 ^ n8734 ;
  assign n26528 = n26524 | n26527 ;
  assign n26529 = n26522 & ~n26528 ;
  assign n26530 = ~n24749 & n26529 ;
  assign n26531 = n10401 ^ n9108 ^ 1'b0 ;
  assign n26532 = ~n26530 & n26531 ;
  assign n26533 = n26532 ^ n898 ^ 1'b0 ;
  assign n26534 = x206 & n2456 ;
  assign n26535 = n3044 & n26534 ;
  assign n26536 = n4873 ^ n1352 ^ n510 ;
  assign n26537 = ( n10478 & n26535 ) | ( n10478 & ~n26536 ) | ( n26535 & ~n26536 ) ;
  assign n26538 = n26537 ^ n22977 ^ 1'b0 ;
  assign n26539 = n19888 ^ n9139 ^ 1'b0 ;
  assign n26540 = ( ~n3070 & n3639 ) | ( ~n3070 & n5309 ) | ( n3639 & n5309 ) ;
  assign n26541 = n1966 & ~n26540 ;
  assign n26542 = ( n4322 & ~n15860 ) | ( n4322 & n17497 ) | ( ~n15860 & n17497 ) ;
  assign n26543 = n26542 ^ n276 ^ 1'b0 ;
  assign n26544 = n26543 ^ n7562 ^ 1'b0 ;
  assign n26545 = n25396 ^ n19985 ^ n14371 ;
  assign n26546 = n21797 | n26545 ;
  assign n26547 = n22226 ^ n5524 ^ n5116 ;
  assign n26549 = ( n2764 & ~n6557 ) | ( n2764 & n6777 ) | ( ~n6557 & n6777 ) ;
  assign n26548 = n3830 | n12952 ;
  assign n26550 = n26549 ^ n26548 ^ 1'b0 ;
  assign n26551 = n7390 | n8671 ;
  assign n26552 = n26551 ^ n17427 ^ 1'b0 ;
  assign n26553 = ~n5905 & n26552 ;
  assign n26554 = ~n1886 & n21496 ;
  assign n26555 = n9097 | n13573 ;
  assign n26556 = n11146 & ~n26555 ;
  assign n26558 = ~n642 & n1301 ;
  assign n26559 = n26558 ^ n5900 ^ 1'b0 ;
  assign n26557 = n8785 & ~n15169 ;
  assign n26560 = n26559 ^ n26557 ^ 1'b0 ;
  assign n26561 = ~n11024 & n26560 ;
  assign n26562 = n26556 & n26561 ;
  assign n26563 = n11157 | n26562 ;
  assign n26564 = n19153 ^ n1750 ^ 1'b0 ;
  assign n26565 = ( n1430 & n5766 ) | ( n1430 & n7117 ) | ( n5766 & n7117 ) ;
  assign n26566 = n26564 & n26565 ;
  assign n26567 = n26566 ^ n10004 ^ 1'b0 ;
  assign n26568 = ~n20035 & n26567 ;
  assign n26569 = n26568 ^ n10152 ^ 1'b0 ;
  assign n26570 = n26563 | n26569 ;
  assign n26571 = n6860 & n23247 ;
  assign n26572 = n26571 ^ n14258 ^ 1'b0 ;
  assign n26573 = n26572 ^ n5486 ^ 1'b0 ;
  assign n26574 = ( n8162 & n20999 ) | ( n8162 & n26573 ) | ( n20999 & n26573 ) ;
  assign n26575 = ( n9289 & ~n10901 ) | ( n9289 & n15120 ) | ( ~n10901 & n15120 ) ;
  assign n26576 = n2075 | n26575 ;
  assign n26577 = n8808 & ~n13807 ;
  assign n26578 = ~n17072 & n26577 ;
  assign n26579 = ( n5671 & n10929 ) | ( n5671 & ~n17742 ) | ( n10929 & ~n17742 ) ;
  assign n26580 = n2241 | n13942 ;
  assign n26581 = n26580 ^ n2361 ^ 1'b0 ;
  assign n26582 = n26581 ^ n18538 ^ 1'b0 ;
  assign n26583 = n6777 | n12699 ;
  assign n26584 = n262 & ~n15820 ;
  assign n26585 = ~n22932 & n26584 ;
  assign n26586 = n10257 & n12084 ;
  assign n26587 = n26586 ^ n1061 ^ 1'b0 ;
  assign n26588 = n4596 | n26587 ;
  assign n26589 = n10827 & ~n26588 ;
  assign n26590 = n3742 & n15254 ;
  assign n26591 = ~n7980 & n26590 ;
  assign n26592 = n14180 ^ x228 ^ 1'b0 ;
  assign n26593 = ~n3488 & n6294 ;
  assign n26594 = n26592 | n26593 ;
  assign n26595 = n26591 & ~n26594 ;
  assign n26596 = ( ~n2680 & n9986 ) | ( ~n2680 & n19953 ) | ( n9986 & n19953 ) ;
  assign n26597 = n14062 ^ x85 ^ 1'b0 ;
  assign n26598 = n14172 ^ n2971 ^ 1'b0 ;
  assign n26599 = n10968 | n26598 ;
  assign n26600 = n22847 ^ n5493 ^ n2593 ;
  assign n26601 = n26600 ^ n11541 ^ 1'b0 ;
  assign n26602 = n22117 & ~n26601 ;
  assign n26603 = n9733 & n24233 ;
  assign n26604 = ~n13188 & n26603 ;
  assign n26605 = ~n26602 & n26604 ;
  assign n26606 = n3591 & ~n15722 ;
  assign n26607 = n6872 ^ n1743 ^ 1'b0 ;
  assign n26608 = n8392 & ~n26607 ;
  assign n26609 = n26608 ^ n8455 ^ n2530 ;
  assign n26610 = n24569 ^ n9520 ^ n873 ;
  assign n26611 = n26610 ^ n2127 ^ 1'b0 ;
  assign n26612 = n26609 | n26611 ;
  assign n26613 = n12946 ^ n8917 ^ 1'b0 ;
  assign n26614 = n26613 ^ n305 ^ 1'b0 ;
  assign n26615 = ( n26606 & n26612 ) | ( n26606 & n26614 ) | ( n26612 & n26614 ) ;
  assign n26616 = n2723 & n10133 ;
  assign n26617 = n26616 ^ n25314 ^ 1'b0 ;
  assign n26618 = ( x244 & n14474 ) | ( x244 & n26617 ) | ( n14474 & n26617 ) ;
  assign n26619 = n22938 ^ n2771 ^ n1391 ;
  assign n26620 = n26619 ^ n5443 ^ 1'b0 ;
  assign n26621 = n2142 | n16325 ;
  assign n26622 = n4450 ^ n4054 ^ 1'b0 ;
  assign n26623 = n26621 & n26622 ;
  assign n26624 = n12500 ^ n5061 ^ 1'b0 ;
  assign n26625 = n22561 ^ n20134 ^ 1'b0 ;
  assign n26626 = ~n10018 & n26625 ;
  assign n26627 = n17898 & ~n26626 ;
  assign n26628 = n9988 | n13624 ;
  assign n26629 = n10371 ^ n7240 ^ 1'b0 ;
  assign n26630 = ~n4311 & n14805 ;
  assign n26631 = n14189 ^ n13718 ^ n360 ;
  assign n26632 = n8882 & ~n26631 ;
  assign n26633 = n25339 ^ n6679 ^ 1'b0 ;
  assign n26634 = n21020 & ~n26633 ;
  assign n26637 = ~x65 & n9319 ;
  assign n26635 = n9379 ^ n2704 ^ 1'b0 ;
  assign n26636 = x218 & n26635 ;
  assign n26638 = n26637 ^ n26636 ^ 1'b0 ;
  assign n26639 = n25184 ^ n14983 ^ n12990 ;
  assign n26640 = n26639 ^ n23310 ^ 1'b0 ;
  assign n26641 = n3880 | n26640 ;
  assign n26642 = n6056 | n26641 ;
  assign n26643 = ( n5659 & n6955 ) | ( n5659 & ~n21562 ) | ( n6955 & ~n21562 ) ;
  assign n26644 = n4412 & n17087 ;
  assign n26645 = ( n15678 & n26643 ) | ( n15678 & n26644 ) | ( n26643 & n26644 ) ;
  assign n26646 = n13526 | n26645 ;
  assign n26647 = ~n23954 & n26216 ;
  assign n26648 = n4987 ^ x0 ^ 1'b0 ;
  assign n26649 = n26648 ^ n16075 ^ n5737 ;
  assign n26650 = n2803 & n19289 ;
  assign n26651 = n18743 | n22452 ;
  assign n26652 = n26650 & ~n26651 ;
  assign n26653 = ( n324 & ~n516 ) | ( n324 & n2828 ) | ( ~n516 & n2828 ) ;
  assign n26654 = n26653 ^ n2952 ^ 1'b0 ;
  assign n26655 = n17754 & ~n26654 ;
  assign n26656 = ( n11248 & ~n17162 ) | ( n11248 & n26655 ) | ( ~n17162 & n26655 ) ;
  assign n26657 = n2092 & ~n26656 ;
  assign n26658 = n26657 ^ n12270 ^ 1'b0 ;
  assign n26659 = n22981 & ~n24206 ;
  assign n26660 = n1793 & ~n26659 ;
  assign n26661 = n17312 ^ n7524 ^ n3000 ;
  assign n26662 = ( n10542 & n19278 ) | ( n10542 & ~n26661 ) | ( n19278 & ~n26661 ) ;
  assign n26663 = n10617 ^ n3096 ^ x244 ;
  assign n26664 = ~n16922 & n21820 ;
  assign n26665 = ~n26663 & n26664 ;
  assign n26666 = n13278 & n25554 ;
  assign n26667 = n5207 & n26666 ;
  assign n26674 = ( n2308 & ~n3460 ) | ( n2308 & n4877 ) | ( ~n3460 & n4877 ) ;
  assign n26668 = n11661 ^ n7252 ^ 1'b0 ;
  assign n26669 = n9052 & ~n26668 ;
  assign n26670 = ~n18575 & n26669 ;
  assign n26671 = n26670 ^ n2630 ^ 1'b0 ;
  assign n26672 = n26671 ^ n8067 ^ 1'b0 ;
  assign n26673 = n7666 & ~n26672 ;
  assign n26675 = n26674 ^ n26673 ^ n8724 ;
  assign n26676 = n1785 ^ x230 ^ 1'b0 ;
  assign n26678 = n2043 | n16288 ;
  assign n26679 = n26678 ^ n16552 ^ 1'b0 ;
  assign n26680 = n1438 & n26679 ;
  assign n26677 = n14157 | n23745 ;
  assign n26681 = n26680 ^ n26677 ^ 1'b0 ;
  assign n26682 = n26681 ^ n11802 ^ n6148 ;
  assign n26683 = ~n13685 & n20051 ;
  assign n26684 = n22535 ^ n21617 ^ 1'b0 ;
  assign n26685 = ( x115 & n5553 ) | ( x115 & ~n14470 ) | ( n5553 & ~n14470 ) ;
  assign n26686 = ~n1074 & n19963 ;
  assign n26687 = ~n4497 & n26686 ;
  assign n26688 = ~n5157 & n26687 ;
  assign n26689 = ( n7846 & ~n15042 ) | ( n7846 & n26688 ) | ( ~n15042 & n26688 ) ;
  assign n26690 = n26689 ^ n3225 ^ 1'b0 ;
  assign n26691 = ~n16095 & n26690 ;
  assign n26692 = n23971 ^ n15922 ^ 1'b0 ;
  assign n26693 = n11498 ^ n4259 ^ 1'b0 ;
  assign n26694 = n3697 & n26693 ;
  assign n26695 = n607 & n26694 ;
  assign n26696 = n26695 ^ n19030 ^ 1'b0 ;
  assign n26697 = n26692 & ~n26696 ;
  assign n26698 = ( n4256 & ~n13720 ) | ( n4256 & n26697 ) | ( ~n13720 & n26697 ) ;
  assign n26699 = ( n11122 & n14786 ) | ( n11122 & ~n26070 ) | ( n14786 & ~n26070 ) ;
  assign n26700 = n26699 ^ n17208 ^ n6249 ;
  assign n26701 = ~n2087 & n16314 ;
  assign n26702 = ( n19494 & n20329 ) | ( n19494 & ~n26701 ) | ( n20329 & ~n26701 ) ;
  assign n26704 = n8205 ^ n3492 ^ n2052 ;
  assign n26705 = n15390 ^ n4435 ^ 1'b0 ;
  assign n26706 = ~n26704 & n26705 ;
  assign n26707 = n26706 ^ n6797 ^ 1'b0 ;
  assign n26708 = n19009 & ~n26707 ;
  assign n26703 = n22918 ^ n6228 ^ n3833 ;
  assign n26709 = n26708 ^ n26703 ^ n23162 ;
  assign n26710 = n4772 & ~n22799 ;
  assign n26711 = n19721 & n26710 ;
  assign n26712 = n3727 & ~n26711 ;
  assign n26713 = n26712 ^ n25740 ^ 1'b0 ;
  assign n26714 = ( n11461 & n18417 ) | ( n11461 & n26614 ) | ( n18417 & n26614 ) ;
  assign n26715 = ( n1510 & ~n9013 ) | ( n1510 & n14857 ) | ( ~n9013 & n14857 ) ;
  assign n26716 = n26483 ^ n23077 ^ n6721 ;
  assign n26717 = n20051 | n26716 ;
  assign n26718 = n26715 | n26717 ;
  assign n26719 = n4977 ^ n2788 ^ 1'b0 ;
  assign n26720 = ( n12401 & n12859 ) | ( n12401 & n26719 ) | ( n12859 & n26719 ) ;
  assign n26721 = n21529 & ~n26720 ;
  assign n26722 = ( ~n9282 & n20617 ) | ( ~n9282 & n26721 ) | ( n20617 & n26721 ) ;
  assign n26723 = ~n7700 & n21187 ;
  assign n26724 = n3739 ^ n3583 ^ n1149 ;
  assign n26725 = n370 & ~n5263 ;
  assign n26726 = n9900 & ~n26725 ;
  assign n26727 = n26724 & n26726 ;
  assign n26728 = n23344 ^ n19816 ^ n11227 ;
  assign n26729 = ~n26727 & n26728 ;
  assign n26730 = n26723 & n26729 ;
  assign n26737 = n5337 | n10546 ;
  assign n26733 = ~n7341 & n22820 ;
  assign n26734 = n26733 ^ n6162 ^ 1'b0 ;
  assign n26731 = n2785 & n8827 ;
  assign n26732 = n26731 ^ n2233 ^ 1'b0 ;
  assign n26735 = n26734 ^ n26732 ^ 1'b0 ;
  assign n26736 = n1088 & n26735 ;
  assign n26738 = n26737 ^ n26736 ^ n7001 ;
  assign n26739 = n17541 | n22606 ;
  assign n26740 = n12302 & ~n26739 ;
  assign n26741 = n14487 & n17384 ;
  assign n26742 = ~n2764 & n26741 ;
  assign n26743 = ( ~x12 & n6043 ) | ( ~x12 & n17970 ) | ( n6043 & n17970 ) ;
  assign n26744 = ( ~n15809 & n17155 ) | ( ~n15809 & n26743 ) | ( n17155 & n26743 ) ;
  assign n26745 = n2399 | n3482 ;
  assign n26746 = ( n6784 & n16098 ) | ( n6784 & n19429 ) | ( n16098 & n19429 ) ;
  assign n26747 = n13850 ^ n2933 ^ 1'b0 ;
  assign n26748 = n26746 & n26747 ;
  assign n26749 = ~n17199 & n20807 ;
  assign n26750 = n26749 ^ n1433 ^ 1'b0 ;
  assign n26752 = n24139 ^ n16238 ^ n8186 ;
  assign n26753 = ( ~n358 & n7462 ) | ( ~n358 & n26752 ) | ( n7462 & n26752 ) ;
  assign n26754 = x62 & ~n26753 ;
  assign n26755 = n26754 ^ n10278 ^ 1'b0 ;
  assign n26751 = x190 & n20302 ;
  assign n26756 = n26755 ^ n26751 ^ 1'b0 ;
  assign n26757 = n17997 ^ n8800 ^ 1'b0 ;
  assign n26758 = n14979 & n26757 ;
  assign n26759 = n19619 & n26012 ;
  assign n26760 = n26759 ^ n1465 ^ 1'b0 ;
  assign n26761 = n26760 ^ n3903 ^ n360 ;
  assign n26767 = n7013 ^ n1689 ^ 1'b0 ;
  assign n26762 = ( n1623 & n15054 ) | ( n1623 & ~n16982 ) | ( n15054 & ~n16982 ) ;
  assign n26763 = ~n10487 & n25763 ;
  assign n26764 = ~n26762 & n26763 ;
  assign n26765 = n1153 & n26764 ;
  assign n26766 = n12993 & ~n26765 ;
  assign n26768 = n26767 ^ n26766 ^ n11077 ;
  assign n26769 = ~n12362 & n24598 ;
  assign n26770 = n26768 & n26769 ;
  assign n26771 = n7371 & ~n8334 ;
  assign n26772 = n12530 ^ n6131 ^ x253 ;
  assign n26773 = n26772 ^ n1874 ^ 1'b0 ;
  assign n26774 = n8119 & ~n15579 ;
  assign n26775 = n3022 & n26774 ;
  assign n26776 = n26775 ^ n23522 ^ 1'b0 ;
  assign n26777 = ~n23215 & n26776 ;
  assign n26778 = n11819 ^ n8793 ^ 1'b0 ;
  assign n26779 = n26778 ^ n15054 ^ n6347 ;
  assign n26780 = n10575 ^ n5299 ^ 1'b0 ;
  assign n26781 = n3228 ^ n2798 ^ 1'b0 ;
  assign n26782 = n26781 ^ n3469 ^ 1'b0 ;
  assign n26783 = n1518 & n26782 ;
  assign n26784 = n10767 & ~n11339 ;
  assign n26785 = ~n3643 & n26784 ;
  assign n26786 = ( n967 & ~n12362 ) | ( n967 & n14018 ) | ( ~n12362 & n14018 ) ;
  assign n26787 = n11032 & n16623 ;
  assign n26788 = n26786 & n26787 ;
  assign n26789 = n6063 ^ n867 ^ 1'b0 ;
  assign n26790 = ~n10440 & n26789 ;
  assign n26791 = n26790 ^ n22060 ^ 1'b0 ;
  assign n26797 = ( n552 & ~n9134 ) | ( n552 & n15539 ) | ( ~n9134 & n15539 ) ;
  assign n26795 = n20160 ^ n11710 ^ n5454 ;
  assign n26792 = n3880 | n16917 ;
  assign n26793 = n26792 ^ n26041 ^ n10419 ;
  assign n26794 = n8716 | n26793 ;
  assign n26796 = n26795 ^ n26794 ^ 1'b0 ;
  assign n26798 = n26797 ^ n26796 ^ n1753 ;
  assign n26799 = ( n4224 & n10866 ) | ( n4224 & ~n17626 ) | ( n10866 & ~n17626 ) ;
  assign n26800 = n21633 ^ n17184 ^ 1'b0 ;
  assign n26801 = n26799 & ~n26800 ;
  assign n26802 = n9931 | n19363 ;
  assign n26803 = n26802 ^ n21716 ^ 1'b0 ;
  assign n26804 = n11146 | n26803 ;
  assign n26805 = ( ~x50 & n9429 ) | ( ~x50 & n10986 ) | ( n9429 & n10986 ) ;
  assign n26806 = n26805 ^ n2630 ^ 1'b0 ;
  assign n26807 = n16064 ^ n11340 ^ 1'b0 ;
  assign n26808 = n24345 | n26807 ;
  assign n26809 = n6474 ^ n3389 ^ 1'b0 ;
  assign n26810 = n23343 & ~n26809 ;
  assign n26811 = n26810 ^ n20889 ^ n5945 ;
  assign n26812 = ~n2225 & n11546 ;
  assign n26813 = n26812 ^ n11868 ^ 1'b0 ;
  assign n26814 = n20561 ^ n8273 ^ n4154 ;
  assign n26815 = n26813 | n26814 ;
  assign n26816 = n1932 & ~n26815 ;
  assign n26817 = n14507 | n26816 ;
  assign n26818 = ( n12323 & ~n19164 ) | ( n12323 & n26817 ) | ( ~n19164 & n26817 ) ;
  assign n26819 = n26811 | n26818 ;
  assign n26820 = ( n3775 & ~n10899 ) | ( n3775 & n20893 ) | ( ~n10899 & n20893 ) ;
  assign n26821 = ~n15468 & n20193 ;
  assign n26822 = ~n26820 & n26821 ;
  assign n26830 = ~n1977 & n9174 ;
  assign n26829 = n5671 | n20160 ;
  assign n26831 = n26830 ^ n26829 ^ 1'b0 ;
  assign n26832 = ( n867 & n6326 ) | ( n867 & ~n19184 ) | ( n6326 & ~n19184 ) ;
  assign n26833 = ( n11907 & n14180 ) | ( n11907 & n26832 ) | ( n14180 & n26832 ) ;
  assign n26834 = ( n19584 & ~n21582 ) | ( n19584 & n26833 ) | ( ~n21582 & n26833 ) ;
  assign n26835 = ~n26831 & n26834 ;
  assign n26823 = n8780 ^ n1074 ^ 1'b0 ;
  assign n26824 = n26823 ^ n16685 ^ n859 ;
  assign n26825 = ~n14866 & n26824 ;
  assign n26826 = n26825 ^ n595 ^ 1'b0 ;
  assign n26827 = ( n8281 & ~n18885 ) | ( n8281 & n26826 ) | ( ~n18885 & n26826 ) ;
  assign n26828 = n10154 & ~n26827 ;
  assign n26836 = n26835 ^ n26828 ^ 1'b0 ;
  assign n26837 = ~n5043 & n23535 ;
  assign n26838 = ~n1311 & n26837 ;
  assign n26839 = n9030 & n11360 ;
  assign n26840 = n22851 ^ n9927 ^ 1'b0 ;
  assign n26841 = n26839 & n26840 ;
  assign n26842 = n19867 ^ n11879 ^ n3337 ;
  assign n26843 = n14686 ^ n7257 ^ n6767 ;
  assign n26844 = n26843 ^ n3328 ^ 1'b0 ;
  assign n26845 = n4410 | n26844 ;
  assign n26856 = ~n11589 & n21459 ;
  assign n26857 = ~n22818 & n26856 ;
  assign n26846 = n3512 & n6630 ;
  assign n26852 = n445 & ~n11574 ;
  assign n26851 = ~n1978 & n6428 ;
  assign n26853 = n26852 ^ n26851 ^ 1'b0 ;
  assign n26847 = ~n9629 & n10978 ;
  assign n26848 = n26847 ^ n8681 ^ 1'b0 ;
  assign n26849 = n26848 ^ n12597 ^ 1'b0 ;
  assign n26850 = n2832 | n26849 ;
  assign n26854 = n26853 ^ n26850 ^ n8171 ;
  assign n26855 = n26846 & ~n26854 ;
  assign n26858 = n26857 ^ n26855 ^ n13309 ;
  assign n26861 = ( n8227 & ~n18924 ) | ( n8227 & n24024 ) | ( ~n18924 & n24024 ) ;
  assign n26859 = n13308 ^ n4383 ^ 1'b0 ;
  assign n26860 = ( n8465 & n11247 ) | ( n8465 & ~n26859 ) | ( n11247 & ~n26859 ) ;
  assign n26862 = n26861 ^ n26860 ^ 1'b0 ;
  assign n26863 = ( n5384 & ~n8517 ) | ( n5384 & n25856 ) | ( ~n8517 & n25856 ) ;
  assign n26866 = n12728 ^ n1088 ^ 1'b0 ;
  assign n26867 = ( n2616 & n17786 ) | ( n2616 & n26866 ) | ( n17786 & n26866 ) ;
  assign n26865 = n19296 ^ n5541 ^ n4818 ;
  assign n26868 = n26867 ^ n26865 ^ n3860 ;
  assign n26864 = n2477 | n4287 ;
  assign n26869 = n26868 ^ n26864 ^ 1'b0 ;
  assign n26870 = n20351 ^ n7243 ^ 1'b0 ;
  assign n26871 = ~n7841 & n9917 ;
  assign n26872 = ( ~n10811 & n18304 ) | ( ~n10811 & n26871 ) | ( n18304 & n26871 ) ;
  assign n26873 = n20487 ^ n9056 ^ 1'b0 ;
  assign n26874 = n3500 & n26873 ;
  assign n26875 = n3375 & ~n25225 ;
  assign n26876 = ~n6938 & n26875 ;
  assign n26877 = ~n12309 & n26876 ;
  assign n26878 = n26877 ^ n12739 ^ 1'b0 ;
  assign n26879 = ~n5894 & n7391 ;
  assign n26880 = n8743 ^ x194 ^ 1'b0 ;
  assign n26881 = ( n17401 & ~n22204 ) | ( n17401 & n26880 ) | ( ~n22204 & n26880 ) ;
  assign n26882 = ( n851 & n5460 ) | ( n851 & ~n26336 ) | ( n5460 & ~n26336 ) ;
  assign n26883 = n21162 ^ n14564 ^ 1'b0 ;
  assign n26884 = n7352 ^ n764 ^ 1'b0 ;
  assign n26885 = n26883 | n26884 ;
  assign n26886 = ( ~n6866 & n9302 ) | ( ~n6866 & n11590 ) | ( n9302 & n11590 ) ;
  assign n26887 = n26886 ^ n480 ^ 1'b0 ;
  assign n26888 = n26885 | n26887 ;
  assign n26889 = x71 & ~n271 ;
  assign n26890 = ~n9804 & n26889 ;
  assign n26891 = n22269 | n26890 ;
  assign n26892 = n26888 & ~n26891 ;
  assign n26893 = n14342 ^ n3633 ^ n1155 ;
  assign n26894 = n3226 | n5557 ;
  assign n26895 = n8334 | n26894 ;
  assign n26896 = n7350 & n26895 ;
  assign n26897 = n16346 | n26896 ;
  assign n26898 = n26897 ^ n1605 ^ 1'b0 ;
  assign n26899 = ~n26893 & n26898 ;
  assign n26900 = ~n13229 & n16903 ;
  assign n26901 = n26900 ^ n24750 ^ 1'b0 ;
  assign n26902 = ( n1427 & n17578 ) | ( n1427 & ~n18661 ) | ( n17578 & ~n18661 ) ;
  assign n26907 = n14034 ^ n4552 ^ n4332 ;
  assign n26908 = ( n400 & n18751 ) | ( n400 & ~n26907 ) | ( n18751 & ~n26907 ) ;
  assign n26903 = n16789 ^ n6832 ^ 1'b0 ;
  assign n26904 = n6476 | n26903 ;
  assign n26905 = n17491 ^ n2277 ^ 1'b0 ;
  assign n26906 = ~n26904 & n26905 ;
  assign n26909 = n26908 ^ n26906 ^ 1'b0 ;
  assign n26910 = ( n2716 & n8066 ) | ( n2716 & n26909 ) | ( n8066 & n26909 ) ;
  assign n26912 = ~n269 & n16844 ;
  assign n26913 = ~n5441 & n26912 ;
  assign n26911 = ( n2106 & ~n3833 ) | ( n2106 & n20143 ) | ( ~n3833 & n20143 ) ;
  assign n26914 = n26913 ^ n26911 ^ 1'b0 ;
  assign n26915 = n1175 & n17854 ;
  assign n26916 = ~n6173 & n26915 ;
  assign n26917 = n4783 | n5276 ;
  assign n26918 = n6833 | n15340 ;
  assign n26919 = n26918 ^ n5660 ^ 1'b0 ;
  assign n26920 = n26919 ^ n21619 ^ n11285 ;
  assign n26921 = ( n26916 & ~n26917 ) | ( n26916 & n26920 ) | ( ~n26917 & n26920 ) ;
  assign n26922 = n16392 ^ n10728 ^ n4762 ;
  assign n26923 = n2066 & ~n9987 ;
  assign n26924 = ~n3837 & n26923 ;
  assign n26925 = n10851 | n26924 ;
  assign n26927 = n1706 & n17565 ;
  assign n26928 = n26927 ^ n14396 ^ n2663 ;
  assign n26926 = n1850 | n24690 ;
  assign n26929 = n26928 ^ n26926 ^ 1'b0 ;
  assign n26930 = n11692 & ~n26929 ;
  assign n26931 = n20057 ^ n8601 ^ n6764 ;
  assign n26932 = n20326 ^ n1390 ^ 1'b0 ;
  assign n26933 = n26931 & n26932 ;
  assign n26934 = n9362 & ~n14603 ;
  assign n26935 = ( n9217 & n26552 ) | ( n9217 & n26934 ) | ( n26552 & n26934 ) ;
  assign n26936 = ( n13903 & n16520 ) | ( n13903 & ~n24345 ) | ( n16520 & ~n24345 ) ;
  assign n26937 = n1954 ^ n1910 ^ 1'b0 ;
  assign n26938 = n26937 ^ n6271 ^ 1'b0 ;
  assign n26939 = ( n735 & n10502 ) | ( n735 & ~n11039 ) | ( n10502 & ~n11039 ) ;
  assign n26940 = n14320 ^ n8316 ^ n6005 ;
  assign n26941 = n26940 ^ n8810 ^ n580 ;
  assign n26942 = ( ~n5915 & n26939 ) | ( ~n5915 & n26941 ) | ( n26939 & n26941 ) ;
  assign n26944 = ( ~n1780 & n4242 ) | ( ~n1780 & n11594 ) | ( n4242 & n11594 ) ;
  assign n26943 = n9142 | n18205 ;
  assign n26945 = n26944 ^ n26943 ^ n14731 ;
  assign n26946 = n17683 ^ n14336 ^ x178 ;
  assign n26947 = n26946 ^ n3325 ^ 1'b0 ;
  assign n26948 = n1240 | n11951 ;
  assign n26949 = n22161 & ~n26948 ;
  assign n26950 = n4211 | n8269 ;
  assign n26951 = n26950 ^ n3792 ^ 1'b0 ;
  assign n26952 = n12989 & n26951 ;
  assign n26953 = n13669 | n26952 ;
  assign n26956 = n5538 ^ n3735 ^ 1'b0 ;
  assign n26954 = n7339 | n9481 ;
  assign n26955 = n26954 ^ n16268 ^ 1'b0 ;
  assign n26957 = n26956 ^ n26955 ^ n4739 ;
  assign n26958 = ( n5356 & n6941 ) | ( n5356 & n22321 ) | ( n6941 & n22321 ) ;
  assign n26959 = ( ~n8551 & n13293 ) | ( ~n8551 & n26958 ) | ( n13293 & n26958 ) ;
  assign n26960 = ( n3061 & n15207 ) | ( n3061 & n26959 ) | ( n15207 & n26959 ) ;
  assign n26961 = n18725 & n26960 ;
  assign n26962 = n21232 & n26961 ;
  assign n26963 = n5596 & n8272 ;
  assign n26964 = n11220 ^ n6347 ^ 1'b0 ;
  assign n26965 = n26964 ^ n18829 ^ n1189 ;
  assign n26966 = ( ~n6150 & n8972 ) | ( ~n6150 & n23605 ) | ( n8972 & n23605 ) ;
  assign n26967 = n17275 ^ n284 ^ 1'b0 ;
  assign n26968 = n8418 ^ x157 ^ 1'b0 ;
  assign n26969 = n26968 ^ n26826 ^ 1'b0 ;
  assign n26970 = ~n1312 & n1753 ;
  assign n26972 = n2220 & n11027 ;
  assign n26973 = n12946 & ~n26972 ;
  assign n26974 = ~n14915 & n26973 ;
  assign n26971 = n2802 | n18084 ;
  assign n26975 = n26974 ^ n26971 ^ 1'b0 ;
  assign n26976 = n26975 ^ n15068 ^ n3832 ;
  assign n26977 = n26976 ^ n18743 ^ n2201 ;
  assign n26978 = n600 & n1372 ;
  assign n26979 = ~n24793 & n26978 ;
  assign n26980 = n9789 ^ n8892 ^ n5251 ;
  assign n26981 = n8204 & n26980 ;
  assign n26982 = ~n26044 & n26981 ;
  assign n26984 = n13012 ^ n9351 ^ n6733 ;
  assign n26983 = n21235 ^ n16959 ^ n469 ;
  assign n26985 = n26984 ^ n26983 ^ n21046 ;
  assign n26986 = ( ~n4744 & n11001 ) | ( ~n4744 & n26985 ) | ( n11001 & n26985 ) ;
  assign n26987 = n3585 | n4979 ;
  assign n26988 = n26986 & ~n26987 ;
  assign n26989 = n2492 | n21995 ;
  assign n26990 = ~n10760 & n23970 ;
  assign n26991 = ( n8333 & n24551 ) | ( n8333 & ~n26990 ) | ( n24551 & ~n26990 ) ;
  assign n26992 = ( n320 & n5577 ) | ( n320 & ~n19352 ) | ( n5577 & ~n19352 ) ;
  assign n26993 = ~n4975 & n26992 ;
  assign n26994 = ( n8851 & n13319 ) | ( n8851 & n26993 ) | ( n13319 & n26993 ) ;
  assign n26995 = n9875 ^ n8739 ^ n3914 ;
  assign n26996 = n7551 | n15941 ;
  assign n26997 = ( n20855 & n26995 ) | ( n20855 & ~n26996 ) | ( n26995 & ~n26996 ) ;
  assign n26998 = n17618 ^ n6204 ^ n2314 ;
  assign n27000 = n19434 ^ n13947 ^ n5720 ;
  assign n26999 = ~x116 & n8317 ;
  assign n27001 = n27000 ^ n26999 ^ n3096 ;
  assign n27002 = n26998 & ~n27001 ;
  assign n27003 = n9660 & n13892 ;
  assign n27004 = ( ~n12488 & n16231 ) | ( ~n12488 & n27003 ) | ( n16231 & n27003 ) ;
  assign n27005 = n3625 | n20085 ;
  assign n27006 = n27005 ^ n23843 ^ 1'b0 ;
  assign n27007 = n1558 & n8148 ;
  assign n27008 = n26464 ^ n18781 ^ n426 ;
  assign n27009 = ( n11524 & n16471 ) | ( n11524 & ~n27008 ) | ( n16471 & ~n27008 ) ;
  assign n27010 = ( n332 & n27007 ) | ( n332 & n27009 ) | ( n27007 & n27009 ) ;
  assign n27011 = ~n12196 & n15174 ;
  assign n27012 = n13129 & n27011 ;
  assign n27013 = n26567 | n27012 ;
  assign n27014 = n27013 ^ n19651 ^ 1'b0 ;
  assign n27015 = ( n5932 & n6626 ) | ( n5932 & n17419 ) | ( n6626 & n17419 ) ;
  assign n27016 = n6227 & ~n27015 ;
  assign n27017 = n27016 ^ n6555 ^ 1'b0 ;
  assign n27018 = n3706 | n27017 ;
  assign n27019 = n1611 | n25780 ;
  assign n27020 = ~n6265 & n14829 ;
  assign n27021 = n27019 & n27020 ;
  assign n27022 = n10078 ^ n4437 ^ 1'b0 ;
  assign n27023 = n15409 | n27022 ;
  assign n27024 = ~n19558 & n27023 ;
  assign n27025 = n27021 & ~n27024 ;
  assign n27027 = n12570 ^ n2104 ^ 1'b0 ;
  assign n27028 = ( n2871 & ~n7898 ) | ( n2871 & n27027 ) | ( ~n7898 & n27027 ) ;
  assign n27026 = n1708 & ~n8456 ;
  assign n27029 = n27028 ^ n27026 ^ 1'b0 ;
  assign n27030 = n7890 | n17935 ;
  assign n27031 = n27030 ^ n14821 ^ 1'b0 ;
  assign n27032 = n14517 ^ n4662 ^ 1'b0 ;
  assign n27033 = n23519 ^ n4745 ^ 1'b0 ;
  assign n27034 = n2155 & ~n27033 ;
  assign n27035 = n19584 & ~n25320 ;
  assign n27036 = ~n4093 & n27035 ;
  assign n27037 = n15084 ^ n1256 ^ 1'b0 ;
  assign n27038 = ( n3605 & n21251 ) | ( n3605 & ~n27037 ) | ( n21251 & ~n27037 ) ;
  assign n27039 = n17243 & n27038 ;
  assign n27040 = ~n6317 & n26583 ;
  assign n27041 = n4190 & n27040 ;
  assign n27042 = n8768 ^ n3114 ^ 1'b0 ;
  assign n27043 = ( ~n6113 & n10511 ) | ( ~n6113 & n13518 ) | ( n10511 & n13518 ) ;
  assign n27044 = n23882 & n27043 ;
  assign n27045 = ~n4100 & n27044 ;
  assign n27046 = n27042 | n27045 ;
  assign n27047 = n27046 ^ n15317 ^ 1'b0 ;
  assign n27048 = ( n1121 & n4359 ) | ( n1121 & ~n12995 ) | ( n4359 & ~n12995 ) ;
  assign n27049 = ~n11000 & n21878 ;
  assign n27050 = n1919 & n27049 ;
  assign n27051 = n27050 ^ n22117 ^ n9122 ;
  assign n27052 = n27051 ^ n23401 ^ n10870 ;
  assign n27053 = n27052 ^ n16110 ^ 1'b0 ;
  assign n27054 = n16826 ^ n14559 ^ 1'b0 ;
  assign n27055 = n27054 ^ n2777 ^ 1'b0 ;
  assign n27056 = ~n7939 & n10998 ;
  assign n27057 = ~n13761 & n27056 ;
  assign n27058 = n27057 ^ n18531 ^ n4356 ;
  assign n27059 = n27058 ^ n3970 ^ 1'b0 ;
  assign n27060 = n27059 ^ n21476 ^ n17073 ;
  assign n27061 = ( n9270 & ~n26567 ) | ( n9270 & n27060 ) | ( ~n26567 & n27060 ) ;
  assign n27077 = ( n3555 & n6056 ) | ( n3555 & n11079 ) | ( n6056 & n11079 ) ;
  assign n27074 = n25552 ^ n22660 ^ n18850 ;
  assign n27075 = n27074 ^ x231 ^ 1'b0 ;
  assign n27076 = ~n4265 & n27075 ;
  assign n27071 = ~n7369 & n19216 ;
  assign n27062 = n11645 ^ n5828 ^ n1532 ;
  assign n27063 = ~n8271 & n27062 ;
  assign n27064 = n2380 & n4255 ;
  assign n27065 = ~n27063 & n27064 ;
  assign n27066 = n17507 ^ n5687 ^ n3614 ;
  assign n27067 = n1440 | n27066 ;
  assign n27068 = n27067 ^ n23754 ^ 1'b0 ;
  assign n27069 = n19905 & n27068 ;
  assign n27070 = n27065 & n27069 ;
  assign n27072 = n27071 ^ n27070 ^ n10786 ;
  assign n27073 = n14272 | n27072 ;
  assign n27078 = n27077 ^ n27076 ^ n27073 ;
  assign n27079 = n5284 ^ n341 ^ 1'b0 ;
  assign n27080 = n10273 & n27079 ;
  assign n27081 = n5746 & n24290 ;
  assign n27082 = n27081 ^ n1108 ^ 1'b0 ;
  assign n27083 = ( n4108 & n12447 ) | ( n4108 & ~n22538 ) | ( n12447 & ~n22538 ) ;
  assign n27084 = n27083 ^ n15550 ^ 1'b0 ;
  assign n27085 = n27082 & n27084 ;
  assign n27086 = n24905 ^ n21506 ^ n3097 ;
  assign n27087 = n6670 & n15694 ;
  assign n27088 = n27086 & ~n27087 ;
  assign n27089 = n27088 ^ n5604 ^ 1'b0 ;
  assign n27090 = n5385 & ~n10468 ;
  assign n27091 = ~n6070 & n27090 ;
  assign n27092 = n22208 ^ n10973 ^ 1'b0 ;
  assign n27093 = ( n441 & n18337 ) | ( n441 & ~n19371 ) | ( n18337 & ~n19371 ) ;
  assign n27094 = n27093 ^ n1838 ^ 1'b0 ;
  assign n27095 = n7009 & n27094 ;
  assign n27096 = ~n27092 & n27095 ;
  assign n27097 = n7196 | n10726 ;
  assign n27098 = n27097 ^ n16049 ^ 1'b0 ;
  assign n27099 = ~n24816 & n27098 ;
  assign n27103 = n257 & ~n17690 ;
  assign n27102 = ~n9389 & n9921 ;
  assign n27104 = n27103 ^ n27102 ^ 1'b0 ;
  assign n27100 = n11644 ^ n4097 ^ 1'b0 ;
  assign n27101 = n27100 ^ n9058 ^ n1168 ;
  assign n27105 = n27104 ^ n27101 ^ n20415 ;
  assign n27106 = n19815 ^ n8798 ^ 1'b0 ;
  assign n27107 = ~n13430 & n27106 ;
  assign n27108 = n24589 ^ n7914 ^ 1'b0 ;
  assign n27109 = n27108 ^ n4306 ^ 1'b0 ;
  assign n27110 = ~n13342 & n27109 ;
  assign n27111 = n27110 ^ n13712 ^ 1'b0 ;
  assign n27112 = ~n14206 & n27111 ;
  assign n27113 = n27107 & n27112 ;
  assign n27114 = n27113 ^ n10482 ^ 1'b0 ;
  assign n27115 = ~n16473 & n27114 ;
  assign n27116 = n18320 ^ n12406 ^ n8049 ;
  assign n27117 = ( n5677 & n12078 ) | ( n5677 & n27116 ) | ( n12078 & n27116 ) ;
  assign n27118 = n13789 ^ n295 ^ x79 ;
  assign n27119 = n27118 ^ n20377 ^ n17960 ;
  assign n27120 = ~n20606 & n27119 ;
  assign n27121 = ~n14465 & n25949 ;
  assign n27122 = ~n6347 & n27121 ;
  assign n27123 = n9014 | n27122 ;
  assign n27124 = n27123 ^ n19462 ^ 1'b0 ;
  assign n27125 = ( n2017 & ~n12232 ) | ( n2017 & n17427 ) | ( ~n12232 & n17427 ) ;
  assign n27126 = n15345 & n21378 ;
  assign n27127 = ~n27125 & n27126 ;
  assign n27128 = ( n9708 & n13667 ) | ( n9708 & ~n18395 ) | ( n13667 & ~n18395 ) ;
  assign n27129 = n15832 & ~n18838 ;
  assign n27130 = n27129 ^ n13457 ^ 1'b0 ;
  assign n27131 = n27128 & ~n27130 ;
  assign n27132 = n14226 & n27131 ;
  assign n27133 = ( n420 & ~n5032 ) | ( n420 & n8137 ) | ( ~n5032 & n8137 ) ;
  assign n27134 = n27133 ^ n16049 ^ 1'b0 ;
  assign n27135 = n2663 & ~n27134 ;
  assign n27136 = n9151 & n21416 ;
  assign n27137 = ( ~n475 & n806 ) | ( ~n475 & n3732 ) | ( n806 & n3732 ) ;
  assign n27138 = n27137 ^ n18913 ^ 1'b0 ;
  assign n27139 = n12296 | n27138 ;
  assign n27140 = n443 | n6420 ;
  assign n27141 = ( n12809 & ~n19990 ) | ( n12809 & n23476 ) | ( ~n19990 & n23476 ) ;
  assign n27142 = n10887 | n27141 ;
  assign n27143 = n27140 & ~n27142 ;
  assign n27144 = ( n1539 & n3883 ) | ( n1539 & ~n17392 ) | ( n3883 & ~n17392 ) ;
  assign n27145 = n9564 ^ n3246 ^ 1'b0 ;
  assign n27146 = n520 & ~n27145 ;
  assign n27147 = ( n15088 & n20961 ) | ( n15088 & n27146 ) | ( n20961 & n27146 ) ;
  assign n27148 = n8666 ^ n632 ^ 1'b0 ;
  assign n27149 = n6387 ^ n3326 ^ 1'b0 ;
  assign n27150 = n27148 & ~n27149 ;
  assign n27151 = n25633 ^ n2683 ^ 1'b0 ;
  assign n27152 = n1874 & n18798 ;
  assign n27153 = ~n27151 & n27152 ;
  assign n27154 = n27153 ^ n18083 ^ n7650 ;
  assign n27155 = n19154 ^ n7493 ^ 1'b0 ;
  assign n27156 = n10734 ^ n7703 ^ 1'b0 ;
  assign n27157 = n10448 ^ n2958 ^ 1'b0 ;
  assign n27158 = n27157 ^ n26472 ^ n23365 ;
  assign n27160 = n17129 ^ n11747 ^ n1975 ;
  assign n27161 = n27160 ^ n6753 ^ 1'b0 ;
  assign n27162 = n2692 | n27161 ;
  assign n27159 = ( n1926 & n7937 ) | ( n1926 & ~n9365 ) | ( n7937 & ~n9365 ) ;
  assign n27163 = n27162 ^ n27159 ^ 1'b0 ;
  assign n27164 = n6869 | n27163 ;
  assign n27165 = n25322 ^ n13295 ^ 1'b0 ;
  assign n27166 = n10228 ^ n7250 ^ 1'b0 ;
  assign n27167 = ~n10243 & n27166 ;
  assign n27168 = ~n8749 & n9499 ;
  assign n27169 = ( ~n13340 & n13579 ) | ( ~n13340 & n27168 ) | ( n13579 & n27168 ) ;
  assign n27170 = ( n3636 & n12462 ) | ( n3636 & n14065 ) | ( n12462 & n14065 ) ;
  assign n27171 = n1029 & ~n9454 ;
  assign n27172 = ~n5620 & n8974 ;
  assign n27173 = n27172 ^ n11990 ^ 1'b0 ;
  assign n27174 = n9665 & ~n10324 ;
  assign n27175 = ~n18339 & n27174 ;
  assign n27176 = n27175 ^ n16462 ^ n12504 ;
  assign n27177 = n2549 | n27176 ;
  assign n27178 = ( n2980 & n13694 ) | ( n2980 & n20616 ) | ( n13694 & n20616 ) ;
  assign n27179 = n2149 ^ n790 ^ 1'b0 ;
  assign n27180 = n5063 & n27179 ;
  assign n27181 = n21083 ^ n16283 ^ n8913 ;
  assign n27182 = ( n10301 & ~n27180 ) | ( n10301 & n27181 ) | ( ~n27180 & n27181 ) ;
  assign n27184 = n7192 ^ n4009 ^ 1'b0 ;
  assign n27185 = n17366 | n27184 ;
  assign n27186 = n10123 & n27185 ;
  assign n27187 = n27186 ^ n19853 ^ 1'b0 ;
  assign n27183 = n4507 ^ n3485 ^ 1'b0 ;
  assign n27188 = n27187 ^ n27183 ^ n7196 ;
  assign n27189 = n9852 | n10841 ;
  assign n27190 = n18990 & ~n27189 ;
  assign n27192 = n25078 ^ n16132 ^ 1'b0 ;
  assign n27193 = n8396 | n27192 ;
  assign n27194 = n27193 ^ n17707 ^ n6777 ;
  assign n27191 = ( ~n1966 & n2364 ) | ( ~n1966 & n7614 ) | ( n2364 & n7614 ) ;
  assign n27195 = n27194 ^ n27191 ^ 1'b0 ;
  assign n27196 = ( x40 & n8307 ) | ( x40 & n24805 ) | ( n8307 & n24805 ) ;
  assign n27197 = n6558 ^ n3006 ^ 1'b0 ;
  assign n27198 = n15357 & ~n27197 ;
  assign n27199 = ~n15335 & n20339 ;
  assign n27200 = x151 & n1705 ;
  assign n27201 = ~n2750 & n27200 ;
  assign n27202 = ( ~x76 & n27199 ) | ( ~x76 & n27201 ) | ( n27199 & n27201 ) ;
  assign n27203 = n11071 | n17060 ;
  assign n27204 = n27202 & ~n27203 ;
  assign n27205 = n8857 ^ n7976 ^ 1'b0 ;
  assign n27206 = n10485 ^ n7922 ^ 1'b0 ;
  assign n27207 = n27206 ^ n17920 ^ n7934 ;
  assign n27208 = n27207 ^ n24138 ^ n17775 ;
  assign n27209 = ~n1745 & n21194 ;
  assign n27210 = ( n1916 & n12547 ) | ( n1916 & ~n21131 ) | ( n12547 & ~n21131 ) ;
  assign n27211 = n25589 ^ n7586 ^ 1'b0 ;
  assign n27212 = n9829 & n27211 ;
  assign n27213 = n7405 & n27212 ;
  assign n27214 = n27213 ^ n12588 ^ 1'b0 ;
  assign n27215 = n27214 ^ n15161 ^ 1'b0 ;
  assign n27216 = n27210 & ~n27215 ;
  assign n27217 = n8859 ^ n7331 ^ 1'b0 ;
  assign n27218 = n13776 | n24966 ;
  assign n27219 = ( ~n3744 & n12931 ) | ( ~n3744 & n15456 ) | ( n12931 & n15456 ) ;
  assign n27220 = ~n6568 & n27219 ;
  assign n27221 = n333 & ~n21865 ;
  assign n27222 = ~n26909 & n27221 ;
  assign n27223 = n18054 ^ n9049 ^ 1'b0 ;
  assign n27224 = n25094 & ~n27223 ;
  assign n27225 = n2061 | n5508 ;
  assign n27226 = n7046 | n27225 ;
  assign n27227 = n7148 & n27226 ;
  assign n27231 = n5271 ^ n4250 ^ n4060 ;
  assign n27232 = ( n4518 & ~n14314 ) | ( n4518 & n27231 ) | ( ~n14314 & n27231 ) ;
  assign n27228 = n18887 ^ n11578 ^ 1'b0 ;
  assign n27229 = ~n5839 & n27228 ;
  assign n27230 = n13135 & n27229 ;
  assign n27233 = n27232 ^ n27230 ^ 1'b0 ;
  assign n27234 = ( n3699 & n5946 ) | ( n3699 & ~n14724 ) | ( n5946 & ~n14724 ) ;
  assign n27235 = n13505 & ~n25787 ;
  assign n27236 = n27235 ^ n15397 ^ 1'b0 ;
  assign n27237 = n27236 ^ n16155 ^ n9918 ;
  assign n27238 = n27237 ^ n3106 ^ n579 ;
  assign n27239 = n27234 & ~n27238 ;
  assign n27240 = n9327 & ~n10353 ;
  assign n27241 = n7867 & ~n8729 ;
  assign n27242 = n27240 & n27241 ;
  assign n27243 = ( x140 & n1552 ) | ( x140 & ~n27242 ) | ( n1552 & ~n27242 ) ;
  assign n27244 = n27243 ^ n6923 ^ 1'b0 ;
  assign n27245 = n4601 & ~n27244 ;
  assign n27246 = n5128 & n25944 ;
  assign n27247 = n27246 ^ n6703 ^ 1'b0 ;
  assign n27248 = n9188 ^ n7803 ^ n3490 ;
  assign n27249 = ( n4769 & n7166 ) | ( n4769 & ~n27248 ) | ( n7166 & ~n27248 ) ;
  assign n27250 = n27249 ^ n12240 ^ n452 ;
  assign n27251 = n27247 & n27250 ;
  assign n27252 = ~n27245 & n27251 ;
  assign n27253 = n26293 | n27252 ;
  assign n27256 = n809 | n8421 ;
  assign n27254 = n12273 | n17218 ;
  assign n27255 = n27254 ^ n22012 ^ 1'b0 ;
  assign n27257 = n27256 ^ n27255 ^ n5407 ;
  assign n27267 = n2279 | n6765 ;
  assign n27268 = n2279 & ~n27267 ;
  assign n27269 = n27268 ^ n5064 ^ n4259 ;
  assign n27258 = n6954 | n13572 ;
  assign n27259 = n27258 ^ n9189 ^ 1'b0 ;
  assign n27262 = n1749 & ~n9685 ;
  assign n27263 = n27262 ^ n3248 ^ 1'b0 ;
  assign n27261 = ~n2850 & n5702 ;
  assign n27264 = n27263 ^ n27261 ^ 1'b0 ;
  assign n27260 = ( n939 & n5025 ) | ( n939 & ~n15337 ) | ( n5025 & ~n15337 ) ;
  assign n27265 = n27264 ^ n27260 ^ 1'b0 ;
  assign n27266 = ~n27259 & n27265 ;
  assign n27270 = n27269 ^ n27266 ^ n17154 ;
  assign n27271 = n20870 | n25894 ;
  assign n27272 = n2841 & ~n27271 ;
  assign n27273 = n2227 & ~n23442 ;
  assign n27274 = n27273 ^ n13147 ^ 1'b0 ;
  assign n27275 = ( n1740 & ~n9451 ) | ( n1740 & n12847 ) | ( ~n9451 & n12847 ) ;
  assign n27276 = n21123 & n27275 ;
  assign n27277 = ( n4445 & n25431 ) | ( n4445 & ~n27276 ) | ( n25431 & ~n27276 ) ;
  assign n27278 = ~n4850 & n5386 ;
  assign n27279 = ~n7270 & n27278 ;
  assign n27280 = ( ~n7248 & n17607 ) | ( ~n7248 & n27279 ) | ( n17607 & n27279 ) ;
  assign n27281 = n11058 ^ n4987 ^ n4617 ;
  assign n27282 = ( n3318 & ~n19485 ) | ( n3318 & n27281 ) | ( ~n19485 & n27281 ) ;
  assign n27283 = n27282 ^ n2333 ^ 1'b0 ;
  assign n27284 = n4867 ^ n2677 ^ 1'b0 ;
  assign n27285 = n10779 & n22700 ;
  assign n27286 = ( n4085 & n7955 ) | ( n4085 & ~n10150 ) | ( n7955 & ~n10150 ) ;
  assign n27288 = n8282 ^ x4 ^ 1'b0 ;
  assign n27289 = n2409 & ~n12579 ;
  assign n27290 = ~x65 & n11659 ;
  assign n27291 = n27289 & n27290 ;
  assign n27292 = ~n27288 & n27291 ;
  assign n27287 = n3070 & n18302 ;
  assign n27293 = n27292 ^ n27287 ^ 1'b0 ;
  assign n27294 = n22538 ^ n18212 ^ 1'b0 ;
  assign n27295 = n27293 & n27294 ;
  assign n27296 = n22089 ^ n893 ^ 1'b0 ;
  assign n27297 = n1924 & n27296 ;
  assign n27298 = n17452 | n18836 ;
  assign n27299 = n12752 | n27298 ;
  assign n27300 = n8740 & n27299 ;
  assign n27301 = n3395 | n23901 ;
  assign n27302 = n27301 ^ n20005 ^ n15616 ;
  assign n27303 = ( n1264 & n3297 ) | ( n1264 & ~n7168 ) | ( n3297 & ~n7168 ) ;
  assign n27304 = ~n2349 & n13145 ;
  assign n27305 = ~n16356 & n27304 ;
  assign n27306 = n21845 ^ n13383 ^ 1'b0 ;
  assign n27307 = n5080 & ~n27306 ;
  assign n27308 = ~n24996 & n27307 ;
  assign n27309 = n5671 | n11963 ;
  assign n27310 = n27309 ^ n10003 ^ 1'b0 ;
  assign n27311 = n10542 | n27310 ;
  assign n27312 = n23931 & ~n27311 ;
  assign n27313 = n10921 & ~n12900 ;
  assign n27314 = n8515 & n27313 ;
  assign n27315 = ~n11215 & n27314 ;
  assign n27316 = n27315 ^ n13708 ^ 1'b0 ;
  assign n27317 = ( x224 & n17385 ) | ( x224 & ~n26042 ) | ( n17385 & ~n26042 ) ;
  assign n27318 = ( n4876 & ~n6252 ) | ( n4876 & n7555 ) | ( ~n6252 & n7555 ) ;
  assign n27319 = n6720 & ~n13488 ;
  assign n27320 = n27319 ^ n16350 ^ 1'b0 ;
  assign n27321 = n27320 ^ n17201 ^ n13632 ;
  assign n27322 = n11859 ^ n10556 ^ 1'b0 ;
  assign n27324 = n5333 ^ n4670 ^ 1'b0 ;
  assign n27325 = n5948 | n27324 ;
  assign n27326 = n15578 | n27325 ;
  assign n27327 = n9726 | n27326 ;
  assign n27323 = ~n10295 & n13461 ;
  assign n27328 = n27327 ^ n27323 ^ 1'b0 ;
  assign n27329 = n18939 ^ n6914 ^ n5209 ;
  assign n27330 = ( ~n8604 & n13588 ) | ( ~n8604 & n27329 ) | ( n13588 & n27329 ) ;
  assign n27331 = ( n7119 & ~n19778 ) | ( n7119 & n24595 ) | ( ~n19778 & n24595 ) ;
  assign n27332 = n8430 | n18046 ;
  assign n27333 = n27332 ^ n17037 ^ 1'b0 ;
  assign n27334 = n19619 ^ n663 ^ 1'b0 ;
  assign n27335 = n21875 ^ n2683 ^ 1'b0 ;
  assign n27336 = n26209 | n27335 ;
  assign n27337 = n27334 | n27336 ;
  assign n27338 = n2328 | n7800 ;
  assign n27339 = n258 & ~n27338 ;
  assign n27340 = n27277 ^ n22405 ^ 1'b0 ;
  assign n27341 = n27339 | n27340 ;
  assign n27342 = n490 & n1903 ;
  assign n27343 = ( n2130 & ~n22639 ) | ( n2130 & n27342 ) | ( ~n22639 & n27342 ) ;
  assign n27344 = n9278 & ~n27343 ;
  assign n27345 = n27344 ^ n24044 ^ 1'b0 ;
  assign n27346 = n9197 ^ n4436 ^ n2661 ;
  assign n27349 = n15279 ^ n13591 ^ 1'b0 ;
  assign n27350 = n27349 ^ n8906 ^ n649 ;
  assign n27347 = n7802 & ~n22616 ;
  assign n27348 = n7042 & n27347 ;
  assign n27351 = n27350 ^ n27348 ^ n25841 ;
  assign n27352 = n3001 & n6886 ;
  assign n27353 = ~n20784 & n23172 ;
  assign n27354 = n27352 & n27353 ;
  assign n27355 = n5961 ^ x202 ^ 1'b0 ;
  assign n27358 = ( n958 & n7261 ) | ( n958 & ~n10896 ) | ( n7261 & ~n10896 ) ;
  assign n27356 = n12037 ^ n10834 ^ 1'b0 ;
  assign n27357 = n7935 & ~n27356 ;
  assign n27359 = n27358 ^ n27357 ^ 1'b0 ;
  assign n27360 = ~x224 & n13310 ;
  assign n27361 = n5205 & n20172 ;
  assign n27362 = n18861 ^ n14994 ^ 1'b0 ;
  assign n27363 = n14583 ^ n1947 ^ 1'b0 ;
  assign n27364 = ~n9276 & n27363 ;
  assign n27365 = n17551 ^ n1795 ^ 1'b0 ;
  assign n27366 = ~n4512 & n23535 ;
  assign n27367 = n27365 & n27366 ;
  assign n27368 = n15290 ^ n11649 ^ 1'b0 ;
  assign n27369 = ~n13299 & n20626 ;
  assign n27370 = n27368 & n27369 ;
  assign n27371 = n16674 ^ n15734 ^ n1737 ;
  assign n27372 = ( n1889 & ~n9371 ) | ( n1889 & n23301 ) | ( ~n9371 & n23301 ) ;
  assign n27373 = ( n18101 & ~n20741 ) | ( n18101 & n27372 ) | ( ~n20741 & n27372 ) ;
  assign n27374 = ( n13421 & n19709 ) | ( n13421 & n27373 ) | ( n19709 & n27373 ) ;
  assign n27376 = n9268 ^ n6150 ^ n2834 ;
  assign n27375 = ( n399 & n12442 ) | ( n399 & n17917 ) | ( n12442 & n17917 ) ;
  assign n27377 = n27376 ^ n27375 ^ n17867 ;
  assign n27380 = n6316 ^ n2793 ^ 1'b0 ;
  assign n27381 = n10761 & n27380 ;
  assign n27378 = n9039 ^ n3534 ^ 1'b0 ;
  assign n27379 = n8850 | n27378 ;
  assign n27382 = n27381 ^ n27379 ^ n3306 ;
  assign n27383 = ~n18976 & n27382 ;
  assign n27384 = ~n1135 & n27383 ;
  assign n27385 = ~n11212 & n17305 ;
  assign n27386 = n949 & n27385 ;
  assign n27387 = n19776 & ~n27386 ;
  assign n27388 = n686 & n2438 ;
  assign n27392 = ( n1321 & ~n6936 ) | ( n1321 & n14843 ) | ( ~n6936 & n14843 ) ;
  assign n27389 = n9278 ^ n5796 ^ 1'b0 ;
  assign n27390 = n13115 ^ n4424 ^ 1'b0 ;
  assign n27391 = n27389 | n27390 ;
  assign n27393 = n27392 ^ n27391 ^ 1'b0 ;
  assign n27394 = n27388 & n27393 ;
  assign n27395 = n19628 ^ n8105 ^ n3133 ;
  assign n27396 = n13665 & ~n27395 ;
  assign n27397 = n27396 ^ n10955 ^ n2613 ;
  assign n27398 = n22391 ^ n22221 ^ 1'b0 ;
  assign n27399 = n9693 ^ n9076 ^ 1'b0 ;
  assign n27400 = ( ~n1127 & n5490 ) | ( ~n1127 & n25388 ) | ( n5490 & n25388 ) ;
  assign n27401 = ( n21487 & ~n21647 ) | ( n21487 & n23494 ) | ( ~n21647 & n23494 ) ;
  assign n27402 = ( n5306 & n27103 ) | ( n5306 & n27401 ) | ( n27103 & n27401 ) ;
  assign n27403 = ~n4351 & n27402 ;
  assign n27404 = ~n27400 & n27403 ;
  assign n27405 = ( ~n1752 & n16101 ) | ( ~n1752 & n27404 ) | ( n16101 & n27404 ) ;
  assign n27406 = n6332 ^ n4471 ^ 1'b0 ;
  assign n27407 = ~n7221 & n27406 ;
  assign n27408 = n17209 & ~n26477 ;
  assign n27409 = n21785 & n27408 ;
  assign n27410 = n19759 | n25779 ;
  assign n27411 = n10509 | n27410 ;
  assign n27412 = n4636 | n6767 ;
  assign n27413 = n2240 & ~n27412 ;
  assign n27414 = ~n259 & n4715 ;
  assign n27415 = n27414 ^ n25174 ^ 1'b0 ;
  assign n27416 = n2586 & ~n27415 ;
  assign n27417 = n27416 ^ n26518 ^ 1'b0 ;
  assign n27418 = n27256 ^ n7605 ^ 1'b0 ;
  assign n27419 = n27417 & ~n27418 ;
  assign n27420 = ~n24865 & n27419 ;
  assign n27421 = n8457 | n27420 ;
  assign n27422 = n27421 ^ n1049 ^ 1'b0 ;
  assign n27423 = n10717 ^ n10474 ^ 1'b0 ;
  assign n27424 = n9500 & ~n27423 ;
  assign n27425 = n27424 ^ n15228 ^ 1'b0 ;
  assign n27426 = n23052 ^ n15394 ^ n5539 ;
  assign n27427 = n27426 ^ n12907 ^ 1'b0 ;
  assign n27428 = n3499 & ~n27427 ;
  assign n27429 = n2440 | n10502 ;
  assign n27430 = ( n14220 & n23607 ) | ( n14220 & ~n27429 ) | ( n23607 & ~n27429 ) ;
  assign n27431 = ( n11865 & n27428 ) | ( n11865 & n27430 ) | ( n27428 & n27430 ) ;
  assign n27432 = n2282 & n10963 ;
  assign n27433 = n27432 ^ n6136 ^ 1'b0 ;
  assign n27434 = ( n12594 & ~n15561 ) | ( n12594 & n16314 ) | ( ~n15561 & n16314 ) ;
  assign n27435 = ( n16555 & ~n27433 ) | ( n16555 & n27434 ) | ( ~n27433 & n27434 ) ;
  assign n27436 = n16409 ^ n4383 ^ 1'b0 ;
  assign n27437 = n3816 | n27436 ;
  assign n27438 = ( n4410 & n26128 ) | ( n4410 & n27437 ) | ( n26128 & n27437 ) ;
  assign n27439 = ~n5697 & n23882 ;
  assign n27440 = n3613 & ~n8727 ;
  assign n27441 = n11794 | n27440 ;
  assign n27442 = n24313 & ~n27441 ;
  assign n27443 = ( n1176 & n3332 ) | ( n1176 & n11768 ) | ( n3332 & n11768 ) ;
  assign n27444 = ~n8648 & n20237 ;
  assign n27445 = n27444 ^ n6923 ^ n2081 ;
  assign n27446 = n5318 | n11129 ;
  assign n27447 = n24919 ^ n14274 ^ n518 ;
  assign n27448 = n27446 & n27447 ;
  assign n27449 = ( ~x174 & n1589 ) | ( ~x174 & n27448 ) | ( n1589 & n27448 ) ;
  assign n27450 = n1961 ^ n879 ^ 1'b0 ;
  assign n27451 = n3715 & n25338 ;
  assign n27453 = n9150 & n24982 ;
  assign n27452 = n24499 ^ n23482 ^ 1'b0 ;
  assign n27454 = n27453 ^ n27452 ^ n15720 ;
  assign n27455 = n15806 | n20805 ;
  assign n27456 = n23458 ^ n22142 ^ n4710 ;
  assign n27457 = n27456 ^ n13127 ^ 1'b0 ;
  assign n27458 = n27457 ^ n25307 ^ n7390 ;
  assign n27459 = n15327 ^ n4886 ^ n4224 ;
  assign n27460 = n3707 | n27459 ;
  assign n27461 = n18978 & ~n27460 ;
  assign n27462 = n6043 | n18449 ;
  assign n27463 = n799 & ~n27462 ;
  assign n27464 = x223 & ~n27463 ;
  assign n27465 = n27461 & n27464 ;
  assign n27466 = n27465 ^ n13484 ^ 1'b0 ;
  assign n27474 = n2704 ^ n2191 ^ n393 ;
  assign n27468 = n7108 & n14452 ;
  assign n27469 = n27468 ^ n397 ^ 1'b0 ;
  assign n27470 = n27469 ^ n4250 ^ n1324 ;
  assign n27471 = n27470 ^ n9463 ^ n4139 ;
  assign n27472 = n18800 ^ n13866 ^ n10816 ;
  assign n27473 = ( n11553 & n27471 ) | ( n11553 & ~n27472 ) | ( n27471 & ~n27472 ) ;
  assign n27467 = ~n16399 & n21900 ;
  assign n27475 = n27474 ^ n27473 ^ n27467 ;
  assign n27476 = ( n918 & n4201 ) | ( n918 & n10284 ) | ( n4201 & n10284 ) ;
  assign n27477 = n3921 & ~n6387 ;
  assign n27478 = n14450 & n27477 ;
  assign n27479 = n24373 & ~n27478 ;
  assign n27480 = ~n27476 & n27479 ;
  assign n27481 = n23896 ^ n14117 ^ n3722 ;
  assign n27482 = n12061 & ~n27481 ;
  assign n27483 = n11857 & n27482 ;
  assign n27484 = ~n432 & n7425 ;
  assign n27485 = n27484 ^ n13012 ^ 1'b0 ;
  assign n27486 = ( n6031 & ~n9510 ) | ( n6031 & n27485 ) | ( ~n9510 & n27485 ) ;
  assign n27487 = n17096 ^ n10954 ^ 1'b0 ;
  assign n27488 = n27487 ^ n8187 ^ 1'b0 ;
  assign n27489 = ( n22127 & n27486 ) | ( n22127 & n27488 ) | ( n27486 & n27488 ) ;
  assign n27490 = n10524 & n21220 ;
  assign n27491 = n27490 ^ n18172 ^ 1'b0 ;
  assign n27492 = n27491 ^ n9188 ^ 1'b0 ;
  assign n27493 = n2925 & n13890 ;
  assign n27494 = n13945 & n27493 ;
  assign n27495 = n1824 & ~n27494 ;
  assign n27496 = ~n9013 & n11938 ;
  assign n27497 = n13771 & n15543 ;
  assign n27498 = ~n27496 & n27497 ;
  assign n27499 = n1374 | n17139 ;
  assign n27500 = n20911 ^ n6107 ^ n4605 ;
  assign n27501 = n4098 & n27500 ;
  assign n27502 = n10903 & ~n19211 ;
  assign n27503 = n12213 & n12973 ;
  assign n27504 = ~n5172 & n27503 ;
  assign n27505 = n25904 ^ n21706 ^ n3647 ;
  assign n27506 = n5736 & ~n17068 ;
  assign n27507 = n27506 ^ n22340 ^ 1'b0 ;
  assign n27508 = n11371 & ~n14341 ;
  assign n27509 = n4954 ^ n4109 ^ n738 ;
  assign n27510 = ( n8332 & ~n9772 ) | ( n8332 & n27509 ) | ( ~n9772 & n27509 ) ;
  assign n27511 = n3894 | n25044 ;
  assign n27512 = n27510 & ~n27511 ;
  assign n27513 = ~n10865 & n15552 ;
  assign n27514 = n27513 ^ n9557 ^ 1'b0 ;
  assign n27515 = ( n1861 & ~n17651 ) | ( n1861 & n24749 ) | ( ~n17651 & n24749 ) ;
  assign n27516 = n5851 & n27515 ;
  assign n27517 = ( ~n8282 & n21322 ) | ( ~n8282 & n27516 ) | ( n21322 & n27516 ) ;
  assign n27522 = ~n18171 & n25369 ;
  assign n27523 = n27522 ^ n5968 ^ 1'b0 ;
  assign n27520 = n10218 | n12005 ;
  assign n27521 = x103 | n27520 ;
  assign n27518 = n11706 ^ n10848 ^ 1'b0 ;
  assign n27519 = n330 | n27518 ;
  assign n27524 = n27523 ^ n27521 ^ n27519 ;
  assign n27525 = n15140 ^ n2913 ^ n1639 ;
  assign n27526 = ( n5060 & n7862 ) | ( n5060 & ~n27525 ) | ( n7862 & ~n27525 ) ;
  assign n27527 = n13993 ^ n8151 ^ n436 ;
  assign n27528 = n11405 ^ n5880 ^ n2748 ;
  assign n27529 = n15794 | n27528 ;
  assign n27530 = x175 & n27529 ;
  assign n27531 = n27527 & n27530 ;
  assign n27532 = n16081 ^ n13275 ^ n12705 ;
  assign n27533 = n2229 & ~n5853 ;
  assign n27534 = n27533 ^ n25453 ^ n21396 ;
  assign n27535 = n9211 & n27534 ;
  assign n27536 = ~n27532 & n27535 ;
  assign n27537 = n10269 ^ n8284 ^ n6595 ;
  assign n27538 = ( ~n405 & n1583 ) | ( ~n405 & n4314 ) | ( n1583 & n4314 ) ;
  assign n27539 = n3819 ^ n2782 ^ 1'b0 ;
  assign n27540 = n2089 | n27539 ;
  assign n27541 = ( n27537 & ~n27538 ) | ( n27537 & n27540 ) | ( ~n27538 & n27540 ) ;
  assign n27542 = x108 & ~n13239 ;
  assign n27543 = n8965 & n27542 ;
  assign n27544 = n27543 ^ n14701 ^ 1'b0 ;
  assign n27545 = n21053 & n27544 ;
  assign n27546 = n7337 & n13741 ;
  assign n27547 = ~n16918 & n27546 ;
  assign n27548 = n20060 ^ n5551 ^ 1'b0 ;
  assign n27549 = n3401 & n27548 ;
  assign n27550 = n27549 ^ n2218 ^ 1'b0 ;
  assign n27551 = ~n27547 & n27550 ;
  assign n27552 = ~n18246 & n27551 ;
  assign n27554 = n5244 & n7026 ;
  assign n27553 = n18530 ^ n3985 ^ 1'b0 ;
  assign n27555 = n27554 ^ n27553 ^ n8560 ;
  assign n27556 = n15570 | n21194 ;
  assign n27557 = n12630 | n27556 ;
  assign n27558 = n27557 ^ n25528 ^ 1'b0 ;
  assign n27559 = n4429 & ~n18892 ;
  assign n27560 = ~n3646 & n18778 ;
  assign n27561 = ( n3696 & ~n20689 ) | ( n3696 & n27560 ) | ( ~n20689 & n27560 ) ;
  assign n27562 = n614 & n7782 ;
  assign n27563 = n27562 ^ n18165 ^ 1'b0 ;
  assign n27564 = ( n2637 & n8790 ) | ( n2637 & n27563 ) | ( n8790 & n27563 ) ;
  assign n27565 = n27564 ^ n23264 ^ n17511 ;
  assign n27566 = n18967 ^ n4686 ^ 1'b0 ;
  assign n27567 = n1920 & ~n27566 ;
  assign n27568 = n18929 & n27567 ;
  assign n27569 = n2065 & n27568 ;
  assign n27570 = ( n388 & n10499 ) | ( n388 & n19369 ) | ( n10499 & n19369 ) ;
  assign n27571 = n1664 & ~n13113 ;
  assign n27572 = n27571 ^ n1933 ^ 1'b0 ;
  assign n27573 = n27570 & n27572 ;
  assign n27576 = n19464 ^ n1641 ^ n703 ;
  assign n27574 = ( n5458 & n8923 ) | ( n5458 & ~n9151 ) | ( n8923 & ~n9151 ) ;
  assign n27575 = n27574 ^ n10540 ^ n9934 ;
  assign n27577 = n27576 ^ n27575 ^ 1'b0 ;
  assign n27578 = n25412 & n27577 ;
  assign n27579 = ~n10041 & n14030 ;
  assign n27580 = n27579 ^ n11422 ^ 1'b0 ;
  assign n27581 = n17198 & ~n21048 ;
  assign n27582 = n9972 & n27581 ;
  assign n27583 = n27582 ^ n25141 ^ n1311 ;
  assign n27584 = ~n3928 & n21727 ;
  assign n27585 = n27584 ^ n2220 ^ 1'b0 ;
  assign n27586 = ( ~n1247 & n11370 ) | ( ~n1247 & n13776 ) | ( n11370 & n13776 ) ;
  assign n27587 = ( n6543 & ~n22921 ) | ( n6543 & n27586 ) | ( ~n22921 & n27586 ) ;
  assign n27588 = ~n17398 & n21728 ;
  assign n27589 = n4318 | n10591 ;
  assign n27590 = n27589 ^ n16163 ^ 1'b0 ;
  assign n27591 = ( n4921 & n10230 ) | ( n4921 & n27590 ) | ( n10230 & n27590 ) ;
  assign n27592 = ( n2328 & ~n9640 ) | ( n2328 & n18266 ) | ( ~n9640 & n18266 ) ;
  assign n27593 = n5937 ^ n1969 ^ 1'b0 ;
  assign n27594 = n8670 & ~n27593 ;
  assign n27595 = n6396 & n27594 ;
  assign n27596 = ~n18373 & n27595 ;
  assign n27597 = n25319 ^ n2624 ^ 1'b0 ;
  assign n27598 = n11454 | n27597 ;
  assign n27599 = n5642 & ~n8111 ;
  assign n27600 = n27599 ^ n11872 ^ 1'b0 ;
  assign n27601 = n21479 & n27600 ;
  assign n27602 = ( n4624 & n11720 ) | ( n4624 & ~n15811 ) | ( n11720 & ~n15811 ) ;
  assign n27603 = ( ~n9218 & n9769 ) | ( ~n9218 & n27602 ) | ( n9769 & n27602 ) ;
  assign n27604 = ~n10580 & n16523 ;
  assign n27605 = n13578 & n27604 ;
  assign n27606 = n19980 | n27605 ;
  assign n27607 = n27606 ^ n5318 ^ 1'b0 ;
  assign n27608 = n27459 ^ n16108 ^ n14684 ;
  assign n27609 = ( n26542 & ~n27607 ) | ( n26542 & n27608 ) | ( ~n27607 & n27608 ) ;
  assign n27610 = n8183 ^ n4941 ^ 1'b0 ;
  assign n27611 = n27610 ^ n19541 ^ 1'b0 ;
  assign n27614 = n26173 ^ n8731 ^ n4979 ;
  assign n27615 = ~n25097 & n27614 ;
  assign n27616 = n25839 & n27615 ;
  assign n27612 = n19709 ^ n4095 ^ 1'b0 ;
  assign n27613 = n7283 | n27612 ;
  assign n27617 = n27616 ^ n27613 ^ 1'b0 ;
  assign n27618 = n3784 | n3858 ;
  assign n27619 = n13412 ^ n12162 ^ 1'b0 ;
  assign n27622 = ( ~n3679 & n4189 ) | ( ~n3679 & n5646 ) | ( n4189 & n5646 ) ;
  assign n27620 = n6406 & n17047 ;
  assign n27621 = n4788 & n27620 ;
  assign n27623 = n27622 ^ n27621 ^ x66 ;
  assign n27624 = n27623 ^ n676 ^ 1'b0 ;
  assign n27625 = ( n27618 & n27619 ) | ( n27618 & ~n27624 ) | ( n27619 & ~n27624 ) ;
  assign n27626 = n19564 ^ n16858 ^ 1'b0 ;
  assign n27627 = ( n5869 & ~n10139 ) | ( n5869 & n26566 ) | ( ~n10139 & n26566 ) ;
  assign n27628 = ( n18703 & ~n19689 ) | ( n18703 & n27627 ) | ( ~n19689 & n27627 ) ;
  assign n27629 = n4292 & ~n7659 ;
  assign n27630 = n2268 & n27629 ;
  assign n27631 = ~n19053 & n27630 ;
  assign n27632 = n27628 & ~n27631 ;
  assign n27633 = n27632 ^ n12624 ^ 1'b0 ;
  assign n27634 = ( ~n4965 & n14120 ) | ( ~n4965 & n25867 ) | ( n14120 & n25867 ) ;
  assign n27635 = n24520 ^ n23189 ^ n8343 ;
  assign n27636 = ~n4680 & n17358 ;
  assign n27637 = ~x0 & n27636 ;
  assign n27638 = n25480 ^ n18741 ^ 1'b0 ;
  assign n27639 = n20411 ^ n19886 ^ 1'b0 ;
  assign n27640 = n24266 & n27639 ;
  assign n27641 = ( n5302 & n12525 ) | ( n5302 & ~n27640 ) | ( n12525 & ~n27640 ) ;
  assign n27642 = n4935 | n8460 ;
  assign n27643 = n27642 ^ n388 ^ 1'b0 ;
  assign n27644 = n3001 | n27643 ;
  assign n27645 = n19216 | n27644 ;
  assign n27646 = ( n10691 & n27641 ) | ( n10691 & ~n27645 ) | ( n27641 & ~n27645 ) ;
  assign n27647 = n17943 ^ n5080 ^ 1'b0 ;
  assign n27648 = ( n1554 & n10956 ) | ( n1554 & n27647 ) | ( n10956 & n27647 ) ;
  assign n27649 = n27648 ^ n8399 ^ x18 ;
  assign n27650 = n27649 ^ n21153 ^ n15699 ;
  assign n27651 = n25928 ^ n1934 ^ 1'b0 ;
  assign n27652 = ( n12606 & ~n24698 ) | ( n12606 & n27651 ) | ( ~n24698 & n27651 ) ;
  assign n27653 = n12179 & ~n15262 ;
  assign n27654 = n27653 ^ n13850 ^ 1'b0 ;
  assign n27655 = n15666 & n27654 ;
  assign n27656 = n13327 | n27655 ;
  assign n27657 = n27656 ^ n455 ^ 1'b0 ;
  assign n27658 = ( n7141 & n20896 ) | ( n7141 & ~n22796 ) | ( n20896 & ~n22796 ) ;
  assign n27659 = n4206 | n27658 ;
  assign n27660 = n19861 | n27659 ;
  assign n27661 = n25188 ^ n23420 ^ 1'b0 ;
  assign n27662 = n2116 | n11131 ;
  assign n27663 = n27662 ^ n4587 ^ 1'b0 ;
  assign n27664 = n8309 & ~n14186 ;
  assign n27665 = n27664 ^ n6847 ^ 1'b0 ;
  assign n27666 = ( ~n25613 & n27663 ) | ( ~n25613 & n27665 ) | ( n27663 & n27665 ) ;
  assign n27667 = n24695 ^ n15057 ^ 1'b0 ;
  assign n27668 = n27667 ^ n22221 ^ n17638 ;
  assign n27669 = ( ~n6787 & n8080 ) | ( ~n6787 & n21284 ) | ( n8080 & n21284 ) ;
  assign n27670 = ~n12907 & n27669 ;
  assign n27671 = n27670 ^ n2773 ^ 1'b0 ;
  assign n27679 = n15972 ^ n7675 ^ 1'b0 ;
  assign n27673 = x11 & ~n6904 ;
  assign n27672 = n10166 | n11279 ;
  assign n27674 = n27673 ^ n27672 ^ 1'b0 ;
  assign n27675 = ~n1440 & n27674 ;
  assign n27676 = n1440 & n27675 ;
  assign n27677 = n3099 | n6884 ;
  assign n27678 = n27676 & ~n27677 ;
  assign n27680 = n27679 ^ n27678 ^ x251 ;
  assign n27681 = n21157 ^ n1743 ^ 1'b0 ;
  assign n27682 = ( n3315 & ~n15432 ) | ( n3315 & n23995 ) | ( ~n15432 & n23995 ) ;
  assign n27683 = n21321 & ~n27682 ;
  assign n27684 = n27683 ^ n14938 ^ 1'b0 ;
  assign n27685 = n16863 | n27684 ;
  assign n27686 = n27681 | n27685 ;
  assign n27687 = n8097 ^ n4619 ^ 1'b0 ;
  assign n27688 = ~n18795 & n27687 ;
  assign n27689 = n27688 ^ n4409 ^ 1'b0 ;
  assign n27690 = n637 & ~n26377 ;
  assign n27691 = n27690 ^ n923 ^ 1'b0 ;
  assign n27692 = ( n15569 & n16018 ) | ( n15569 & n27691 ) | ( n16018 & n27691 ) ;
  assign n27693 = n11166 & ~n23314 ;
  assign n27694 = n27693 ^ n10849 ^ 1'b0 ;
  assign n27695 = n14708 | n18459 ;
  assign n27696 = n15123 & ~n27695 ;
  assign n27697 = ( n4963 & ~n23771 ) | ( n4963 & n27696 ) | ( ~n23771 & n27696 ) ;
  assign n27698 = n27697 ^ n770 ^ 1'b0 ;
  assign n27699 = n25429 ^ n18900 ^ n2595 ;
  assign n27700 = n8116 ^ n4454 ^ 1'b0 ;
  assign n27701 = n8974 ^ n1658 ^ 1'b0 ;
  assign n27702 = n1381 & n27701 ;
  assign n27703 = ~n27700 & n27702 ;
  assign n27704 = n7922 ^ n4823 ^ 1'b0 ;
  assign n27705 = ( n27699 & n27703 ) | ( n27699 & n27704 ) | ( n27703 & n27704 ) ;
  assign n27706 = ~n13593 & n18814 ;
  assign n27707 = ~n14899 & n27706 ;
  assign n27708 = x65 & n27707 ;
  assign n27709 = ( n19174 & n21285 ) | ( n19174 & ~n27708 ) | ( n21285 & ~n27708 ) ;
  assign n27710 = ( n2274 & n6355 ) | ( n2274 & n27709 ) | ( n6355 & n27709 ) ;
  assign n27711 = n18025 | n27710 ;
  assign n27712 = n12323 | n14297 ;
  assign n27713 = n8787 | n27712 ;
  assign n27714 = n27713 ^ n8698 ^ n4912 ;
  assign n27715 = ( n3384 & n4334 ) | ( n3384 & ~n4841 ) | ( n4334 & ~n4841 ) ;
  assign n27716 = n14791 & n15913 ;
  assign n27717 = n27715 & ~n27716 ;
  assign n27718 = ~n1646 & n27717 ;
  assign n27719 = n27718 ^ n20583 ^ n12576 ;
  assign n27720 = n21352 ^ n13785 ^ n8004 ;
  assign n27721 = ~n26528 & n27720 ;
  assign n27722 = n14309 & n27721 ;
  assign n27723 = n20786 ^ n6358 ^ 1'b0 ;
  assign n27724 = ~n27722 & n27723 ;
  assign n27725 = n27724 ^ n27619 ^ 1'b0 ;
  assign n27726 = n10631 ^ n2281 ^ 1'b0 ;
  assign n27727 = n4199 & n27726 ;
  assign n27728 = n26681 ^ n18863 ^ 1'b0 ;
  assign n27729 = n15590 ^ n6192 ^ 1'b0 ;
  assign n27730 = n12404 & ~n27729 ;
  assign n27731 = n15036 ^ x85 ^ 1'b0 ;
  assign n27732 = ( n716 & ~n12266 ) | ( n716 & n21004 ) | ( ~n12266 & n21004 ) ;
  assign n27733 = n27732 ^ n22030 ^ n15170 ;
  assign n27734 = n12738 ^ n12237 ^ n2774 ;
  assign n27735 = n19433 ^ n8452 ^ 1'b0 ;
  assign n27736 = n10524 & ~n27735 ;
  assign n27737 = ( n23612 & n27734 ) | ( n23612 & n27736 ) | ( n27734 & n27736 ) ;
  assign n27738 = n17392 ^ n13740 ^ n7462 ;
  assign n27739 = n26219 ^ n14098 ^ 1'b0 ;
  assign n27740 = n27738 & ~n27739 ;
  assign n27741 = n27740 ^ n16611 ^ 1'b0 ;
  assign n27742 = n14102 | n27741 ;
  assign n27743 = n2561 & n5765 ;
  assign n27744 = n6460 & n11591 ;
  assign n27745 = n4694 ^ x82 ^ 1'b0 ;
  assign n27746 = ~n14622 & n27745 ;
  assign n27747 = n12399 & n27746 ;
  assign n27748 = n27744 & ~n27747 ;
  assign n27749 = n18924 & n27748 ;
  assign n27751 = n6159 ^ n3009 ^ n1067 ;
  assign n27750 = n3883 | n10688 ;
  assign n27752 = n27751 ^ n27750 ^ 1'b0 ;
  assign n27753 = ( n2645 & n3254 ) | ( n2645 & n27752 ) | ( n3254 & n27752 ) ;
  assign n27754 = n524 & ~n27753 ;
  assign n27755 = ~n9414 & n27754 ;
  assign n27756 = ( n9378 & n25496 ) | ( n9378 & n27540 ) | ( n25496 & n27540 ) ;
  assign n27757 = n452 ^ n354 ^ 1'b0 ;
  assign n27758 = ~n6456 & n27757 ;
  assign n27759 = n10723 ^ n9594 ^ n7788 ;
  assign n27760 = n27759 ^ n18169 ^ 1'b0 ;
  assign n27761 = n3335 | n27760 ;
  assign n27762 = ( n8607 & n27758 ) | ( n8607 & ~n27761 ) | ( n27758 & ~n27761 ) ;
  assign n27763 = ( ~n9365 & n16484 ) | ( ~n9365 & n21682 ) | ( n16484 & n21682 ) ;
  assign n27766 = n2993 & ~n10684 ;
  assign n27764 = n16164 & ~n19840 ;
  assign n27765 = n2649 & n27764 ;
  assign n27767 = n27766 ^ n27765 ^ 1'b0 ;
  assign n27768 = n25630 | n27767 ;
  assign n27769 = n27478 ^ n22246 ^ n21348 ;
  assign n27770 = n19509 ^ n15827 ^ 1'b0 ;
  assign n27771 = n20115 ^ n6705 ^ n2043 ;
  assign n27772 = n27771 ^ n13340 ^ 1'b0 ;
  assign n27773 = n2223 | n18327 ;
  assign n27774 = n3264 & ~n27773 ;
  assign n27775 = n27774 ^ n20392 ^ n16699 ;
  assign n27776 = n962 | n10880 ;
  assign n27777 = n1107 | n27776 ;
  assign n27778 = n27777 ^ n26952 ^ n17773 ;
  assign n27779 = ~n27775 & n27778 ;
  assign n27780 = x55 | n8705 ;
  assign n27781 = n3530 | n21703 ;
  assign n27782 = n27781 ^ n22798 ^ 1'b0 ;
  assign n27783 = n2041 & n15842 ;
  assign n27784 = ( n17081 & ~n26414 ) | ( n17081 & n27783 ) | ( ~n26414 & n27783 ) ;
  assign n27785 = ( n1120 & n17652 ) | ( n1120 & n27784 ) | ( n17652 & n27784 ) ;
  assign n27786 = n16495 ^ n413 ^ 1'b0 ;
  assign n27787 = n7285 & n15668 ;
  assign n27788 = ~n5716 & n27787 ;
  assign n27789 = n18027 ^ n3167 ^ 1'b0 ;
  assign n27790 = n27788 | n27789 ;
  assign n27791 = n6870 ^ n2156 ^ 1'b0 ;
  assign n27792 = n12162 & ~n27791 ;
  assign n27793 = ~n9053 & n27792 ;
  assign n27794 = n24610 | n27793 ;
  assign n27795 = ( n11247 & n27790 ) | ( n11247 & ~n27794 ) | ( n27790 & ~n27794 ) ;
  assign n27796 = n10774 ^ n5460 ^ 1'b0 ;
  assign n27797 = n24267 & ~n27796 ;
  assign n27798 = n14664 ^ n5100 ^ 1'b0 ;
  assign n27799 = x156 & ~n27798 ;
  assign n27800 = n9143 ^ n2531 ^ 1'b0 ;
  assign n27801 = n25759 | n27800 ;
  assign n27802 = n27801 ^ n7752 ^ 1'b0 ;
  assign n27803 = n14786 & ~n27802 ;
  assign n27804 = n27799 & ~n27803 ;
  assign n27807 = ~n12709 & n17327 ;
  assign n27808 = n23490 & n27807 ;
  assign n27805 = n6636 ^ n4905 ^ 1'b0 ;
  assign n27806 = n294 & ~n27805 ;
  assign n27809 = n27808 ^ n27806 ^ 1'b0 ;
  assign n27810 = n1287 & n17023 ;
  assign n27811 = ~n23805 & n27810 ;
  assign n27812 = n1379 | n3856 ;
  assign n27813 = n5500 & ~n27812 ;
  assign n27814 = ~n3042 & n27813 ;
  assign n27815 = n21856 ^ n4435 ^ 1'b0 ;
  assign n27816 = ~n3623 & n27815 ;
  assign n27817 = n2465 & n14874 ;
  assign n27818 = ( n17600 & n18538 ) | ( n17600 & n27817 ) | ( n18538 & n27817 ) ;
  assign n27819 = n980 & n9109 ;
  assign n27820 = ~n2466 & n27819 ;
  assign n27821 = ( n14464 & n18602 ) | ( n14464 & ~n27820 ) | ( n18602 & ~n27820 ) ;
  assign n27822 = n25361 & n27821 ;
  assign n27823 = n12202 ^ n5496 ^ n4029 ;
  assign n27824 = n8776 & ~n27823 ;
  assign n27825 = n2532 ^ n402 ^ 1'b0 ;
  assign n27826 = n3034 | n27825 ;
  assign n27827 = n27826 ^ n19770 ^ 1'b0 ;
  assign n27828 = n27827 ^ n25536 ^ n22125 ;
  assign n27829 = n27828 ^ n26605 ^ 1'b0 ;
  assign n27830 = n24673 & n26974 ;
  assign n27831 = ~n13167 & n18424 ;
  assign n27832 = n17572 | n20453 ;
  assign n27833 = n8972 | n27832 ;
  assign n27834 = n27833 ^ n2386 ^ 1'b0 ;
  assign n27835 = n3120 & n17887 ;
  assign n27836 = n27835 ^ n4975 ^ 1'b0 ;
  assign n27837 = ( n15119 & ~n18169 ) | ( n15119 & n18284 ) | ( ~n18169 & n18284 ) ;
  assign n27838 = ~n2945 & n27837 ;
  assign n27839 = n24751 ^ n10339 ^ n4527 ;
  assign n27840 = n19278 ^ n16167 ^ 1'b0 ;
  assign n27841 = ~n26192 & n27840 ;
  assign n27842 = ( n2961 & ~n6394 ) | ( n2961 & n7815 ) | ( ~n6394 & n7815 ) ;
  assign n27843 = n23167 | n27842 ;
  assign n27844 = ( n4376 & n16778 ) | ( n4376 & ~n18140 ) | ( n16778 & ~n18140 ) ;
  assign n27845 = n27844 ^ n5990 ^ 1'b0 ;
  assign n27846 = n1884 & ~n20462 ;
  assign n27847 = n27846 ^ n24620 ^ n9626 ;
  assign n27848 = n2812 | n17044 ;
  assign n27849 = n27848 ^ n4206 ^ 1'b0 ;
  assign n27850 = n4532 ^ n4507 ^ x133 ;
  assign n27851 = ~n27849 & n27850 ;
  assign n27852 = ~n19579 & n27851 ;
  assign n27853 = n9188 ^ n4488 ^ 1'b0 ;
  assign n27854 = n8543 ^ n5947 ^ n1643 ;
  assign n27855 = ( n4618 & n11112 ) | ( n4618 & n27854 ) | ( n11112 & n27854 ) ;
  assign n27856 = n27855 ^ n10361 ^ n4659 ;
  assign n27857 = n9377 ^ n5385 ^ n1494 ;
  assign n27858 = n27857 ^ n16784 ^ n6967 ;
  assign n27859 = ~n15731 & n27858 ;
  assign n27860 = n8906 & ~n23279 ;
  assign n27861 = ~n481 & n27860 ;
  assign n27862 = n7952 | n14648 ;
  assign n27863 = n5208 | n27862 ;
  assign n27864 = n11789 | n27863 ;
  assign n27865 = n27864 ^ n18886 ^ 1'b0 ;
  assign n27866 = n2620 & n27865 ;
  assign n27867 = ~n1334 & n27515 ;
  assign n27868 = n4959 ^ n4820 ^ 1'b0 ;
  assign n27869 = n16847 ^ n9739 ^ n7081 ;
  assign n27870 = ( n8289 & ~n27868 ) | ( n8289 & n27869 ) | ( ~n27868 & n27869 ) ;
  assign n27871 = n17707 ^ n15758 ^ n6332 ;
  assign n27872 = n10688 | n17401 ;
  assign n27873 = n27872 ^ n18195 ^ n15572 ;
  assign n27876 = ~n609 & n6390 ;
  assign n27877 = ~n1887 & n27876 ;
  assign n27878 = ( n1118 & n8711 ) | ( n1118 & n27877 ) | ( n8711 & n27877 ) ;
  assign n27879 = n27878 ^ n12542 ^ n10342 ;
  assign n27880 = n27879 ^ n10964 ^ 1'b0 ;
  assign n27874 = n2160 ^ n820 ^ 1'b0 ;
  assign n27875 = n12423 | n27874 ;
  assign n27881 = n27880 ^ n27875 ^ n5871 ;
  assign n27884 = x67 & ~n2388 ;
  assign n27885 = n27884 ^ n4954 ^ 1'b0 ;
  assign n27882 = ( ~n7689 & n8171 ) | ( ~n7689 & n8706 ) | ( n8171 & n8706 ) ;
  assign n27883 = n27882 ^ n6216 ^ 1'b0 ;
  assign n27886 = n27885 ^ n27883 ^ 1'b0 ;
  assign n27887 = n27881 & ~n27886 ;
  assign n27888 = n24479 ^ n3420 ^ 1'b0 ;
  assign n27889 = n17224 ^ n1607 ^ 1'b0 ;
  assign n27890 = ( n17035 & n27888 ) | ( n17035 & ~n27889 ) | ( n27888 & ~n27889 ) ;
  assign n27891 = ~n5262 & n6580 ;
  assign n27892 = n8133 | n27891 ;
  assign n27893 = n9218 & n18563 ;
  assign n27894 = n10761 & n15506 ;
  assign n27895 = n27894 ^ n26600 ^ 1'b0 ;
  assign n27896 = n27893 | n27895 ;
  assign n27897 = x254 ^ x246 ^ 1'b0 ;
  assign n27898 = n4368 & ~n26329 ;
  assign n27899 = x209 & ~n5574 ;
  assign n27900 = n17563 ^ n17145 ^ n6470 ;
  assign n27901 = n27899 | n27900 ;
  assign n27902 = n8251 & ~n27901 ;
  assign n27903 = ( n1414 & ~n17525 ) | ( n1414 & n19434 ) | ( ~n17525 & n19434 ) ;
  assign n27904 = n12061 ^ n593 ^ 1'b0 ;
  assign n27905 = ( n20209 & n27903 ) | ( n20209 & ~n27904 ) | ( n27903 & ~n27904 ) ;
  assign n27909 = ~n2788 & n5154 ;
  assign n27910 = n27909 ^ n12481 ^ 1'b0 ;
  assign n27906 = n3930 ^ n2978 ^ n2507 ;
  assign n27907 = n27906 ^ n9182 ^ 1'b0 ;
  assign n27908 = n6917 | n27907 ;
  assign n27911 = n27910 ^ n27908 ^ n20110 ;
  assign n27912 = n12167 & n19957 ;
  assign n27913 = n22065 | n27912 ;
  assign n27914 = n27913 ^ n23921 ^ 1'b0 ;
  assign n27915 = n9150 ^ n7185 ^ 1'b0 ;
  assign n27916 = n15372 | n27915 ;
  assign n27917 = ( ~n12622 & n26911 ) | ( ~n12622 & n27916 ) | ( n26911 & n27916 ) ;
  assign n27918 = n18161 ^ n7223 ^ 1'b0 ;
  assign n27919 = n22593 ^ n15662 ^ n14760 ;
  assign n27920 = n2586 & ~n23022 ;
  assign n27921 = n18354 ^ n8033 ^ x223 ;
  assign n27922 = ~n15763 & n18446 ;
  assign n27923 = ~n27921 & n27922 ;
  assign n27924 = n23518 ^ n16359 ^ 1'b0 ;
  assign n27925 = ~n2093 & n27924 ;
  assign n27926 = n19602 ^ n5470 ^ 1'b0 ;
  assign n27929 = n3863 ^ n3245 ^ 1'b0 ;
  assign n27930 = n5063 & n27929 ;
  assign n27927 = n19253 & ~n23946 ;
  assign n27928 = ~n24434 & n27927 ;
  assign n27931 = n27930 ^ n27928 ^ n26475 ;
  assign n27932 = n13894 ^ n12571 ^ n9501 ;
  assign n27933 = n19756 ^ n19379 ^ 1'b0 ;
  assign n27934 = n22214 | n27933 ;
  assign n27935 = ( ~n341 & n21515 ) | ( ~n341 & n25129 ) | ( n21515 & n25129 ) ;
  assign n27936 = ( n14890 & n19507 ) | ( n14890 & ~n27935 ) | ( n19507 & ~n27935 ) ;
  assign n27937 = n3031 ^ n1297 ^ 1'b0 ;
  assign n27938 = n12866 & ~n27937 ;
  assign n27939 = n27938 ^ n7391 ^ 1'b0 ;
  assign n27940 = n27939 ^ n2040 ^ n637 ;
  assign n27941 = ( n21968 & n27936 ) | ( n21968 & ~n27940 ) | ( n27936 & ~n27940 ) ;
  assign n27942 = n27941 ^ n17515 ^ 1'b0 ;
  assign n27943 = n21396 ^ n11500 ^ 1'b0 ;
  assign n27944 = n930 | n10220 ;
  assign n27945 = n7943 | n27944 ;
  assign n27946 = n12166 ^ n7441 ^ 1'b0 ;
  assign n27947 = n27946 ^ n23921 ^ 1'b0 ;
  assign n27948 = n27947 ^ n19313 ^ 1'b0 ;
  assign n27949 = n27948 ^ n19989 ^ n11546 ;
  assign n27950 = n21094 ^ n14095 ^ n5005 ;
  assign n27951 = n1539 & ~n21141 ;
  assign n27952 = n21141 & n27951 ;
  assign n27953 = n18356 ^ n1870 ^ 1'b0 ;
  assign n27954 = n27952 & n27953 ;
  assign n27955 = n8492 & n8775 ;
  assign n27956 = n27955 ^ n19630 ^ 1'b0 ;
  assign n27957 = n7447 ^ n5989 ^ 1'b0 ;
  assign n27958 = n22847 ^ n18388 ^ n8041 ;
  assign n27959 = n2108 & n5286 ;
  assign n27960 = n27959 ^ n21403 ^ 1'b0 ;
  assign n27961 = n1098 | n12230 ;
  assign n27962 = n21083 & ~n27961 ;
  assign n27963 = n27962 ^ n26088 ^ 1'b0 ;
  assign n27964 = n13788 & ~n27963 ;
  assign n27973 = ( ~n5795 & n7068 ) | ( ~n5795 & n19253 ) | ( n7068 & n19253 ) ;
  assign n27965 = ( n1948 & n3182 ) | ( n1948 & n25313 ) | ( n3182 & n25313 ) ;
  assign n27966 = n27965 ^ n4394 ^ 1'b0 ;
  assign n27967 = ~n6220 & n27966 ;
  assign n27968 = n19193 ^ n13888 ^ n12605 ;
  assign n27969 = n27968 ^ n12549 ^ n7050 ;
  assign n27970 = n27969 ^ n325 ^ 1'b0 ;
  assign n27971 = n27967 & n27970 ;
  assign n27972 = ~n331 & n27971 ;
  assign n27974 = n27973 ^ n27972 ^ 1'b0 ;
  assign n27975 = n22485 | n27974 ;
  assign n27976 = n23164 ^ n9569 ^ n7626 ;
  assign n27977 = n7358 | n16241 ;
  assign n27978 = n24792 ^ n14427 ^ 1'b0 ;
  assign n27979 = ~n4708 & n27978 ;
  assign n27980 = ~n24064 & n27979 ;
  assign n27981 = n5261 | n17068 ;
  assign n27982 = n27981 ^ n6732 ^ 1'b0 ;
  assign n27983 = n25821 & n27982 ;
  assign n27984 = n27983 ^ n3966 ^ 1'b0 ;
  assign n27985 = n17723 ^ n7356 ^ 1'b0 ;
  assign n27986 = n27984 & ~n27985 ;
  assign n27987 = n27986 ^ n13342 ^ 1'b0 ;
  assign n27988 = n4844 | n27987 ;
  assign n27989 = n27988 ^ n404 ^ 1'b0 ;
  assign n27990 = n14462 | n14892 ;
  assign n27991 = n27990 ^ n3499 ^ 1'b0 ;
  assign n27992 = n27989 & n27991 ;
  assign n27993 = ( n6796 & n17064 ) | ( n6796 & n21876 ) | ( n17064 & n21876 ) ;
  assign n27994 = ( n6453 & n12775 ) | ( n6453 & ~n27993 ) | ( n12775 & ~n27993 ) ;
  assign n27995 = n21198 ^ n16531 ^ n3872 ;
  assign n27996 = n8946 ^ n8433 ^ n1040 ;
  assign n27997 = n27996 ^ n23406 ^ 1'b0 ;
  assign n27998 = n27995 & ~n27997 ;
  assign n27999 = n27998 ^ n8187 ^ 1'b0 ;
  assign n28000 = ~n18451 & n27999 ;
  assign n28001 = ~n16922 & n19914 ;
  assign n28002 = n17095 ^ n15360 ^ n11753 ;
  assign n28003 = n15829 ^ n10466 ^ n1826 ;
  assign n28005 = n6041 | n26916 ;
  assign n28004 = ~n11157 & n13850 ;
  assign n28006 = n28005 ^ n28004 ^ 1'b0 ;
  assign n28007 = ( n14476 & ~n28003 ) | ( n14476 & n28006 ) | ( ~n28003 & n28006 ) ;
  assign n28008 = ( n3953 & n18498 ) | ( n3953 & n28007 ) | ( n18498 & n28007 ) ;
  assign n28010 = n9394 ^ x94 ^ 1'b0 ;
  assign n28009 = n11619 ^ n9146 ^ 1'b0 ;
  assign n28011 = n28010 ^ n28009 ^ n18373 ;
  assign n28012 = n27651 ^ n2100 ^ 1'b0 ;
  assign n28013 = n28011 & n28012 ;
  assign n28014 = ( n2864 & n9232 ) | ( n2864 & ~n26145 ) | ( n9232 & ~n26145 ) ;
  assign n28015 = n28014 ^ n23817 ^ 1'b0 ;
  assign n28016 = ~n20351 & n28015 ;
  assign n28017 = n28016 ^ n22631 ^ 1'b0 ;
  assign n28018 = ~n20625 & n28017 ;
  assign n28019 = ( n3246 & n4499 ) | ( n3246 & ~n13423 ) | ( n4499 & ~n13423 ) ;
  assign n28020 = n15153 ^ n14192 ^ n6733 ;
  assign n28021 = n18845 ^ n14155 ^ 1'b0 ;
  assign n28022 = ( n3016 & ~n5741 ) | ( n3016 & n5823 ) | ( ~n5741 & n5823 ) ;
  assign n28023 = n18223 ^ n17441 ^ 1'b0 ;
  assign n28024 = n28022 | n28023 ;
  assign n28025 = n19759 ^ n4075 ^ 1'b0 ;
  assign n28026 = ~n4583 & n28025 ;
  assign n28027 = n22846 ^ n3283 ^ 1'b0 ;
  assign n28028 = n24663 & n28027 ;
  assign n28029 = n7859 & n28028 ;
  assign n28030 = ( n21234 & n28026 ) | ( n21234 & n28029 ) | ( n28026 & n28029 ) ;
  assign n28031 = ( ~n17867 & n28024 ) | ( ~n17867 & n28030 ) | ( n28024 & n28030 ) ;
  assign n28032 = n25773 ^ n22987 ^ n10267 ;
  assign n28033 = n21934 ^ n11447 ^ 1'b0 ;
  assign n28034 = n413 & ~n1446 ;
  assign n28035 = n7981 | n28034 ;
  assign n28036 = n28035 ^ n3781 ^ 1'b0 ;
  assign n28037 = ( n1511 & n11302 ) | ( n1511 & n28036 ) | ( n11302 & n28036 ) ;
  assign n28038 = ~n16355 & n24917 ;
  assign n28039 = n28037 & n28038 ;
  assign n28040 = ~n4788 & n9232 ;
  assign n28041 = n28040 ^ n6495 ^ 1'b0 ;
  assign n28042 = n28041 ^ n16357 ^ 1'b0 ;
  assign n28043 = n28042 ^ n16540 ^ 1'b0 ;
  assign n28044 = n11631 ^ n7360 ^ n4180 ;
  assign n28045 = n28044 ^ n27496 ^ n9111 ;
  assign n28046 = ( n3026 & n6216 ) | ( n3026 & n7611 ) | ( n6216 & n7611 ) ;
  assign n28048 = ( n4790 & ~n11862 ) | ( n4790 & n14059 ) | ( ~n11862 & n14059 ) ;
  assign n28047 = n23040 & n26955 ;
  assign n28049 = n28048 ^ n28047 ^ 1'b0 ;
  assign n28050 = n6611 & n8724 ;
  assign n28051 = n28050 ^ n7220 ^ 1'b0 ;
  assign n28052 = n18888 ^ n10151 ^ 1'b0 ;
  assign n28053 = ~n5753 & n28052 ;
  assign n28054 = n2335 | n5264 ;
  assign n28055 = n28053 | n28054 ;
  assign n28056 = n17507 & n28055 ;
  assign n28057 = ~n17783 & n28056 ;
  assign n28058 = n2839 & n15680 ;
  assign n28059 = ~n28057 & n28058 ;
  assign n28060 = x147 & n15456 ;
  assign n28061 = n15757 & n28060 ;
  assign n28062 = ~n6037 & n28061 ;
  assign n28063 = n8652 & ~n13871 ;
  assign n28064 = ~n9191 & n28063 ;
  assign n28065 = n3463 & ~n6985 ;
  assign n28066 = n28065 ^ n22394 ^ n10648 ;
  assign n28067 = n28066 ^ n5346 ^ 1'b0 ;
  assign n28068 = n586 | n28067 ;
  assign n28069 = n28068 ^ n10172 ^ 1'b0 ;
  assign n28070 = n20209 ^ n17130 ^ n1054 ;
  assign n28071 = n21030 ^ n11332 ^ 1'b0 ;
  assign n28072 = ~n8366 & n25323 ;
  assign n28073 = n21716 & n28072 ;
  assign n28074 = ( n4148 & ~n10634 ) | ( n4148 & n23460 ) | ( ~n10634 & n23460 ) ;
  assign n28075 = n28074 ^ n24237 ^ 1'b0 ;
  assign n28076 = ( n1983 & ~n4190 ) | ( n1983 & n11515 ) | ( ~n4190 & n11515 ) ;
  assign n28077 = n15654 ^ n2205 ^ 1'b0 ;
  assign n28078 = n9078 & n26305 ;
  assign n28081 = n5553 & ~n7926 ;
  assign n28079 = n13755 ^ n2811 ^ 1'b0 ;
  assign n28080 = n13317 & n28079 ;
  assign n28082 = n28081 ^ n28080 ^ 1'b0 ;
  assign n28083 = n13812 | n28082 ;
  assign n28084 = n14606 | n28083 ;
  assign n28085 = n10278 | n21678 ;
  assign n28089 = n1418 & ~n10173 ;
  assign n28086 = ~n2903 & n8730 ;
  assign n28087 = n4260 & n28086 ;
  assign n28088 = n7873 | n28087 ;
  assign n28090 = n28089 ^ n28088 ^ 1'b0 ;
  assign n28091 = n9578 | n28090 ;
  assign n28092 = n8908 | n28091 ;
  assign n28093 = ( n4851 & n8008 ) | ( n4851 & ~n28092 ) | ( n8008 & ~n28092 ) ;
  assign n28094 = n7064 ^ n5838 ^ 1'b0 ;
  assign n28095 = ~n22305 & n28094 ;
  assign n28096 = n28095 ^ n22094 ^ 1'b0 ;
  assign n28098 = n7916 & n9149 ;
  assign n28097 = n6071 & ~n14821 ;
  assign n28099 = n28098 ^ n28097 ^ 1'b0 ;
  assign n28100 = ~n9664 & n28099 ;
  assign n28101 = n11903 ^ n7046 ^ 1'b0 ;
  assign n28102 = ~n4287 & n28101 ;
  assign n28103 = ~n17618 & n21980 ;
  assign n28104 = n28103 ^ n18085 ^ n16865 ;
  assign n28105 = ( n3484 & ~n11478 ) | ( n3484 & n28104 ) | ( ~n11478 & n28104 ) ;
  assign n28107 = n20533 ^ n4544 ^ n374 ;
  assign n28108 = n2504 & n28107 ;
  assign n28109 = n8337 ^ n4087 ^ n2218 ;
  assign n28110 = n28108 & n28109 ;
  assign n28111 = n10014 & n28110 ;
  assign n28106 = n15871 ^ n6722 ^ n1879 ;
  assign n28112 = n28111 ^ n28106 ^ n25028 ;
  assign n28113 = n19461 ^ n10595 ^ n1836 ;
  assign n28114 = n28113 ^ n4590 ^ n1652 ;
  assign n28115 = n22725 ^ n7223 ^ n4209 ;
  assign n28116 = n397 & ~n28115 ;
  assign n28117 = n9899 & n28116 ;
  assign n28118 = n2918 ^ n1484 ^ 1'b0 ;
  assign n28119 = n23134 & ~n28118 ;
  assign n28120 = n28113 & n28119 ;
  assign n28121 = ~n9127 & n25494 ;
  assign n28122 = n1617 & n28121 ;
  assign n28123 = n7481 & ~n21231 ;
  assign n28124 = n23452 & n28123 ;
  assign n28125 = ( n4554 & ~n15599 ) | ( n4554 & n15764 ) | ( ~n15599 & n15764 ) ;
  assign n28128 = n10216 ^ n9258 ^ 1'b0 ;
  assign n28129 = n872 & n28128 ;
  assign n28126 = n6379 ^ n1659 ^ 1'b0 ;
  assign n28127 = ~n26907 & n28126 ;
  assign n28130 = n28129 ^ n28127 ^ 1'b0 ;
  assign n28131 = ( n4734 & n8008 ) | ( n4734 & ~n24408 ) | ( n8008 & ~n24408 ) ;
  assign n28132 = ~n12753 & n23457 ;
  assign n28133 = n24255 ^ n22991 ^ n8011 ;
  assign n28134 = ( ~n28131 & n28132 ) | ( ~n28131 & n28133 ) | ( n28132 & n28133 ) ;
  assign n28135 = n6295 ^ n1903 ^ 1'b0 ;
  assign n28136 = n2232 | n28135 ;
  assign n28137 = ( ~n9588 & n23255 ) | ( ~n9588 & n28136 ) | ( n23255 & n28136 ) ;
  assign n28138 = ( n2731 & n11414 ) | ( n2731 & n20164 ) | ( n11414 & n20164 ) ;
  assign n28139 = n28138 ^ n15839 ^ n13953 ;
  assign n28140 = n17004 & ~n28120 ;
  assign n28141 = n1695 & n28140 ;
  assign n28142 = x69 | n14173 ;
  assign n28143 = n28142 ^ n20511 ^ 1'b0 ;
  assign n28144 = ~n16183 & n28143 ;
  assign n28145 = n28144 ^ n24451 ^ 1'b0 ;
  assign n28146 = n24706 ^ n24500 ^ 1'b0 ;
  assign n28147 = n2205 | n28146 ;
  assign n28148 = n20283 ^ n12304 ^ 1'b0 ;
  assign n28149 = ( n8331 & n17976 ) | ( n8331 & ~n28148 ) | ( n17976 & ~n28148 ) ;
  assign n28152 = n20139 ^ n3995 ^ n1524 ;
  assign n28150 = ( ~n1380 & n14870 ) | ( ~n1380 & n27140 ) | ( n14870 & n27140 ) ;
  assign n28151 = n28150 ^ n12329 ^ 1'b0 ;
  assign n28153 = n28152 ^ n28151 ^ 1'b0 ;
  assign n28154 = n22970 & ~n28153 ;
  assign n28155 = n261 & ~n13270 ;
  assign n28156 = n14894 & n28155 ;
  assign n28157 = n28156 ^ n18098 ^ n7212 ;
  assign n28158 = ( ~n10036 & n11796 ) | ( ~n10036 & n24162 ) | ( n11796 & n24162 ) ;
  assign n28159 = ( n1735 & n7670 ) | ( n1735 & ~n17908 ) | ( n7670 & ~n17908 ) ;
  assign n28160 = n28158 & n28159 ;
  assign n28172 = n1283 | n5380 ;
  assign n28173 = n4298 | n28172 ;
  assign n28170 = n21642 ^ n8299 ^ 1'b0 ;
  assign n28171 = ( n1629 & n12692 ) | ( n1629 & ~n28170 ) | ( n12692 & ~n28170 ) ;
  assign n28161 = n2994 & n8537 ;
  assign n28162 = n28161 ^ n16806 ^ n11492 ;
  assign n28164 = n14721 ^ n6560 ^ n4104 ;
  assign n28163 = n21097 & n22449 ;
  assign n28165 = n28164 ^ n28163 ^ 1'b0 ;
  assign n28166 = ~n1057 & n3737 ;
  assign n28167 = ( n2514 & n8172 ) | ( n2514 & ~n16228 ) | ( n8172 & ~n16228 ) ;
  assign n28168 = ( n7232 & ~n28166 ) | ( n7232 & n28167 ) | ( ~n28166 & n28167 ) ;
  assign n28169 = ( n28162 & ~n28165 ) | ( n28162 & n28168 ) | ( ~n28165 & n28168 ) ;
  assign n28174 = n28173 ^ n28171 ^ n28169 ;
  assign n28175 = n18040 ^ n6640 ^ n3880 ;
  assign n28176 = n28175 ^ n7361 ^ 1'b0 ;
  assign n28177 = ( n19414 & ~n19857 ) | ( n19414 & n28176 ) | ( ~n19857 & n28176 ) ;
  assign n28178 = n8940 | n14807 ;
  assign n28179 = n28177 & ~n28178 ;
  assign n28187 = n23477 ^ n10277 ^ n8233 ;
  assign n28188 = n10225 | n28187 ;
  assign n28180 = ~n7236 & n12527 ;
  assign n28181 = ~n5286 & n28180 ;
  assign n28182 = n7542 & ~n16409 ;
  assign n28183 = n1945 | n6612 ;
  assign n28184 = n28183 ^ n23618 ^ 1'b0 ;
  assign n28185 = n28182 & ~n28184 ;
  assign n28186 = n28181 & n28185 ;
  assign n28189 = n28188 ^ n28186 ^ n7500 ;
  assign n28190 = ~n28179 & n28189 ;
  assign n28191 = n6625 & ~n7401 ;
  assign n28192 = n28191 ^ n5693 ^ n5201 ;
  assign n28193 = n27956 | n28192 ;
  assign n28194 = n17678 | n28193 ;
  assign n28195 = ~n11863 & n12649 ;
  assign n28200 = n12492 ^ n8373 ^ n5458 ;
  assign n28196 = ( n8357 & n14136 ) | ( n8357 & ~n16199 ) | ( n14136 & ~n16199 ) ;
  assign n28197 = n6395 & n28196 ;
  assign n28198 = n28197 ^ n10774 ^ 1'b0 ;
  assign n28199 = n28198 ^ n1963 ^ 1'b0 ;
  assign n28201 = n28200 ^ n28199 ^ 1'b0 ;
  assign n28202 = n3994 & n16662 ;
  assign n28203 = ~n13163 & n28202 ;
  assign n28204 = n24417 & ~n28203 ;
  assign n28205 = ~n8133 & n16665 ;
  assign n28206 = n1791 & n28205 ;
  assign n28207 = n28206 ^ n9790 ^ 1'b0 ;
  assign n28208 = ( n28201 & n28204 ) | ( n28201 & n28207 ) | ( n28204 & n28207 ) ;
  assign n28209 = x230 & ~n16838 ;
  assign n28210 = n14328 & n28209 ;
  assign n28211 = ( ~n12906 & n17494 ) | ( ~n12906 & n28210 ) | ( n17494 & n28210 ) ;
  assign n28212 = ( n3209 & ~n11676 ) | ( n3209 & n14494 ) | ( ~n11676 & n14494 ) ;
  assign n28213 = n4179 & ~n28212 ;
  assign n28214 = n14584 & n21973 ;
  assign n28215 = n17302 & n28214 ;
  assign n28216 = n12631 & n15279 ;
  assign n28217 = n15270 ^ n9700 ^ n3157 ;
  assign n28221 = ~n2771 & n14992 ;
  assign n28222 = n28221 ^ n3909 ^ 1'b0 ;
  assign n28218 = n5935 | n21420 ;
  assign n28219 = n14283 ^ n7744 ^ 1'b0 ;
  assign n28220 = ~n28218 & n28219 ;
  assign n28223 = n28222 ^ n28220 ^ n20777 ;
  assign n28224 = n12536 ^ n769 ^ 1'b0 ;
  assign n28225 = n3001 | n28224 ;
  assign n28226 = n28225 ^ n26775 ^ 1'b0 ;
  assign n28227 = ~n28223 & n28226 ;
  assign n28228 = n3195 & ~n18459 ;
  assign n28229 = n28228 ^ n10290 ^ 1'b0 ;
  assign n28230 = n27430 | n28229 ;
  assign n28231 = n2062 | n28230 ;
  assign n28232 = n8461 & ~n28231 ;
  assign n28233 = n7742 ^ n3901 ^ 1'b0 ;
  assign n28234 = n8209 & ~n11445 ;
  assign n28235 = n4530 & ~n6124 ;
  assign n28236 = n28235 ^ n11958 ^ 1'b0 ;
  assign n28237 = n6488 & ~n9642 ;
  assign n28238 = ~n7741 & n28237 ;
  assign n28239 = n28238 ^ n459 ^ 1'b0 ;
  assign n28240 = n28236 & ~n28239 ;
  assign n28241 = ~n15835 & n28240 ;
  assign n28242 = n10284 & ~n16268 ;
  assign n28243 = n28242 ^ n918 ^ 1'b0 ;
  assign n28244 = n4783 | n5324 ;
  assign n28245 = n25165 ^ n15344 ^ 1'b0 ;
  assign n28246 = n21536 | n28245 ;
  assign n28247 = ( n7108 & n9116 ) | ( n7108 & n21629 ) | ( n9116 & n21629 ) ;
  assign n28248 = n28246 | n28247 ;
  assign n28249 = ( n28243 & n28244 ) | ( n28243 & ~n28248 ) | ( n28244 & ~n28248 ) ;
  assign n28250 = x14 & ~n7627 ;
  assign n28251 = n22702 & ~n28250 ;
  assign n28252 = ~n13297 & n28251 ;
  assign n28253 = n28252 ^ n6690 ^ n640 ;
  assign n28255 = ( ~n1753 & n14902 ) | ( ~n1753 & n15230 ) | ( n14902 & n15230 ) ;
  assign n28256 = n28255 ^ n15625 ^ n8697 ;
  assign n28254 = n11560 & n23130 ;
  assign n28257 = n28256 ^ n28254 ^ 1'b0 ;
  assign n28258 = n1422 | n2800 ;
  assign n28259 = n26609 & ~n28258 ;
  assign n28260 = n9470 ^ n2721 ^ 1'b0 ;
  assign n28261 = n21741 | n28260 ;
  assign n28262 = n21905 | n28261 ;
  assign n28263 = n3182 | n28262 ;
  assign n28264 = n28263 ^ n11457 ^ n1057 ;
  assign n28265 = n12845 ^ n9524 ^ n6199 ;
  assign n28266 = ( n20830 & n23465 ) | ( n20830 & ~n28265 ) | ( n23465 & ~n28265 ) ;
  assign n28267 = n9637 | n15351 ;
  assign n28268 = n6672 & n12474 ;
  assign n28269 = n28268 ^ n4890 ^ 1'b0 ;
  assign n28270 = n11451 ^ n6460 ^ 1'b0 ;
  assign n28271 = n16759 ^ n2512 ^ n1545 ;
  assign n28272 = n28270 | n28271 ;
  assign n28273 = n12533 & ~n23376 ;
  assign n28274 = n28273 ^ n4779 ^ 1'b0 ;
  assign n28275 = n28274 ^ n27729 ^ 1'b0 ;
  assign n28276 = n28275 ^ n20807 ^ 1'b0 ;
  assign n28278 = n1541 | n10243 ;
  assign n28279 = n3614 | n28278 ;
  assign n28280 = ~n27079 & n28279 ;
  assign n28277 = ( ~n4749 & n13382 ) | ( ~n4749 & n20742 ) | ( n13382 & n20742 ) ;
  assign n28281 = n28280 ^ n28277 ^ n9286 ;
  assign n28282 = ( x80 & x122 ) | ( x80 & ~n7391 ) | ( x122 & ~n7391 ) ;
  assign n28283 = n4727 & ~n12222 ;
  assign n28284 = n1087 & n28283 ;
  assign n28285 = n28284 ^ n26323 ^ n6341 ;
  assign n28286 = n782 & n5697 ;
  assign n28287 = ( n11623 & n16115 ) | ( n11623 & n28286 ) | ( n16115 & n28286 ) ;
  assign n28288 = n28287 ^ n18671 ^ 1'b0 ;
  assign n28289 = n16181 & ~n26720 ;
  assign n28290 = ~n17071 & n28289 ;
  assign n28291 = n9767 & n19226 ;
  assign n28292 = n9239 & n28291 ;
  assign n28293 = ( n5408 & n12988 ) | ( n5408 & n13693 ) | ( n12988 & n13693 ) ;
  assign n28294 = ( n1298 & n2760 ) | ( n1298 & n7238 ) | ( n2760 & n7238 ) ;
  assign n28295 = ~n4711 & n8253 ;
  assign n28296 = ( ~n5326 & n11251 ) | ( ~n5326 & n28295 ) | ( n11251 & n28295 ) ;
  assign n28297 = ( n7122 & n10400 ) | ( n7122 & ~n14573 ) | ( n10400 & ~n14573 ) ;
  assign n28298 = ( n12013 & ~n28296 ) | ( n12013 & n28297 ) | ( ~n28296 & n28297 ) ;
  assign n28299 = n22926 ^ n4652 ^ n1586 ;
  assign n28300 = n28299 ^ n12430 ^ x86 ;
  assign n28301 = n26680 ^ n18229 ^ 1'b0 ;
  assign n28302 = n28301 ^ n23563 ^ 1'b0 ;
  assign n28303 = n24725 ^ n7884 ^ 1'b0 ;
  assign n28304 = n8515 & n28303 ;
  assign n28305 = n12550 ^ n8483 ^ n5341 ;
  assign n28306 = ~n11124 & n28305 ;
  assign n28307 = n28306 ^ n15285 ^ 1'b0 ;
  assign n28308 = ~n28304 & n28307 ;
  assign n28309 = ( x237 & n6365 ) | ( x237 & ~n6725 ) | ( n6365 & ~n6725 ) ;
  assign n28310 = n13743 ^ n12806 ^ 1'b0 ;
  assign n28311 = n18750 | n28310 ;
  assign n28312 = n4304 | n28311 ;
  assign n28313 = n7904 & n11766 ;
  assign n28314 = n28313 ^ n14815 ^ n842 ;
  assign n28315 = n3675 ^ n3251 ^ n3118 ;
  assign n28316 = n28315 ^ n13623 ^ 1'b0 ;
  assign n28318 = ~n14266 & n17463 ;
  assign n28317 = x33 & n19377 ;
  assign n28319 = n28318 ^ n28317 ^ 1'b0 ;
  assign n28320 = n16128 & n19256 ;
  assign n28321 = n15067 ^ n7980 ^ 1'b0 ;
  assign n28322 = ~n28320 & n28321 ;
  assign n28323 = ~n702 & n1909 ;
  assign n28324 = n11213 & ~n20721 ;
  assign n28325 = n28324 ^ n4346 ^ 1'b0 ;
  assign n28326 = n28323 & n28325 ;
  assign n28327 = ( n1629 & n8156 ) | ( n1629 & n21251 ) | ( n8156 & n21251 ) ;
  assign n28328 = n28327 ^ n10308 ^ n9931 ;
  assign n28333 = n2520 & n5408 ;
  assign n28334 = n10735 & n28333 ;
  assign n28329 = n5924 ^ n2501 ^ 1'b0 ;
  assign n28330 = n10577 & n28329 ;
  assign n28331 = ( n9742 & ~n11853 ) | ( n9742 & n28330 ) | ( ~n11853 & n28330 ) ;
  assign n28332 = ~n18887 & n28331 ;
  assign n28335 = n28334 ^ n28332 ^ 1'b0 ;
  assign n28336 = n19195 & ~n28335 ;
  assign n28337 = ( n6778 & ~n11591 ) | ( n6778 & n13486 ) | ( ~n11591 & n13486 ) ;
  assign n28338 = n26954 ^ n5384 ^ 1'b0 ;
  assign n28339 = n7216 & ~n28338 ;
  assign n28340 = ~n16791 & n28339 ;
  assign n28341 = ( n27093 & n28337 ) | ( n27093 & n28340 ) | ( n28337 & n28340 ) ;
  assign n28342 = n1178 | n28341 ;
  assign n28343 = n28341 & ~n28342 ;
  assign n28344 = n27478 ^ n22246 ^ 1'b0 ;
  assign n28345 = ( n9699 & ~n17614 ) | ( n9699 & n28344 ) | ( ~n17614 & n28344 ) ;
  assign n28346 = ( n7126 & ~n28343 ) | ( n7126 & n28345 ) | ( ~n28343 & n28345 ) ;
  assign n28347 = ( n9357 & n17060 ) | ( n9357 & ~n23335 ) | ( n17060 & ~n23335 ) ;
  assign n28348 = n3717 & ~n28347 ;
  assign n28349 = n28348 ^ n5144 ^ 1'b0 ;
  assign n28350 = ( n14896 & n18414 ) | ( n14896 & ~n24233 ) | ( n18414 & ~n24233 ) ;
  assign n28351 = n20554 ^ n8234 ^ 1'b0 ;
  assign n28352 = n23845 | n28351 ;
  assign n28353 = ~n28350 & n28352 ;
  assign n28354 = n11998 ^ n4004 ^ 1'b0 ;
  assign n28355 = n24120 & ~n28354 ;
  assign n28356 = ~n19485 & n28355 ;
  assign n28357 = ~n5795 & n28356 ;
  assign n28358 = ( n6911 & ~n20582 ) | ( n6911 & n23812 ) | ( ~n20582 & n23812 ) ;
  assign n28359 = ( n14848 & n17851 ) | ( n14848 & ~n28358 ) | ( n17851 & ~n28358 ) ;
  assign n28360 = n14848 ^ n7158 ^ 1'b0 ;
  assign n28361 = n2847 | n28360 ;
  assign n28362 = n10409 ^ n6673 ^ 1'b0 ;
  assign n28363 = ~n28361 & n28362 ;
  assign n28364 = ~n455 & n28363 ;
  assign n28365 = ~n4008 & n28364 ;
  assign n28366 = n2595 & n28365 ;
  assign n28367 = n28366 ^ n9273 ^ 1'b0 ;
  assign n28368 = ~n3760 & n16894 ;
  assign n28369 = n28368 ^ n22595 ^ 1'b0 ;
  assign n28370 = n12881 ^ n11257 ^ 1'b0 ;
  assign n28376 = n14029 ^ n4369 ^ n3042 ;
  assign n28371 = n22068 ^ n17976 ^ 1'b0 ;
  assign n28372 = n7705 | n20007 ;
  assign n28373 = n9608 & ~n28372 ;
  assign n28374 = n2714 | n28373 ;
  assign n28375 = n28371 & ~n28374 ;
  assign n28377 = n28376 ^ n28375 ^ x159 ;
  assign n28378 = ~n3817 & n6184 ;
  assign n28379 = n3946 | n4101 ;
  assign n28380 = n28379 ^ n1766 ^ 1'b0 ;
  assign n28381 = n28378 | n28380 ;
  assign n28382 = n28381 ^ n2412 ^ 1'b0 ;
  assign n28383 = ( n7395 & n18651 ) | ( n7395 & n28382 ) | ( n18651 & n28382 ) ;
  assign n28384 = ( n10230 & n16686 ) | ( n10230 & ~n28383 ) | ( n16686 & ~n28383 ) ;
  assign n28385 = ( ~n10623 & n28377 ) | ( ~n10623 & n28384 ) | ( n28377 & n28384 ) ;
  assign n28386 = n5436 & n15659 ;
  assign n28387 = ~n5251 & n28386 ;
  assign n28388 = n16989 ^ n6252 ^ 1'b0 ;
  assign n28389 = ( n23817 & n28387 ) | ( n23817 & n28388 ) | ( n28387 & n28388 ) ;
  assign n28390 = n23472 ^ n12814 ^ n11181 ;
  assign n28391 = ( n1438 & n4328 ) | ( n1438 & ~n4423 ) | ( n4328 & ~n4423 ) ;
  assign n28392 = ( n8756 & n16479 ) | ( n8756 & n28391 ) | ( n16479 & n28391 ) ;
  assign n28393 = n21827 & n28392 ;
  assign n28396 = n4301 | n20046 ;
  assign n28397 = n12914 | n28396 ;
  assign n28394 = n7370 ^ n3754 ^ 1'b0 ;
  assign n28395 = ( n12033 & ~n15564 ) | ( n12033 & n28394 ) | ( ~n15564 & n28394 ) ;
  assign n28398 = n28397 ^ n28395 ^ 1'b0 ;
  assign n28399 = ( n1868 & n9919 ) | ( n1868 & n22517 ) | ( n9919 & n22517 ) ;
  assign n28400 = n11965 | n23081 ;
  assign n28401 = n13923 | n28400 ;
  assign n28402 = ( n963 & n17232 ) | ( n963 & n28401 ) | ( n17232 & n28401 ) ;
  assign n28403 = n16028 ^ n1868 ^ n1049 ;
  assign n28404 = ( n3149 & n19723 ) | ( n3149 & ~n28403 ) | ( n19723 & ~n28403 ) ;
  assign n28405 = n1475 & n23864 ;
  assign n28406 = ~n11518 & n28405 ;
  assign n28408 = ( n1352 & n6502 ) | ( n1352 & n7602 ) | ( n6502 & n7602 ) ;
  assign n28407 = ( n5663 & ~n7156 ) | ( n5663 & n7300 ) | ( ~n7156 & n7300 ) ;
  assign n28409 = n28408 ^ n28407 ^ n1933 ;
  assign n28410 = ( n22844 & ~n24099 ) | ( n22844 & n26951 ) | ( ~n24099 & n26951 ) ;
  assign n28411 = n8437 ^ n5251 ^ 1'b0 ;
  assign n28412 = ( n3637 & n9675 ) | ( n3637 & n28411 ) | ( n9675 & n28411 ) ;
  assign n28413 = n22802 ^ n21209 ^ 1'b0 ;
  assign n28414 = n8374 & n28413 ;
  assign n28415 = n28414 ^ n3874 ^ 1'b0 ;
  assign n28416 = n10418 ^ n9632 ^ n9498 ;
  assign n28417 = ( n8795 & n21219 ) | ( n8795 & ~n28416 ) | ( n21219 & ~n28416 ) ;
  assign n28418 = ( ~n6872 & n28415 ) | ( ~n6872 & n28417 ) | ( n28415 & n28417 ) ;
  assign n28419 = n1695 | n23054 ;
  assign n28420 = n28419 ^ n3356 ^ 1'b0 ;
  assign n28421 = n28420 ^ n6986 ^ 1'b0 ;
  assign n28422 = n26623 ^ n22387 ^ 1'b0 ;
  assign n28423 = n28421 & ~n28422 ;
  assign n28424 = n6030 & n18463 ;
  assign n28425 = n22121 ^ n1468 ^ n814 ;
  assign n28426 = n19171 ^ n18926 ^ n5910 ;
  assign n28427 = n332 & ~n1356 ;
  assign n28428 = n1356 & n28427 ;
  assign n28429 = n804 & n2160 ;
  assign n28430 = ~n2160 & n28429 ;
  assign n28431 = n12573 & ~n28430 ;
  assign n28432 = n28428 & n28431 ;
  assign n28433 = n28432 ^ n21371 ^ 1'b0 ;
  assign n28434 = n20038 & n28433 ;
  assign n28435 = n2937 ^ n1370 ^ 1'b0 ;
  assign n28436 = n22043 & ~n28435 ;
  assign n28442 = n9984 ^ n9742 ^ 1'b0 ;
  assign n28443 = n11150 | n28442 ;
  assign n28437 = ( n763 & n2849 ) | ( n763 & n14116 ) | ( n2849 & n14116 ) ;
  assign n28438 = ~n11853 & n28437 ;
  assign n28439 = n28438 ^ n21776 ^ 1'b0 ;
  assign n28440 = ( n5737 & ~n9188 ) | ( n5737 & n22360 ) | ( ~n9188 & n22360 ) ;
  assign n28441 = n28439 & n28440 ;
  assign n28444 = n28443 ^ n28441 ^ 1'b0 ;
  assign n28445 = n10211 | n28444 ;
  assign n28446 = n2997 & ~n18981 ;
  assign n28447 = n23084 | n28446 ;
  assign n28448 = n20517 & n28447 ;
  assign n28449 = n3801 & n28448 ;
  assign n28450 = n3442 | n5704 ;
  assign n28451 = n7559 & ~n28450 ;
  assign n28452 = n537 | n4581 ;
  assign n28453 = n28452 ^ x154 ^ 1'b0 ;
  assign n28454 = n28451 & ~n28453 ;
  assign n28455 = n26332 ^ n20141 ^ 1'b0 ;
  assign n28456 = ~n689 & n11113 ;
  assign n28457 = ~n21322 & n28456 ;
  assign n28458 = n4644 | n28457 ;
  assign n28459 = n28458 ^ n4516 ^ 1'b0 ;
  assign n28461 = n23978 ^ n15859 ^ n3484 ;
  assign n28460 = n9249 & ~n21611 ;
  assign n28462 = n28461 ^ n28460 ^ 1'b0 ;
  assign n28463 = n5289 | n9082 ;
  assign n28464 = n16100 | n28463 ;
  assign n28465 = n28464 ^ n14722 ^ n3840 ;
  assign n28466 = n12631 ^ n2450 ^ 1'b0 ;
  assign n28467 = ~n27116 & n28466 ;
  assign n28468 = n14798 & n28467 ;
  assign n28469 = n28468 ^ n16385 ^ 1'b0 ;
  assign n28470 = n14277 & n23180 ;
  assign n28471 = ~n28469 & n28470 ;
  assign n28473 = ~n13160 & n22925 ;
  assign n28474 = ( n2016 & n15938 ) | ( n2016 & n28473 ) | ( n15938 & n28473 ) ;
  assign n28472 = ~n7313 & n9052 ;
  assign n28475 = n28474 ^ n28472 ^ 1'b0 ;
  assign n28476 = ~n3254 & n28247 ;
  assign n28477 = ~n22397 & n28476 ;
  assign n28478 = n5795 & n23988 ;
  assign n28479 = n28478 ^ n9160 ^ n6683 ;
  assign n28480 = ( ~n10702 & n10858 ) | ( ~n10702 & n28479 ) | ( n10858 & n28479 ) ;
  assign n28481 = n28188 ^ n4995 ^ 1'b0 ;
  assign n28482 = n27611 ^ n8947 ^ 1'b0 ;
  assign n28483 = ~n28481 & n28482 ;
  assign n28484 = n8218 | n12852 ;
  assign n28485 = n2191 & n27071 ;
  assign n28486 = n28485 ^ n21077 ^ 1'b0 ;
  assign n28487 = n25002 ^ n2616 ^ 1'b0 ;
  assign n28488 = n28486 & ~n28487 ;
  assign n28489 = ~x66 & n28488 ;
  assign n28490 = ~n21892 & n28489 ;
  assign n28491 = n5442 & ~n17976 ;
  assign n28492 = n3903 & n28491 ;
  assign n28493 = ( ~n8377 & n8607 ) | ( ~n8377 & n28492 ) | ( n8607 & n28492 ) ;
  assign n28494 = n28493 ^ n2425 ^ 1'b0 ;
  assign n28495 = n18252 | n28494 ;
  assign n28496 = n28495 ^ n20170 ^ 1'b0 ;
  assign n28497 = n25662 ^ n23970 ^ n6895 ;
  assign n28498 = n10240 ^ n9951 ^ n7416 ;
  assign n28499 = n17901 ^ n17171 ^ n2093 ;
  assign n28500 = n28499 ^ n8307 ^ 1'b0 ;
  assign n28501 = n28500 ^ n3437 ^ 1'b0 ;
  assign n28502 = n22129 | n24986 ;
  assign n28503 = n28502 ^ n28162 ^ 1'b0 ;
  assign n28504 = n26079 ^ n16904 ^ 1'b0 ;
  assign n28505 = n14733 & n28504 ;
  assign n28506 = n28505 ^ n19061 ^ 1'b0 ;
  assign n28510 = n11122 ^ n1510 ^ 1'b0 ;
  assign n28511 = ~n7879 & n28510 ;
  assign n28509 = n9199 | n22488 ;
  assign n28512 = n28511 ^ n28509 ^ 1'b0 ;
  assign n28507 = n1581 & n18556 ;
  assign n28508 = n20745 & n28507 ;
  assign n28513 = n28512 ^ n28508 ^ n22899 ;
  assign n28514 = ( ~n3026 & n6370 ) | ( ~n3026 & n13282 ) | ( n6370 & n13282 ) ;
  assign n28515 = ~n3996 & n28514 ;
  assign n28516 = n28515 ^ n12462 ^ 1'b0 ;
  assign n28526 = ( n1438 & ~n7650 ) | ( n1438 & n13986 ) | ( ~n7650 & n13986 ) ;
  assign n28525 = ~n10722 & n15567 ;
  assign n28527 = n28526 ^ n28525 ^ 1'b0 ;
  assign n28518 = n12562 ^ n10079 ^ n9794 ;
  assign n28517 = ~n261 & n12915 ;
  assign n28519 = n28518 ^ n28517 ^ 1'b0 ;
  assign n28520 = n28519 ^ n22840 ^ n3320 ;
  assign n28521 = ~n4540 & n28520 ;
  assign n28522 = ~n2864 & n10514 ;
  assign n28523 = n28522 ^ n24125 ^ 1'b0 ;
  assign n28524 = n28521 & ~n28523 ;
  assign n28528 = n28527 ^ n28524 ^ 1'b0 ;
  assign n28529 = n17417 | n28528 ;
  assign n28530 = n28529 ^ n11536 ^ 1'b0 ;
  assign n28531 = n21158 | n22987 ;
  assign n28535 = ( n10863 & n14421 ) | ( n10863 & ~n19925 ) | ( n14421 & ~n19925 ) ;
  assign n28532 = n11409 ^ n5740 ^ n1192 ;
  assign n28533 = n28532 ^ n21397 ^ 1'b0 ;
  assign n28534 = ~n26026 & n28533 ;
  assign n28536 = n28535 ^ n28534 ^ n16399 ;
  assign n28537 = n23235 & n28536 ;
  assign n28538 = n13417 ^ n5947 ^ n2340 ;
  assign n28539 = n28538 ^ n20972 ^ 1'b0 ;
  assign n28540 = x205 & ~n4538 ;
  assign n28541 = n17723 & n28540 ;
  assign n28546 = n955 & ~n2468 ;
  assign n28547 = n28546 ^ n10284 ^ 1'b0 ;
  assign n28545 = ( x5 & n11857 ) | ( x5 & n14237 ) | ( n11857 & n14237 ) ;
  assign n28542 = n3058 | n3202 ;
  assign n28543 = n28542 ^ n6369 ^ 1'b0 ;
  assign n28544 = n17183 & ~n28543 ;
  assign n28548 = n28547 ^ n28545 ^ n28544 ;
  assign n28549 = ( ~n26512 & n28541 ) | ( ~n26512 & n28548 ) | ( n28541 & n28548 ) ;
  assign n28550 = n14717 ^ n13341 ^ n6618 ;
  assign n28551 = n13516 & n20791 ;
  assign n28552 = n11303 ^ n6231 ^ 1'b0 ;
  assign n28553 = n28551 | n28552 ;
  assign n28555 = n9211 | n10157 ;
  assign n28554 = n13666 & ~n20019 ;
  assign n28556 = n28555 ^ n28554 ^ 1'b0 ;
  assign n28557 = n9963 ^ n6085 ^ 1'b0 ;
  assign n28558 = n28557 ^ n6833 ^ 1'b0 ;
  assign n28559 = n28558 ^ n13683 ^ n13234 ;
  assign n28560 = n28559 ^ n4283 ^ n1108 ;
  assign n28561 = n19238 ^ n6763 ^ 1'b0 ;
  assign n28562 = ~n23740 & n28561 ;
  assign n28563 = ~n7108 & n28562 ;
  assign n28564 = n28563 ^ n6349 ^ 1'b0 ;
  assign n28565 = n16145 ^ n15676 ^ n2347 ;
  assign n28566 = ( n4005 & n10895 ) | ( n4005 & n28565 ) | ( n10895 & n28565 ) ;
  assign n28567 = n18461 ^ n9771 ^ 1'b0 ;
  assign n28568 = n17444 ^ n15333 ^ 1'b0 ;
  assign n28569 = n7842 ^ n2045 ^ 1'b0 ;
  assign n28570 = ~n2582 & n28569 ;
  assign n28571 = n9458 ^ n8223 ^ n5780 ;
  assign n28572 = ( n10173 & ~n17276 ) | ( n10173 & n28571 ) | ( ~n17276 & n28571 ) ;
  assign n28573 = n18457 ^ n4284 ^ n3803 ;
  assign n28574 = n28573 ^ n20965 ^ 1'b0 ;
  assign n28575 = n28574 ^ n14816 ^ n5781 ;
  assign n28576 = n6782 | n18942 ;
  assign n28577 = n2428 & ~n28576 ;
  assign n28578 = n8008 | n20447 ;
  assign n28579 = n28577 | n28578 ;
  assign n28580 = n28355 | n28579 ;
  assign n28581 = n25597 ^ n9295 ^ n6331 ;
  assign n28582 = n28581 ^ n9129 ^ 1'b0 ;
  assign n28583 = n27700 ^ n9932 ^ n1153 ;
  assign n28584 = n28582 & n28583 ;
  assign n28585 = n28584 ^ n1487 ^ 1'b0 ;
  assign n28586 = n28585 ^ n13689 ^ 1'b0 ;
  assign n28587 = ( n9757 & ~n16590 ) | ( n9757 & n27425 ) | ( ~n16590 & n27425 ) ;
  assign n28589 = n13349 ^ n5110 ^ n2677 ;
  assign n28588 = n2555 & n26545 ;
  assign n28590 = n28589 ^ n28588 ^ n6852 ;
  assign n28591 = n1209 & n20876 ;
  assign n28592 = n400 & n13082 ;
  assign n28593 = n28592 ^ n3856 ^ 1'b0 ;
  assign n28594 = n28581 ^ n8498 ^ n5926 ;
  assign n28595 = n22390 & ~n28594 ;
  assign n28596 = n28595 ^ n13639 ^ 1'b0 ;
  assign n28597 = n25563 & ~n28596 ;
  assign n28598 = n28597 ^ n9087 ^ 1'b0 ;
  assign n28599 = n15506 ^ n7968 ^ n5823 ;
  assign n28600 = n28599 ^ n14228 ^ 1'b0 ;
  assign n28601 = n4876 & ~n6533 ;
  assign n28602 = n28601 ^ n28523 ^ 1'b0 ;
  assign n28603 = n10411 ^ n944 ^ 1'b0 ;
  assign n28604 = n28603 ^ n9824 ^ 1'b0 ;
  assign n28605 = ~n4820 & n28604 ;
  assign n28606 = n26312 ^ n23701 ^ 1'b0 ;
  assign n28607 = n18550 & ~n28606 ;
  assign n28608 = n28607 ^ n18292 ^ 1'b0 ;
  assign n28609 = ~n17824 & n28608 ;
  assign n28610 = n28609 ^ n26538 ^ 1'b0 ;
  assign n28612 = n5236 | n14621 ;
  assign n28611 = n27766 ^ n22605 ^ n7296 ;
  assign n28613 = n28612 ^ n28611 ^ n2643 ;
  assign n28614 = ( n431 & n3141 ) | ( n431 & n6931 ) | ( n3141 & n6931 ) ;
  assign n28615 = n3123 ^ n2234 ^ x159 ;
  assign n28616 = n28615 ^ n18049 ^ 1'b0 ;
  assign n28617 = ~n28614 & n28616 ;
  assign n28620 = ( ~n4502 & n6782 ) | ( ~n4502 & n9096 ) | ( n6782 & n9096 ) ;
  assign n28621 = n28620 ^ n15791 ^ n5112 ;
  assign n28618 = ( n7649 & ~n11376 ) | ( n7649 & n15345 ) | ( ~n11376 & n15345 ) ;
  assign n28619 = n19787 & n28618 ;
  assign n28622 = n28621 ^ n28619 ^ 1'b0 ;
  assign n28623 = n24444 ^ n11001 ^ 1'b0 ;
  assign n28624 = ~n28622 & n28623 ;
  assign n28625 = n14618 & n25498 ;
  assign n28626 = n21809 & ~n28625 ;
  assign n28627 = n4707 & n28626 ;
  assign n28628 = n2070 & ~n16047 ;
  assign n28629 = n8869 & n28628 ;
  assign n28630 = n704 & n8201 ;
  assign n28631 = n28630 ^ n1805 ^ 1'b0 ;
  assign n28632 = ~n20280 & n21431 ;
  assign n28633 = n28632 ^ n3491 ^ n1056 ;
  assign n28634 = n28319 & n28633 ;
  assign n28635 = n22512 & ~n24303 ;
  assign n28636 = ( n1624 & n6115 ) | ( n1624 & ~n27825 ) | ( n6115 & ~n27825 ) ;
  assign n28637 = n27930 & n28636 ;
  assign n28638 = n28637 ^ n5328 ^ 1'b0 ;
  assign n28639 = x151 & n28638 ;
  assign n28640 = ( n1192 & ~n1669 ) | ( n1192 & n12461 ) | ( ~n1669 & n12461 ) ;
  assign n28641 = n28640 ^ n6184 ^ n796 ;
  assign n28642 = ~n13390 & n28641 ;
  assign n28643 = n28642 ^ n11693 ^ 1'b0 ;
  assign n28644 = n28643 ^ n5201 ^ 1'b0 ;
  assign n28645 = n28639 & n28644 ;
  assign n28646 = ~n1754 & n3931 ;
  assign n28647 = n28646 ^ n3110 ^ 1'b0 ;
  assign n28648 = n28647 ^ n17787 ^ 1'b0 ;
  assign n28649 = ( n3254 & n4315 ) | ( n3254 & ~n6088 ) | ( n4315 & ~n6088 ) ;
  assign n28650 = n13621 | n28649 ;
  assign n28651 = n28650 ^ n16010 ^ 1'b0 ;
  assign n28652 = n2455 & n28651 ;
  assign n28653 = n7392 | n28652 ;
  assign n28654 = n28653 ^ n18853 ^ 1'b0 ;
  assign n28655 = n26199 ^ n8594 ^ 1'b0 ;
  assign n28656 = n7919 & ~n28655 ;
  assign n28657 = n28656 ^ n26034 ^ x66 ;
  assign n28658 = n21810 ^ n20754 ^ n3360 ;
  assign n28659 = n28658 ^ n3488 ^ 1'b0 ;
  assign n28660 = n2665 & n28659 ;
  assign n28661 = n27089 & ~n28660 ;
  assign n28662 = ~x24 & n28661 ;
  assign n28663 = n17088 ^ n3508 ^ n421 ;
  assign n28664 = n1900 ^ x36 ^ 1'b0 ;
  assign n28665 = n28664 ^ n19832 ^ n12973 ;
  assign n28666 = n12061 ^ n9465 ^ 1'b0 ;
  assign n28667 = n20256 | n28666 ;
  assign n28668 = n28665 | n28667 ;
  assign n28669 = n17961 | n28668 ;
  assign n28670 = n12570 ^ n3750 ^ 1'b0 ;
  assign n28671 = n7732 & n11762 ;
  assign n28672 = ( n5504 & ~n8156 ) | ( n5504 & n28671 ) | ( ~n8156 & n28671 ) ;
  assign n28673 = ~n5994 & n7633 ;
  assign n28674 = ~n26182 & n28673 ;
  assign n28675 = n28674 ^ n10472 ^ n2906 ;
  assign n28677 = n8598 | n23761 ;
  assign n28678 = n3802 & ~n28677 ;
  assign n28679 = n8819 & ~n28678 ;
  assign n28680 = ~n15244 & n28679 ;
  assign n28676 = n2338 & ~n24040 ;
  assign n28681 = n28680 ^ n28676 ^ n21322 ;
  assign n28682 = n3375 ^ n1102 ^ 1'b0 ;
  assign n28683 = n8904 | n13421 ;
  assign n28684 = ~n6068 & n23519 ;
  assign n28685 = n8253 & ~n13386 ;
  assign n28686 = n7343 & ~n28685 ;
  assign n28687 = ( n4763 & n5743 ) | ( n4763 & ~n28686 ) | ( n5743 & ~n28686 ) ;
  assign n28688 = n23991 ^ n10364 ^ 1'b0 ;
  assign n28689 = n28687 | n28688 ;
  assign n28690 = n8678 & ~n14963 ;
  assign n28691 = n28690 ^ n9151 ^ 1'b0 ;
  assign n28692 = ~n1988 & n22277 ;
  assign n28693 = ~n14995 & n28692 ;
  assign n28694 = n5452 ^ n4309 ^ 1'b0 ;
  assign n28695 = n12741 & n28694 ;
  assign n28696 = n28695 ^ n15359 ^ 1'b0 ;
  assign n28697 = ~n28693 & n28696 ;
  assign n28698 = n28697 ^ n22206 ^ n8638 ;
  assign n28706 = ~n2229 & n5709 ;
  assign n28702 = n21317 | n28177 ;
  assign n28703 = n17218 ^ n12861 ^ 1'b0 ;
  assign n28704 = ~n28702 & n28703 ;
  assign n28701 = n12031 & n24609 ;
  assign n28705 = n28704 ^ n28701 ^ 1'b0 ;
  assign n28699 = n18829 | n25844 ;
  assign n28700 = n5514 & n28699 ;
  assign n28707 = n28706 ^ n28705 ^ n28700 ;
  assign n28708 = n9536 ^ n3636 ^ 1'b0 ;
  assign n28709 = n22153 | n28708 ;
  assign n28710 = n3309 & ~n9189 ;
  assign n28711 = n28457 ^ n24022 ^ 1'b0 ;
  assign n28712 = n11371 | n28711 ;
  assign n28713 = ( n10546 & ~n26018 ) | ( n10546 & n28712 ) | ( ~n26018 & n28712 ) ;
  assign n28714 = ( ~n11684 & n28710 ) | ( ~n11684 & n28713 ) | ( n28710 & n28713 ) ;
  assign n28715 = n24735 ^ n17723 ^ 1'b0 ;
  assign n28716 = ( ~n4198 & n5430 ) | ( ~n4198 & n5473 ) | ( n5430 & n5473 ) ;
  assign n28717 = n5540 | n9469 ;
  assign n28718 = ( ~n5238 & n28716 ) | ( ~n5238 & n28717 ) | ( n28716 & n28717 ) ;
  assign n28719 = n1518 & n25587 ;
  assign n28720 = n28719 ^ n6973 ^ 1'b0 ;
  assign n28721 = n7666 & n18550 ;
  assign n28722 = n28721 ^ n13157 ^ 1'b0 ;
  assign n28723 = n1796 | n28722 ;
  assign n28724 = n12701 & ~n28723 ;
  assign n28726 = ( n2789 & n8280 ) | ( n2789 & n8628 ) | ( n8280 & n8628 ) ;
  assign n28725 = n1359 & n6117 ;
  assign n28727 = n28726 ^ n28725 ^ 1'b0 ;
  assign n28728 = n28727 ^ n18028 ^ n7507 ;
  assign n28729 = ~n12756 & n28728 ;
  assign n28730 = n16421 & ~n26568 ;
  assign n28731 = ~n18283 & n28730 ;
  assign n28734 = ( n3275 & n4739 ) | ( n3275 & ~n22286 ) | ( n4739 & ~n22286 ) ;
  assign n28732 = ~n14672 & n15174 ;
  assign n28733 = n20536 & n28732 ;
  assign n28735 = n28734 ^ n28733 ^ 1'b0 ;
  assign n28736 = ~n17295 & n28735 ;
  assign n28737 = n2739 & ~n13721 ;
  assign n28738 = n28737 ^ n13283 ^ 1'b0 ;
  assign n28739 = n28738 ^ n5302 ^ 1'b0 ;
  assign n28740 = ( n9472 & ~n20995 ) | ( n9472 & n26830 ) | ( ~n20995 & n26830 ) ;
  assign n28741 = n18800 ^ n2722 ^ 1'b0 ;
  assign n28742 = ~n28740 & n28741 ;
  assign n28743 = n4062 & ~n15191 ;
  assign n28744 = ~n9561 & n28743 ;
  assign n28745 = ( n352 & n24275 ) | ( n352 & n27488 ) | ( n24275 & n27488 ) ;
  assign n28746 = ~n6163 & n10043 ;
  assign n28747 = n6163 & n28746 ;
  assign n28748 = n19005 | n28747 ;
  assign n28749 = n19005 & ~n28748 ;
  assign n28750 = n24927 | n28749 ;
  assign n28751 = n6294 & ~n28750 ;
  assign n28752 = ( n280 & n20604 ) | ( n280 & ~n28751 ) | ( n20604 & ~n28751 ) ;
  assign n28753 = n16480 ^ n14265 ^ n11492 ;
  assign n28754 = n25054 ^ n6653 ^ 1'b0 ;
  assign n28755 = ~n28753 & n28754 ;
  assign n28756 = ~n8568 & n14766 ;
  assign n28757 = n28756 ^ n3757 ^ 1'b0 ;
  assign n28758 = n7201 & ~n9294 ;
  assign n28759 = n518 & n28758 ;
  assign n28760 = n21606 | n28759 ;
  assign n28761 = n28757 & ~n28760 ;
  assign n28762 = n28761 ^ n2380 ^ 1'b0 ;
  assign n28763 = n27290 & ~n28762 ;
  assign n28764 = n23022 ^ n16841 ^ n6408 ;
  assign n28765 = ( n5589 & n8087 ) | ( n5589 & n8604 ) | ( n8087 & n8604 ) ;
  assign n28766 = n2101 & n2814 ;
  assign n28767 = ~n13924 & n28766 ;
  assign n28770 = n20468 ^ x156 ^ 1'b0 ;
  assign n28768 = n26130 ^ n11033 ^ n3846 ;
  assign n28769 = n17565 & ~n28768 ;
  assign n28771 = n28770 ^ n28769 ^ 1'b0 ;
  assign n28772 = n28771 ^ n2377 ^ 1'b0 ;
  assign n28773 = ( ~n9907 & n28767 ) | ( ~n9907 & n28772 ) | ( n28767 & n28772 ) ;
  assign n28774 = ( ~n28764 & n28765 ) | ( ~n28764 & n28773 ) | ( n28765 & n28773 ) ;
  assign n28776 = n6984 | n7694 ;
  assign n28777 = n7817 | n28776 ;
  assign n28778 = ( ~n3858 & n10841 ) | ( ~n3858 & n28777 ) | ( n10841 & n28777 ) ;
  assign n28775 = n6045 & n22595 ;
  assign n28779 = n28778 ^ n28775 ^ n13421 ;
  assign n28780 = n16885 ^ n4516 ^ 1'b0 ;
  assign n28781 = ( ~n2084 & n5647 ) | ( ~n2084 & n6428 ) | ( n5647 & n6428 ) ;
  assign n28782 = n19628 & n28781 ;
  assign n28783 = n28782 ^ n18921 ^ 1'b0 ;
  assign n28784 = ~n10707 & n28783 ;
  assign n28785 = n19827 ^ n7781 ^ 1'b0 ;
  assign n28786 = n12730 & ~n15455 ;
  assign n28787 = n28786 ^ n6216 ^ 1'b0 ;
  assign n28788 = n28787 ^ n16895 ^ n1832 ;
  assign n28789 = ~x212 & n28788 ;
  assign n28791 = n15415 ^ n12504 ^ 1'b0 ;
  assign n28790 = n2268 & ~n18234 ;
  assign n28792 = n28791 ^ n28790 ^ 1'b0 ;
  assign n28793 = n17119 & n28792 ;
  assign n28794 = n19062 ^ x122 ^ 1'b0 ;
  assign n28801 = n21187 ^ n13256 ^ 1'b0 ;
  assign n28798 = n12653 & n19098 ;
  assign n28799 = n28798 ^ n8262 ^ 1'b0 ;
  assign n28800 = ( n1311 & n5309 ) | ( n1311 & n28799 ) | ( n5309 & n28799 ) ;
  assign n28795 = n26185 ^ n22912 ^ 1'b0 ;
  assign n28796 = n23709 & n28795 ;
  assign n28797 = n13232 & n28796 ;
  assign n28802 = n28801 ^ n28800 ^ n28797 ;
  assign n28803 = n6058 & ~n6941 ;
  assign n28804 = n964 & n28803 ;
  assign n28805 = n28804 ^ n14365 ^ n8657 ;
  assign n28806 = ( ~n12563 & n19648 ) | ( ~n12563 & n25805 ) | ( n19648 & n25805 ) ;
  assign n28807 = n10903 & ~n28806 ;
  assign n28808 = ~n15898 & n23878 ;
  assign n28809 = n17626 & n28808 ;
  assign n28810 = n16520 ^ n446 ^ 1'b0 ;
  assign n28811 = n28810 ^ n3887 ^ 1'b0 ;
  assign n28812 = n19401 & n19474 ;
  assign n28813 = n6398 & n7444 ;
  assign n28814 = n28813 ^ n23107 ^ n4656 ;
  assign n28815 = n4037 | n4600 ;
  assign n28816 = n7431 & ~n28815 ;
  assign n28817 = n28816 ^ n21403 ^ 1'b0 ;
  assign n28819 = n885 & n12469 ;
  assign n28818 = n3318 ^ n2878 ^ 1'b0 ;
  assign n28820 = n28819 ^ n28818 ^ n7314 ;
  assign n28821 = n11332 & n18330 ;
  assign n28822 = n10550 ^ n3432 ^ 1'b0 ;
  assign n28823 = n1912 | n28822 ;
  assign n28824 = n28823 ^ n26650 ^ 1'b0 ;
  assign n28825 = n3855 | n22303 ;
  assign n28826 = ~n14568 & n14768 ;
  assign n28827 = n28826 ^ n640 ^ 1'b0 ;
  assign n28828 = ( ~n10159 & n28825 ) | ( ~n10159 & n28827 ) | ( n28825 & n28827 ) ;
  assign n28829 = n24366 ^ n21238 ^ 1'b0 ;
  assign n28830 = n26816 | n28829 ;
  assign n28831 = n10317 ^ x19 ^ 1'b0 ;
  assign n28832 = n11443 & n28831 ;
  assign n28833 = n28832 ^ n18322 ^ 1'b0 ;
  assign n28834 = ~n7688 & n28833 ;
  assign n28835 = n28834 ^ n24685 ^ n16609 ;
  assign n28836 = n24301 ^ n10741 ^ 1'b0 ;
  assign n28837 = n6035 & n11724 ;
  assign n28838 = n24058 ^ n11075 ^ 1'b0 ;
  assign n28839 = n14126 & n18230 ;
  assign n28840 = ~n7015 & n28839 ;
  assign n28841 = n822 & ~n11024 ;
  assign n28842 = ~n7046 & n28841 ;
  assign n28843 = n28842 ^ n2009 ^ 1'b0 ;
  assign n28844 = ( n6912 & n7700 ) | ( n6912 & ~n14640 ) | ( n7700 & ~n14640 ) ;
  assign n28845 = ( n3855 & n5060 ) | ( n3855 & ~n8041 ) | ( n5060 & ~n8041 ) ;
  assign n28846 = n8041 & ~n17489 ;
  assign n28847 = ( n27433 & ~n28845 ) | ( n27433 & n28846 ) | ( ~n28845 & n28846 ) ;
  assign n28848 = n28847 ^ n7857 ^ 1'b0 ;
  assign n28849 = n24457 & ~n28848 ;
  assign n28853 = ~n3070 & n8262 ;
  assign n28854 = n9965 ^ n7285 ^ 1'b0 ;
  assign n28855 = n28853 | n28854 ;
  assign n28850 = ( ~n13181 & n19417 ) | ( ~n13181 & n21034 ) | ( n19417 & n21034 ) ;
  assign n28851 = n28850 ^ n9178 ^ 1'b0 ;
  assign n28852 = n3962 & n28851 ;
  assign n28856 = n28855 ^ n28852 ^ 1'b0 ;
  assign n28857 = n21582 ^ n15985 ^ 1'b0 ;
  assign n28858 = ~n2929 & n16414 ;
  assign n28859 = n28857 & n28858 ;
  assign n28860 = n23055 | n28859 ;
  assign n28861 = ( x215 & ~x222 ) | ( x215 & n1078 ) | ( ~x222 & n1078 ) ;
  assign n28862 = ~n6625 & n28861 ;
  assign n28863 = n28862 ^ n3521 ^ 1'b0 ;
  assign n28864 = n25204 ^ n5736 ^ 1'b0 ;
  assign n28865 = n18264 & ~n28864 ;
  assign n28866 = n1645 & n28865 ;
  assign n28867 = ~n26218 & n28866 ;
  assign n28868 = n28863 & n28867 ;
  assign n28869 = n28868 ^ n8558 ^ 1'b0 ;
  assign n28870 = n20905 ^ n2006 ^ 1'b0 ;
  assign n28871 = x119 & n10537 ;
  assign n28872 = n28870 & n28871 ;
  assign n28873 = n22929 ^ n8468 ^ n6694 ;
  assign n28874 = n1917 & n5122 ;
  assign n28875 = x137 & n5500 ;
  assign n28876 = ~n28874 & n28875 ;
  assign n28877 = ( ~n7323 & n14079 ) | ( ~n7323 & n18330 ) | ( n14079 & n18330 ) ;
  assign n28878 = n9634 & n10079 ;
  assign n28879 = n28878 ^ n9803 ^ 1'b0 ;
  assign n28880 = n28879 ^ n14292 ^ 1'b0 ;
  assign n28881 = ~n28877 & n28880 ;
  assign n28882 = ~n28876 & n28881 ;
  assign n28883 = n20077 ^ n3082 ^ 1'b0 ;
  assign n28884 = ( ~n1898 & n7327 ) | ( ~n1898 & n10562 ) | ( n7327 & n10562 ) ;
  assign n28885 = n28884 ^ n3208 ^ 1'b0 ;
  assign n28886 = ~n20112 & n28885 ;
  assign n28887 = n18466 ^ n8828 ^ n5424 ;
  assign n28888 = n28887 ^ n1342 ^ 1'b0 ;
  assign n28889 = n27619 | n28888 ;
  assign n28890 = n19192 & n26795 ;
  assign n28891 = n28890 ^ n4627 ^ 1'b0 ;
  assign n28892 = n18984 & ~n24088 ;
  assign n28893 = ~n23953 & n28892 ;
  assign n28894 = n18531 ^ n17068 ^ n10639 ;
  assign n28895 = n28894 ^ n8268 ^ 1'b0 ;
  assign n28896 = n16959 | n28895 ;
  assign n28897 = n28896 ^ n14590 ^ n10416 ;
  assign n28898 = n28897 ^ n27281 ^ n2586 ;
  assign n28899 = n16733 & ~n21269 ;
  assign n28900 = ~n6912 & n28899 ;
  assign n28901 = n13283 | n28900 ;
  assign n28902 = ( n6586 & ~n12383 ) | ( n6586 & n13673 ) | ( ~n12383 & n13673 ) ;
  assign n28903 = n28902 ^ n23215 ^ n15486 ;
  assign n28904 = n11281 ^ n3429 ^ n1097 ;
  assign n28905 = ( n13795 & n28363 ) | ( n13795 & n28904 ) | ( n28363 & n28904 ) ;
  assign n28906 = n28905 ^ n13408 ^ 1'b0 ;
  assign n28907 = n3156 & ~n13882 ;
  assign n28908 = ~n13540 & n28907 ;
  assign n28909 = n28908 ^ n11350 ^ 1'b0 ;
  assign n28910 = n13207 | n15820 ;
  assign n28911 = ( n11747 & n13778 ) | ( n11747 & n18570 ) | ( n13778 & n18570 ) ;
  assign n28921 = n11732 ^ x138 ^ 1'b0 ;
  assign n28912 = ( n13296 & n14817 ) | ( n13296 & ~n23285 ) | ( n14817 & ~n23285 ) ;
  assign n28913 = n12023 ^ n1035 ^ 1'b0 ;
  assign n28914 = n26734 | n28913 ;
  assign n28915 = n25338 ^ n4471 ^ 1'b0 ;
  assign n28916 = ~n28914 & n28915 ;
  assign n28917 = ~n16141 & n28916 ;
  assign n28918 = n28912 & n28917 ;
  assign n28919 = n9169 | n28918 ;
  assign n28920 = n28919 ^ n26199 ^ 1'b0 ;
  assign n28922 = n28921 ^ n28920 ^ n7307 ;
  assign n28926 = ( ~n6551 & n7403 ) | ( ~n6551 & n11677 ) | ( n7403 & n11677 ) ;
  assign n28924 = n964 & ~n3805 ;
  assign n28923 = n1912 & ~n20814 ;
  assign n28925 = n28924 ^ n28923 ^ 1'b0 ;
  assign n28927 = n28926 ^ n28925 ^ n16507 ;
  assign n28928 = ( x191 & ~n11512 ) | ( x191 & n15425 ) | ( ~n11512 & n15425 ) ;
  assign n28929 = n28928 ^ n13776 ^ n13510 ;
  assign n28932 = n22133 ^ n9016 ^ 1'b0 ;
  assign n28930 = n7452 ^ n6780 ^ 1'b0 ;
  assign n28931 = ~n22605 & n28930 ;
  assign n28933 = n28932 ^ n28931 ^ 1'b0 ;
  assign n28934 = n24231 & n28933 ;
  assign n28935 = n18067 | n20300 ;
  assign n28936 = n910 | n28935 ;
  assign n28937 = n17628 ^ n6324 ^ 1'b0 ;
  assign n28938 = ~n6495 & n28937 ;
  assign n28939 = ( n3459 & ~n6011 ) | ( n3459 & n21749 ) | ( ~n6011 & n21749 ) ;
  assign n28940 = ( n3116 & n7240 ) | ( n3116 & ~n7573 ) | ( n7240 & ~n7573 ) ;
  assign n28941 = ( x54 & n1919 ) | ( x54 & n4466 ) | ( n1919 & n4466 ) ;
  assign n28942 = n2860 & n17470 ;
  assign n28943 = n28942 ^ n8982 ^ 1'b0 ;
  assign n28944 = n17350 | n19689 ;
  assign n28945 = ( n12516 & n18595 ) | ( n12516 & n28944 ) | ( n18595 & n28944 ) ;
  assign n28946 = n4077 & n22025 ;
  assign n28947 = n28946 ^ n19587 ^ 1'b0 ;
  assign n28948 = ~n3122 & n4719 ;
  assign n28949 = n28948 ^ n6113 ^ 1'b0 ;
  assign n28950 = ( n3029 & ~n9636 ) | ( n3029 & n28949 ) | ( ~n9636 & n28949 ) ;
  assign n28951 = n22053 | n28950 ;
  assign n28952 = n28947 & ~n28951 ;
  assign n28953 = n13724 | n27120 ;
  assign n28954 = n4573 & n17561 ;
  assign n28955 = n28954 ^ n9588 ^ x98 ;
  assign n28956 = n23087 ^ n13570 ^ n3430 ;
  assign n28957 = n18059 ^ n455 ^ 1'b0 ;
  assign n28958 = ~n6733 & n28957 ;
  assign n28959 = ( ~n3466 & n3627 ) | ( ~n3466 & n3713 ) | ( n3627 & n3713 ) ;
  assign n28960 = n24343 | n28959 ;
  assign n28961 = n28960 ^ n15333 ^ 1'b0 ;
  assign n28962 = n20727 ^ n12832 ^ 1'b0 ;
  assign n28963 = n11795 & n28962 ;
  assign n28964 = ( n2113 & n28961 ) | ( n2113 & n28963 ) | ( n28961 & n28963 ) ;
  assign n28965 = n10653 & n15526 ;
  assign n28966 = n28024 ^ n15347 ^ 1'b0 ;
  assign n28967 = n912 & ~n28966 ;
  assign n28968 = n9449 ^ n3056 ^ 1'b0 ;
  assign n28969 = n16034 ^ n3435 ^ 1'b0 ;
  assign n28970 = ~n4068 & n28969 ;
  assign n28971 = n912 & n28970 ;
  assign n28972 = n28971 ^ n13450 ^ 1'b0 ;
  assign n28973 = n333 & ~n28972 ;
  assign n28974 = n28973 ^ n20328 ^ 1'b0 ;
  assign n28975 = ( n28967 & n28968 ) | ( n28967 & n28974 ) | ( n28968 & n28974 ) ;
  assign n28979 = ( n2113 & n6414 ) | ( n2113 & n21244 ) | ( n6414 & n21244 ) ;
  assign n28980 = n28979 ^ n1191 ^ 1'b0 ;
  assign n28977 = n1468 & ~n12308 ;
  assign n28978 = n4006 & n28977 ;
  assign n28976 = n663 & n15744 ;
  assign n28981 = n28980 ^ n28978 ^ n28976 ;
  assign n28982 = n2033 & ~n7248 ;
  assign n28983 = n8106 & n28982 ;
  assign n28984 = n28983 ^ n16810 ^ 1'b0 ;
  assign n28992 = n8495 ^ n8127 ^ n6626 ;
  assign n28993 = n18535 ^ n9137 ^ n5331 ;
  assign n28994 = ~n28992 & n28993 ;
  assign n28985 = n1022 | n9406 ;
  assign n28986 = ~n5146 & n12905 ;
  assign n28987 = n23313 & n28986 ;
  assign n28988 = ( n3303 & n11339 ) | ( n3303 & ~n28987 ) | ( n11339 & ~n28987 ) ;
  assign n28989 = n2861 & n28988 ;
  assign n28990 = n28989 ^ n13274 ^ 1'b0 ;
  assign n28991 = n28985 & n28990 ;
  assign n28995 = n28994 ^ n28991 ^ 1'b0 ;
  assign n28996 = n4249 & ~n4670 ;
  assign n28997 = n4217 & ~n22246 ;
  assign n28998 = n28997 ^ n17071 ^ 1'b0 ;
  assign n28999 = n28998 ^ n22167 ^ n4108 ;
  assign n29000 = ( n939 & ~n5675 ) | ( n939 & n16112 ) | ( ~n5675 & n16112 ) ;
  assign n29001 = n13000 & ~n29000 ;
  assign n29006 = n24307 ^ n18891 ^ 1'b0 ;
  assign n29007 = n3521 | n29006 ;
  assign n29005 = x28 & n24391 ;
  assign n29008 = n29007 ^ n29005 ^ n3699 ;
  assign n29009 = n29008 ^ n7731 ^ 1'b0 ;
  assign n29002 = ( ~n8177 & n12767 ) | ( ~n8177 & n19432 ) | ( n12767 & n19432 ) ;
  assign n29003 = ( ~n14689 & n15009 ) | ( ~n14689 & n29002 ) | ( n15009 & n29002 ) ;
  assign n29004 = ( n16449 & n20885 ) | ( n16449 & n29003 ) | ( n20885 & n29003 ) ;
  assign n29010 = n29009 ^ n29004 ^ n12343 ;
  assign n29011 = x114 & n6824 ;
  assign n29012 = n29011 ^ n14802 ^ x59 ;
  assign n29013 = n20937 ^ n18249 ^ n11368 ;
  assign n29014 = n26288 ^ n23383 ^ n14891 ;
  assign n29015 = ~n21378 & n23406 ;
  assign n29016 = ~n2530 & n29015 ;
  assign n29017 = n5228 | n7784 ;
  assign n29018 = n4987 & ~n29017 ;
  assign n29019 = n29018 ^ n10536 ^ 1'b0 ;
  assign n29020 = n25148 ^ n2853 ^ 1'b0 ;
  assign n29021 = n26916 & n29020 ;
  assign n29022 = ( n14146 & n15360 ) | ( n14146 & ~n24564 ) | ( n15360 & ~n24564 ) ;
  assign n29024 = n2390 & n8495 ;
  assign n29023 = x103 & n12581 ;
  assign n29025 = n29024 ^ n29023 ^ 1'b0 ;
  assign n29026 = n29025 ^ n28201 ^ n19711 ;
  assign n29027 = n29026 ^ n27373 ^ 1'b0 ;
  assign n29028 = n13558 & n16456 ;
  assign n29029 = n8667 ^ n3801 ^ n1359 ;
  assign n29030 = ( ~n4335 & n10280 ) | ( ~n4335 & n29029 ) | ( n10280 & n29029 ) ;
  assign n29031 = ~n14050 & n29030 ;
  assign n29034 = n20350 ^ n16148 ^ 1'b0 ;
  assign n29035 = n18174 | n29034 ;
  assign n29036 = n962 | n29035 ;
  assign n29032 = n11930 | n18885 ;
  assign n29033 = n29032 ^ n1971 ^ 1'b0 ;
  assign n29037 = n29036 ^ n29033 ^ n12604 ;
  assign n29038 = n3984 & ~n25295 ;
  assign n29039 = n13557 | n27889 ;
  assign n29040 = ~n4064 & n11868 ;
  assign n29041 = ( n10377 & n14886 ) | ( n10377 & n22617 ) | ( n14886 & n22617 ) ;
  assign n29042 = ( n2345 & n29040 ) | ( n2345 & ~n29041 ) | ( n29040 & ~n29041 ) ;
  assign n29043 = n23852 ^ n12570 ^ 1'b0 ;
  assign n29044 = n18266 | n21489 ;
  assign n29045 = n5132 ^ n2406 ^ 1'b0 ;
  assign n29046 = n5201 & n29045 ;
  assign n29047 = ( ~n18128 & n28087 ) | ( ~n18128 & n29046 ) | ( n28087 & n29046 ) ;
  assign n29048 = ~n3675 & n12152 ;
  assign n29050 = n23562 ^ n9704 ^ n6045 ;
  assign n29051 = n14774 & ~n29050 ;
  assign n29052 = ~n3823 & n29051 ;
  assign n29049 = n23608 ^ n12891 ^ 1'b0 ;
  assign n29053 = n29052 ^ n29049 ^ 1'b0 ;
  assign n29054 = n29053 ^ n25538 ^ n10078 ;
  assign n29055 = n17081 ^ n16952 ^ 1'b0 ;
  assign n29056 = n17012 & n29055 ;
  assign n29057 = n26527 & n29056 ;
  assign n29058 = n2614 | n23626 ;
  assign n29059 = n29058 ^ n16316 ^ 1'b0 ;
  assign n29060 = ( ~n1764 & n8073 ) | ( ~n1764 & n19149 ) | ( n8073 & n19149 ) ;
  assign n29061 = n27496 & ~n29060 ;
  assign n29062 = n29061 ^ n15041 ^ 1'b0 ;
  assign n29067 = n14873 ^ n2858 ^ 1'b0 ;
  assign n29066 = ( n1607 & n18770 ) | ( n1607 & n26984 ) | ( n18770 & n26984 ) ;
  assign n29063 = ~n4284 & n23761 ;
  assign n29064 = n29063 ^ n19758 ^ n12012 ;
  assign n29065 = n8230 | n29064 ;
  assign n29068 = n29067 ^ n29066 ^ n29065 ;
  assign n29069 = n22467 & ~n29068 ;
  assign n29070 = ( n6928 & n8574 ) | ( n6928 & n9499 ) | ( n8574 & n9499 ) ;
  assign n29071 = n29070 ^ n8357 ^ 1'b0 ;
  assign n29072 = n29071 ^ n26875 ^ n675 ;
  assign n29073 = ( n17314 & ~n23378 ) | ( n17314 & n23717 ) | ( ~n23378 & n23717 ) ;
  assign n29074 = ~x14 & n12421 ;
  assign n29075 = n29074 ^ n1078 ^ 1'b0 ;
  assign n29078 = n5710 & ~n18467 ;
  assign n29079 = n29078 ^ n6840 ^ 1'b0 ;
  assign n29076 = n18281 ^ n3377 ^ 1'b0 ;
  assign n29077 = n29076 ^ n15011 ^ 1'b0 ;
  assign n29080 = n29079 ^ n29077 ^ 1'b0 ;
  assign n29081 = ~n29075 & n29080 ;
  assign n29082 = n29081 ^ n22479 ^ n8872 ;
  assign n29084 = n1588 ^ n1484 ^ 1'b0 ;
  assign n29083 = n14798 & n25717 ;
  assign n29085 = n29084 ^ n29083 ^ 1'b0 ;
  assign n29086 = n29085 ^ n25986 ^ n3791 ;
  assign n29087 = n5485 ^ x115 ^ 1'b0 ;
  assign n29088 = n29087 ^ n6545 ^ 1'b0 ;
  assign n29089 = x21 & ~n29088 ;
  assign n29090 = n29089 ^ n6435 ^ n1446 ;
  assign n29091 = ( n27187 & n27430 ) | ( n27187 & ~n29090 ) | ( n27430 & ~n29090 ) ;
  assign n29092 = n7183 ^ n2117 ^ n363 ;
  assign n29093 = n11647 & ~n29092 ;
  assign n29094 = ~n13684 & n29093 ;
  assign n29095 = ( ~n15911 & n18294 ) | ( ~n15911 & n29094 ) | ( n18294 & n29094 ) ;
  assign n29096 = n5025 & n11632 ;
  assign n29097 = n4242 | n29096 ;
  assign n29098 = n29097 ^ n5965 ^ 1'b0 ;
  assign n29099 = ( n12638 & n29095 ) | ( n12638 & ~n29098 ) | ( n29095 & ~n29098 ) ;
  assign n29100 = n28765 ^ n11129 ^ 1'b0 ;
  assign n29101 = n9120 & ~n29100 ;
  assign n29102 = n23329 ^ n2665 ^ 1'b0 ;
  assign n29104 = n2194 | n11153 ;
  assign n29103 = ( n3557 & n8239 ) | ( n3557 & ~n18895 ) | ( n8239 & ~n18895 ) ;
  assign n29105 = n29104 ^ n29103 ^ 1'b0 ;
  assign n29106 = n29105 ^ n14981 ^ 1'b0 ;
  assign n29107 = n8250 & n29106 ;
  assign n29108 = n17310 ^ n10841 ^ 1'b0 ;
  assign n29109 = n29108 ^ n11190 ^ 1'b0 ;
  assign n29110 = n9228 & ~n10688 ;
  assign n29111 = n18254 & n29110 ;
  assign n29112 = n29111 ^ n16788 ^ 1'b0 ;
  assign n29113 = ~n27622 & n29112 ;
  assign n29114 = n2585 & ~n4703 ;
  assign n29115 = ~n29113 & n29114 ;
  assign n29116 = n29115 ^ n11507 ^ n9921 ;
  assign n29117 = n8367 ^ n3116 ^ 1'b0 ;
  assign n29118 = n29117 ^ n4443 ^ 1'b0 ;
  assign n29119 = n8898 & n29118 ;
  assign n29120 = n10125 & n29119 ;
  assign n29121 = n15320 ^ n2006 ^ 1'b0 ;
  assign n29122 = n29121 ^ n7671 ^ 1'b0 ;
  assign n29123 = n2615 & ~n7288 ;
  assign n29124 = n17971 & n29123 ;
  assign n29125 = n29124 ^ n21581 ^ n18717 ;
  assign n29126 = ~n6017 & n23992 ;
  assign n29127 = n29125 & n29126 ;
  assign n29128 = n26187 ^ n5148 ^ n2246 ;
  assign n29129 = ( n757 & ~n7270 ) | ( n757 & n8063 ) | ( ~n7270 & n8063 ) ;
  assign n29130 = n29129 ^ n16270 ^ n3444 ;
  assign n29131 = ( n5076 & n21430 ) | ( n5076 & n29130 ) | ( n21430 & n29130 ) ;
  assign n29132 = n8703 & n21893 ;
  assign n29133 = n17267 & n29132 ;
  assign n29134 = ( ~n315 & n5440 ) | ( ~n315 & n20410 ) | ( n5440 & n20410 ) ;
  assign n29135 = n13097 ^ n5177 ^ n268 ;
  assign n29136 = ( x134 & ~n25480 ) | ( x134 & n26848 ) | ( ~n25480 & n26848 ) ;
  assign n29137 = ~n19832 & n25395 ;
  assign n29138 = n10204 & n29137 ;
  assign n29139 = n29136 | n29138 ;
  assign n29140 = n29139 ^ n615 ^ 1'b0 ;
  assign n29141 = n6186 & ~n15841 ;
  assign n29142 = n13713 ^ n6286 ^ 1'b0 ;
  assign n29144 = n8496 ^ n4996 ^ n4095 ;
  assign n29143 = ( x56 & n12829 ) | ( x56 & ~n19523 ) | ( n12829 & ~n19523 ) ;
  assign n29145 = n29144 ^ n29143 ^ n8942 ;
  assign n29146 = ~n2786 & n19109 ;
  assign n29147 = n28375 ^ n14622 ^ n262 ;
  assign n29148 = n4540 & n14086 ;
  assign n29149 = n29148 ^ n13794 ^ 1'b0 ;
  assign n29150 = n29149 ^ n13351 ^ 1'b0 ;
  assign n29151 = n7968 | n10995 ;
  assign n29152 = n26284 | n29151 ;
  assign n29153 = ( n2076 & n7055 ) | ( n2076 & ~n14607 ) | ( n7055 & ~n14607 ) ;
  assign n29154 = ( ~n1304 & n8709 ) | ( ~n1304 & n19020 ) | ( n8709 & n19020 ) ;
  assign n29155 = n29154 ^ n20711 ^ 1'b0 ;
  assign n29156 = n29153 & n29155 ;
  assign n29157 = ( ~n6729 & n11224 ) | ( ~n6729 & n16004 ) | ( n11224 & n16004 ) ;
  assign n29158 = n9987 | n29157 ;
  assign n29159 = n29156 | n29158 ;
  assign n29160 = n7206 ^ n6493 ^ 1'b0 ;
  assign n29161 = ~n5157 & n29160 ;
  assign n29162 = n22724 ^ n8931 ^ 1'b0 ;
  assign n29163 = ~n2697 & n29162 ;
  assign n29165 = n6991 ^ n3114 ^ 1'b0 ;
  assign n29164 = n16559 | n23780 ;
  assign n29166 = n29165 ^ n29164 ^ 1'b0 ;
  assign n29167 = ( ~n24088 & n24494 ) | ( ~n24088 & n29166 ) | ( n24494 & n29166 ) ;
  assign n29168 = ( ~n29161 & n29163 ) | ( ~n29161 & n29167 ) | ( n29163 & n29167 ) ;
  assign n29169 = n8225 | n17890 ;
  assign n29170 = n29169 ^ n7334 ^ 1'b0 ;
  assign n29171 = n29170 ^ n25740 ^ n2696 ;
  assign n29172 = n29171 ^ n16453 ^ n2031 ;
  assign n29173 = n29172 ^ n14741 ^ n7052 ;
  assign n29174 = ( ~n10399 & n13687 ) | ( ~n10399 & n29173 ) | ( n13687 & n29173 ) ;
  assign n29175 = n8418 | n9186 ;
  assign n29176 = ~n8333 & n29175 ;
  assign n29177 = n7527 & ~n29176 ;
  assign n29178 = n29177 ^ n7355 ^ 1'b0 ;
  assign n29179 = n19556 | n29178 ;
  assign n29183 = n29108 ^ n11740 ^ 1'b0 ;
  assign n29180 = ~n9457 & n12184 ;
  assign n29181 = n29180 ^ n15375 ^ 1'b0 ;
  assign n29182 = ~n16458 & n29181 ;
  assign n29184 = n29183 ^ n29182 ^ 1'b0 ;
  assign n29187 = ( ~n1518 & n3309 ) | ( ~n1518 & n25170 ) | ( n3309 & n25170 ) ;
  assign n29185 = n10013 ^ n4826 ^ n1621 ;
  assign n29186 = ( n19303 & n20688 ) | ( n19303 & ~n29185 ) | ( n20688 & ~n29185 ) ;
  assign n29188 = n29187 ^ n29186 ^ n25135 ;
  assign n29190 = ~n24163 & n28639 ;
  assign n29189 = ~n22431 & n24818 ;
  assign n29191 = n29190 ^ n29189 ^ 1'b0 ;
  assign n29192 = n24759 ^ n22113 ^ n4575 ;
  assign n29193 = ( n533 & n591 ) | ( n533 & ~n16356 ) | ( n591 & ~n16356 ) ;
  assign n29194 = n13238 | n19950 ;
  assign n29195 = n23626 | n29194 ;
  assign n29196 = n12312 | n29195 ;
  assign n29197 = n29196 ^ n15313 ^ n4906 ;
  assign n29198 = ~n7453 & n9966 ;
  assign n29199 = n29197 & n29198 ;
  assign n29200 = ~n8243 & n24237 ;
  assign n29201 = ( ~n6800 & n18471 ) | ( ~n6800 & n28261 ) | ( n18471 & n28261 ) ;
  assign n29202 = ~n9933 & n28204 ;
  assign n29203 = n9541 | n11177 ;
  assign n29204 = n1850 & ~n29203 ;
  assign n29210 = n7969 & ~n23739 ;
  assign n29211 = n19775 & n29210 ;
  assign n29206 = n24589 ^ n24401 ^ 1'b0 ;
  assign n29207 = n29206 ^ n23008 ^ n9389 ;
  assign n29205 = ~n1607 & n14543 ;
  assign n29208 = n29207 ^ n29205 ^ 1'b0 ;
  assign n29209 = ~n2063 & n29208 ;
  assign n29212 = n29211 ^ n29209 ^ 1'b0 ;
  assign n29213 = n7123 & ~n29212 ;
  assign n29214 = n29213 ^ n19925 ^ 1'b0 ;
  assign n29215 = n13556 ^ n6091 ^ 1'b0 ;
  assign n29216 = n7213 & ~n29215 ;
  assign n29217 = n29216 ^ n637 ^ 1'b0 ;
  assign n29218 = n8577 & n25628 ;
  assign n29219 = n29218 ^ n6630 ^ 1'b0 ;
  assign n29220 = n6136 | n29219 ;
  assign n29221 = n29217 | n29220 ;
  assign n29222 = n18643 ^ n4340 ^ 1'b0 ;
  assign n29224 = n9468 ^ n2945 ^ 1'b0 ;
  assign n29225 = n7151 & ~n29224 ;
  assign n29226 = ~n8120 & n29225 ;
  assign n29223 = n1199 | n5240 ;
  assign n29227 = n29226 ^ n29223 ^ 1'b0 ;
  assign n29228 = n20602 | n29108 ;
  assign n29230 = n24266 ^ n11385 ^ 1'b0 ;
  assign n29231 = n14515 & n29230 ;
  assign n29229 = n15561 & n25627 ;
  assign n29232 = n29231 ^ n29229 ^ 1'b0 ;
  assign n29233 = n28740 ^ n27201 ^ n18218 ;
  assign n29234 = ( ~n8306 & n10049 ) | ( ~n8306 & n12418 ) | ( n10049 & n12418 ) ;
  assign n29235 = n25526 ^ n393 ^ 1'b0 ;
  assign n29236 = n21970 ^ n9816 ^ 1'b0 ;
  assign n29237 = n16371 & ~n29236 ;
  assign n29238 = n8992 & ~n29237 ;
  assign n29239 = n5449 & n9479 ;
  assign n29240 = ~n506 & n29239 ;
  assign n29241 = n29240 ^ n24681 ^ n16459 ;
  assign n29242 = ~n21584 & n21897 ;
  assign n29243 = n29242 ^ n23679 ^ n7519 ;
  assign n29244 = n12428 ^ n5236 ^ 1'b0 ;
  assign n29245 = ~n3672 & n29244 ;
  assign n29246 = n11416 & n15953 ;
  assign n29247 = n23486 & ~n29246 ;
  assign n29248 = ~n29245 & n29247 ;
  assign n29249 = n11179 | n23687 ;
  assign n29250 = n29249 ^ n7524 ^ 1'b0 ;
  assign n29251 = n532 | n29250 ;
  assign n29252 = n15153 & n21497 ;
  assign n29253 = n5470 | n29252 ;
  assign n29254 = n15518 ^ n9494 ^ n6798 ;
  assign n29255 = n24983 ^ n12090 ^ 1'b0 ;
  assign n29256 = n29254 & ~n29255 ;
  assign n29258 = n26165 ^ n4552 ^ 1'b0 ;
  assign n29259 = x168 & ~n29258 ;
  assign n29257 = ~n8027 & n10423 ;
  assign n29260 = n29259 ^ n29257 ^ 1'b0 ;
  assign n29267 = ~n5947 & n7792 ;
  assign n29268 = n19857 & n29267 ;
  assign n29269 = n17186 & ~n29268 ;
  assign n29270 = n29269 ^ n13539 ^ 1'b0 ;
  assign n29261 = n4560 ^ n2367 ^ 1'b0 ;
  assign n29262 = n29261 ^ n7323 ^ 1'b0 ;
  assign n29263 = n29262 ^ n23430 ^ n8458 ;
  assign n29264 = n29263 ^ n11378 ^ n5722 ;
  assign n29265 = n29264 ^ n3375 ^ n2542 ;
  assign n29266 = n10674 | n29265 ;
  assign n29271 = n29270 ^ n29266 ^ 1'b0 ;
  assign n29272 = n3902 ^ n1672 ^ n1229 ;
  assign n29273 = n16203 ^ n5620 ^ 1'b0 ;
  assign n29274 = n29273 ^ n2091 ^ 1'b0 ;
  assign n29275 = n14944 | n19508 ;
  assign n29276 = ~n6121 & n28286 ;
  assign n29277 = ~n9798 & n29276 ;
  assign n29278 = n2398 & n3532 ;
  assign n29279 = ( n7491 & n25740 ) | ( n7491 & ~n29278 ) | ( n25740 & ~n29278 ) ;
  assign n29280 = n3012 | n29279 ;
  assign n29281 = n23358 | n29280 ;
  assign n29282 = n3256 | n11454 ;
  assign n29283 = n21393 | n22808 ;
  assign n29284 = ( n3315 & n8169 ) | ( n3315 & n13835 ) | ( n8169 & n13835 ) ;
  assign n29285 = n6868 | n15651 ;
  assign n29286 = n11064 | n29285 ;
  assign n29287 = n21157 & n29286 ;
  assign n29288 = ~n8367 & n18390 ;
  assign n29289 = n17312 ^ n9195 ^ n8584 ;
  assign n29290 = n29289 ^ n9492 ^ n683 ;
  assign n29291 = n13771 & ~n29290 ;
  assign n29292 = n25810 & n29291 ;
  assign n29293 = ( ~n5447 & n11565 ) | ( ~n5447 & n15673 ) | ( n11565 & n15673 ) ;
  assign n29294 = n15056 ^ n6387 ^ 1'b0 ;
  assign n29295 = ~n4062 & n29294 ;
  assign n29296 = ( n13875 & ~n29293 ) | ( n13875 & n29295 ) | ( ~n29293 & n29295 ) ;
  assign n29297 = ( n4343 & n11334 ) | ( n4343 & n20611 ) | ( n11334 & n20611 ) ;
  assign n29298 = n29297 ^ n10310 ^ 1'b0 ;
  assign n29299 = n29296 & n29298 ;
  assign n29300 = n4704 ^ n1759 ^ n952 ;
  assign n29301 = ( n9131 & ~n10340 ) | ( n9131 & n22457 ) | ( ~n10340 & n22457 ) ;
  assign n29302 = n29301 ^ n25020 ^ n7142 ;
  assign n29311 = n13037 ^ n9934 ^ 1'b0 ;
  assign n29312 = n2628 | n29311 ;
  assign n29313 = n29312 ^ n20675 ^ 1'b0 ;
  assign n29307 = n12859 ^ n2613 ^ 1'b0 ;
  assign n29308 = n22170 | n29307 ;
  assign n29303 = n26332 ^ n3052 ^ 1'b0 ;
  assign n29304 = n10001 & n29303 ;
  assign n29305 = ( x147 & n19229 ) | ( x147 & ~n29304 ) | ( n19229 & ~n29304 ) ;
  assign n29306 = n12094 | n29305 ;
  assign n29309 = n29308 ^ n29306 ^ n13814 ;
  assign n29310 = ~n7154 & n29309 ;
  assign n29314 = n29313 ^ n29310 ^ 1'b0 ;
  assign n29315 = x146 & ~n10427 ;
  assign n29316 = n29315 ^ n1133 ^ 1'b0 ;
  assign n29317 = ( n1075 & n10294 ) | ( n1075 & ~n19478 ) | ( n10294 & ~n19478 ) ;
  assign n29318 = n29317 ^ n28709 ^ n19963 ;
  assign n29319 = n9199 ^ n6061 ^ n2152 ;
  assign n29324 = ( ~n4168 & n8031 ) | ( ~n4168 & n8175 ) | ( n8031 & n8175 ) ;
  assign n29325 = n29324 ^ n21791 ^ n8361 ;
  assign n29320 = ( n3401 & n8976 ) | ( n3401 & ~n11737 ) | ( n8976 & ~n11737 ) ;
  assign n29321 = n13334 ^ n5843 ^ x96 ;
  assign n29322 = n29320 & ~n29321 ;
  assign n29323 = ~n6515 & n29322 ;
  assign n29326 = n29325 ^ n29323 ^ 1'b0 ;
  assign n29327 = n29326 ^ n10811 ^ 1'b0 ;
  assign n29328 = n14323 | n14443 ;
  assign n29329 = n29328 ^ n27175 ^ 1'b0 ;
  assign n29330 = n29329 ^ n19112 ^ 1'b0 ;
  assign n29331 = n1623 & n15502 ;
  assign n29332 = ~n3249 & n29331 ;
  assign n29333 = n8625 & ~n29332 ;
  assign n29334 = n10615 & n29333 ;
  assign n29335 = n27458 | n29334 ;
  assign n29336 = n29330 | n29335 ;
  assign n29337 = n17897 ^ n9076 ^ 1'b0 ;
  assign n29338 = ( n17154 & ~n23393 ) | ( n17154 & n29337 ) | ( ~n23393 & n29337 ) ;
  assign n29339 = ( n1367 & n2513 ) | ( n1367 & n7696 ) | ( n2513 & n7696 ) ;
  assign n29340 = n8315 & ~n29339 ;
  assign n29341 = n2155 & n29340 ;
  assign n29342 = n5592 | n17970 ;
  assign n29343 = n27780 ^ n3000 ^ 1'b0 ;
  assign n29344 = n25003 & n29343 ;
  assign n29345 = n29344 ^ n23073 ^ n5853 ;
  assign n29346 = n6941 | n7170 ;
  assign n29347 = ~n6409 & n21478 ;
  assign n29348 = n29347 ^ n15113 ^ 1'b0 ;
  assign n29349 = ( n23991 & ~n29346 ) | ( n23991 & n29348 ) | ( ~n29346 & n29348 ) ;
  assign n29350 = n29349 ^ n28166 ^ n24504 ;
  assign n29351 = n24040 ^ n3112 ^ 1'b0 ;
  assign n29352 = n29351 ^ n3613 ^ n3382 ;
  assign n29359 = ~n9422 & n13995 ;
  assign n29353 = n9291 ^ n4250 ^ 1'b0 ;
  assign n29355 = n4109 | n8155 ;
  assign n29354 = n22904 ^ n10571 ^ n8013 ;
  assign n29356 = n29355 ^ n29354 ^ 1'b0 ;
  assign n29357 = n29353 & n29356 ;
  assign n29358 = n3826 | n29357 ;
  assign n29360 = n29359 ^ n29358 ^ 1'b0 ;
  assign n29361 = n26358 & n29360 ;
  assign n29362 = n19776 ^ n17408 ^ 1'b0 ;
  assign n29363 = n17256 | n29362 ;
  assign n29364 = n11649 | n29363 ;
  assign n29365 = ( ~n5466 & n8851 ) | ( ~n5466 & n12502 ) | ( n8851 & n12502 ) ;
  assign n29366 = n29365 ^ n23419 ^ n2261 ;
  assign n29367 = ~n3891 & n10461 ;
  assign n29368 = n5556 & n29367 ;
  assign n29369 = n25433 & ~n29368 ;
  assign n29370 = ~n2428 & n9414 ;
  assign n29371 = n29370 ^ n18345 ^ 1'b0 ;
  assign n29372 = n28874 & ~n29371 ;
  assign n29373 = n19898 & n29372 ;
  assign n29374 = ( ~n892 & n8119 ) | ( ~n892 & n18657 ) | ( n8119 & n18657 ) ;
  assign n29375 = n14205 ^ n8406 ^ 1'b0 ;
  assign n29376 = n29374 | n29375 ;
  assign n29377 = n10991 ^ n2615 ^ 1'b0 ;
  assign n29378 = n5138 & ~n29377 ;
  assign n29379 = ( ~n9025 & n29376 ) | ( ~n9025 & n29378 ) | ( n29376 & n29378 ) ;
  assign n29382 = n23387 ^ n10945 ^ 1'b0 ;
  assign n29383 = n7490 | n29382 ;
  assign n29380 = ( n6218 & n19429 ) | ( n6218 & ~n21224 ) | ( n19429 & ~n21224 ) ;
  assign n29381 = ( ~n8345 & n11248 ) | ( ~n8345 & n29380 ) | ( n11248 & n29380 ) ;
  assign n29384 = n29383 ^ n29381 ^ n6348 ;
  assign n29385 = n12735 ^ n6178 ^ 1'b0 ;
  assign n29386 = x114 & ~n29385 ;
  assign n29388 = ( n15959 & ~n24540 ) | ( n15959 & n27600 ) | ( ~n24540 & n27600 ) ;
  assign n29387 = n21166 & ~n27091 ;
  assign n29389 = n29388 ^ n29387 ^ 1'b0 ;
  assign n29390 = n7048 & n12795 ;
  assign n29391 = ~n17629 & n29390 ;
  assign n29392 = n29222 & ~n29391 ;
  assign n29393 = n29389 & n29392 ;
  assign n29394 = n19182 ^ n15168 ^ 1'b0 ;
  assign n29395 = n10841 & n24029 ;
  assign n29396 = ~n12190 & n19059 ;
  assign n29397 = n29395 | n29396 ;
  assign n29398 = ( n3343 & ~n16447 ) | ( n3343 & n29397 ) | ( ~n16447 & n29397 ) ;
  assign n29399 = n25909 ^ n13635 ^ n3644 ;
  assign n29400 = n4360 & n19577 ;
  assign n29401 = n8171 & n29400 ;
  assign n29402 = n3689 & ~n14310 ;
  assign n29403 = n18639 ^ n4601 ^ n318 ;
  assign n29404 = ( ~n16802 & n28771 ) | ( ~n16802 & n29403 ) | ( n28771 & n29403 ) ;
  assign n29405 = n1120 | n4455 ;
  assign n29406 = ( ~n3260 & n28458 ) | ( ~n3260 & n29405 ) | ( n28458 & n29405 ) ;
  assign n29407 = ( ~n2575 & n7566 ) | ( ~n2575 & n14138 ) | ( n7566 & n14138 ) ;
  assign n29408 = n7511 & ~n29407 ;
  assign n29409 = n29408 ^ n6863 ^ 1'b0 ;
  assign n29410 = ( n4112 & n21628 ) | ( n4112 & n29409 ) | ( n21628 & n29409 ) ;
  assign n29411 = n29410 ^ n15607 ^ n3996 ;
  assign n29412 = n11070 ^ n450 ^ 1'b0 ;
  assign n29413 = n1605 & ~n29412 ;
  assign n29414 = n3984 ^ n1983 ^ 1'b0 ;
  assign n29415 = n29413 | n29414 ;
  assign n29416 = ( n1573 & ~n3598 ) | ( n1573 & n5034 ) | ( ~n3598 & n5034 ) ;
  assign n29417 = n29416 ^ n9608 ^ n5602 ;
  assign n29418 = n29415 & n29417 ;
  assign n29419 = n15327 & n15879 ;
  assign n29420 = n7943 & n28394 ;
  assign n29421 = n4524 | n8689 ;
  assign n29422 = ~n1810 & n29421 ;
  assign n29423 = n29422 ^ n12130 ^ 1'b0 ;
  assign n29424 = n6808 | n29423 ;
  assign n29425 = n459 & ~n1024 ;
  assign n29426 = n29425 ^ n1664 ^ 1'b0 ;
  assign n29427 = n8019 ^ n1932 ^ 1'b0 ;
  assign n29428 = ~n29426 & n29427 ;
  assign n29429 = ~n7127 & n29428 ;
  assign n29430 = n2153 | n5592 ;
  assign n29431 = n410 & ~n29430 ;
  assign n29432 = ~n3227 & n16500 ;
  assign n29433 = ~n3835 & n29432 ;
  assign n29434 = n29431 & n29433 ;
  assign n29435 = n22973 ^ n14793 ^ 1'b0 ;
  assign n29436 = n3174 & n24361 ;
  assign n29437 = n29436 ^ n23498 ^ 1'b0 ;
  assign n29438 = n19647 & n29437 ;
  assign n29439 = n16993 ^ n627 ^ 1'b0 ;
  assign n29440 = ( n820 & n7261 ) | ( n820 & n29439 ) | ( n7261 & n29439 ) ;
  assign n29442 = n1385 & n4127 ;
  assign n29443 = ~n1358 & n29442 ;
  assign n29444 = n29443 ^ n6428 ^ n1475 ;
  assign n29441 = n22084 | n28277 ;
  assign n29445 = n29444 ^ n29441 ^ 1'b0 ;
  assign n29449 = n1135 & ~n9306 ;
  assign n29450 = n29449 ^ n13806 ^ 1'b0 ;
  assign n29451 = n19099 & n21431 ;
  assign n29452 = n29450 & n29451 ;
  assign n29446 = ( ~n6150 & n9900 ) | ( ~n6150 & n19834 ) | ( n9900 & n19834 ) ;
  assign n29447 = n29446 ^ n7232 ^ 1'b0 ;
  assign n29448 = ~n1051 & n29447 ;
  assign n29453 = n29452 ^ n29448 ^ 1'b0 ;
  assign n29454 = n8685 | n12161 ;
  assign n29455 = n29454 ^ n10777 ^ 1'b0 ;
  assign n29456 = ( n5266 & n25000 ) | ( n5266 & n29455 ) | ( n25000 & n29455 ) ;
  assign n29457 = n2730 ^ n2486 ^ 1'b0 ;
  assign n29458 = n29456 & ~n29457 ;
  assign n29459 = n15129 & n20763 ;
  assign n29460 = n29459 ^ n25769 ^ 1'b0 ;
  assign n29461 = n29460 ^ n15713 ^ 1'b0 ;
  assign n29462 = n7937 | n29461 ;
  assign n29463 = n29462 ^ n6076 ^ 1'b0 ;
  assign n29464 = n14007 & n29463 ;
  assign n29465 = ( n6707 & n8826 ) | ( n6707 & ~n12575 ) | ( n8826 & ~n12575 ) ;
  assign n29466 = n29465 ^ n3504 ^ n2361 ;
  assign n29467 = ( n6342 & n28549 ) | ( n6342 & n29466 ) | ( n28549 & n29466 ) ;
  assign n29468 = n11564 & n28323 ;
  assign n29469 = n8422 | n21412 ;
  assign n29470 = n17079 | n28327 ;
  assign n29471 = n4553 ^ n3796 ^ 1'b0 ;
  assign n29472 = n7227 & ~n29471 ;
  assign n29473 = ( n9966 & ~n12404 ) | ( n9966 & n23040 ) | ( ~n12404 & n23040 ) ;
  assign n29474 = n4257 & n29473 ;
  assign n29475 = ~n21751 & n25661 ;
  assign n29476 = n29475 ^ n18955 ^ 1'b0 ;
  assign n29477 = ( n29472 & n29474 ) | ( n29472 & n29476 ) | ( n29474 & n29476 ) ;
  assign n29478 = n26966 ^ n10617 ^ n3156 ;
  assign n29479 = ( n26188 & n27710 ) | ( n26188 & ~n29478 ) | ( n27710 & ~n29478 ) ;
  assign n29480 = n18619 & ~n29096 ;
  assign n29481 = ~n11342 & n29480 ;
  assign n29482 = n11363 ^ n2767 ^ 1'b0 ;
  assign n29483 = ~n8422 & n29482 ;
  assign n29484 = n5951 & n10007 ;
  assign n29485 = n29484 ^ n4284 ^ 1'b0 ;
  assign n29486 = n29485 ^ n10723 ^ 1'b0 ;
  assign n29487 = n29483 & ~n29486 ;
  assign n29488 = ~n3456 & n17568 ;
  assign n29489 = n29488 ^ n1084 ^ 1'b0 ;
  assign n29490 = n7158 | n29489 ;
  assign n29491 = n20321 & ~n28087 ;
  assign n29492 = n13023 & n29491 ;
  assign n29495 = ~n3264 & n4289 ;
  assign n29496 = n29495 ^ n6124 ^ 1'b0 ;
  assign n29493 = n14620 ^ n2213 ^ 1'b0 ;
  assign n29494 = ~n812 & n29493 ;
  assign n29497 = n29496 ^ n29494 ^ n12163 ;
  assign n29498 = n5965 & n28010 ;
  assign n29499 = n29498 ^ n18061 ^ 1'b0 ;
  assign n29500 = n12894 ^ n8973 ^ 1'b0 ;
  assign n29501 = n1733 & n12487 ;
  assign n29502 = n29501 ^ n25102 ^ n1217 ;
  assign n29503 = n598 | n29502 ;
  assign n29504 = n3518 | n27070 ;
  assign n29505 = n3122 & ~n29504 ;
  assign n29507 = n7983 | n11124 ;
  assign n29508 = n13305 | n29507 ;
  assign n29506 = ~n19893 & n20763 ;
  assign n29509 = n29508 ^ n29506 ^ 1'b0 ;
  assign n29510 = n2442 & n12946 ;
  assign n29511 = n29510 ^ n16831 ^ n4986 ;
  assign n29512 = ( ~n4501 & n5849 ) | ( ~n4501 & n29511 ) | ( n5849 & n29511 ) ;
  assign n29513 = n3994 ^ n659 ^ 1'b0 ;
  assign n29514 = ~n17136 & n29513 ;
  assign n29515 = ( ~n1309 & n8839 ) | ( ~n1309 & n29514 ) | ( n8839 & n29514 ) ;
  assign n29516 = n25552 & ~n29515 ;
  assign n29517 = n29516 ^ n26805 ^ 1'b0 ;
  assign n29518 = ~n2911 & n14518 ;
  assign n29519 = n1211 & n29518 ;
  assign n29520 = n22479 ^ n10018 ^ n2791 ;
  assign n29521 = n4160 & n29520 ;
  assign n29522 = n29519 & n29521 ;
  assign n29523 = n20826 ^ n10229 ^ n9043 ;
  assign n29524 = ( n4916 & n15525 ) | ( n4916 & n23739 ) | ( n15525 & n23739 ) ;
  assign n29525 = ~n10973 & n29524 ;
  assign n29526 = n28947 ^ n4822 ^ x171 ;
  assign n29528 = n272 | n7771 ;
  assign n29529 = n29528 ^ n2124 ^ 1'b0 ;
  assign n29530 = n29529 ^ n3498 ^ 1'b0 ;
  assign n29531 = n6390 & n29530 ;
  assign n29527 = n3974 & n18934 ;
  assign n29532 = n29531 ^ n29527 ^ 1'b0 ;
  assign n29533 = n18928 ^ n8234 ^ 1'b0 ;
  assign n29534 = ( n4749 & ~n14366 ) | ( n4749 & n29533 ) | ( ~n14366 & n29533 ) ;
  assign n29535 = n2004 & n11263 ;
  assign n29536 = n29535 ^ n5166 ^ 1'b0 ;
  assign n29537 = n29534 & ~n29536 ;
  assign n29538 = n29537 ^ n20459 ^ 1'b0 ;
  assign n29539 = n3561 & ~n21194 ;
  assign n29540 = n29539 ^ n3804 ^ 1'b0 ;
  assign n29541 = n19206 ^ n15491 ^ 1'b0 ;
  assign n29542 = n29540 & ~n29541 ;
  assign n29543 = n22333 & ~n27057 ;
  assign n29544 = n29543 ^ n15491 ^ 1'b0 ;
  assign n29545 = x246 & n18668 ;
  assign n29546 = n29545 ^ n657 ^ 1'b0 ;
  assign n29547 = n12229 ^ n9052 ^ n3901 ;
  assign n29548 = ( ~n3061 & n29546 ) | ( ~n3061 & n29547 ) | ( n29546 & n29547 ) ;
  assign n29549 = n29548 ^ n26896 ^ n14308 ;
  assign n29550 = n14133 & n24735 ;
  assign n29551 = n29550 ^ n3358 ^ 1'b0 ;
  assign n29552 = n12076 ^ n262 ^ x110 ;
  assign n29553 = n29552 ^ n22006 ^ 1'b0 ;
  assign n29554 = n3863 & n29553 ;
  assign n29558 = n15214 ^ n2753 ^ 1'b0 ;
  assign n29555 = n8330 ^ n1359 ^ 1'b0 ;
  assign n29556 = ~n3170 & n29555 ;
  assign n29557 = n29556 ^ n1487 ^ 1'b0 ;
  assign n29559 = n29558 ^ n29557 ^ n2791 ;
  assign n29563 = ~n6140 & n22216 ;
  assign n29560 = n13354 ^ n13168 ^ 1'b0 ;
  assign n29561 = n7389 ^ n2630 ^ 1'b0 ;
  assign n29562 = n29560 | n29561 ;
  assign n29564 = n29563 ^ n29562 ^ 1'b0 ;
  assign n29565 = n15029 & ~n18961 ;
  assign n29566 = ~n16035 & n29565 ;
  assign n29571 = n17351 ^ n12478 ^ 1'b0 ;
  assign n29567 = n4481 | n18449 ;
  assign n29568 = n4053 & ~n29567 ;
  assign n29569 = n1643 | n29568 ;
  assign n29570 = n29569 ^ n24182 ^ 1'b0 ;
  assign n29572 = n29571 ^ n29570 ^ 1'b0 ;
  assign n29573 = n29566 | n29572 ;
  assign n29574 = ( n9160 & n12612 ) | ( n9160 & ~n29573 ) | ( n12612 & ~n29573 ) ;
  assign n29575 = n18751 ^ n17120 ^ n9521 ;
  assign n29576 = ( n5819 & n7920 ) | ( n5819 & n14715 ) | ( n7920 & n14715 ) ;
  assign n29577 = n29576 ^ n8873 ^ n5126 ;
  assign n29578 = n29577 ^ n27028 ^ 1'b0 ;
  assign n29579 = n5789 ^ n2705 ^ 1'b0 ;
  assign n29580 = ( n8902 & n15989 ) | ( n8902 & n29579 ) | ( n15989 & n29579 ) ;
  assign n29581 = n25751 ^ n3027 ^ 1'b0 ;
  assign n29582 = n29580 & ~n29581 ;
  assign n29583 = n24383 ^ n11343 ^ n8919 ;
  assign n29584 = n9298 | n29583 ;
  assign n29585 = n4346 & ~n29584 ;
  assign n29586 = ( ~n4089 & n8780 ) | ( ~n4089 & n20548 ) | ( n8780 & n20548 ) ;
  assign n29587 = ~n19005 & n29586 ;
  assign n29588 = n9341 ^ n8566 ^ 1'b0 ;
  assign n29589 = n2957 & ~n29588 ;
  assign n29590 = n29589 ^ n574 ^ 1'b0 ;
  assign n29591 = ~n29587 & n29590 ;
  assign n29596 = n10997 ^ n3331 ^ 1'b0 ;
  assign n29592 = n1924 & ~n6721 ;
  assign n29593 = n29592 ^ n3902 ^ 1'b0 ;
  assign n29594 = n1346 | n29593 ;
  assign n29595 = n29594 ^ n3787 ^ 1'b0 ;
  assign n29597 = n29596 ^ n29595 ^ 1'b0 ;
  assign n29598 = ( n3281 & ~n13531 ) | ( n3281 & n21382 ) | ( ~n13531 & n21382 ) ;
  assign n29599 = n12121 | n18208 ;
  assign n29600 = n13391 & n29599 ;
  assign n29601 = ~n29598 & n29600 ;
  assign n29602 = n12118 | n26556 ;
  assign n29605 = n3074 | n6372 ;
  assign n29606 = n4061 & n29605 ;
  assign n29607 = ~n14613 & n29606 ;
  assign n29603 = n6242 & ~n26986 ;
  assign n29604 = n19223 & n29603 ;
  assign n29608 = n29607 ^ n29604 ^ n16727 ;
  assign n29609 = ( n2666 & n18388 ) | ( n2666 & n23593 ) | ( n18388 & n23593 ) ;
  assign n29610 = ( n357 & ~n19431 ) | ( n357 & n29593 ) | ( ~n19431 & n29593 ) ;
  assign n29611 = n13907 ^ n10098 ^ 1'b0 ;
  assign n29612 = n24476 | n29611 ;
  assign n29613 = ~n6480 & n29612 ;
  assign n29614 = n24444 ^ n20063 ^ n2638 ;
  assign n29615 = n6523 | n10396 ;
  assign n29616 = n14848 | n29615 ;
  assign n29617 = n29616 ^ n5183 ^ 1'b0 ;
  assign n29618 = n11898 ^ n10595 ^ n8070 ;
  assign n29619 = ~n18920 & n29618 ;
  assign n29620 = ~n26631 & n29619 ;
  assign n29621 = n23929 ^ n8734 ^ n2410 ;
  assign n29622 = ( n6574 & n15794 ) | ( n6574 & n29621 ) | ( n15794 & n29621 ) ;
  assign n29623 = n24443 ^ n22586 ^ n11323 ;
  assign n29624 = n12312 | n13352 ;
  assign n29625 = n29624 ^ n15348 ^ 1'b0 ;
  assign n29626 = n3502 & n29625 ;
  assign n29627 = n23564 ^ n7252 ^ x47 ;
  assign n29628 = n15717 & n29627 ;
  assign n29629 = n26833 ^ n2247 ^ 1'b0 ;
  assign n29630 = n22398 & ~n29629 ;
  assign n29631 = n29630 ^ n27498 ^ 1'b0 ;
  assign n29632 = n29628 | n29631 ;
  assign n29633 = x119 & n20015 ;
  assign n29634 = n29633 ^ n2447 ^ 1'b0 ;
  assign n29635 = n5458 & ~n11165 ;
  assign n29636 = ~n29634 & n29635 ;
  assign n29637 = n18664 ^ n12459 ^ 1'b0 ;
  assign n29638 = n29636 | n29637 ;
  assign n29639 = n16023 | n17439 ;
  assign n29640 = n29249 | n29639 ;
  assign n29641 = x91 & ~n423 ;
  assign n29642 = ~n2456 & n29641 ;
  assign n29643 = n8747 ^ n5506 ^ n3814 ;
  assign n29644 = ( n11543 & n29642 ) | ( n11543 & n29643 ) | ( n29642 & n29643 ) ;
  assign n29647 = ~n6952 & n7257 ;
  assign n29646 = n20782 ^ n7217 ^ 1'b0 ;
  assign n29645 = n19628 ^ n15116 ^ n5733 ;
  assign n29648 = n29647 ^ n29646 ^ n29645 ;
  assign n29649 = n5523 & n7206 ;
  assign n29650 = n28440 ^ n27012 ^ n5642 ;
  assign n29651 = n7363 ^ n1006 ^ 1'b0 ;
  assign n29652 = n1066 | n29651 ;
  assign n29653 = n20814 ^ n15835 ^ 1'b0 ;
  assign n29654 = n29652 | n29653 ;
  assign n29655 = ~n861 & n5949 ;
  assign n29656 = n29655 ^ n25465 ^ 1'b0 ;
  assign n29657 = n29654 | n29656 ;
  assign n29658 = n11357 | n29657 ;
  assign n29659 = n29658 ^ n26900 ^ 1'b0 ;
  assign n29660 = ~n5754 & n25405 ;
  assign n29661 = n6090 | n22206 ;
  assign n29662 = ( n9658 & ~n29660 ) | ( n9658 & n29661 ) | ( ~n29660 & n29661 ) ;
  assign n29663 = n12766 ^ n1061 ^ 1'b0 ;
  assign n29664 = n16289 | n29663 ;
  assign n29665 = n3460 & ~n29664 ;
  assign n29666 = ~n3127 & n29665 ;
  assign n29667 = ~n930 & n2131 ;
  assign n29668 = n29667 ^ n14789 ^ 1'b0 ;
  assign n29669 = ( n1307 & n4253 ) | ( n1307 & ~n5833 ) | ( n4253 & ~n5833 ) ;
  assign n29670 = n29669 ^ n18440 ^ n12766 ;
  assign n29671 = n16789 ^ n8842 ^ n4023 ;
  assign n29672 = n5026 | n16327 ;
  assign n29673 = ( n16883 & n25228 ) | ( n16883 & n29672 ) | ( n25228 & n29672 ) ;
  assign n29674 = n5322 & n18721 ;
  assign n29675 = n25171 ^ n16547 ^ n8159 ;
  assign n29676 = ( ~n2847 & n29674 ) | ( ~n2847 & n29675 ) | ( n29674 & n29675 ) ;
  assign n29677 = n7364 ^ x110 ^ 1'b0 ;
  assign n29678 = n7478 & ~n29677 ;
  assign n29679 = n28775 & n29678 ;
  assign n29680 = n29679 ^ n22302 ^ 1'b0 ;
  assign n29681 = ( ~n5130 & n12383 ) | ( ~n5130 & n15868 ) | ( n12383 & n15868 ) ;
  assign n29682 = n4318 & n29681 ;
  assign n29683 = n29680 & n29682 ;
  assign n29684 = n4206 ^ n2295 ^ 1'b0 ;
  assign n29685 = n21798 & n29684 ;
  assign n29686 = ~n14193 & n29685 ;
  assign n29687 = n4674 | n29686 ;
  assign n29688 = n29687 ^ n4060 ^ 1'b0 ;
  assign n29689 = n5003 & n11546 ;
  assign n29690 = ~n29688 & n29689 ;
  assign n29691 = ( n523 & n12429 ) | ( n523 & n29690 ) | ( n12429 & n29690 ) ;
  assign n29692 = n29691 ^ n17064 ^ n3465 ;
  assign n29693 = n3012 | n13571 ;
  assign n29694 = n29693 ^ n17635 ^ n2225 ;
  assign n29695 = n17933 ^ n12546 ^ 1'b0 ;
  assign n29696 = ~n1526 & n9654 ;
  assign n29697 = ( n20012 & n29053 ) | ( n20012 & n29696 ) | ( n29053 & n29696 ) ;
  assign n29698 = n28074 ^ n16600 ^ x129 ;
  assign n29699 = n14634 & ~n15314 ;
  assign n29700 = n29699 ^ n27283 ^ 1'b0 ;
  assign n29701 = n15828 | n29700 ;
  assign n29702 = n6229 ^ n2548 ^ 1'b0 ;
  assign n29703 = ~n3462 & n29702 ;
  assign n29704 = ~n10776 & n26944 ;
  assign n29705 = ~n29703 & n29704 ;
  assign n29707 = n2303 ^ n2225 ^ 1'b0 ;
  assign n29708 = ~n9018 & n29707 ;
  assign n29709 = n29708 ^ n7513 ^ n2822 ;
  assign n29706 = n9150 & ~n9997 ;
  assign n29710 = n29709 ^ n29706 ^ 1'b0 ;
  assign n29711 = n29710 ^ n24792 ^ 1'b0 ;
  assign n29714 = ( n5504 & n10976 ) | ( n5504 & n15187 ) | ( n10976 & n15187 ) ;
  assign n29712 = n8067 ^ n392 ^ 1'b0 ;
  assign n29713 = n6096 & n29712 ;
  assign n29715 = n29714 ^ n29713 ^ n6258 ;
  assign n29716 = n17014 ^ n6823 ^ 1'b0 ;
  assign n29717 = n18457 ^ n1889 ^ 1'b0 ;
  assign n29718 = n5816 & ~n21105 ;
  assign n29719 = n16685 ^ n13474 ^ n4646 ;
  assign n29720 = ( n4072 & n9956 ) | ( n4072 & ~n29719 ) | ( n9956 & ~n29719 ) ;
  assign n29721 = ~n11091 & n18795 ;
  assign n29722 = ( n5294 & n14430 ) | ( n5294 & ~n21274 ) | ( n14430 & ~n21274 ) ;
  assign n29723 = n7500 | n29707 ;
  assign n29724 = ~n12554 & n27086 ;
  assign n29725 = n1039 & n29724 ;
  assign n29726 = n6146 ^ n734 ^ 1'b0 ;
  assign n29727 = n29726 ^ n18672 ^ n1681 ;
  assign n29728 = ~n15919 & n29727 ;
  assign n29729 = n18638 & n29728 ;
  assign n29730 = n20379 ^ n3147 ^ 1'b0 ;
  assign n29731 = n340 | n7300 ;
  assign n29732 = n29731 ^ n7108 ^ 1'b0 ;
  assign n29733 = n29732 ^ n24461 ^ 1'b0 ;
  assign n29734 = ( n3829 & n4949 ) | ( n3829 & ~n13039 ) | ( n4949 & ~n13039 ) ;
  assign n29735 = n20321 & n29734 ;
  assign n29736 = n7518 & ~n24919 ;
  assign n29737 = ~n23073 & n29736 ;
  assign n29738 = n15362 ^ n9398 ^ n6150 ;
  assign n29739 = n29738 ^ n20655 ^ 1'b0 ;
  assign n29740 = ~n17431 & n29739 ;
  assign n29741 = n6586 & n13478 ;
  assign n29743 = n15627 ^ n6966 ^ 1'b0 ;
  assign n29742 = n9387 | n16427 ;
  assign n29744 = n29743 ^ n29742 ^ 1'b0 ;
  assign n29745 = n6427 & ~n12780 ;
  assign n29746 = n3511 | n7187 ;
  assign n29747 = n12221 & ~n29746 ;
  assign n29748 = ( ~n7372 & n9072 ) | ( ~n7372 & n10315 ) | ( n9072 & n10315 ) ;
  assign n29749 = n29748 ^ n21866 ^ 1'b0 ;
  assign n29750 = n22238 | n29749 ;
  assign n29751 = n5923 & n18862 ;
  assign n29752 = n656 & n3566 ;
  assign n29753 = ~n3583 & n29752 ;
  assign n29754 = n19373 ^ n12038 ^ 1'b0 ;
  assign n29755 = ~n29753 & n29754 ;
  assign n29756 = ( ~n2171 & n18847 ) | ( ~n2171 & n29050 ) | ( n18847 & n29050 ) ;
  assign n29757 = n1454 & n20333 ;
  assign n29758 = n27654 ^ n17154 ^ 1'b0 ;
  assign n29759 = n5277 | n12461 ;
  assign n29760 = n2365 | n29759 ;
  assign n29761 = n1977 | n29760 ;
  assign n29762 = ( n8870 & ~n18378 ) | ( n8870 & n29761 ) | ( ~n18378 & n29761 ) ;
  assign n29763 = n29359 ^ n2321 ^ 1'b0 ;
  assign n29764 = n25854 ^ n22488 ^ 1'b0 ;
  assign n29765 = n15112 ^ n7087 ^ n3029 ;
  assign n29766 = ~n15989 & n29765 ;
  assign n29767 = n12274 | n29766 ;
  assign n29768 = n11449 | n14297 ;
  assign n29769 = n9113 | n17932 ;
  assign n29770 = n29769 ^ n7959 ^ 1'b0 ;
  assign n29771 = ~n29768 & n29770 ;
  assign n29772 = n5135 ^ n1035 ^ 1'b0 ;
  assign n29773 = n3493 & n29772 ;
  assign n29774 = ~n4244 & n29773 ;
  assign n29775 = ~n8984 & n29774 ;
  assign n29776 = ~n8990 & n24916 ;
  assign n29777 = n29776 ^ n11568 ^ 1'b0 ;
  assign n29778 = n24894 ^ n12699 ^ n9182 ;
  assign n29779 = n21927 | n29778 ;
  assign n29780 = n15173 | n29779 ;
  assign n29781 = n29780 ^ n25342 ^ n2036 ;
  assign n29782 = n5990 & n20182 ;
  assign n29783 = ( ~x95 & n20285 ) | ( ~x95 & n29782 ) | ( n20285 & n29782 ) ;
  assign n29784 = n4749 | n23716 ;
  assign n29785 = n9544 & n17812 ;
  assign n29786 = ~n29784 & n29785 ;
  assign n29787 = n9994 ^ n3101 ^ 1'b0 ;
  assign n29788 = n24150 ^ n15551 ^ n5100 ;
  assign n29789 = ( n23913 & ~n29787 ) | ( n23913 & n29788 ) | ( ~n29787 & n29788 ) ;
  assign n29790 = n11536 | n29789 ;
  assign n29791 = n29790 ^ n16810 ^ 1'b0 ;
  assign n29792 = ~n9076 & n23301 ;
  assign n29793 = n5718 & n29792 ;
  assign n29794 = ~n29791 & n29793 ;
  assign n29795 = n23457 & n27028 ;
  assign n29796 = n6546 | n29795 ;
  assign n29797 = n27365 ^ n17761 ^ n3301 ;
  assign n29798 = n1191 & n14318 ;
  assign n29799 = n29798 ^ n4117 ^ 1'b0 ;
  assign n29800 = n444 & n6148 ;
  assign n29801 = ~n444 & n29800 ;
  assign n29802 = ~n2208 & n9482 ;
  assign n29803 = n2208 & n29802 ;
  assign n29804 = n29801 | n29803 ;
  assign n29805 = n29804 ^ n10233 ^ 1'b0 ;
  assign n29806 = n18442 & n29805 ;
  assign n29807 = ~n29799 & n29806 ;
  assign n29808 = n29807 ^ n21424 ^ n9003 ;
  assign n29809 = ( n503 & n1401 ) | ( n503 & n10644 ) | ( n1401 & n10644 ) ;
  assign n29810 = n8657 | n29809 ;
  assign n29811 = n21963 | n29810 ;
  assign n29812 = n20303 ^ x11 ^ 1'b0 ;
  assign n29813 = n14283 | n29812 ;
  assign n29814 = ~n916 & n10133 ;
  assign n29815 = n29814 ^ n9591 ^ 1'b0 ;
  assign n29816 = n18911 & ~n29815 ;
  assign n29817 = ~n21001 & n29816 ;
  assign n29818 = n18873 ^ n5839 ^ 1'b0 ;
  assign n29824 = n14617 ^ n6832 ^ n392 ;
  assign n29825 = n29824 ^ n16294 ^ n9472 ;
  assign n29819 = n2319 | n7920 ;
  assign n29820 = n29819 ^ n8484 ^ 1'b0 ;
  assign n29821 = ~n742 & n27614 ;
  assign n29822 = n409 & n29821 ;
  assign n29823 = n29820 | n29822 ;
  assign n29826 = n29825 ^ n29823 ^ 1'b0 ;
  assign n29827 = n1998 | n11476 ;
  assign n29828 = n29827 ^ n4497 ^ 1'b0 ;
  assign n29829 = ( ~x54 & n5509 ) | ( ~x54 & n29828 ) | ( n5509 & n29828 ) ;
  assign n29830 = ~n9894 & n21236 ;
  assign n29831 = ~n9691 & n29830 ;
  assign n29832 = n20717 ^ n5514 ^ n1374 ;
  assign n29833 = n29832 ^ n14226 ^ n8450 ;
  assign n29834 = n12426 & ~n29833 ;
  assign n29835 = n6005 & n29834 ;
  assign n29836 = n29835 ^ n14001 ^ n6169 ;
  assign n29837 = ( n23017 & n29831 ) | ( n23017 & n29836 ) | ( n29831 & n29836 ) ;
  assign n29838 = n1075 & n29837 ;
  assign n29840 = n29784 ^ n10243 ^ 1'b0 ;
  assign n29839 = n22881 ^ n15161 ^ n2156 ;
  assign n29841 = n29840 ^ n29839 ^ n27452 ;
  assign n29842 = n7172 ^ n4705 ^ n3680 ;
  assign n29843 = n13674 | n29842 ;
  assign n29844 = n23564 & ~n29843 ;
  assign n29845 = n8898 & n17830 ;
  assign n29846 = n29844 & n29845 ;
  assign n29847 = ~n11035 & n13764 ;
  assign n29848 = n7862 ^ n6907 ^ 1'b0 ;
  assign n29849 = ( n14790 & ~n20358 ) | ( n14790 & n29848 ) | ( ~n20358 & n29848 ) ;
  assign n29850 = n29849 ^ n21890 ^ n11995 ;
  assign n29851 = n23608 ^ n15654 ^ n11244 ;
  assign n29852 = ~n17077 & n22492 ;
  assign n29853 = n29851 & n29852 ;
  assign n29854 = n15348 ^ n12106 ^ 1'b0 ;
  assign n29855 = ( n17908 & n19446 ) | ( n17908 & n23910 ) | ( n19446 & n23910 ) ;
  assign n29860 = n8510 & n12356 ;
  assign n29857 = n16300 ^ n8506 ^ 1'b0 ;
  assign n29858 = n1533 & n29857 ;
  assign n29859 = n29858 ^ n24052 ^ n3442 ;
  assign n29856 = n24963 ^ n1294 ^ 1'b0 ;
  assign n29861 = n29860 ^ n29859 ^ n29856 ;
  assign n29862 = n12947 | n16214 ;
  assign n29863 = n12265 & ~n29862 ;
  assign n29864 = n29863 ^ n13660 ^ n8050 ;
  assign n29865 = n18061 | n29864 ;
  assign n29866 = n5216 & ~n18103 ;
  assign n29867 = ~n15174 & n29866 ;
  assign n29868 = n29867 ^ n16473 ^ n13052 ;
  assign n29869 = ~n9298 & n29868 ;
  assign n29870 = n29869 ^ n3200 ^ 1'b0 ;
  assign n29871 = n13145 ^ n11816 ^ n543 ;
  assign n29872 = n24844 ^ n23909 ^ 1'b0 ;
  assign n29873 = n27015 | n29872 ;
  assign n29874 = n29871 | n29873 ;
  assign n29875 = ~n16325 & n29874 ;
  assign n29876 = ~n23642 & n26681 ;
  assign n29877 = n2812 & ~n19182 ;
  assign n29878 = ~n14341 & n29877 ;
  assign n29879 = n28057 ^ n19957 ^ n7107 ;
  assign n29880 = n8309 & ~n10657 ;
  assign n29881 = n4272 ^ n1149 ^ 1'b0 ;
  assign n29882 = n21698 ^ n5950 ^ 1'b0 ;
  assign n29883 = n7420 | n29882 ;
  assign n29884 = ( ~n979 & n2824 ) | ( ~n979 & n14214 ) | ( n2824 & n14214 ) ;
  assign n29885 = ( ~n10623 & n25819 ) | ( ~n10623 & n29884 ) | ( n25819 & n29884 ) ;
  assign n29886 = n20731 ^ n19463 ^ 1'b0 ;
  assign n29887 = n10239 ^ n3550 ^ 1'b0 ;
  assign n29888 = n10209 ^ n7496 ^ 1'b0 ;
  assign n29889 = n29887 | n29888 ;
  assign n29890 = n1943 | n3254 ;
  assign n29891 = n29890 ^ n6472 ^ 1'b0 ;
  assign n29892 = ( n15776 & ~n26797 ) | ( n15776 & n29891 ) | ( ~n26797 & n29891 ) ;
  assign n29893 = n21494 & ~n26711 ;
  assign n29894 = n29893 ^ n14485 ^ 1'b0 ;
  assign n29895 = n24324 | n29894 ;
  assign n29897 = n9016 ^ n5357 ^ 1'b0 ;
  assign n29898 = ~n2124 & n29897 ;
  assign n29896 = n29070 ^ n3275 ^ 1'b0 ;
  assign n29899 = n29898 ^ n29896 ^ n3600 ;
  assign n29900 = n20160 ^ n6163 ^ 1'b0 ;
  assign n29901 = ~n9322 & n29900 ;
  assign n29902 = n29901 ^ x108 ^ 1'b0 ;
  assign n29903 = n29902 ^ n27302 ^ 1'b0 ;
  assign n29904 = n29899 & ~n29903 ;
  assign n29905 = n28104 ^ n9184 ^ 1'b0 ;
  assign n29906 = n12837 | n29905 ;
  assign n29907 = n29906 ^ n15249 ^ n1726 ;
  assign n29908 = n14457 ^ n5791 ^ n352 ;
  assign n29909 = ( n10223 & ~n10433 ) | ( n10223 & n29908 ) | ( ~n10433 & n29908 ) ;
  assign n29910 = n11138 ^ n8352 ^ n1279 ;
  assign n29911 = n29910 ^ n25284 ^ n8201 ;
  assign n29912 = n29911 ^ n12668 ^ 1'b0 ;
  assign n29913 = n15902 & ~n29912 ;
  assign n29914 = ( n6478 & ~n14180 ) | ( n6478 & n20305 ) | ( ~n14180 & n20305 ) ;
  assign n29915 = n29914 ^ n5285 ^ n1315 ;
  assign n29916 = n29915 ^ n12081 ^ 1'b0 ;
  assign n29917 = n9023 | n29916 ;
  assign n29918 = n17109 ^ n3753 ^ 1'b0 ;
  assign n29919 = n3675 | n29918 ;
  assign n29920 = n19030 & n29919 ;
  assign n29926 = n5368 & ~n10930 ;
  assign n29927 = n29926 ^ n9792 ^ 1'b0 ;
  assign n29921 = n26609 ^ n12467 ^ 1'b0 ;
  assign n29922 = ( ~n7725 & n24684 ) | ( ~n7725 & n29921 ) | ( n24684 & n29921 ) ;
  assign n29923 = n21759 & ~n29922 ;
  assign n29924 = ~n20668 & n29923 ;
  assign n29925 = n29924 ^ n3378 ^ 1'b0 ;
  assign n29928 = n29927 ^ n29925 ^ n21538 ;
  assign n29929 = n20438 ^ n17205 ^ 1'b0 ;
  assign n29930 = n29245 ^ n14847 ^ 1'b0 ;
  assign n29931 = ( n28014 & n29929 ) | ( n28014 & n29930 ) | ( n29929 & n29930 ) ;
  assign n29932 = n8567 & n15728 ;
  assign n29933 = n29932 ^ n22812 ^ n14443 ;
  assign n29934 = n29933 ^ n18571 ^ n18191 ;
  assign n29935 = n4363 & ~n25596 ;
  assign n29936 = ~n10970 & n29935 ;
  assign n29941 = n17847 | n18777 ;
  assign n29938 = n3909 | n15753 ;
  assign n29939 = n9452 & ~n29938 ;
  assign n29937 = n23901 ^ n23075 ^ n334 ;
  assign n29940 = n29939 ^ n29937 ^ n16504 ;
  assign n29942 = n29941 ^ n29940 ^ 1'b0 ;
  assign n29943 = ( n10684 & n21943 ) | ( n10684 & n29643 ) | ( n21943 & n29643 ) ;
  assign n29944 = n21189 & ~n29943 ;
  assign n29945 = n22353 & n29944 ;
  assign n29946 = n3611 & ~n16058 ;
  assign n29947 = n27457 & ~n29946 ;
  assign n29948 = n29947 ^ n5494 ^ 1'b0 ;
  assign n29949 = n7300 ^ n4202 ^ 1'b0 ;
  assign n29950 = n27724 ^ n15675 ^ 1'b0 ;
  assign n29951 = n29949 & n29950 ;
  assign n29952 = n23074 ^ n10489 ^ n4198 ;
  assign n29953 = n21470 ^ n13929 ^ 1'b0 ;
  assign n29954 = ~n2216 & n29953 ;
  assign n29955 = ( x199 & n28384 ) | ( x199 & n29954 ) | ( n28384 & n29954 ) ;
  assign n29958 = n5674 & n11345 ;
  assign n29959 = ~n9141 & n29958 ;
  assign n29956 = n13932 ^ n1482 ^ 1'b0 ;
  assign n29957 = ~n9546 & n29956 ;
  assign n29960 = n29959 ^ n29957 ^ 1'b0 ;
  assign n29961 = n19368 ^ n18253 ^ 1'b0 ;
  assign n29962 = ( ~n16754 & n18284 ) | ( ~n16754 & n29961 ) | ( n18284 & n29961 ) ;
  assign n29963 = ~n2061 & n29765 ;
  assign n29965 = n5462 ^ n2457 ^ 1'b0 ;
  assign n29964 = n3652 & ~n6687 ;
  assign n29966 = n29965 ^ n29964 ^ 1'b0 ;
  assign n29967 = n10109 & ~n29966 ;
  assign n29968 = n29963 & n29967 ;
  assign n29969 = n7905 | n19706 ;
  assign n29970 = ~n12542 & n29969 ;
  assign n29977 = n21077 ^ n16136 ^ n2687 ;
  assign n29974 = n4856 & ~n13359 ;
  assign n29975 = ~n20545 & n29974 ;
  assign n29976 = n29975 ^ n8133 ^ 1'b0 ;
  assign n29971 = n9902 ^ n2470 ^ 1'b0 ;
  assign n29972 = n8637 ^ n4552 ^ 1'b0 ;
  assign n29973 = ( n13873 & n29971 ) | ( n13873 & n29972 ) | ( n29971 & n29972 ) ;
  assign n29978 = n29977 ^ n29976 ^ n29973 ;
  assign n29979 = n2684 | n3148 ;
  assign n29980 = n26339 | n29979 ;
  assign n29981 = n8210 & n22473 ;
  assign n29982 = ( n10091 & n18770 ) | ( n10091 & ~n27176 ) | ( n18770 & ~n27176 ) ;
  assign n29983 = ( n2558 & n8133 ) | ( n2558 & ~n11108 ) | ( n8133 & ~n11108 ) ;
  assign n29984 = n8423 | n29983 ;
  assign n29985 = n29984 ^ n11539 ^ 1'b0 ;
  assign n29986 = n18682 ^ n2691 ^ x43 ;
  assign n29987 = ~n23589 & n29986 ;
  assign n29988 = n4466 & n29987 ;
  assign n29989 = ( ~n5722 & n29985 ) | ( ~n5722 & n29988 ) | ( n29985 & n29988 ) ;
  assign n29990 = ~n23001 & n28506 ;
  assign n29991 = n29990 ^ n8282 ^ 1'b0 ;
  assign n29992 = n9857 ^ n7163 ^ 1'b0 ;
  assign n29993 = n19089 ^ n17611 ^ n10926 ;
  assign n29994 = n17465 ^ n3063 ^ 1'b0 ;
  assign n29995 = n10324 ^ n9116 ^ 1'b0 ;
  assign n29996 = ( n3502 & n29994 ) | ( n3502 & ~n29995 ) | ( n29994 & ~n29995 ) ;
  assign n29997 = n15838 & n22662 ;
  assign n29998 = ( ~n16542 & n20410 ) | ( ~n16542 & n23289 ) | ( n20410 & n23289 ) ;
  assign n30002 = n12351 & ~n21944 ;
  assign n30003 = ( n6048 & n9662 ) | ( n6048 & n30002 ) | ( n9662 & n30002 ) ;
  assign n29999 = n5221 & n10822 ;
  assign n30000 = ~n27669 & n29999 ;
  assign n30001 = n30000 ^ n17733 ^ n739 ;
  assign n30004 = n30003 ^ n30001 ^ 1'b0 ;
  assign n30005 = n2620 & n7602 ;
  assign n30006 = n30005 ^ n16348 ^ 1'b0 ;
  assign n30007 = n30006 ^ n8336 ^ 1'b0 ;
  assign n30008 = ~n2741 & n13822 ;
  assign n30009 = n30008 ^ n12270 ^ 1'b0 ;
  assign n30010 = n12000 & ~n30009 ;
  assign n30011 = n30010 ^ n14973 ^ n10281 ;
  assign n30012 = n22571 ^ n20858 ^ n14233 ;
  assign n30013 = ( ~n11564 & n12181 ) | ( ~n11564 & n14564 ) | ( n12181 & n14564 ) ;
  assign n30014 = n722 & n1871 ;
  assign n30016 = n14833 ^ n5044 ^ n1854 ;
  assign n30015 = n26853 ^ n23783 ^ n10502 ;
  assign n30017 = n30016 ^ n30015 ^ 1'b0 ;
  assign n30018 = ( n20161 & ~n23636 ) | ( n20161 & n28307 ) | ( ~n23636 & n28307 ) ;
  assign n30019 = ( n1916 & ~n4147 ) | ( n1916 & n27246 ) | ( ~n4147 & n27246 ) ;
  assign n30020 = n6463 & ~n7649 ;
  assign n30021 = n26560 ^ n11734 ^ 1'b0 ;
  assign n30022 = n30020 | n30021 ;
  assign n30023 = x84 & n30022 ;
  assign n30024 = ( n4255 & n30019 ) | ( n4255 & n30023 ) | ( n30019 & n30023 ) ;
  assign n30025 = x58 & n13870 ;
  assign n30026 = ( ~x154 & n742 ) | ( ~x154 & n7916 ) | ( n742 & n7916 ) ;
  assign n30027 = n30026 ^ n9938 ^ 1'b0 ;
  assign n30028 = n23703 & ~n30027 ;
  assign n30029 = ~n2525 & n30028 ;
  assign n30030 = n30029 ^ n26753 ^ 1'b0 ;
  assign n30031 = n8904 & ~n30030 ;
  assign n30032 = n30031 ^ n10290 ^ 1'b0 ;
  assign n30033 = n30025 & ~n30032 ;
  assign n30034 = n7999 | n25697 ;
  assign n30035 = n11384 ^ n932 ^ 1'b0 ;
  assign n30036 = n21335 ^ n18040 ^ n17734 ;
  assign n30037 = ( n1736 & n13522 ) | ( n1736 & ~n24120 ) | ( n13522 & ~n24120 ) ;
  assign n30038 = n9568 | n30037 ;
  assign n30039 = n27392 ^ n20487 ^ n17529 ;
  assign n30040 = ( ~n9634 & n18667 ) | ( ~n9634 & n28565 ) | ( n18667 & n28565 ) ;
  assign n30041 = n30040 ^ n7421 ^ n3264 ;
  assign n30042 = n6414 & ~n22878 ;
  assign n30043 = n30042 ^ n16900 ^ n10695 ;
  assign n30045 = ~n8635 & n11820 ;
  assign n30046 = n4171 & n30045 ;
  assign n30044 = n645 | n5493 ;
  assign n30047 = n30046 ^ n30044 ^ n24150 ;
  assign n30050 = n6740 ^ n6622 ^ n952 ;
  assign n30051 = n30050 ^ n17291 ^ 1'b0 ;
  assign n30052 = n1874 & ~n30051 ;
  assign n30053 = n30052 ^ n15927 ^ n1643 ;
  assign n30054 = n29616 & n30053 ;
  assign n30055 = n17626 & n30054 ;
  assign n30048 = n9754 ^ n8730 ^ n4036 ;
  assign n30049 = ( n7622 & n15485 ) | ( n7622 & ~n30048 ) | ( n15485 & ~n30048 ) ;
  assign n30056 = n30055 ^ n30049 ^ 1'b0 ;
  assign n30057 = ~n13521 & n16512 ;
  assign n30058 = n30057 ^ n18462 ^ 1'b0 ;
  assign n30059 = n30058 ^ n5452 ^ n4239 ;
  assign n30060 = n7797 ^ n4741 ^ 1'b0 ;
  assign n30061 = ( n6156 & n14244 ) | ( n6156 & n21983 ) | ( n14244 & n21983 ) ;
  assign n30062 = n15720 ^ n14624 ^ n13833 ;
  assign n30063 = n30062 ^ n18054 ^ n10405 ;
  assign n30064 = n22003 ^ n3309 ^ 1'b0 ;
  assign n30065 = ~n12591 & n15779 ;
  assign n30066 = n30065 ^ n14370 ^ 1'b0 ;
  assign n30067 = n3140 & n3999 ;
  assign n30068 = n12566 & n30067 ;
  assign n30069 = n30068 ^ n7412 ^ 1'b0 ;
  assign n30070 = x112 & n30069 ;
  assign n30071 = n17678 ^ n11332 ^ 1'b0 ;
  assign n30072 = ~n21711 & n30071 ;
  assign n30073 = n30072 ^ n22172 ^ n21141 ;
  assign n30076 = n3226 ^ n2999 ^ 1'b0 ;
  assign n30077 = n8465 | n30076 ;
  assign n30078 = n3722 | n30077 ;
  assign n30079 = n30078 ^ n9056 ^ 1'b0 ;
  assign n30080 = n30079 ^ n10274 ^ 1'b0 ;
  assign n30074 = n3888 ^ x179 ^ 1'b0 ;
  assign n30075 = ~n23440 & n30074 ;
  assign n30081 = n30080 ^ n30075 ^ 1'b0 ;
  assign n30082 = n6666 | n16605 ;
  assign n30083 = n28816 ^ n4446 ^ 1'b0 ;
  assign n30084 = ~n15566 & n30083 ;
  assign n30085 = n30084 ^ n14771 ^ 1'b0 ;
  assign n30086 = n4627 & n30085 ;
  assign n30087 = n17800 ^ n16789 ^ 1'b0 ;
  assign n30088 = n17079 | n30087 ;
  assign n30089 = n30086 & ~n30088 ;
  assign n30090 = n30089 ^ n29301 ^ 1'b0 ;
  assign n30091 = n524 & ~n7642 ;
  assign n30092 = n30091 ^ n1290 ^ 1'b0 ;
  assign n30093 = n25917 ^ n5770 ^ 1'b0 ;
  assign n30094 = ( n544 & n22050 ) | ( n544 & n30093 ) | ( n22050 & n30093 ) ;
  assign n30095 = n11116 ^ n9499 ^ 1'b0 ;
  assign n30096 = n2008 & n30095 ;
  assign n30097 = ( n16054 & n23386 ) | ( n16054 & n30096 ) | ( n23386 & n30096 ) ;
  assign n30098 = n17818 ^ n5872 ^ 1'b0 ;
  assign n30099 = n24520 | n30098 ;
  assign n30100 = n8838 & n15685 ;
  assign n30101 = n30100 ^ n9255 ^ 1'b0 ;
  assign n30102 = n30101 ^ n5126 ^ 1'b0 ;
  assign n30103 = n11891 ^ n7750 ^ n3713 ;
  assign n30104 = ( ~x114 & n3629 ) | ( ~x114 & n30103 ) | ( n3629 & n30103 ) ;
  assign n30106 = ~n18929 & n27669 ;
  assign n30107 = n30106 ^ n1635 ^ 1'b0 ;
  assign n30105 = n8335 | n22963 ;
  assign n30108 = n30107 ^ n30105 ^ 1'b0 ;
  assign n30109 = ( ~n30102 & n30104 ) | ( ~n30102 & n30108 ) | ( n30104 & n30108 ) ;
  assign n30110 = ( n12421 & ~n14146 ) | ( n12421 & n14708 ) | ( ~n14146 & n14708 ) ;
  assign n30111 = n30110 ^ n6886 ^ 1'b0 ;
  assign n30112 = ( ~n4249 & n7600 ) | ( ~n4249 & n15983 ) | ( n7600 & n15983 ) ;
  assign n30113 = n30112 ^ n19965 ^ n14065 ;
  assign n30114 = ~n7255 & n18535 ;
  assign n30115 = n18774 ^ n9079 ^ 1'b0 ;
  assign n30116 = n6097 & n30115 ;
  assign n30117 = n4190 | n8915 ;
  assign n30118 = n30117 ^ n17062 ^ 1'b0 ;
  assign n30119 = ~n25105 & n30118 ;
  assign n30120 = ~n30116 & n30119 ;
  assign n30121 = n793 & ~n30120 ;
  assign n30122 = n17358 ^ n12109 ^ 1'b0 ;
  assign n30123 = n15732 | n30122 ;
  assign n30124 = n20814 ^ n10553 ^ n2991 ;
  assign n30125 = n2343 & n30124 ;
  assign n30126 = ( x207 & n937 ) | ( x207 & n6582 ) | ( n937 & n6582 ) ;
  assign n30127 = ( ~n4659 & n28048 ) | ( ~n4659 & n30126 ) | ( n28048 & n30126 ) ;
  assign n30128 = n3219 | n30127 ;
  assign n30129 = n11382 ^ x79 ^ 1'b0 ;
  assign n30130 = n6083 & n30129 ;
  assign n30131 = ~n9927 & n30130 ;
  assign n30132 = n30131 ^ n17370 ^ 1'b0 ;
  assign n30133 = x84 & n27995 ;
  assign n30134 = ~n25604 & n30133 ;
  assign n30135 = n4591 | n12868 ;
  assign n30136 = x3 & ~n30135 ;
  assign n30137 = n30136 ^ n18320 ^ 1'b0 ;
  assign n30138 = n28380 | n30137 ;
  assign n30139 = n26984 ^ n25136 ^ 1'b0 ;
  assign n30140 = ( ~n2177 & n7480 ) | ( ~n2177 & n12866 ) | ( n7480 & n12866 ) ;
  assign n30141 = ~n8870 & n30140 ;
  assign n30142 = n7398 & n30141 ;
  assign n30143 = ( ~n5364 & n8188 ) | ( ~n5364 & n10621 ) | ( n8188 & n10621 ) ;
  assign n30144 = n30143 ^ n16990 ^ x111 ;
  assign n30145 = n30144 ^ n8916 ^ x58 ;
  assign n30146 = n26177 ^ n18484 ^ 1'b0 ;
  assign n30147 = n3907 & ~n30146 ;
  assign n30148 = n2978 & ~n7401 ;
  assign n30149 = n30148 ^ n1543 ^ 1'b0 ;
  assign n30150 = ( ~n27758 & n29195 ) | ( ~n27758 & n30149 ) | ( n29195 & n30149 ) ;
  assign n30151 = n6781 & ~n30150 ;
  assign n30152 = n30151 ^ n27921 ^ 1'b0 ;
  assign n30153 = n17997 ^ n2160 ^ 1'b0 ;
  assign n30154 = n1822 & ~n30153 ;
  assign n30155 = ~n9508 & n30154 ;
  assign n30156 = ( n12389 & n14940 ) | ( n12389 & ~n30155 ) | ( n14940 & ~n30155 ) ;
  assign n30157 = ( ~n6512 & n17399 ) | ( ~n6512 & n26536 ) | ( n17399 & n26536 ) ;
  assign n30158 = ( n3227 & ~n15767 ) | ( n3227 & n30157 ) | ( ~n15767 & n30157 ) ;
  assign n30159 = n8809 & n16444 ;
  assign n30160 = n15335 ^ n13234 ^ n5909 ;
  assign n30161 = n15851 & n30160 ;
  assign n30162 = n22535 & n30161 ;
  assign n30163 = n30162 ^ n20881 ^ 1'b0 ;
  assign n30164 = n9341 & n30163 ;
  assign n30165 = ~n28426 & n30164 ;
  assign n30166 = n13163 & ~n18876 ;
  assign n30167 = n6053 & ~n14913 ;
  assign n30168 = n30166 & n30167 ;
  assign n30169 = n7165 & n30168 ;
  assign n30170 = n29070 ^ n28699 ^ 1'b0 ;
  assign n30171 = n24670 | n30170 ;
  assign n30173 = n6897 ^ n3249 ^ n1723 ;
  assign n30172 = n10472 ^ n9666 ^ n3727 ;
  assign n30174 = n30173 ^ n30172 ^ n5539 ;
  assign n30175 = n30174 ^ n23844 ^ n14917 ;
  assign n30176 = n28414 ^ n1749 ^ n471 ;
  assign n30177 = n30176 ^ n18506 ^ n18157 ;
  assign n30178 = n30177 ^ n18892 ^ 1'b0 ;
  assign n30179 = n23946 ^ n7763 ^ n5662 ;
  assign n30180 = n30179 ^ n19024 ^ 1'b0 ;
  assign n30181 = x72 | n8537 ;
  assign n30182 = n30181 ^ n16759 ^ 1'b0 ;
  assign n30183 = n10490 & n30182 ;
  assign n30184 = n343 & ~n21054 ;
  assign n30185 = n10779 ^ n9875 ^ n6725 ;
  assign n30186 = n8769 & n17117 ;
  assign n30187 = ~n6795 & n23456 ;
  assign n30188 = ~n6625 & n30187 ;
  assign n30189 = n11551 ^ n2519 ^ n1907 ;
  assign n30190 = ( n10834 & ~n12620 ) | ( n10834 & n30189 ) | ( ~n12620 & n30189 ) ;
  assign n30191 = n24759 & ~n30190 ;
  assign n30192 = n30191 ^ n413 ^ 1'b0 ;
  assign n30193 = ( n23432 & ~n30188 ) | ( n23432 & n30192 ) | ( ~n30188 & n30192 ) ;
  assign n30194 = n25112 ^ n2163 ^ 1'b0 ;
  assign n30195 = n2399 & ~n30194 ;
  assign n30196 = n30195 ^ n19531 ^ 1'b0 ;
  assign n30197 = ( n4310 & n6457 ) | ( n4310 & n23040 ) | ( n6457 & n23040 ) ;
  assign n30198 = n30197 ^ n4075 ^ n2086 ;
  assign n30199 = n30198 ^ n10738 ^ 1'b0 ;
  assign n30200 = n20888 & ~n30199 ;
  assign n30205 = n9855 ^ n2492 ^ 1'b0 ;
  assign n30206 = n6279 | n30205 ;
  assign n30201 = n1684 & n19703 ;
  assign n30202 = ~n17689 & n30201 ;
  assign n30203 = n30202 ^ n23543 ^ 1'b0 ;
  assign n30204 = n16999 & n30203 ;
  assign n30207 = n30206 ^ n30204 ^ 1'b0 ;
  assign n30208 = n4268 | n30207 ;
  assign n30210 = n7529 & ~n10932 ;
  assign n30209 = n6442 ^ n5021 ^ n1086 ;
  assign n30211 = n30210 ^ n30209 ^ n2743 ;
  assign n30212 = n14099 ^ n10955 ^ n1102 ;
  assign n30213 = n7167 & ~n10171 ;
  assign n30214 = ~n15615 & n30213 ;
  assign n30215 = n5570 | n30214 ;
  assign n30216 = n22744 ^ n15784 ^ 1'b0 ;
  assign n30217 = n20884 | n30216 ;
  assign n30218 = n12959 & ~n30217 ;
  assign n30219 = n30218 ^ n23745 ^ 1'b0 ;
  assign n30220 = n16115 ^ n8023 ^ n5506 ;
  assign n30221 = n17412 & n30220 ;
  assign n30222 = n22037 ^ n3422 ^ 1'b0 ;
  assign n30223 = n30222 ^ n14351 ^ 1'b0 ;
  assign n30229 = ( n3205 & ~n6368 ) | ( n3205 & n10181 ) | ( ~n6368 & n10181 ) ;
  assign n30228 = n4536 ^ n1191 ^ 1'b0 ;
  assign n30230 = n30229 ^ n30228 ^ 1'b0 ;
  assign n30231 = n3621 & ~n30230 ;
  assign n30232 = n30231 ^ n12194 ^ 1'b0 ;
  assign n30224 = n8462 ^ n2774 ^ 1'b0 ;
  assign n30225 = n14990 ^ n14243 ^ 1'b0 ;
  assign n30226 = n30224 | n30225 ;
  assign n30227 = n18361 & ~n30226 ;
  assign n30233 = n30232 ^ n30227 ^ 1'b0 ;
  assign n30234 = n7181 ^ n923 ^ 1'b0 ;
  assign n30235 = n18164 & n30234 ;
  assign n30236 = n15405 ^ n11588 ^ n8325 ;
  assign n30237 = n15645 ^ n289 ^ 1'b0 ;
  assign n30238 = n30237 ^ n23055 ^ 1'b0 ;
  assign n30239 = n30238 ^ n10721 ^ n5006 ;
  assign n30240 = ( ~n19836 & n23162 ) | ( ~n19836 & n25399 ) | ( n23162 & n25399 ) ;
  assign n30241 = n30240 ^ n9244 ^ 1'b0 ;
  assign n30242 = n15301 | n17084 ;
  assign n30243 = ( n6076 & ~n9647 ) | ( n6076 & n12359 ) | ( ~n9647 & n12359 ) ;
  assign n30244 = ( ~n30241 & n30242 ) | ( ~n30241 & n30243 ) | ( n30242 & n30243 ) ;
  assign n30245 = n24276 ^ n16510 ^ 1'b0 ;
  assign n30246 = n27610 & n30245 ;
  assign n30247 = x235 & n6739 ;
  assign n30248 = n30247 ^ n7534 ^ 1'b0 ;
  assign n30249 = n27392 ^ n23986 ^ n11383 ;
  assign n30250 = n332 & n15244 ;
  assign n30251 = ~n25492 & n30250 ;
  assign n30252 = n26693 | n29280 ;
  assign n30254 = n4008 | n11584 ;
  assign n30255 = n30254 ^ n5766 ^ 1'b0 ;
  assign n30256 = n1418 | n24690 ;
  assign n30257 = n30255 & ~n30256 ;
  assign n30253 = ( n4465 & n28188 ) | ( n4465 & ~n29849 ) | ( n28188 & ~n29849 ) ;
  assign n30258 = n30257 ^ n30253 ^ 1'b0 ;
  assign n30259 = n30258 ^ n16669 ^ n9259 ;
  assign n30260 = x80 & ~n2347 ;
  assign n30261 = n30260 ^ n13239 ^ n1920 ;
  assign n30262 = n8192 & n29071 ;
  assign n30263 = ~n9376 & n14197 ;
  assign n30264 = n8964 & n30263 ;
  assign n30265 = n11536 | n30042 ;
  assign n30266 = n30264 & n30265 ;
  assign n30267 = ~n1029 & n17763 ;
  assign n30270 = n10571 | n15860 ;
  assign n30271 = n30270 ^ n28959 ^ n3061 ;
  assign n30268 = n7388 ^ n3392 ^ 1'b0 ;
  assign n30269 = n30268 ^ n18880 ^ n4786 ;
  assign n30272 = n30271 ^ n30269 ^ n3097 ;
  assign n30273 = n27263 ^ n1819 ^ 1'b0 ;
  assign n30274 = n13341 | n16926 ;
  assign n30275 = n23612 ^ n8726 ^ n8666 ;
  assign n30276 = n27625 | n30275 ;
  assign n30277 = n26886 & ~n30276 ;
  assign n30278 = n977 | n4809 ;
  assign n30279 = n30278 ^ n21273 ^ n21229 ;
  assign n30280 = n25754 | n30279 ;
  assign n30281 = n30280 ^ n3125 ^ 1'b0 ;
  assign n30282 = n17656 ^ n9693 ^ n4283 ;
  assign n30283 = ( n16294 & ~n17813 ) | ( n16294 & n26823 ) | ( ~n17813 & n26823 ) ;
  assign n30284 = n30283 ^ n26355 ^ n22864 ;
  assign n30285 = n6862 & ~n27279 ;
  assign n30286 = ~n26040 & n30285 ;
  assign n30287 = n30286 ^ n17294 ^ 1'b0 ;
  assign n30288 = n8715 & ~n10430 ;
  assign n30289 = n30288 ^ n3012 ^ 1'b0 ;
  assign n30290 = n30289 ^ n15533 ^ 1'b0 ;
  assign n30291 = n8939 & ~n30290 ;
  assign n30292 = n16362 & n21348 ;
  assign n30293 = n19862 ^ n12739 ^ n6821 ;
  assign n30294 = n8504 | n14016 ;
  assign n30295 = ( n6691 & n11197 ) | ( n6691 & ~n11224 ) | ( n11197 & ~n11224 ) ;
  assign n30296 = ~n4850 & n30295 ;
  assign n30297 = ~n30294 & n30296 ;
  assign n30298 = ( n30292 & n30293 ) | ( n30292 & ~n30297 ) | ( n30293 & ~n30297 ) ;
  assign n30299 = ~n9306 & n29206 ;
  assign n30300 = ~n19836 & n30299 ;
  assign n30301 = n30300 ^ n26797 ^ 1'b0 ;
  assign n30302 = ~n4419 & n6064 ;
  assign n30303 = n479 | n6856 ;
  assign n30304 = n23760 | n30303 ;
  assign n30305 = n10552 & ~n30304 ;
  assign n30306 = n1646 & n16453 ;
  assign n30307 = n30305 & n30306 ;
  assign n30313 = ( n4289 & n10287 ) | ( n4289 & n24837 ) | ( n10287 & n24837 ) ;
  assign n30308 = n15686 ^ n13610 ^ 1'b0 ;
  assign n30309 = n30308 ^ n26875 ^ 1'b0 ;
  assign n30310 = n6602 | n18944 ;
  assign n30311 = n20649 & n30310 ;
  assign n30312 = n30309 & ~n30311 ;
  assign n30314 = n30313 ^ n30312 ^ 1'b0 ;
  assign n30317 = n12135 | n20605 ;
  assign n30318 = n18838 | n30317 ;
  assign n30315 = ( ~n6540 & n11476 ) | ( ~n6540 & n13702 ) | ( n11476 & n13702 ) ;
  assign n30316 = n19371 & ~n30315 ;
  assign n30319 = n30318 ^ n30316 ^ 1'b0 ;
  assign n30320 = n15959 ^ x74 ^ 1'b0 ;
  assign n30321 = n21097 ^ n11501 ^ 1'b0 ;
  assign n30323 = n28704 ^ n22528 ^ n8762 ;
  assign n30322 = ~n11475 & n28756 ;
  assign n30324 = n30323 ^ n30322 ^ 1'b0 ;
  assign n30325 = n30324 ^ n29173 ^ n22821 ;
  assign n30326 = n5977 | n8427 ;
  assign n30327 = n30326 ^ n20941 ^ 1'b0 ;
  assign n30328 = n939 & ~n16277 ;
  assign n30329 = ~n18159 & n30328 ;
  assign n30330 = n30329 ^ n15660 ^ 1'b0 ;
  assign n30331 = n30327 & ~n30330 ;
  assign n30332 = n8601 | n21016 ;
  assign n30333 = n4893 & ~n30332 ;
  assign n30334 = n16744 & ~n22923 ;
  assign n30335 = ( ~n10144 & n23129 ) | ( ~n10144 & n23930 ) | ( n23129 & n23930 ) ;
  assign n30336 = n30335 ^ n5371 ^ n5212 ;
  assign n30337 = ~n22210 & n23249 ;
  assign n30338 = n30337 ^ n28005 ^ 1'b0 ;
  assign n30339 = n14870 ^ n6911 ^ 1'b0 ;
  assign n30340 = ( n21683 & ~n30338 ) | ( n21683 & n30339 ) | ( ~n30338 & n30339 ) ;
  assign n30341 = n30336 | n30340 ;
  assign n30342 = n6594 ^ n1654 ^ 1'b0 ;
  assign n30343 = n30342 ^ n7488 ^ 1'b0 ;
  assign n30344 = n20397 | n30343 ;
  assign n30345 = n3770 & ~n13824 ;
  assign n30346 = n30345 ^ n5681 ^ 1'b0 ;
  assign n30347 = n7032 & n30346 ;
  assign n30348 = ~n23722 & n30347 ;
  assign n30349 = ( x70 & n30068 ) | ( x70 & ~n30348 ) | ( n30068 & ~n30348 ) ;
  assign n30350 = n19061 ^ n9242 ^ 1'b0 ;
  assign n30351 = ( n3945 & n5356 ) | ( n3945 & ~n30350 ) | ( n5356 & ~n30350 ) ;
  assign n30352 = ~n2531 & n8375 ;
  assign n30353 = n30351 & n30352 ;
  assign n30354 = n30353 ^ n6139 ^ 1'b0 ;
  assign n30355 = ~n1049 & n11181 ;
  assign n30356 = n30355 ^ n19128 ^ 1'b0 ;
  assign n30357 = ( n4454 & ~n8817 ) | ( n4454 & n14657 ) | ( ~n8817 & n14657 ) ;
  assign n30358 = ~n2401 & n30357 ;
  assign n30359 = n30358 ^ n8014 ^ 1'b0 ;
  assign n30360 = n30359 ^ n9421 ^ n3930 ;
  assign n30361 = ( n9705 & n16834 ) | ( n9705 & n23972 ) | ( n16834 & n23972 ) ;
  assign n30362 = n12364 ^ n449 ^ 1'b0 ;
  assign n30363 = n19152 | n30362 ;
  assign n30364 = n30361 & ~n30363 ;
  assign n30365 = n4807 ^ n4053 ^ n2960 ;
  assign n30366 = n30365 ^ n18143 ^ n1403 ;
  assign n30367 = n30366 ^ n9603 ^ x169 ;
  assign n30368 = n30367 ^ n14424 ^ 1'b0 ;
  assign n30369 = n14945 | n30368 ;
  assign n30370 = n27334 ^ n8786 ^ 1'b0 ;
  assign n30371 = ( n4155 & n23077 ) | ( n4155 & n30370 ) | ( n23077 & n30370 ) ;
  assign n30372 = n24157 & ~n30371 ;
  assign n30373 = n30369 & n30372 ;
  assign n30374 = n16336 ^ n877 ^ 1'b0 ;
  assign n30375 = n30374 ^ n23612 ^ n18565 ;
  assign n30376 = n13071 ^ n4053 ^ 1'b0 ;
  assign n30377 = ( x100 & n27968 ) | ( x100 & n30376 ) | ( n27968 & n30376 ) ;
  assign n30378 = n11806 ^ n10000 ^ 1'b0 ;
  assign n30381 = n3520 | n5642 ;
  assign n30380 = n15842 & ~n22134 ;
  assign n30382 = n30381 ^ n30380 ^ n6041 ;
  assign n30383 = n30382 ^ n2952 ^ 1'b0 ;
  assign n30384 = n3463 & n30383 ;
  assign n30379 = n5353 ^ n1318 ^ 1'b0 ;
  assign n30385 = n30384 ^ n30379 ^ 1'b0 ;
  assign n30386 = n30385 ^ n22840 ^ n19503 ;
  assign n30387 = n4777 & n23413 ;
  assign n30388 = n30387 ^ n20844 ^ 1'b0 ;
  assign n30389 = n7616 ^ n3411 ^ 1'b0 ;
  assign n30390 = n2009 | n30389 ;
  assign n30391 = ~n2614 & n4688 ;
  assign n30392 = ~n2382 & n30391 ;
  assign n30393 = ( n758 & ~n22057 ) | ( n758 & n30392 ) | ( ~n22057 & n30392 ) ;
  assign n30394 = n30393 ^ n2152 ^ 1'b0 ;
  assign n30395 = ( n13066 & n19149 ) | ( n13066 & ~n30394 ) | ( n19149 & ~n30394 ) ;
  assign n30396 = n21654 ^ n5017 ^ 1'b0 ;
  assign n30397 = n28998 ^ n6479 ^ n4766 ;
  assign n30398 = n11449 | n30397 ;
  assign n30399 = n30398 ^ n11062 ^ 1'b0 ;
  assign n30400 = n30399 ^ n29249 ^ 1'b0 ;
  assign n30401 = ~n18508 & n30400 ;
  assign n30402 = n19940 ^ n5126 ^ 1'b0 ;
  assign n30403 = n8969 & ~n30402 ;
  assign n30404 = n30403 ^ n11376 ^ 1'b0 ;
  assign n30405 = n18017 ^ n8317 ^ 1'b0 ;
  assign n30406 = n30404 & n30405 ;
  assign n30407 = n3605 & ~n11500 ;
  assign n30408 = n30407 ^ n19512 ^ n16481 ;
  assign n30409 = n30408 ^ n28985 ^ 1'b0 ;
  assign n30410 = ~n25533 & n30409 ;
  assign n30411 = n13096 ^ n7826 ^ 1'b0 ;
  assign n30412 = n30411 ^ n301 ^ 1'b0 ;
  assign n30413 = n9447 | n30412 ;
  assign n30414 = n367 & n18919 ;
  assign n30415 = n30413 & n30414 ;
  assign n30416 = n15154 | n17141 ;
  assign n30417 = ~n20784 & n23178 ;
  assign n30419 = n21046 ^ n12532 ^ 1'b0 ;
  assign n30418 = x130 & ~n4707 ;
  assign n30420 = n30419 ^ n30418 ^ 1'b0 ;
  assign n30421 = ~n737 & n30420 ;
  assign n30422 = n9612 | n20410 ;
  assign n30423 = n18770 & n19650 ;
  assign n30424 = n30423 ^ n22478 ^ 1'b0 ;
  assign n30425 = ( n3579 & ~n13832 ) | ( n3579 & n28761 ) | ( ~n13832 & n28761 ) ;
  assign n30426 = n20475 | n30425 ;
  assign n30427 = n25346 & ~n30426 ;
  assign n30428 = n8581 | n30427 ;
  assign n30429 = n30428 ^ n9505 ^ 1'b0 ;
  assign n30430 = n12304 | n14135 ;
  assign n30431 = n30430 ^ n3821 ^ 1'b0 ;
  assign n30432 = n29703 ^ n17954 ^ 1'b0 ;
  assign n30433 = n30432 ^ n8272 ^ 1'b0 ;
  assign n30434 = ~n30431 & n30433 ;
  assign n30435 = n4510 & n19945 ;
  assign n30436 = n30435 ^ n17446 ^ n17040 ;
  assign n30437 = n1273 & ~n30436 ;
  assign n30438 = n30437 ^ n19172 ^ 1'b0 ;
  assign n30439 = n25642 | n30438 ;
  assign n30440 = n30439 ^ n28037 ^ n16030 ;
  assign n30441 = ( n8418 & n15805 ) | ( n8418 & ~n30440 ) | ( n15805 & ~n30440 ) ;
  assign n30442 = n15815 ^ n15011 ^ n9228 ;
  assign n30443 = n30442 ^ n5741 ^ 1'b0 ;
  assign n30444 = n1735 & n12900 ;
  assign n30445 = n30444 ^ n12406 ^ 1'b0 ;
  assign n30446 = n9596 ^ n4986 ^ 1'b0 ;
  assign n30447 = n30445 | n30446 ;
  assign n30448 = ( ~n1516 & n26646 ) | ( ~n1516 & n30447 ) | ( n26646 & n30447 ) ;
  assign n30449 = ~n1226 & n13687 ;
  assign n30450 = n30449 ^ n9508 ^ 1'b0 ;
  assign n30451 = n7031 | n12613 ;
  assign n30452 = n477 | n30451 ;
  assign n30454 = ~n2422 & n5442 ;
  assign n30455 = n30454 ^ n8634 ^ 1'b0 ;
  assign n30456 = n30455 ^ n4629 ^ 1'b0 ;
  assign n30453 = n7296 | n28272 ;
  assign n30457 = n30456 ^ n30453 ^ 1'b0 ;
  assign n30458 = n21118 & ~n27985 ;
  assign n30459 = ( ~n5535 & n30219 ) | ( ~n5535 & n30458 ) | ( n30219 & n30458 ) ;
  assign n30460 = ( ~x246 & n6336 ) | ( ~x246 & n8555 ) | ( n6336 & n8555 ) ;
  assign n30461 = ~n11293 & n19648 ;
  assign n30462 = n30460 & n30461 ;
  assign n30463 = n2338 & n5815 ;
  assign n30464 = n30462 & n30463 ;
  assign n30465 = n19093 ^ n14369 ^ 1'b0 ;
  assign n30466 = ( n686 & n9413 ) | ( n686 & n28887 ) | ( n9413 & n28887 ) ;
  assign n30467 = n30466 ^ n6976 ^ 1'b0 ;
  assign n30468 = n12977 & ~n30467 ;
  assign n30469 = ( x212 & n5205 ) | ( x212 & ~n30468 ) | ( n5205 & ~n30468 ) ;
  assign n30470 = n2782 | n13388 ;
  assign n30471 = n30470 ^ n21192 ^ n4799 ;
  assign n30472 = ( n7505 & n8276 ) | ( n7505 & ~n21087 ) | ( n8276 & ~n21087 ) ;
  assign n30473 = n9334 ^ n2947 ^ 1'b0 ;
  assign n30474 = n13713 ^ n3921 ^ 1'b0 ;
  assign n30475 = n7579 & n30474 ;
  assign n30476 = ~n23992 & n30475 ;
  assign n30477 = n3273 | n25104 ;
  assign n30478 = n29195 | n30477 ;
  assign n30479 = n30478 ^ n22088 ^ 1'b0 ;
  assign n30480 = n16459 ^ n13590 ^ n1438 ;
  assign n30481 = n363 & n29927 ;
  assign n30482 = n19368 ^ n7173 ^ 1'b0 ;
  assign n30483 = n782 & n30482 ;
  assign n30484 = n30483 ^ n11460 ^ n6328 ;
  assign n30485 = n27027 ^ n3546 ^ n2036 ;
  assign n30486 = n1137 | n30485 ;
  assign n30487 = n9373 ^ n7436 ^ n3106 ;
  assign n30488 = ( ~n2761 & n14518 ) | ( ~n2761 & n14685 ) | ( n14518 & n14685 ) ;
  assign n30489 = ( ~n4715 & n12705 ) | ( ~n4715 & n30488 ) | ( n12705 & n30488 ) ;
  assign n30490 = n10622 & n12400 ;
  assign n30491 = ~n28930 & n30490 ;
  assign n30492 = n4626 | n18327 ;
  assign n30493 = n30491 & ~n30492 ;
  assign n30494 = ~n23173 & n30493 ;
  assign n30495 = n4077 | n28336 ;
  assign n30496 = n24938 ^ n21671 ^ n4180 ;
  assign n30497 = n26257 ^ n19424 ^ n7051 ;
  assign n30498 = ( ~n4457 & n15967 ) | ( ~n4457 & n30497 ) | ( n15967 & n30497 ) ;
  assign n30499 = ~n17097 & n22162 ;
  assign n30500 = ( n18530 & n28618 ) | ( n18530 & n30499 ) | ( n28618 & n30499 ) ;
  assign n30501 = n19610 ^ n1417 ^ 1'b0 ;
  assign n30502 = ~n11227 & n30501 ;
  assign n30503 = n3361 & n30502 ;
  assign n30504 = ~n1666 & n30503 ;
  assign n30505 = n15163 | n20754 ;
  assign n30506 = n30505 ^ n19401 ^ 1'b0 ;
  assign n30507 = n18385 ^ n2606 ^ n947 ;
  assign n30508 = n30507 ^ n881 ^ 1'b0 ;
  assign n30509 = n21251 ^ n18349 ^ 1'b0 ;
  assign n30510 = n30509 ^ n19947 ^ n10464 ;
  assign n30511 = n14957 | n30510 ;
  assign n30512 = n11804 & ~n30511 ;
  assign n30513 = n26175 ^ n25899 ^ 1'b0 ;
  assign n30520 = n10049 | n11002 ;
  assign n30521 = n2103 | n30520 ;
  assign n30514 = n2945 & ~n11179 ;
  assign n30515 = ~n12984 & n30514 ;
  assign n30516 = n4457 | n12924 ;
  assign n30517 = n6396 | n30516 ;
  assign n30518 = ~n30515 & n30517 ;
  assign n30519 = n30518 ^ x194 ^ 1'b0 ;
  assign n30522 = n30521 ^ n30519 ^ n12569 ;
  assign n30523 = n11605 ^ n10631 ^ 1'b0 ;
  assign n30524 = n13585 & n17808 ;
  assign n30525 = ~n30523 & n30524 ;
  assign n30526 = n18639 | n30525 ;
  assign n30527 = n6705 & ~n30526 ;
  assign n30528 = n30527 ^ n11347 ^ 1'b0 ;
  assign n30529 = n14210 ^ n4023 ^ 1'b0 ;
  assign n30530 = n30529 ^ n27079 ^ n9450 ;
  assign n30533 = n23980 ^ n593 ^ 1'b0 ;
  assign n30534 = n26291 & ~n30533 ;
  assign n30535 = n22332 & ~n30534 ;
  assign n30536 = n13376 ^ n8345 ^ n5082 ;
  assign n30537 = n3585 | n30536 ;
  assign n30538 = n30535 | n30537 ;
  assign n30531 = n14362 & ~n24848 ;
  assign n30532 = ~n14624 & n30531 ;
  assign n30539 = n30538 ^ n30532 ^ 1'b0 ;
  assign n30540 = ~n4713 & n26291 ;
  assign n30541 = n16838 | n17576 ;
  assign n30542 = n14818 | n30541 ;
  assign n30543 = n30542 ^ n7353 ^ 1'b0 ;
  assign n30544 = ~n5406 & n14218 ;
  assign n30545 = n5681 & ~n22345 ;
  assign n30546 = n305 & n14620 ;
  assign n30547 = ( ~n20615 & n28005 ) | ( ~n20615 & n30546 ) | ( n28005 & n30546 ) ;
  assign n30548 = x10 | n30547 ;
  assign n30549 = n29454 | n30548 ;
  assign n30550 = ( n22340 & n30545 ) | ( n22340 & n30549 ) | ( n30545 & n30549 ) ;
  assign n30551 = ~n271 & n13466 ;
  assign n30552 = n30551 ^ n11221 ^ 1'b0 ;
  assign n30553 = n14173 ^ n7709 ^ 1'b0 ;
  assign n30554 = n27446 & n30553 ;
  assign n30555 = n29186 ^ n22374 ^ n18380 ;
  assign n30556 = n24570 ^ n21410 ^ 1'b0 ;
  assign n30557 = n7944 | n30556 ;
  assign n30558 = n14697 ^ n10800 ^ 1'b0 ;
  assign n30559 = n19929 ^ n17252 ^ 1'b0 ;
  assign n30560 = n16148 & n30559 ;
  assign n30561 = n21449 ^ n365 ^ 1'b0 ;
  assign n30562 = n944 & ~n7268 ;
  assign n30563 = n30562 ^ n1896 ^ 1'b0 ;
  assign n30564 = ( n10976 & ~n26540 ) | ( n10976 & n30563 ) | ( ~n26540 & n30563 ) ;
  assign n30565 = ( n16976 & ~n28331 ) | ( n16976 & n30564 ) | ( ~n28331 & n30564 ) ;
  assign n30566 = ( n4480 & ~n15817 ) | ( n4480 & n30462 ) | ( ~n15817 & n30462 ) ;
  assign n30567 = n12784 ^ n9082 ^ n5926 ;
  assign n30568 = ( n22168 & n29391 ) | ( n22168 & n30567 ) | ( n29391 & n30567 ) ;
  assign n30569 = ~n6869 & n7994 ;
  assign n30570 = ~n13297 & n30569 ;
  assign n30571 = n3894 & ~n18390 ;
  assign n30572 = n30571 ^ n1108 ^ n301 ;
  assign n30573 = n28804 ^ n338 ^ 1'b0 ;
  assign n30574 = n14224 | n22338 ;
  assign n30575 = n30573 & ~n30574 ;
  assign n30576 = ( ~n18035 & n28131 ) | ( ~n18035 & n30575 ) | ( n28131 & n30575 ) ;
  assign n30577 = n14745 ^ n12832 ^ n8598 ;
  assign n30581 = n16690 ^ n13529 ^ n8091 ;
  assign n30578 = n5117 | n5381 ;
  assign n30579 = n30578 ^ n3371 ^ 1'b0 ;
  assign n30580 = n3634 & n30579 ;
  assign n30582 = n30581 ^ n30580 ^ n12430 ;
  assign n30584 = n9613 | n14975 ;
  assign n30585 = n30584 ^ n2858 ^ 1'b0 ;
  assign n30583 = ~n5499 & n15143 ;
  assign n30586 = n30585 ^ n30583 ^ 1'b0 ;
  assign n30587 = n5272 & n29732 ;
  assign n30588 = n1868 & n30587 ;
  assign n30589 = x102 & n2620 ;
  assign n30590 = n7234 & n30589 ;
  assign n30595 = n23472 ^ n22593 ^ 1'b0 ;
  assign n30596 = n13655 & n30595 ;
  assign n30591 = n10913 ^ n2944 ^ 1'b0 ;
  assign n30592 = n30591 ^ n26504 ^ 1'b0 ;
  assign n30593 = n22971 | n30592 ;
  assign n30594 = n12481 & ~n30593 ;
  assign n30597 = n30596 ^ n30594 ^ 1'b0 ;
  assign n30598 = n29221 ^ n19297 ^ 1'b0 ;
  assign n30599 = ( n370 & n2116 ) | ( n370 & n16541 ) | ( n2116 & n16541 ) ;
  assign n30600 = n21244 ^ n20420 ^ n5522 ;
  assign n30601 = n16492 & n30600 ;
  assign n30602 = ~n11219 & n30601 ;
  assign n30603 = n30602 ^ n4995 ^ 1'b0 ;
  assign n30604 = n7014 & n30603 ;
  assign n30605 = n4701 ^ n1674 ^ n962 ;
  assign n30606 = ( n946 & n30604 ) | ( n946 & ~n30605 ) | ( n30604 & ~n30605 ) ;
  assign n30607 = n19157 ^ n17157 ^ 1'b0 ;
  assign n30608 = n367 & ~n30607 ;
  assign n30609 = n22324 ^ n8613 ^ 1'b0 ;
  assign n30610 = ~n24002 & n30609 ;
  assign n30611 = n30267 ^ n11831 ^ 1'b0 ;
  assign n30612 = n15091 & n30611 ;
  assign n30613 = ( n8178 & n11572 ) | ( n8178 & n29261 ) | ( n11572 & n29261 ) ;
  assign n30614 = n21785 ^ n3804 ^ 1'b0 ;
  assign n30615 = n28131 & n30614 ;
  assign n30619 = n698 | n18341 ;
  assign n30620 = n25862 & ~n30619 ;
  assign n30616 = n14154 & ~n18043 ;
  assign n30617 = n1752 & n30616 ;
  assign n30618 = n2419 & ~n30617 ;
  assign n30621 = n30620 ^ n30618 ^ 1'b0 ;
  assign n30622 = n27222 ^ n7226 ^ 1'b0 ;
  assign n30623 = n11193 & ~n28270 ;
  assign n30624 = n30623 ^ n3521 ^ 1'b0 ;
  assign n30625 = n8969 & n12900 ;
  assign n30626 = n30625 ^ n2905 ^ 1'b0 ;
  assign n30627 = n8093 & ~n21071 ;
  assign n30628 = n30626 & ~n30627 ;
  assign n30629 = n24759 & ~n26648 ;
  assign n30630 = n30629 ^ n27614 ^ 1'b0 ;
  assign n30631 = n30630 ^ n9420 ^ 1'b0 ;
  assign n30632 = ~n12104 & n30631 ;
  assign n30633 = n30632 ^ n21625 ^ n4745 ;
  assign n30636 = ( n12522 & n24900 ) | ( n12522 & ~n29395 ) | ( n24900 & ~n29395 ) ;
  assign n30637 = n30636 ^ n23251 ^ n8201 ;
  assign n30634 = x11 & n13672 ;
  assign n30635 = n30634 ^ n4187 ^ 1'b0 ;
  assign n30638 = n30637 ^ n30635 ^ n16674 ;
  assign n30639 = n2124 | n4513 ;
  assign n30640 = ~n3149 & n25427 ;
  assign n30641 = n4374 & ~n22702 ;
  assign n30642 = n25179 ^ n12276 ^ 1'b0 ;
  assign n30643 = n8330 ^ n8176 ^ 1'b0 ;
  assign n30644 = n11225 & ~n30643 ;
  assign n30645 = ( n1422 & n2875 ) | ( n1422 & ~n21830 ) | ( n2875 & ~n21830 ) ;
  assign n30646 = ~n3432 & n30645 ;
  assign n30647 = n30646 ^ n3744 ^ 1'b0 ;
  assign n30648 = n15153 ^ n4553 ^ 1'b0 ;
  assign n30649 = ( n4232 & n30647 ) | ( n4232 & n30648 ) | ( n30647 & n30648 ) ;
  assign n30650 = n12066 ^ n9319 ^ 1'b0 ;
  assign n30651 = ( n5349 & n9981 ) | ( n5349 & ~n10047 ) | ( n9981 & ~n10047 ) ;
  assign n30652 = n30651 ^ n8568 ^ n1689 ;
  assign n30653 = ( n3184 & n8052 ) | ( n3184 & n9816 ) | ( n8052 & n9816 ) ;
  assign n30654 = ~n17571 & n30411 ;
  assign n30655 = n30654 ^ n19282 ^ 1'b0 ;
  assign n30656 = n10626 ^ n7254 ^ 1'b0 ;
  assign n30661 = n16568 ^ n11199 ^ 1'b0 ;
  assign n30662 = n8652 | n30661 ;
  assign n30657 = n11566 ^ n11031 ^ n5803 ;
  assign n30658 = ~x106 & n30657 ;
  assign n30659 = ~n256 & n30658 ;
  assign n30660 = n30659 ^ n28106 ^ n18751 ;
  assign n30663 = n30662 ^ n30660 ^ 1'b0 ;
  assign n30664 = ( n2413 & n8254 ) | ( n2413 & n13514 ) | ( n8254 & n13514 ) ;
  assign n30665 = n13223 & n25256 ;
  assign n30666 = ~n8066 & n30665 ;
  assign n30667 = n30666 ^ n12977 ^ 1'b0 ;
  assign n30668 = n30664 | n30667 ;
  assign n30669 = n26942 & ~n30668 ;
  assign n30670 = n5367 & n30669 ;
  assign n30671 = n22888 ^ n8241 ^ n7493 ;
  assign n30672 = n15462 & ~n19569 ;
  assign n30673 = n30671 & n30672 ;
  assign n30674 = ( n4993 & n14109 ) | ( n4993 & ~n30673 ) | ( n14109 & ~n30673 ) ;
  assign n30675 = n18666 ^ n1521 ^ n1239 ;
  assign n30676 = n30675 ^ n22025 ^ n2702 ;
  assign n30677 = ~n1782 & n23805 ;
  assign n30678 = ~n2325 & n30677 ;
  assign n30679 = ( n2321 & n2930 ) | ( n2321 & n4076 ) | ( n2930 & n4076 ) ;
  assign n30680 = n30679 ^ n22594 ^ 1'b0 ;
  assign n30681 = n9391 & ~n30680 ;
  assign n30682 = n3665 & n4575 ;
  assign n30683 = n2790 & n30682 ;
  assign n30684 = n4513 & ~n25941 ;
  assign n30685 = n9851 & n10418 ;
  assign n30686 = n548 | n11078 ;
  assign n30687 = ~n4983 & n18619 ;
  assign n30688 = n30687 ^ n4841 ^ 1'b0 ;
  assign n30689 = n4494 | n30688 ;
  assign n30690 = n30689 ^ n29576 ^ n9912 ;
  assign n30691 = ~n3363 & n7196 ;
  assign n30692 = n3363 & n30691 ;
  assign n30693 = ~n820 & n2155 ;
  assign n30694 = n820 & n30693 ;
  assign n30697 = n5256 | n10060 ;
  assign n30698 = n18534 ^ n11149 ^ 1'b0 ;
  assign n30699 = ~n7458 & n30698 ;
  assign n30700 = ( n6807 & n28756 ) | ( n6807 & n30699 ) | ( n28756 & n30699 ) ;
  assign n30701 = ( n23042 & ~n30697 ) | ( n23042 & n30700 ) | ( ~n30697 & n30700 ) ;
  assign n30702 = n30701 ^ n5470 ^ 1'b0 ;
  assign n30703 = n11006 & ~n30702 ;
  assign n30704 = n30703 ^ n20008 ^ 1'b0 ;
  assign n30695 = n15155 & ~n23949 ;
  assign n30696 = n30695 ^ n27288 ^ n16233 ;
  assign n30705 = n30704 ^ n30696 ^ 1'b0 ;
  assign n30706 = ( ~n30692 & n30694 ) | ( ~n30692 & n30705 ) | ( n30694 & n30705 ) ;
  assign n30707 = n13238 ^ n9876 ^ n7308 ;
  assign n30708 = ( n4720 & n7936 ) | ( n4720 & ~n30707 ) | ( n7936 & ~n30707 ) ;
  assign n30709 = n867 | n30708 ;
  assign n30710 = n4353 & ~n30709 ;
  assign n30711 = n9147 | n30710 ;
  assign n30712 = n21292 ^ n1099 ^ 1'b0 ;
  assign n30713 = ~n10686 & n30712 ;
  assign n30714 = n17881 ^ n10004 ^ 1'b0 ;
  assign n30715 = ( n16779 & n21818 ) | ( n16779 & ~n30714 ) | ( n21818 & ~n30714 ) ;
  assign n30716 = n15753 ^ n15717 ^ 1'b0 ;
  assign n30717 = n30715 & n30716 ;
  assign n30718 = n30717 ^ n9757 ^ n9405 ;
  assign n30719 = n3643 & ~n26250 ;
  assign n30720 = n30719 ^ n17657 ^ n8734 ;
  assign n30721 = n15845 ^ n15478 ^ n5302 ;
  assign n30723 = n12047 ^ n4724 ^ n1284 ;
  assign n30722 = n29265 ^ n3918 ^ 1'b0 ;
  assign n30724 = n30723 ^ n30722 ^ n3323 ;
  assign n30725 = n24403 ^ n10532 ^ n9255 ;
  assign n30726 = ( n6101 & n15621 ) | ( n6101 & ~n28300 ) | ( n15621 & ~n28300 ) ;
  assign n30727 = n1541 ^ n289 ^ 1'b0 ;
  assign n30728 = ( ~n7515 & n8488 ) | ( ~n7515 & n28200 ) | ( n8488 & n28200 ) ;
  assign n30729 = n29917 ^ n9378 ^ 1'b0 ;
  assign n30730 = n30728 & ~n30729 ;
  assign n30731 = ( n5574 & ~n8958 ) | ( n5574 & n16238 ) | ( ~n8958 & n16238 ) ;
  assign n30732 = ~n7452 & n30731 ;
  assign n30733 = n21228 & n30732 ;
  assign n30734 = n30733 ^ n20289 ^ n11044 ;
  assign n30735 = ( n1773 & n13289 ) | ( n1773 & ~n16003 ) | ( n13289 & ~n16003 ) ;
  assign n30736 = ( n8502 & n10953 ) | ( n8502 & ~n30735 ) | ( n10953 & ~n30735 ) ;
  assign n30737 = n30736 ^ n26648 ^ n12967 ;
  assign n30738 = n25148 ^ n3009 ^ 1'b0 ;
  assign n30739 = n30738 ^ n7011 ^ n5316 ;
  assign n30740 = n30737 & n30739 ;
  assign n30741 = ~n7276 & n22560 ;
  assign n30742 = ~n14856 & n17635 ;
  assign n30743 = n30741 & n30742 ;
  assign n30744 = n23614 ^ n18247 ^ n8122 ;
  assign n30745 = n22885 ^ n9911 ^ n6551 ;
  assign n30746 = n29932 ^ n8769 ^ n2306 ;
  assign n30747 = ~n7932 & n14452 ;
  assign n30748 = n30747 ^ n29090 ^ 1'b0 ;
  assign n30749 = n18559 ^ n3246 ^ 1'b0 ;
  assign n30750 = n11666 ^ n5383 ^ 1'b0 ;
  assign n30751 = n5909 ^ n5500 ^ n4036 ;
  assign n30754 = n20115 ^ n2887 ^ 1'b0 ;
  assign n30752 = n7698 ^ n4552 ^ 1'b0 ;
  assign n30753 = n4138 & n30752 ;
  assign n30755 = n30754 ^ n30753 ^ 1'b0 ;
  assign n30756 = n7688 ^ n1264 ^ 1'b0 ;
  assign n30757 = n11543 & n12000 ;
  assign n30758 = n30757 ^ n19508 ^ 1'b0 ;
  assign n30759 = n21333 & ~n22131 ;
  assign n30760 = n30759 ^ n7256 ^ 1'b0 ;
  assign n30761 = n5205 & ~n7812 ;
  assign n30762 = n30761 ^ n30132 ^ 1'b0 ;
  assign n30763 = n21752 ^ n21513 ^ 1'b0 ;
  assign n30764 = ~n17803 & n30763 ;
  assign n30765 = ( ~n7201 & n9145 ) | ( ~n7201 & n12491 ) | ( n9145 & n12491 ) ;
  assign n30766 = n30765 ^ n28018 ^ n5482 ;
  assign n30767 = n26504 ^ n11823 ^ 1'b0 ;
  assign n30768 = x147 & n27247 ;
  assign n30769 = ~n22878 & n30768 ;
  assign n30770 = n19650 ^ n16964 ^ n9583 ;
  assign n30771 = n11231 & ~n12721 ;
  assign n30772 = n30771 ^ n6593 ^ 1'b0 ;
  assign n30773 = n30770 & n30772 ;
  assign n30774 = n27116 & n30773 ;
  assign n30775 = ~n5300 & n8294 ;
  assign n30776 = n30775 ^ n6807 ^ 1'b0 ;
  assign n30777 = ( n2796 & ~n15556 ) | ( n2796 & n30776 ) | ( ~n15556 & n30776 ) ;
  assign n30778 = n30777 ^ n24247 ^ 1'b0 ;
  assign n30779 = ~n30774 & n30778 ;
  assign n30780 = n20123 & n22141 ;
  assign n30781 = ( n4538 & n19845 ) | ( n4538 & n30780 ) | ( n19845 & n30780 ) ;
  assign n30782 = ( ~n4648 & n28397 ) | ( ~n4648 & n30781 ) | ( n28397 & n30781 ) ;
  assign n30783 = ~n13155 & n22133 ;
  assign n30784 = ~n4137 & n9626 ;
  assign n30785 = n11118 & ~n29833 ;
  assign n30786 = ~n30784 & n30785 ;
  assign n30787 = n30786 ^ n22301 ^ n17312 ;
  assign n30788 = ( n8120 & ~n19770 ) | ( n8120 & n27850 ) | ( ~n19770 & n27850 ) ;
  assign n30789 = n23075 & n30788 ;
  assign n30794 = n7579 & ~n17058 ;
  assign n30795 = n3623 & n30794 ;
  assign n30790 = n1037 & n6253 ;
  assign n30791 = n11413 & n30790 ;
  assign n30792 = n10709 | n30791 ;
  assign n30793 = n15088 | n30792 ;
  assign n30796 = n30795 ^ n30793 ^ 1'b0 ;
  assign n30797 = n28167 ^ n18140 ^ n13251 ;
  assign n30799 = n15389 ^ n10007 ^ 1'b0 ;
  assign n30798 = n1855 | n15649 ;
  assign n30800 = n30799 ^ n30798 ^ 1'b0 ;
  assign n30801 = n22214 ^ n12746 ^ 1'b0 ;
  assign n30802 = n30800 | n30801 ;
  assign n30803 = n8122 & n17246 ;
  assign n30804 = n19514 ^ n16352 ^ n14385 ;
  assign n30805 = n15873 & n30293 ;
  assign n30806 = ( n18749 & ~n30804 ) | ( n18749 & n30805 ) | ( ~n30804 & n30805 ) ;
  assign n30807 = ( n1093 & n11045 ) | ( n1093 & n13722 ) | ( n11045 & n13722 ) ;
  assign n30808 = ( ~n1863 & n2592 ) | ( ~n1863 & n24431 ) | ( n2592 & n24431 ) ;
  assign n30809 = n30808 ^ n4917 ^ 1'b0 ;
  assign n30810 = ( n6967 & ~n30807 ) | ( n6967 & n30809 ) | ( ~n30807 & n30809 ) ;
  assign n30811 = n20664 ^ n17134 ^ n2563 ;
  assign n30812 = ~n9432 & n28548 ;
  assign n30813 = ~n9252 & n30812 ;
  assign n30814 = n10284 | n11715 ;
  assign n30815 = n11536 ^ n3962 ^ 1'b0 ;
  assign n30816 = n15743 | n30815 ;
  assign n30817 = n30814 | n30816 ;
  assign n30818 = ( n14445 & ~n22616 ) | ( n14445 & n30817 ) | ( ~n22616 & n30817 ) ;
  assign n30819 = n637 & ~n12385 ;
  assign n30820 = n11942 | n30819 ;
  assign n30821 = n30818 | n30820 ;
  assign n30822 = ( n8872 & n18435 ) | ( n8872 & n28884 ) | ( n18435 & n28884 ) ;
  assign n30823 = n27864 ^ n19411 ^ 1'b0 ;
  assign n30824 = n1803 | n3392 ;
  assign n30825 = n30824 ^ n16132 ^ x58 ;
  assign n30826 = n2263 & n30825 ;
  assign n30827 = n9994 ^ n693 ^ 1'b0 ;
  assign n30828 = n30494 ^ n30010 ^ n6978 ;
  assign n30829 = ( ~n15727 & n22868 ) | ( ~n15727 & n22948 ) | ( n22868 & n22948 ) ;
  assign n30830 = n9812 & n23843 ;
  assign n30831 = n30830 ^ n15983 ^ 1'b0 ;
  assign n30834 = n5301 & ~n29421 ;
  assign n30832 = ~n1438 & n9141 ;
  assign n30833 = n30832 ^ n16037 ^ 1'b0 ;
  assign n30835 = n30834 ^ n30833 ^ 1'b0 ;
  assign n30836 = ~n22734 & n30835 ;
  assign n30837 = n23494 ^ n11390 ^ 1'b0 ;
  assign n30838 = n19951 ^ n4925 ^ 1'b0 ;
  assign n30839 = n30838 ^ n11872 ^ 1'b0 ;
  assign n30840 = n392 & ~n30839 ;
  assign n30841 = ( n17204 & n26914 ) | ( n17204 & ~n30840 ) | ( n26914 & ~n30840 ) ;
  assign n30844 = n2608 & n25352 ;
  assign n30845 = ~n3356 & n30844 ;
  assign n30843 = ~n8051 & n25274 ;
  assign n30846 = n30845 ^ n30843 ^ 1'b0 ;
  assign n30842 = n8031 & n13851 ;
  assign n30847 = n30846 ^ n30842 ^ 1'b0 ;
  assign n30848 = ~n8312 & n17850 ;
  assign n30849 = n12554 & n30848 ;
  assign n30850 = n16710 & ~n29891 ;
  assign n30851 = n30850 ^ n4313 ^ 1'b0 ;
  assign n30852 = n2946 | n30851 ;
  assign n30853 = n30852 ^ n11796 ^ 1'b0 ;
  assign n30854 = n22726 ^ n19662 ^ 1'b0 ;
  assign n30855 = ~n1108 & n2675 ;
  assign n30856 = n30855 ^ n8390 ^ 1'b0 ;
  assign n30857 = n6037 & ~n30856 ;
  assign n30858 = ~n7903 & n30857 ;
  assign n30859 = n30858 ^ n24052 ^ n5093 ;
  assign n30860 = n28985 ^ n6105 ^ 1'b0 ;
  assign n30861 = n643 & ~n30860 ;
  assign n30862 = n30861 ^ n19743 ^ n4513 ;
  assign n30863 = ~n3675 & n14995 ;
  assign n30864 = ~n11368 & n30863 ;
  assign n30865 = n30864 ^ n17803 ^ n2444 ;
  assign n30866 = n8883 ^ n8323 ^ n3614 ;
  assign n30867 = n4254 & ~n30866 ;
  assign n30868 = n30867 ^ n5259 ^ 1'b0 ;
  assign n30869 = n30868 ^ n14774 ^ n2583 ;
  assign n30870 = n1026 & n14091 ;
  assign n30871 = n1409 | n7087 ;
  assign n30872 = n30870 | n30871 ;
  assign n30873 = n19691 ^ n5488 ^ 1'b0 ;
  assign n30874 = n15228 & n30873 ;
  assign n30875 = n19874 ^ n7342 ^ 1'b0 ;
  assign n30877 = n2048 & ~n18989 ;
  assign n30878 = n6687 & n30877 ;
  assign n30876 = n10922 ^ n6374 ^ 1'b0 ;
  assign n30879 = n30878 ^ n30876 ^ n7531 ;
  assign n30880 = ( ~n3175 & n11364 ) | ( ~n3175 & n30879 ) | ( n11364 & n30879 ) ;
  assign n30881 = n10770 ^ n872 ^ 1'b0 ;
  assign n30882 = ~n12879 & n30881 ;
  assign n30883 = ( n1827 & n2399 ) | ( n1827 & n2508 ) | ( n2399 & n2508 ) ;
  assign n30884 = n30883 ^ n16429 ^ 1'b0 ;
  assign n30885 = n5430 & n30884 ;
  assign n30886 = n19127 ^ n10139 ^ n2154 ;
  assign n30887 = ( n30882 & ~n30885 ) | ( n30882 & n30886 ) | ( ~n30885 & n30886 ) ;
  assign n30888 = n13086 ^ n11886 ^ 1'b0 ;
  assign n30889 = n29844 ^ n23057 ^ n3983 ;
  assign n30892 = n5874 ^ n4898 ^ n1476 ;
  assign n30890 = n14474 ^ n3799 ^ 1'b0 ;
  assign n30891 = n2611 & n30890 ;
  assign n30893 = n30892 ^ n30891 ^ 1'b0 ;
  assign n30894 = n13011 & n29446 ;
  assign n30895 = n7619 & n30894 ;
  assign n30897 = n24602 ^ n4119 ^ 1'b0 ;
  assign n30896 = n6798 | n7905 ;
  assign n30898 = n30897 ^ n30896 ^ 1'b0 ;
  assign n30901 = ( n3083 & ~n4062 ) | ( n3083 & n7367 ) | ( ~n4062 & n7367 ) ;
  assign n30902 = ( n5109 & n9870 ) | ( n5109 & n30901 ) | ( n9870 & n30901 ) ;
  assign n30899 = n2989 & n7482 ;
  assign n30900 = n413 & n30899 ;
  assign n30903 = n30902 ^ n30900 ^ 1'b0 ;
  assign n30904 = ~n11813 & n30903 ;
  assign n30905 = n8704 & n20377 ;
  assign n30906 = ~n15258 & n15334 ;
  assign n30907 = n30906 ^ n3218 ^ 1'b0 ;
  assign n30908 = n21278 | n22171 ;
  assign n30909 = n30907 & n30908 ;
  assign n30910 = n30909 ^ n19711 ^ 1'b0 ;
  assign n30911 = n30910 ^ n24394 ^ 1'b0 ;
  assign n30912 = ~n5274 & n30911 ;
  assign n30913 = n5729 | n5731 ;
  assign n30914 = n30913 ^ n24519 ^ 1'b0 ;
  assign n30915 = n1384 & ~n30914 ;
  assign n30916 = ( n15405 & ~n17971 ) | ( n15405 & n26244 ) | ( ~n17971 & n26244 ) ;
  assign n30917 = n30916 ^ n13488 ^ n9780 ;
  assign n30918 = n30915 & ~n30917 ;
  assign n30919 = n23837 & n30918 ;
  assign n30920 = n18531 ^ n8036 ^ 1'b0 ;
  assign n30921 = n30920 ^ n16203 ^ n3910 ;
  assign n30922 = n27289 ^ n10947 ^ 1'b0 ;
  assign n30923 = ~n20767 & n30922 ;
  assign n30924 = n30923 ^ n14247 ^ n8960 ;
  assign n30930 = n6802 ^ n4779 ^ n3811 ;
  assign n30931 = n28107 & ~n30930 ;
  assign n30925 = n2229 & ~n14979 ;
  assign n30926 = n3338 | n30925 ;
  assign n30927 = n14652 & ~n30926 ;
  assign n30928 = n11903 & ~n25736 ;
  assign n30929 = n30927 & n30928 ;
  assign n30932 = n30931 ^ n30929 ^ n29840 ;
  assign n30933 = n11356 ^ n6897 ^ n2411 ;
  assign n30934 = n20074 ^ n8757 ^ 1'b0 ;
  assign n30935 = ( n1331 & ~n7452 ) | ( n1331 & n19902 ) | ( ~n7452 & n19902 ) ;
  assign n30936 = n1108 & ~n30935 ;
  assign n30937 = n30936 ^ n19822 ^ 1'b0 ;
  assign n30938 = n8177 & n29326 ;
  assign n30939 = n30938 ^ n5485 ^ 1'b0 ;
  assign n30940 = ~n3088 & n3594 ;
  assign n30941 = n30940 ^ n16826 ^ n6297 ;
  assign n30942 = ( n6188 & n30939 ) | ( n6188 & ~n30941 ) | ( n30939 & ~n30941 ) ;
  assign n30943 = n6646 ^ n6145 ^ 1'b0 ;
  assign n30944 = n9961 & ~n24324 ;
  assign n30945 = ( n10457 & ~n30943 ) | ( n10457 & n30944 ) | ( ~n30943 & n30944 ) ;
  assign n30946 = n11953 ^ n7049 ^ 1'b0 ;
  assign n30947 = n9470 & ~n17842 ;
  assign n30948 = n30947 ^ n9234 ^ 1'b0 ;
  assign n30949 = ~n8768 & n16612 ;
  assign n30950 = n30948 & n30949 ;
  assign n30951 = n19125 & ~n26929 ;
  assign n30952 = ~n2450 & n30951 ;
  assign n30953 = ( ~n8103 & n10214 ) | ( ~n8103 & n16048 ) | ( n10214 & n16048 ) ;
  assign n30954 = n7217 ^ n4965 ^ 1'b0 ;
  assign n30955 = n5373 & n30954 ;
  assign n30956 = ( n1915 & n2191 ) | ( n1915 & ~n6299 ) | ( n2191 & ~n6299 ) ;
  assign n30957 = n30956 ^ n25695 ^ n20377 ;
  assign n30958 = n436 & n12278 ;
  assign n30959 = n30958 ^ n8316 ^ 1'b0 ;
  assign n30960 = n30959 ^ n26916 ^ x200 ;
  assign n30961 = n24901 & ~n30960 ;
  assign n30962 = n1745 ^ n398 ^ x129 ;
  assign n30963 = n27539 ^ n14924 ^ 1'b0 ;
  assign n30964 = ~n30962 & n30963 ;
  assign n30965 = n30964 ^ n9083 ^ 1'b0 ;
  assign n30966 = ~n11964 & n30965 ;
  assign n30967 = ~n30961 & n30966 ;
  assign n30968 = n27247 ^ n4156 ^ n542 ;
  assign n30969 = ( n8344 & ~n11088 ) | ( n8344 & n30319 ) | ( ~n11088 & n30319 ) ;
  assign n30970 = n16733 & ~n22374 ;
  assign n30971 = x89 & n2475 ;
  assign n30972 = n2367 & n30971 ;
  assign n30973 = n9756 | n30972 ;
  assign n30974 = n7515 | n30973 ;
  assign n30975 = n10047 & ~n20605 ;
  assign n30976 = ( n7815 & n30974 ) | ( n7815 & n30975 ) | ( n30974 & n30975 ) ;
  assign n30977 = n4675 & ~n30976 ;
  assign n30978 = n30977 ^ n27734 ^ 1'b0 ;
  assign n30979 = n5250 | n14056 ;
  assign n30980 = n30979 ^ n9580 ^ 1'b0 ;
  assign n30981 = n26946 ^ n21264 ^ n19257 ;
  assign n30982 = n9764 ^ n8324 ^ 1'b0 ;
  assign n30983 = n30982 ^ n23928 ^ n8125 ;
  assign n30984 = n5081 | n26902 ;
  assign n30985 = n20028 & ~n30984 ;
  assign n30986 = n22130 ^ n19950 ^ n1497 ;
  assign n30987 = n30986 ^ n13909 ^ n7475 ;
  assign n30988 = n11853 | n21601 ;
  assign n30989 = n5132 & ~n30988 ;
  assign n30990 = n30989 ^ n21948 ^ 1'b0 ;
  assign n30991 = ( n15484 & ~n30987 ) | ( n15484 & n30990 ) | ( ~n30987 & n30990 ) ;
  assign n30992 = n10043 | n22431 ;
  assign n30993 = n355 & ~n13438 ;
  assign n30994 = ~n1270 & n30993 ;
  assign n30995 = n30994 ^ n4577 ^ 1'b0 ;
  assign n30996 = n12249 & ~n30995 ;
  assign n30997 = ( n18730 & n18765 ) | ( n18730 & n30996 ) | ( n18765 & n30996 ) ;
  assign n30998 = n20123 ^ n8125 ^ 1'b0 ;
  assign n30999 = ( ~n992 & n6186 ) | ( ~n992 & n26297 ) | ( n6186 & n26297 ) ;
  assign n31000 = n12421 ^ n5637 ^ 1'b0 ;
  assign n31001 = n20660 | n31000 ;
  assign n31002 = ( ~x56 & n21282 ) | ( ~x56 & n22374 ) | ( n21282 & n22374 ) ;
  assign n31003 = n8368 ^ n2883 ^ 1'b0 ;
  assign n31004 = n4644 & n31003 ;
  assign n31005 = n18351 & ~n31004 ;
  assign n31006 = n9232 ^ n8902 ^ n633 ;
  assign n31007 = n31006 ^ n5060 ^ 1'b0 ;
  assign n31008 = n5376 | n23476 ;
  assign n31009 = n31008 ^ n21453 ^ 1'b0 ;
  assign n31010 = n31009 ^ n8597 ^ n7664 ;
  assign n31011 = n15357 & n31010 ;
  assign n31012 = ~n16822 & n31011 ;
  assign n31013 = n31012 ^ n18582 ^ 1'b0 ;
  assign n31014 = n28109 ^ n18774 ^ n3709 ;
  assign n31015 = n31014 ^ n7170 ^ 1'b0 ;
  assign n31016 = n5455 ^ n3633 ^ 1'b0 ;
  assign n31017 = n31015 & n31016 ;
  assign n31018 = ( n5539 & ~n14409 ) | ( n5539 & n20904 ) | ( ~n14409 & n20904 ) ;
  assign n31019 = x185 & n31018 ;
  assign n31026 = ( x122 & n7574 ) | ( x122 & n13414 ) | ( n7574 & n13414 ) ;
  assign n31020 = n15212 ^ n9294 ^ 1'b0 ;
  assign n31021 = ( n2846 & ~n6101 ) | ( n2846 & n31020 ) | ( ~n6101 & n31020 ) ;
  assign n31022 = n6870 & n20245 ;
  assign n31023 = ~n31021 & n31022 ;
  assign n31024 = n5360 | n31023 ;
  assign n31025 = n20410 | n31024 ;
  assign n31027 = n31026 ^ n31025 ^ n6204 ;
  assign n31029 = n29707 ^ n26472 ^ n21313 ;
  assign n31028 = n10597 & ~n16288 ;
  assign n31030 = n31029 ^ n31028 ^ 1'b0 ;
  assign n31031 = ~n1009 & n17224 ;
  assign n31032 = n11383 ^ n6000 ^ n4564 ;
  assign n31033 = n31032 ^ n24394 ^ 1'b0 ;
  assign n31034 = n31031 & n31033 ;
  assign n31035 = n481 & ~n8621 ;
  assign n31036 = n31035 ^ n329 ^ 1'b0 ;
  assign n31037 = n25854 ^ n7180 ^ 1'b0 ;
  assign n31038 = n27074 & ~n31037 ;
  assign n31039 = n31036 & n31038 ;
  assign n31040 = ~n19574 & n25369 ;
  assign n31041 = n31040 ^ n2573 ^ 1'b0 ;
  assign n31042 = ( n379 & n881 ) | ( n379 & ~n10760 ) | ( n881 & ~n10760 ) ;
  assign n31043 = n13675 & n31042 ;
  assign n31044 = ~x167 & n31043 ;
  assign n31045 = ~n31041 & n31044 ;
  assign n31046 = n2036 & ~n16667 ;
  assign n31047 = n11727 & n31046 ;
  assign n31048 = n19261 ^ n15805 ^ 1'b0 ;
  assign n31049 = ~n31047 & n31048 ;
  assign n31050 = n2336 & n10722 ;
  assign n31051 = ( ~n8276 & n31049 ) | ( ~n8276 & n31050 ) | ( n31049 & n31050 ) ;
  assign n31052 = n8943 ^ n5157 ^ 1'b0 ;
  assign n31053 = n3256 & ~n4571 ;
  assign n31054 = n31053 ^ n21122 ^ n11069 ;
  assign n31055 = n31054 ^ n9087 ^ 1'b0 ;
  assign n31056 = ( n26096 & n31052 ) | ( n26096 & ~n31055 ) | ( n31052 & ~n31055 ) ;
  assign n31057 = ~n6047 & n14486 ;
  assign n31058 = n12063 | n31057 ;
  assign n31059 = n4319 & ~n31058 ;
  assign n31060 = x200 & n21028 ;
  assign n31061 = n31060 ^ n17999 ^ n11579 ;
  assign n31062 = ~n8411 & n27578 ;
  assign n31063 = ~n31061 & n31062 ;
  assign n31064 = ( ~n4870 & n5662 ) | ( ~n4870 & n22256 ) | ( n5662 & n22256 ) ;
  assign n31065 = n31064 ^ n12952 ^ 1'b0 ;
  assign n31066 = n31065 ^ n3469 ^ n3200 ;
  assign n31067 = n4516 ^ n1569 ^ 1'b0 ;
  assign n31069 = ~n5384 & n8359 ;
  assign n31068 = n19193 | n28743 ;
  assign n31070 = n31069 ^ n31068 ^ 1'b0 ;
  assign n31071 = ( n1753 & n13854 ) | ( n1753 & n16982 ) | ( n13854 & n16982 ) ;
  assign n31072 = ( n10579 & ~n21863 ) | ( n10579 & n31071 ) | ( ~n21863 & n31071 ) ;
  assign n31073 = n4138 & n6634 ;
  assign n31074 = n31073 ^ n21099 ^ n20445 ;
  assign n31075 = n8560 | n10655 ;
  assign n31076 = ( x98 & n1701 ) | ( x98 & n10702 ) | ( n1701 & n10702 ) ;
  assign n31077 = n11096 & ~n18763 ;
  assign n31078 = n31076 & n31077 ;
  assign n31079 = n8791 & ~n18493 ;
  assign n31080 = n31079 ^ n4342 ^ 1'b0 ;
  assign n31081 = n4998 & n17961 ;
  assign n31082 = n14331 ^ n2319 ^ 1'b0 ;
  assign n31083 = n15173 & ~n31082 ;
  assign n31084 = ~n6240 & n31083 ;
  assign n31085 = n6848 & n31084 ;
  assign n31086 = n17881 | n31085 ;
  assign n31087 = n31086 ^ n12363 ^ 1'b0 ;
  assign n31088 = ~n3433 & n24049 ;
  assign n31089 = ~n31087 & n31088 ;
  assign n31090 = n25413 ^ n1221 ^ 1'b0 ;
  assign n31091 = n9320 & n31090 ;
  assign n31092 = ( n3952 & n24670 ) | ( n3952 & n31091 ) | ( n24670 & n31091 ) ;
  assign n31093 = ( n6133 & n9061 ) | ( n6133 & n10183 ) | ( n9061 & n10183 ) ;
  assign n31094 = n31093 ^ n18233 ^ n11669 ;
  assign n31095 = ~n4996 & n14275 ;
  assign n31096 = n5589 | n17723 ;
  assign n31097 = n31096 ^ n12837 ^ 1'b0 ;
  assign n31098 = n29625 & ~n31097 ;
  assign n31099 = n31098 ^ n7367 ^ 1'b0 ;
  assign n31100 = n31099 ^ n13963 ^ 1'b0 ;
  assign n31101 = ~n19530 & n29534 ;
  assign n31102 = n30701 & n31101 ;
  assign n31103 = ~n7217 & n10152 ;
  assign n31104 = n31103 ^ n24208 ^ 1'b0 ;
  assign n31105 = ~n8588 & n31104 ;
  assign n31106 = n4912 & ~n9746 ;
  assign n31107 = ~n16179 & n31106 ;
  assign n31108 = n3666 & n7786 ;
  assign n31109 = n31108 ^ n8369 ^ 1'b0 ;
  assign n31110 = n31109 ^ n864 ^ 1'b0 ;
  assign n31111 = n31107 & n31110 ;
  assign n31112 = n10846 & n31111 ;
  assign n31113 = n10109 & ~n24717 ;
  assign n31114 = ~n22098 & n31113 ;
  assign n31115 = n5046 | n24719 ;
  assign n31116 = n8960 | n31115 ;
  assign n31117 = n3387 & n15240 ;
  assign n31118 = n10078 ^ n6188 ^ 1'b0 ;
  assign n31119 = n28716 & n31118 ;
  assign n31120 = n31119 ^ n15388 ^ n5744 ;
  assign n31121 = ( n19501 & n31117 ) | ( n19501 & n31120 ) | ( n31117 & n31120 ) ;
  assign n31123 = n4359 & n6480 ;
  assign n31122 = ~n19445 & n21042 ;
  assign n31124 = n31123 ^ n31122 ^ 1'b0 ;
  assign n31125 = n30483 ^ n19421 ^ 1'b0 ;
  assign n31126 = ~n31124 & n31125 ;
  assign n31127 = ( n15630 & n29591 ) | ( n15630 & n31126 ) | ( n29591 & n31126 ) ;
  assign n31128 = n14522 ^ n8793 ^ 1'b0 ;
  assign n31129 = n31128 ^ n14806 ^ n12446 ;
  assign n31130 = n10555 ^ n4107 ^ 1'b0 ;
  assign n31131 = n2966 & ~n13698 ;
  assign n31132 = n13915 ^ n12186 ^ 1'b0 ;
  assign n31133 = n3191 & n31132 ;
  assign n31134 = ( ~n1483 & n10517 ) | ( ~n1483 & n19815 ) | ( n10517 & n19815 ) ;
  assign n31135 = n13593 | n31134 ;
  assign n31136 = n31133 | n31135 ;
  assign n31137 = ~n13999 & n29809 ;
  assign n31138 = n18842 ^ n11070 ^ 1'b0 ;
  assign n31139 = n1776 | n31138 ;
  assign n31140 = n20404 ^ n9981 ^ 1'b0 ;
  assign n31141 = ~n1906 & n31140 ;
  assign n31142 = n31139 & ~n31141 ;
  assign n31143 = n24803 & n31142 ;
  assign n31144 = ~n21987 & n31143 ;
  assign n31145 = ( n2977 & n15728 ) | ( n2977 & ~n26375 ) | ( n15728 & ~n26375 ) ;
  assign n31146 = ~n16890 & n31145 ;
  assign n31147 = n31146 ^ n14927 ^ 1'b0 ;
  assign n31151 = n28846 ^ n15054 ^ n12832 ;
  assign n31150 = n23910 & n25861 ;
  assign n31152 = n31151 ^ n31150 ^ 1'b0 ;
  assign n31148 = n10405 ^ n8478 ^ n1634 ;
  assign n31149 = n8170 | n31148 ;
  assign n31153 = n31152 ^ n31149 ^ 1'b0 ;
  assign n31155 = n13760 ^ n5044 ^ n3872 ;
  assign n31154 = n12418 ^ n2841 ^ 1'b0 ;
  assign n31156 = n31155 ^ n31154 ^ n14579 ;
  assign n31157 = n17505 ^ n17410 ^ n4890 ;
  assign n31158 = n5126 & n11907 ;
  assign n31159 = n31158 ^ n24254 ^ n2165 ;
  assign n31160 = n4413 ^ n2823 ^ 1'b0 ;
  assign n31161 = n3173 & n31160 ;
  assign n31162 = ~n1438 & n31161 ;
  assign n31163 = ( n9024 & n11765 ) | ( n9024 & n24397 ) | ( n11765 & n24397 ) ;
  assign n31164 = n6108 & ~n31163 ;
  assign n31165 = n8291 ^ n6984 ^ 1'b0 ;
  assign n31166 = ( n6237 & n12277 ) | ( n6237 & n31165 ) | ( n12277 & n31165 ) ;
  assign n31167 = ( ~n10957 & n22047 ) | ( ~n10957 & n31166 ) | ( n22047 & n31166 ) ;
  assign n31168 = n31167 ^ n12356 ^ 1'b0 ;
  assign n31169 = ( n9458 & n26096 ) | ( n9458 & n27937 ) | ( n26096 & n27937 ) ;
  assign n31170 = n31168 | n31169 ;
  assign n31171 = n31164 & ~n31170 ;
  assign n31172 = ( n1537 & ~n8916 ) | ( n1537 & n9432 ) | ( ~n8916 & n9432 ) ;
  assign n31173 = n11776 ^ n9552 ^ n5522 ;
  assign n31174 = n7306 & n30770 ;
  assign n31175 = n31174 ^ n16198 ^ 1'b0 ;
  assign n31176 = n30320 ^ n25018 ^ 1'b0 ;
  assign n31177 = n31175 | n31176 ;
  assign n31178 = ( n13107 & n13814 ) | ( n13107 & n23352 ) | ( n13814 & n23352 ) ;
  assign n31179 = n7079 & ~n31178 ;
  assign n31180 = n13841 & n31179 ;
  assign n31181 = ( n413 & n7151 ) | ( n413 & ~n31180 ) | ( n7151 & ~n31180 ) ;
  assign n31182 = ( n9401 & ~n21624 ) | ( n9401 & n31181 ) | ( ~n21624 & n31181 ) ;
  assign n31185 = n19438 & ~n20266 ;
  assign n31186 = ~x180 & n31185 ;
  assign n31187 = n6699 & ~n31186 ;
  assign n31188 = n31187 ^ n8676 ^ 1'b0 ;
  assign n31183 = ( n8247 & ~n10529 ) | ( n8247 & n28810 ) | ( ~n10529 & n28810 ) ;
  assign n31184 = ~n11478 & n31183 ;
  assign n31189 = n31188 ^ n31184 ^ 1'b0 ;
  assign n31190 = n31189 ^ n19098 ^ n15559 ;
  assign n31191 = n6624 & ~n29729 ;
  assign n31192 = n702 | n20679 ;
  assign n31193 = n31192 ^ n8477 ^ 1'b0 ;
  assign n31194 = ~n29538 & n31193 ;
  assign n31195 = ~n13066 & n31194 ;
  assign n31196 = n1535 ^ n707 ^ 1'b0 ;
  assign n31197 = ( x65 & n12219 ) | ( x65 & ~n19359 ) | ( n12219 & ~n19359 ) ;
  assign n31205 = n9050 ^ n1104 ^ 1'b0 ;
  assign n31203 = n18924 | n19931 ;
  assign n31204 = n31203 ^ n18063 ^ 1'b0 ;
  assign n31198 = ( ~n5438 & n10283 ) | ( ~n5438 & n19674 ) | ( n10283 & n19674 ) ;
  assign n31199 = n30559 ^ n12480 ^ n9595 ;
  assign n31200 = ( n3034 & n7841 ) | ( n3034 & ~n31199 ) | ( n7841 & ~n31199 ) ;
  assign n31201 = ~n31198 & n31200 ;
  assign n31202 = n31201 ^ n27849 ^ 1'b0 ;
  assign n31206 = n31205 ^ n31204 ^ n31202 ;
  assign n31207 = ~n799 & n30554 ;
  assign n31208 = n31207 ^ n8019 ^ 1'b0 ;
  assign n31209 = ( ~n3411 & n6672 ) | ( ~n3411 & n7551 ) | ( n6672 & n7551 ) ;
  assign n31210 = n23979 | n31209 ;
  assign n31211 = n5526 & n7790 ;
  assign n31212 = ~n24275 & n31211 ;
  assign n31213 = n12205 ^ n7827 ^ n5538 ;
  assign n31214 = n10251 & ~n21562 ;
  assign n31215 = n31214 ^ n21581 ^ 1'b0 ;
  assign n31216 = ( n4958 & n31213 ) | ( n4958 & ~n31215 ) | ( n31213 & ~n31215 ) ;
  assign n31217 = n5970 & ~n31216 ;
  assign n31218 = ~n21413 & n31217 ;
  assign n31221 = n24240 ^ n22301 ^ n13177 ;
  assign n31219 = n24885 ^ n6697 ^ 1'b0 ;
  assign n31220 = n26868 & ~n31219 ;
  assign n31222 = n31221 ^ n31220 ^ n14075 ;
  assign n31223 = n1421 & n24299 ;
  assign n31224 = n2191 | n10204 ;
  assign n31225 = n31224 ^ n28596 ^ n414 ;
  assign n31226 = n19446 ^ n12771 ^ n3437 ;
  assign n31227 = n31226 ^ n3638 ^ 1'b0 ;
  assign n31228 = n9549 | n28685 ;
  assign n31229 = n24257 & n24299 ;
  assign n31230 = n31229 ^ n19255 ^ 1'b0 ;
  assign n31231 = ~n31228 & n31230 ;
  assign n31232 = ~n31227 & n31231 ;
  assign n31233 = n2954 & ~n3804 ;
  assign n31234 = n31233 ^ n998 ^ 1'b0 ;
  assign n31235 = n31234 ^ n10813 ^ n4575 ;
  assign n31239 = n6502 & n9347 ;
  assign n31240 = ~n693 & n31239 ;
  assign n31237 = n857 | n2084 ;
  assign n31238 = n31237 ^ n7169 ^ 1'b0 ;
  assign n31241 = n31240 ^ n31238 ^ n14721 ;
  assign n31242 = n31241 ^ n5561 ^ 1'b0 ;
  assign n31243 = n31242 ^ n12121 ^ n10793 ;
  assign n31236 = ( n4287 & ~n6821 ) | ( n4287 & n9521 ) | ( ~n6821 & n9521 ) ;
  assign n31244 = n31243 ^ n31236 ^ 1'b0 ;
  assign n31245 = n15970 | n31244 ;
  assign n31246 = n31245 ^ n13466 ^ 1'b0 ;
  assign n31247 = n25985 ^ n14789 ^ n6854 ;
  assign n31249 = n7562 ^ n3206 ^ n3009 ;
  assign n31248 = n4255 | n16705 ;
  assign n31250 = n31249 ^ n31248 ^ 1'b0 ;
  assign n31251 = ( n3872 & n4848 ) | ( n3872 & n15254 ) | ( n4848 & n15254 ) ;
  assign n31252 = ( n2422 & ~n28166 ) | ( n2422 & n31251 ) | ( ~n28166 & n31251 ) ;
  assign n31253 = ( n2843 & n7127 ) | ( n2843 & ~n31252 ) | ( n7127 & ~n31252 ) ;
  assign n31254 = n7856 | n31253 ;
  assign n31255 = n31254 ^ n26522 ^ 1'b0 ;
  assign n31256 = ~n7843 & n31255 ;
  assign n31257 = n690 & n17306 ;
  assign n31258 = n3466 ^ n855 ^ 1'b0 ;
  assign n31259 = ~n11778 & n31258 ;
  assign n31260 = ~n23777 & n31259 ;
  assign n31261 = ~n24373 & n31260 ;
  assign n31262 = ( ~n27889 & n31243 ) | ( ~n27889 & n31261 ) | ( n31243 & n31261 ) ;
  assign n31263 = n28877 ^ n7689 ^ n5261 ;
  assign n31264 = n31263 ^ n22034 ^ 1'b0 ;
  assign n31265 = n2638 & n31264 ;
  assign n31266 = n24413 ^ n11857 ^ 1'b0 ;
  assign n31267 = ~n2151 & n31266 ;
  assign n31271 = n2624 & ~n7254 ;
  assign n31269 = x107 & n13760 ;
  assign n31270 = n31269 ^ n10442 ^ 1'b0 ;
  assign n31268 = n22933 | n24192 ;
  assign n31272 = n31271 ^ n31270 ^ n31268 ;
  assign n31273 = n7396 & n31037 ;
  assign n31274 = n31273 ^ n16699 ^ n15961 ;
  assign n31275 = n10788 | n11913 ;
  assign n31276 = n31275 ^ n3982 ^ 1'b0 ;
  assign n31277 = n31276 ^ n27851 ^ n24067 ;
  assign n31278 = n31277 ^ n10004 ^ 1'b0 ;
  assign n31279 = ( ~n4573 & n29304 ) | ( ~n4573 & n31278 ) | ( n29304 & n31278 ) ;
  assign n31280 = ( n17958 & n18032 ) | ( n17958 & ~n18106 ) | ( n18032 & ~n18106 ) ;
  assign n31286 = n30255 ^ n4769 ^ n3264 ;
  assign n31285 = n18330 ^ n16213 ^ n6626 ;
  assign n31287 = n31286 ^ n31285 ^ 1'b0 ;
  assign n31281 = ~n1578 & n7073 ;
  assign n31282 = n26026 ^ n7412 ^ 1'b0 ;
  assign n31283 = n31281 | n31282 ;
  assign n31284 = n10305 & ~n31283 ;
  assign n31288 = n31287 ^ n31284 ^ 1'b0 ;
  assign n31289 = n17671 ^ n806 ^ 1'b0 ;
  assign n31290 = n8433 | n31289 ;
  assign n31291 = n27043 ^ n26944 ^ n4382 ;
  assign n31292 = n31291 ^ n23661 ^ 1'b0 ;
  assign n31293 = n31290 | n31292 ;
  assign n31294 = n13768 ^ n5909 ^ 1'b0 ;
  assign n31295 = n5337 ^ n733 ^ 1'b0 ;
  assign n31296 = n31295 ^ n4023 ^ 1'b0 ;
  assign n31297 = n13499 ^ n468 ^ 1'b0 ;
  assign n31298 = n9603 & n31297 ;
  assign n31299 = n10860 ^ n9252 ^ 1'b0 ;
  assign n31300 = n3736 & ~n31299 ;
  assign n31301 = n31298 & n31300 ;
  assign n31302 = n31296 & n31301 ;
  assign n31303 = n10223 & n16555 ;
  assign n31304 = n976 & n31303 ;
  assign n31305 = n31304 ^ n23691 ^ 1'b0 ;
  assign n31306 = n4552 | n5795 ;
  assign n31307 = n584 & n11606 ;
  assign n31308 = n31307 ^ n28196 ^ n20237 ;
  assign n31309 = n15054 ^ n2267 ^ 1'b0 ;
  assign n31310 = ~n2220 & n31309 ;
  assign n31311 = ~n15335 & n23880 ;
  assign n31312 = n31311 ^ n4708 ^ 1'b0 ;
  assign n31313 = ( n3032 & ~n17329 ) | ( n3032 & n18084 ) | ( ~n17329 & n18084 ) ;
  assign n31314 = n26142 ^ n1344 ^ 1'b0 ;
  assign n31315 = n4535 & n11332 ;
  assign n31316 = n17509 ^ n14458 ^ 1'b0 ;
  assign n31317 = ( n31314 & n31315 ) | ( n31314 & n31316 ) | ( n31315 & n31316 ) ;
  assign n31318 = ~n5300 & n6060 ;
  assign n31319 = n31318 ^ n10400 ^ n9391 ;
  assign n31320 = n31319 ^ n11357 ^ 1'b0 ;
  assign n31321 = n14658 & ~n16258 ;
  assign n31322 = n31321 ^ n12015 ^ 1'b0 ;
  assign n31323 = n19236 ^ n7138 ^ 1'b0 ;
  assign n31324 = ( n31320 & n31322 ) | ( n31320 & ~n31323 ) | ( n31322 & ~n31323 ) ;
  assign n31326 = ~n6323 & n25385 ;
  assign n31325 = n11940 ^ n8574 ^ x228 ;
  assign n31327 = n31326 ^ n31325 ^ 1'b0 ;
  assign n31328 = ~n7049 & n31327 ;
  assign n31329 = n3604 | n26540 ;
  assign n31330 = n455 & n17743 ;
  assign n31331 = n31330 ^ n16317 ^ 1'b0 ;
  assign n31332 = n293 & ~n31331 ;
  assign n31333 = n18854 & n31332 ;
  assign n31334 = ( n11925 & ~n13380 ) | ( n11925 & n30046 ) | ( ~n13380 & n30046 ) ;
  assign n31335 = n31334 ^ n11079 ^ 1'b0 ;
  assign n31336 = n15281 ^ n6247 ^ n4952 ;
  assign n31337 = n11294 | n31336 ;
  assign n31338 = ~n1345 & n4585 ;
  assign n31339 = n31338 ^ n4881 ^ 1'b0 ;
  assign n31340 = n31337 | n31339 ;
  assign n31341 = ( n1037 & n4490 ) | ( n1037 & ~n7947 ) | ( n4490 & ~n7947 ) ;
  assign n31342 = ~n2924 & n31341 ;
  assign n31343 = n21354 ^ n19981 ^ 1'b0 ;
  assign n31344 = ~n9997 & n31343 ;
  assign n31345 = n31344 ^ n15067 ^ 1'b0 ;
  assign n31346 = n24619 ^ n16058 ^ n12327 ;
  assign n31347 = n31346 ^ n13777 ^ n2365 ;
  assign n31348 = n31347 ^ n12031 ^ 1'b0 ;
  assign n31349 = n18774 & ~n31348 ;
  assign n31350 = ( n1493 & ~n25070 ) | ( n1493 & n27263 ) | ( ~n25070 & n27263 ) ;
  assign n31351 = n11173 & ~n16616 ;
  assign n31352 = n31351 ^ n9655 ^ 1'b0 ;
  assign n31353 = n18634 | n31352 ;
  assign n31354 = n31352 & ~n31353 ;
  assign n31355 = n1867 & ~n31354 ;
  assign n31356 = ~n31350 & n31355 ;
  assign n31357 = n1081 & ~n7489 ;
  assign n31358 = n27704 & n31357 ;
  assign n31359 = n17442 ^ n2075 ^ n1360 ;
  assign n31360 = ( ~n1435 & n28806 ) | ( ~n1435 & n31359 ) | ( n28806 & n31359 ) ;
  assign n31361 = n31360 ^ n23110 ^ n15809 ;
  assign n31362 = n18178 ^ n1900 ^ 1'b0 ;
  assign n31363 = n31361 & n31362 ;
  assign n31364 = ( n14714 & ~n25951 ) | ( n14714 & n31363 ) | ( ~n25951 & n31363 ) ;
  assign n31365 = n14695 ^ n10678 ^ n3627 ;
  assign n31366 = ~n5905 & n30513 ;
  assign n31367 = ~n31365 & n31366 ;
  assign n31368 = n10769 ^ n4171 ^ 1'b0 ;
  assign n31369 = ~n413 & n31368 ;
  assign n31370 = n31369 ^ n6266 ^ 1'b0 ;
  assign n31371 = n17572 & n31370 ;
  assign n31372 = n14022 & ~n31371 ;
  assign n31373 = n19169 ^ n9580 ^ n3436 ;
  assign n31374 = ~n17386 & n31373 ;
  assign n31375 = n31374 ^ n7878 ^ 1'b0 ;
  assign n31376 = x67 | n31375 ;
  assign n31377 = n31376 ^ n14780 ^ 1'b0 ;
  assign n31378 = ( ~n5221 & n17614 ) | ( ~n5221 & n23784 ) | ( n17614 & n23784 ) ;
  assign n31379 = ( ~n3579 & n9746 ) | ( ~n3579 & n20749 ) | ( n9746 & n20749 ) ;
  assign n31380 = n31379 ^ n17120 ^ n9595 ;
  assign n31381 = n6331 | n31380 ;
  assign n31382 = n16230 ^ n6531 ^ 1'b0 ;
  assign n31383 = n2398 & n31382 ;
  assign n31384 = n20423 ^ n8470 ^ 1'b0 ;
  assign n31385 = n5125 | n31384 ;
  assign n31386 = n12031 | n31385 ;
  assign n31387 = n31383 & n31386 ;
  assign n31388 = n1884 & n31387 ;
  assign n31389 = n16662 & n23373 ;
  assign n31390 = n31389 ^ n10181 ^ 1'b0 ;
  assign n31391 = n31390 ^ x84 ^ 1'b0 ;
  assign n31392 = n31388 | n31391 ;
  assign n31393 = n13679 ^ n7537 ^ 1'b0 ;
  assign n31394 = n12335 & ~n31393 ;
  assign n31395 = ~n7089 & n31394 ;
  assign n31396 = ~n3160 & n31395 ;
  assign n31397 = n14098 ^ n11058 ^ 1'b0 ;
  assign n31398 = n19982 ^ n3742 ^ 1'b0 ;
  assign n31399 = n15864 | n31398 ;
  assign n31402 = n757 | n12479 ;
  assign n31403 = n31402 ^ n27930 ^ n5125 ;
  assign n31400 = n14737 ^ n10911 ^ n2131 ;
  assign n31401 = n31400 ^ n23472 ^ n17883 ;
  assign n31404 = n31403 ^ n31401 ^ n23076 ;
  assign n31405 = ( n1909 & n6479 ) | ( n1909 & ~n31404 ) | ( n6479 & ~n31404 ) ;
  assign n31406 = ( n2914 & ~n7058 ) | ( n2914 & n13566 ) | ( ~n7058 & n13566 ) ;
  assign n31407 = ( n1934 & n29258 ) | ( n1934 & n31406 ) | ( n29258 & n31406 ) ;
  assign n31408 = n31407 ^ n20281 ^ n3823 ;
  assign n31410 = ( n3503 & n6533 ) | ( n3503 & n12384 ) | ( n6533 & n12384 ) ;
  assign n31411 = n3937 & ~n31410 ;
  assign n31412 = ~n1901 & n31411 ;
  assign n31413 = n26968 & ~n31412 ;
  assign n31409 = n17681 & n27990 ;
  assign n31414 = n31413 ^ n31409 ^ 1'b0 ;
  assign n31415 = n7207 | n16782 ;
  assign n31416 = n31415 ^ n7356 ^ 1'b0 ;
  assign n31417 = n16319 ^ n8842 ^ n3687 ;
  assign n31418 = n31417 ^ n20508 ^ 1'b0 ;
  assign n31419 = x109 & ~n31418 ;
  assign n31420 = n1273 & n14848 ;
  assign n31421 = n31420 ^ n23001 ^ n20573 ;
  assign n31422 = n21862 ^ n20377 ^ n7178 ;
  assign n31423 = n14212 ^ n12000 ^ 1'b0 ;
  assign n31424 = n2254 | n22805 ;
  assign n31425 = ( ~n5080 & n9484 ) | ( ~n5080 & n12646 ) | ( n9484 & n12646 ) ;
  assign n31426 = n31425 ^ n9361 ^ 1'b0 ;
  assign n31427 = n31424 & ~n31426 ;
  assign n31428 = n3444 | n21305 ;
  assign n31429 = n31428 ^ n28773 ^ n5251 ;
  assign n31430 = n17958 ^ n5367 ^ 1'b0 ;
  assign n31431 = n31430 ^ n2182 ^ 1'b0 ;
  assign n31432 = n5902 & ~n6659 ;
  assign n31433 = n6145 ^ n5926 ^ 1'b0 ;
  assign n31434 = n31433 ^ n14715 ^ n7115 ;
  assign n31435 = n12143 & ~n31434 ;
  assign n31436 = n31435 ^ x159 ^ 1'b0 ;
  assign n31437 = ~n11865 & n31436 ;
  assign n31438 = n31437 ^ n29154 ^ n12970 ;
  assign n31439 = n277 & n9994 ;
  assign n31440 = n31439 ^ n8520 ^ 1'b0 ;
  assign n31441 = n15143 & ~n31440 ;
  assign n31442 = n31441 ^ n19540 ^ 1'b0 ;
  assign n31443 = n3048 & n31442 ;
  assign n31444 = ( n9789 & n17493 ) | ( n9789 & ~n21936 ) | ( n17493 & ~n21936 ) ;
  assign n31449 = n9448 ^ n7635 ^ 1'b0 ;
  assign n31450 = n23612 | n31449 ;
  assign n31446 = n17500 ^ n8936 ^ n435 ;
  assign n31445 = n11008 & ~n18769 ;
  assign n31447 = n31446 ^ n31445 ^ 1'b0 ;
  assign n31448 = n25777 & ~n31447 ;
  assign n31451 = n31450 ^ n31448 ^ 1'b0 ;
  assign n31452 = n11089 ^ n9016 ^ 1'b0 ;
  assign n31453 = n9379 | n10851 ;
  assign n31454 = n7785 | n18084 ;
  assign n31455 = n4789 & ~n31454 ;
  assign n31459 = ~n3219 & n19304 ;
  assign n31457 = n19953 ^ n3573 ^ n2935 ;
  assign n31456 = n12135 ^ n10741 ^ 1'b0 ;
  assign n31458 = n31457 ^ n31456 ^ n1995 ;
  assign n31460 = n31459 ^ n31458 ^ n25974 ;
  assign n31461 = n21555 ^ n4536 ^ 1'b0 ;
  assign n31462 = ( ~n25419 & n28089 ) | ( ~n25419 & n31461 ) | ( n28089 & n31461 ) ;
  assign n31463 = ( ~n17764 & n18331 ) | ( ~n17764 & n24324 ) | ( n18331 & n24324 ) ;
  assign n31464 = n31463 ^ n16231 ^ n1482 ;
  assign n31465 = ( n6304 & n26148 ) | ( n6304 & n27947 ) | ( n26148 & n27947 ) ;
  assign n31466 = n22526 & n30204 ;
  assign n31467 = n31466 ^ n4757 ^ 1'b0 ;
  assign n31468 = ( n5191 & n12479 ) | ( n5191 & ~n16403 ) | ( n12479 & ~n16403 ) ;
  assign n31469 = n24523 | n31468 ;
  assign n31470 = n10878 ^ n1461 ^ 1'b0 ;
  assign n31471 = ~n5724 & n16154 ;
  assign n31472 = n6964 & n31471 ;
  assign n31475 = ( ~n4394 & n14511 ) | ( ~n4394 & n26192 ) | ( n14511 & n26192 ) ;
  assign n31473 = n21795 ^ n8024 ^ n7633 ;
  assign n31474 = n31473 ^ n17323 ^ n1736 ;
  assign n31476 = n31475 ^ n31474 ^ 1'b0 ;
  assign n31477 = n5341 & ~n31476 ;
  assign n31480 = ~n3697 & n25170 ;
  assign n31478 = n9433 & ~n27204 ;
  assign n31479 = n21111 & n31478 ;
  assign n31481 = n31480 ^ n31479 ^ 1'b0 ;
  assign n31482 = ~n13225 & n27388 ;
  assign n31483 = ~n1574 & n31482 ;
  assign n31484 = n4338 | n28014 ;
  assign n31485 = n31484 ^ n15795 ^ 1'b0 ;
  assign n31486 = ( ~n9405 & n27540 ) | ( ~n9405 & n31485 ) | ( n27540 & n31485 ) ;
  assign n31487 = n2694 ^ n1155 ^ 1'b0 ;
  assign n31488 = n31487 ^ n19982 ^ 1'b0 ;
  assign n31489 = ~n11782 & n31488 ;
  assign n31490 = ( n3810 & n4890 ) | ( n3810 & n14491 ) | ( n4890 & n14491 ) ;
  assign n31491 = n17921 & n31490 ;
  assign n31492 = ~n1662 & n31491 ;
  assign n31493 = n10945 ^ n297 ^ 1'b0 ;
  assign n31494 = n31492 | n31493 ;
  assign n31495 = n31489 & n31494 ;
  assign n31496 = n29596 ^ n19655 ^ n4113 ;
  assign n31497 = n6538 | n19525 ;
  assign n31498 = ( n8568 & n31496 ) | ( n8568 & n31497 ) | ( n31496 & n31497 ) ;
  assign n31502 = ( ~n3970 & n5207 ) | ( ~n3970 & n26866 ) | ( n5207 & n26866 ) ;
  assign n31500 = n12895 ^ n1808 ^ 1'b0 ;
  assign n31501 = n31500 ^ n18759 ^ 1'b0 ;
  assign n31499 = n26408 ^ n1385 ^ 1'b0 ;
  assign n31503 = n31502 ^ n31501 ^ n31499 ;
  assign n31504 = ( ~n1080 & n25482 ) | ( ~n1080 & n29426 ) | ( n25482 & n29426 ) ;
  assign n31505 = n26015 | n31504 ;
  assign n31506 = n15414 | n31505 ;
  assign n31507 = n31506 ^ n7970 ^ 1'b0 ;
  assign n31511 = n15237 ^ n4986 ^ 1'b0 ;
  assign n31512 = n12900 & n31511 ;
  assign n31508 = ( n676 & n20904 ) | ( n676 & n22096 ) | ( n20904 & n22096 ) ;
  assign n31509 = n12229 & ~n31508 ;
  assign n31510 = n31509 ^ n468 ^ 1'b0 ;
  assign n31513 = n31512 ^ n31510 ^ n5418 ;
  assign n31514 = n4575 | n12849 ;
  assign n31515 = n31514 ^ n31076 ^ n17787 ;
  assign n31516 = n26619 & ~n31515 ;
  assign n31517 = n31516 ^ n22989 ^ 1'b0 ;
  assign n31519 = ( n2795 & ~n7110 ) | ( n2795 & n18273 ) | ( ~n7110 & n18273 ) ;
  assign n31518 = ~n8754 & n12551 ;
  assign n31520 = n31519 ^ n31518 ^ 1'b0 ;
  assign n31521 = ~n28536 & n31520 ;
  assign n31522 = n31521 ^ n9394 ^ 1'b0 ;
  assign n31523 = n1108 | n9455 ;
  assign n31524 = ~n9175 & n31523 ;
  assign n31525 = ( n21169 & ~n31304 ) | ( n21169 & n31524 ) | ( ~n31304 & n31524 ) ;
  assign n31526 = n15263 ^ n7782 ^ 1'b0 ;
  assign n31527 = ~n29171 & n31526 ;
  assign n31528 = n12876 & ~n17846 ;
  assign n31529 = n31528 ^ n1716 ^ 1'b0 ;
  assign n31530 = n31529 ^ n29756 ^ 1'b0 ;
  assign n31531 = n2388 | n31530 ;
  assign n31532 = n7870 ^ n528 ^ 1'b0 ;
  assign n31533 = n17729 ^ n12331 ^ n2702 ;
  assign n31534 = ~n31532 & n31533 ;
  assign n31535 = n31531 & n31534 ;
  assign n31536 = n5641 & n13025 ;
  assign n31537 = n31536 ^ n29454 ^ 1'b0 ;
  assign n31538 = ~n2783 & n12266 ;
  assign n31539 = n31538 ^ n28473 ^ 1'b0 ;
  assign n31540 = n17890 ^ n5236 ^ 1'b0 ;
  assign n31541 = n10464 & ~n31540 ;
  assign n31542 = n7098 | n10056 ;
  assign n31543 = n2263 & ~n31542 ;
  assign n31544 = n25027 & ~n31543 ;
  assign n31545 = ( n31539 & n31541 ) | ( n31539 & n31544 ) | ( n31541 & n31544 ) ;
  assign n31546 = x11 & n31545 ;
  assign n31547 = n31546 ^ n16084 ^ 1'b0 ;
  assign n31548 = n12459 | n24712 ;
  assign n31549 = n31548 ^ n15272 ^ 1'b0 ;
  assign n31550 = n8568 | n13621 ;
  assign n31555 = ( n2544 & n11275 ) | ( n2544 & n18244 ) | ( n11275 & n18244 ) ;
  assign n31556 = n352 | n17692 ;
  assign n31557 = n31555 & ~n31556 ;
  assign n31551 = n15651 | n21286 ;
  assign n31552 = n18638 ^ n17685 ^ 1'b0 ;
  assign n31553 = n31551 & ~n31552 ;
  assign n31554 = ~n19614 & n31553 ;
  assign n31558 = n31557 ^ n31554 ^ 1'b0 ;
  assign n31559 = n3941 ^ n636 ^ n353 ;
  assign n31560 = n31559 ^ n25939 ^ n20310 ;
  assign n31561 = ( n5660 & n17147 ) | ( n5660 & n31560 ) | ( n17147 & n31560 ) ;
  assign n31564 = ~n4606 & n29713 ;
  assign n31565 = n31564 ^ n13365 ^ 1'b0 ;
  assign n31562 = n2155 & n27576 ;
  assign n31563 = n4796 & n31562 ;
  assign n31566 = n31565 ^ n31563 ^ 1'b0 ;
  assign n31571 = ( n5972 & n6864 ) | ( n5972 & ~n10049 ) | ( n6864 & ~n10049 ) ;
  assign n31568 = n9601 ^ n615 ^ 1'b0 ;
  assign n31569 = n31568 ^ n15351 ^ n11821 ;
  assign n31567 = n10630 & ~n27509 ;
  assign n31570 = n31569 ^ n31567 ^ 1'b0 ;
  assign n31572 = n31571 ^ n31570 ^ n21552 ;
  assign n31574 = n4944 & ~n5799 ;
  assign n31575 = n31574 ^ n10599 ^ 1'b0 ;
  assign n31573 = n20130 ^ n12654 ^ 1'b0 ;
  assign n31576 = n31575 ^ n31573 ^ n11419 ;
  assign n31577 = n10739 ^ n1173 ^ 1'b0 ;
  assign n31578 = ~n361 & n13143 ;
  assign n31579 = n5791 & n31578 ;
  assign n31580 = n31577 & ~n31579 ;
  assign n31581 = n7755 & n31580 ;
  assign n31582 = n17568 ^ n9432 ^ 1'b0 ;
  assign n31583 = n19468 | n31582 ;
  assign n31584 = n13938 ^ n11233 ^ 1'b0 ;
  assign n31585 = ~n1390 & n31584 ;
  assign n31586 = ~n17623 & n31585 ;
  assign n31587 = n31586 ^ n21358 ^ 1'b0 ;
  assign n31588 = n8191 & ~n12601 ;
  assign n31589 = n31588 ^ n1986 ^ 1'b0 ;
  assign n31590 = n14161 ^ n285 ^ 1'b0 ;
  assign n31591 = n31589 & ~n31590 ;
  assign n31592 = n31591 ^ n17322 ^ n1365 ;
  assign n31593 = ( n31379 & n31587 ) | ( n31379 & ~n31592 ) | ( n31587 & ~n31592 ) ;
  assign n31594 = n7183 & ~n12313 ;
  assign n31595 = n17681 & ~n31594 ;
  assign n31598 = n19130 ^ n9394 ^ 1'b0 ;
  assign n31599 = ~n11287 & n31598 ;
  assign n31596 = ~n10723 & n12570 ;
  assign n31597 = n3828 & n31596 ;
  assign n31600 = n31599 ^ n31597 ^ 1'b0 ;
  assign n31601 = n19831 | n31600 ;
  assign n31602 = n31601 ^ n1911 ^ 1'b0 ;
  assign n31603 = n13673 | n15523 ;
  assign n31604 = n31603 ^ n2669 ^ 1'b0 ;
  assign n31605 = n23664 ^ n19635 ^ n13694 ;
  assign n31607 = n9725 & n12269 ;
  assign n31608 = n31607 ^ n3120 ^ 1'b0 ;
  assign n31609 = n24161 | n31608 ;
  assign n31610 = n12968 & ~n31609 ;
  assign n31611 = n31610 ^ n12736 ^ n10144 ;
  assign n31606 = n10671 ^ n5665 ^ n1164 ;
  assign n31612 = n31611 ^ n31606 ^ n23549 ;
  assign n31613 = n11738 & ~n31612 ;
  assign n31614 = ~n1932 & n31613 ;
  assign n31615 = n31614 ^ n16126 ^ n5146 ;
  assign n31616 = n12960 ^ n11296 ^ 1'b0 ;
  assign n31617 = n31616 ^ n21178 ^ n2843 ;
  assign n31618 = n2205 | n11885 ;
  assign n31619 = n1016 & ~n31618 ;
  assign n31620 = n21395 & ~n31619 ;
  assign n31621 = ~n6804 & n31620 ;
  assign n31622 = n4060 & n22806 ;
  assign n31623 = n30144 ^ n25376 ^ 1'b0 ;
  assign n31624 = n17945 & n31623 ;
  assign n31625 = n31624 ^ n25334 ^ 1'b0 ;
  assign n31626 = n2036 & ~n31625 ;
  assign n31627 = ( n31621 & ~n31622 ) | ( n31621 & n31626 ) | ( ~n31622 & n31626 ) ;
  assign n31628 = ~n5932 & n20626 ;
  assign n31629 = n31628 ^ n12709 ^ 1'b0 ;
  assign n31631 = n17754 ^ n17529 ^ n8343 ;
  assign n31632 = ( n7213 & n10192 ) | ( n7213 & n14081 ) | ( n10192 & n14081 ) ;
  assign n31633 = ( n15904 & n29782 ) | ( n15904 & n31632 ) | ( n29782 & n31632 ) ;
  assign n31634 = ( n17114 & n31631 ) | ( n17114 & ~n31633 ) | ( n31631 & ~n31633 ) ;
  assign n31630 = ~n6744 & n11549 ;
  assign n31635 = n31634 ^ n31630 ^ 1'b0 ;
  assign n31636 = ~n10353 & n15486 ;
  assign n31637 = n31636 ^ n1743 ^ 1'b0 ;
  assign n31638 = ( n26992 & ~n30573 ) | ( n26992 & n31637 ) | ( ~n30573 & n31637 ) ;
  assign n31639 = n31638 ^ n7622 ^ 1'b0 ;
  assign n31640 = n19227 ^ n14753 ^ n8306 ;
  assign n31641 = n7625 & n15749 ;
  assign n31642 = ( n9576 & n13624 ) | ( n9576 & n18098 ) | ( n13624 & n18098 ) ;
  assign n31643 = n31642 ^ n25242 ^ 1'b0 ;
  assign n31644 = n31643 ^ n8151 ^ n6153 ;
  assign n31645 = n13187 ^ n3690 ^ n761 ;
  assign n31646 = ( ~n22658 & n31644 ) | ( ~n22658 & n31645 ) | ( n31644 & n31645 ) ;
  assign n31647 = n7750 | n16534 ;
  assign n31648 = n31647 ^ n832 ^ 1'b0 ;
  assign n31649 = ~n14058 & n31648 ;
  assign n31650 = n19963 ^ n7194 ^ n6295 ;
  assign n31651 = n6340 | n20183 ;
  assign n31652 = n14972 | n31651 ;
  assign n31653 = ~n28901 & n31652 ;
  assign n31654 = ~n18664 & n31653 ;
  assign n31655 = ( x44 & ~n31650 ) | ( x44 & n31654 ) | ( ~n31650 & n31654 ) ;
  assign n31656 = n17068 ^ n5916 ^ 1'b0 ;
  assign n31657 = n5777 ^ n2775 ^ 1'b0 ;
  assign n31658 = n31657 ^ n20715 ^ 1'b0 ;
  assign n31659 = n5374 & ~n6606 ;
  assign n31660 = n20923 & n31659 ;
  assign n31661 = n31660 ^ n13158 ^ n7209 ;
  assign n31662 = n19556 | n31661 ;
  assign n31663 = n31662 ^ n31634 ^ 1'b0 ;
  assign n31664 = n28361 ^ n5279 ^ 1'b0 ;
  assign n31665 = ~n3099 & n31664 ;
  assign n31666 = n31665 ^ n26757 ^ n20269 ;
  assign n31667 = n24248 & n27663 ;
  assign n31668 = n31667 ^ n14632 ^ 1'b0 ;
  assign n31669 = n3180 & n25831 ;
  assign n31670 = n31669 ^ n7447 ^ 1'b0 ;
  assign n31671 = ( n31666 & n31668 ) | ( n31666 & n31670 ) | ( n31668 & n31670 ) ;
  assign n31672 = n14177 & ~n22694 ;
  assign n31673 = n31672 ^ n3769 ^ 1'b0 ;
  assign n31676 = n4932 & n13624 ;
  assign n31677 = n31676 ^ n6969 ^ 1'b0 ;
  assign n31674 = n29515 ^ n18070 ^ 1'b0 ;
  assign n31675 = n6156 | n31674 ;
  assign n31678 = n31677 ^ n31675 ^ n7475 ;
  assign n31679 = n31678 ^ n21703 ^ 1'b0 ;
  assign n31680 = n19945 ^ n15663 ^ 1'b0 ;
  assign n31684 = n936 & ~n3985 ;
  assign n31685 = n31684 ^ n10938 ^ 1'b0 ;
  assign n31686 = n10769 & ~n31685 ;
  assign n31681 = n14007 ^ n7004 ^ n2197 ;
  assign n31682 = n31681 ^ n26489 ^ n4267 ;
  assign n31683 = ( ~n2476 & n8290 ) | ( ~n2476 & n31682 ) | ( n8290 & n31682 ) ;
  assign n31687 = n31686 ^ n31683 ^ n14325 ;
  assign n31689 = x110 & ~n16195 ;
  assign n31690 = n31689 ^ n11332 ^ 1'b0 ;
  assign n31688 = n4016 & ~n12410 ;
  assign n31691 = n31690 ^ n31688 ^ 1'b0 ;
  assign n31692 = n600 & ~n3894 ;
  assign n31693 = n3894 & n31692 ;
  assign n31694 = x179 & ~n31693 ;
  assign n31695 = ~x179 & n31694 ;
  assign n31696 = n7386 & ~n31695 ;
  assign n31697 = ~n7386 & n31696 ;
  assign n31698 = n5504 & ~n31697 ;
  assign n31699 = n31698 ^ n11826 ^ 1'b0 ;
  assign n31700 = n1083 & ~n14415 ;
  assign n31701 = n31700 ^ n1211 ^ 1'b0 ;
  assign n31702 = n5760 & n7777 ;
  assign n31703 = ~n5809 & n31702 ;
  assign n31704 = ( n6396 & ~n12163 ) | ( n6396 & n31703 ) | ( ~n12163 & n31703 ) ;
  assign n31705 = ( ~n20130 & n20591 ) | ( ~n20130 & n31704 ) | ( n20591 & n31704 ) ;
  assign n31706 = n13305 & n31705 ;
  assign n31707 = n30228 ^ n4700 ^ 1'b0 ;
  assign n31708 = ~n11457 & n31707 ;
  assign n31709 = ( n16758 & n18054 ) | ( n16758 & ~n31708 ) | ( n18054 & ~n31708 ) ;
  assign n31710 = n31709 ^ n13483 ^ n3154 ;
  assign n31711 = ( x35 & ~n31706 ) | ( x35 & n31710 ) | ( ~n31706 & n31710 ) ;
  assign n31712 = ( n22483 & ~n26472 ) | ( n22483 & n31569 ) | ( ~n26472 & n31569 ) ;
  assign n31713 = n8715 ^ n4771 ^ n4557 ;
  assign n31714 = n28519 ^ n9581 ^ 1'b0 ;
  assign n31715 = n31713 & ~n31714 ;
  assign n31716 = ~n24444 & n31715 ;
  assign n31717 = n4306 | n6617 ;
  assign n31718 = n31717 ^ n5303 ^ 1'b0 ;
  assign n31719 = n9965 ^ n785 ^ 1'b0 ;
  assign n31720 = n28851 & n31719 ;
  assign n31721 = n22643 ^ n20701 ^ 1'b0 ;
  assign n31722 = n24336 ^ n2542 ^ 1'b0 ;
  assign n31723 = ( n16444 & n31612 ) | ( n16444 & ~n31722 ) | ( n31612 & ~n31722 ) ;
  assign n31724 = n4097 & ~n17404 ;
  assign n31725 = n24599 & n31724 ;
  assign n31726 = n24694 ^ n9825 ^ 1'b0 ;
  assign n31727 = n31726 ^ n16748 ^ 1'b0 ;
  assign n31728 = ( n9056 & n16640 ) | ( n9056 & ~n18318 ) | ( n16640 & ~n18318 ) ;
  assign n31729 = n26486 | n31728 ;
  assign n31730 = n31727 | n31729 ;
  assign n31731 = n9218 & ~n28265 ;
  assign n31732 = n3889 ^ n2400 ^ 1'b0 ;
  assign n31733 = n31731 & n31732 ;
  assign n31735 = n19674 & n20182 ;
  assign n31736 = n9369 & n31735 ;
  assign n31734 = n5585 | n10329 ;
  assign n31737 = n31736 ^ n31734 ^ 1'b0 ;
  assign n31738 = n2194 & n31737 ;
  assign n31739 = n15626 ^ n790 ^ 1'b0 ;
  assign n31740 = n15985 | n31739 ;
  assign n31741 = ~n543 & n6945 ;
  assign n31742 = n20185 & ~n24543 ;
  assign n31743 = ( n6945 & n12998 ) | ( n6945 & ~n18920 ) | ( n12998 & ~n18920 ) ;
  assign n31744 = n31743 ^ n30458 ^ n9852 ;
  assign n31745 = ~n11565 & n16777 ;
  assign n31746 = n31745 ^ n16357 ^ n15362 ;
  assign n31747 = n13478 & n31746 ;
  assign n31748 = n24894 ^ n13349 ^ n3794 ;
  assign n31749 = ( n6466 & n26527 ) | ( n6466 & ~n31748 ) | ( n26527 & ~n31748 ) ;
  assign n31750 = n31749 ^ n25175 ^ n21680 ;
  assign n31751 = n21949 & ~n30994 ;
  assign n31752 = n31751 ^ n617 ^ 1'b0 ;
  assign n31757 = n16119 ^ n8817 ^ n5144 ;
  assign n31758 = ~n16352 & n31757 ;
  assign n31759 = n31758 ^ n23035 ^ 1'b0 ;
  assign n31756 = ( n3764 & n8994 ) | ( n3764 & ~n28308 ) | ( n8994 & ~n28308 ) ;
  assign n31753 = n31588 ^ n13001 ^ 1'b0 ;
  assign n31754 = n23215 | n31753 ;
  assign n31755 = n31754 ^ n23867 ^ 1'b0 ;
  assign n31760 = n31759 ^ n31756 ^ n31755 ;
  assign n31761 = n31760 ^ n12645 ^ 1'b0 ;
  assign n31762 = n27864 & ~n31761 ;
  assign n31763 = n30525 ^ n5378 ^ 1'b0 ;
  assign n31766 = ~n1267 & n22654 ;
  assign n31767 = ~n14432 & n31766 ;
  assign n31764 = n23563 | n31224 ;
  assign n31765 = n18355 & ~n31764 ;
  assign n31768 = n31767 ^ n31765 ^ n753 ;
  assign n31769 = ( ~n8893 & n9309 ) | ( ~n8893 & n31768 ) | ( n9309 & n31768 ) ;
  assign n31770 = ~n4198 & n8369 ;
  assign n31771 = n11891 ^ n1616 ^ 1'b0 ;
  assign n31772 = n31770 & ~n31771 ;
  assign n31773 = n3166 & n31772 ;
  assign n31774 = n31773 ^ n24403 ^ 1'b0 ;
  assign n31775 = n14247 | n15717 ;
  assign n31776 = n31775 ^ n18490 ^ n2939 ;
  assign n31777 = n17573 & ~n24344 ;
  assign n31778 = n31777 ^ n16981 ^ 1'b0 ;
  assign n31779 = n21179 & n31778 ;
  assign n31780 = n14592 ^ n3860 ^ 1'b0 ;
  assign n31781 = n1427 & ~n31780 ;
  assign n31782 = n31781 ^ x153 ^ 1'b0 ;
  assign n31783 = n8739 & n31782 ;
  assign n31784 = ~n31779 & n31783 ;
  assign n31785 = ( n3187 & n23371 ) | ( n3187 & n24949 ) | ( n23371 & n24949 ) ;
  assign n31786 = n1385 & n6369 ;
  assign n31787 = ~n31785 & n31786 ;
  assign n31790 = n24358 ^ n19865 ^ n9556 ;
  assign n31788 = ( n4461 & n5318 ) | ( n4461 & n6339 ) | ( n5318 & n6339 ) ;
  assign n31789 = n4079 & ~n31788 ;
  assign n31791 = n31790 ^ n31789 ^ 1'b0 ;
  assign n31792 = n855 ^ x12 ^ 1'b0 ;
  assign n31793 = n5916 & ~n31792 ;
  assign n31794 = ( ~n10005 & n14251 ) | ( ~n10005 & n31793 ) | ( n14251 & n31793 ) ;
  assign n31795 = n31794 ^ n2783 ^ 1'b0 ;
  assign n31796 = n8921 & ~n31795 ;
  assign n31797 = n31796 ^ n13735 ^ 1'b0 ;
  assign n31798 = n31791 & n31797 ;
  assign n31801 = n21382 ^ n11703 ^ n2179 ;
  assign n31799 = n18354 ^ n6739 ^ 1'b0 ;
  assign n31800 = ~n2635 & n31799 ;
  assign n31802 = n31801 ^ n31800 ^ n25666 ;
  assign n31803 = n15799 & n26693 ;
  assign n31804 = n26903 & n31803 ;
  assign n31805 = n31804 ^ n5153 ^ n5109 ;
  assign n31806 = ( n5891 & n19070 ) | ( n5891 & n31805 ) | ( n19070 & n31805 ) ;
  assign n31807 = ( n1354 & ~n10452 ) | ( n1354 & n17618 ) | ( ~n10452 & n17618 ) ;
  assign n31808 = n31807 ^ n21777 ^ n15335 ;
  assign n31809 = ~n3272 & n17597 ;
  assign n31810 = ( x51 & n6868 ) | ( x51 & ~n9124 ) | ( n6868 & ~n9124 ) ;
  assign n31811 = n939 | n12960 ;
  assign n31812 = n31811 ^ n7815 ^ 1'b0 ;
  assign n31813 = ~n10000 & n31812 ;
  assign n31814 = n10819 & ~n31813 ;
  assign n31815 = ~n5842 & n6479 ;
  assign n31816 = n31815 ^ n9989 ^ 1'b0 ;
  assign n31817 = n12572 & n31816 ;
  assign n31818 = n20376 & n31817 ;
  assign n31819 = n28196 & ~n31818 ;
  assign n31820 = n989 & n31819 ;
  assign n31821 = ( n11631 & n20316 ) | ( n11631 & ~n31820 ) | ( n20316 & ~n31820 ) ;
  assign n31822 = n3640 | n6211 ;
  assign n31823 = n2042 | n31822 ;
  assign n31824 = ( n4575 & ~n24922 ) | ( n4575 & n31823 ) | ( ~n24922 & n31823 ) ;
  assign n31825 = n31824 ^ n22678 ^ n4902 ;
  assign n31826 = n2576 & ~n11741 ;
  assign n31827 = n31826 ^ n10793 ^ 1'b0 ;
  assign n31828 = n305 & ~n6520 ;
  assign n31829 = ( x162 & n4152 ) | ( x162 & n9302 ) | ( n4152 & n9302 ) ;
  assign n31830 = n7987 & n31829 ;
  assign n31831 = n22796 & n31830 ;
  assign n31832 = n4838 & ~n31831 ;
  assign n31833 = n31832 ^ n18329 ^ n5880 ;
  assign n31834 = n14087 ^ n8844 ^ n480 ;
  assign n31835 = ( n20009 & n31833 ) | ( n20009 & n31834 ) | ( n31833 & n31834 ) ;
  assign n31836 = n7921 & ~n31835 ;
  assign n31837 = n17493 ^ n10653 ^ n6935 ;
  assign n31838 = n31837 ^ n22170 ^ n9019 ;
  assign n31839 = n14636 & ~n31838 ;
  assign n31840 = ~n17477 & n31839 ;
  assign n31841 = n6554 ^ n3271 ^ 1'b0 ;
  assign n31842 = ~n16987 & n31841 ;
  assign n31843 = n8517 & ~n31832 ;
  assign n31844 = ~n31842 & n31843 ;
  assign n31845 = n14077 ^ n3112 ^ n793 ;
  assign n31846 = n417 & n31845 ;
  assign n31847 = n10012 | n29426 ;
  assign n31848 = n30543 ^ n21635 ^ n9455 ;
  assign n31849 = n6118 | n11349 ;
  assign n31850 = ( n6211 & ~n8269 ) | ( n6211 & n17758 ) | ( ~n8269 & n17758 ) ;
  assign n31851 = n27607 ^ n5341 ^ 1'b0 ;
  assign n31852 = n31850 | n31851 ;
  assign n31853 = n26998 & ~n28042 ;
  assign n31854 = n31515 ^ n18906 ^ 1'b0 ;
  assign n31857 = n13379 & n17802 ;
  assign n31855 = n7119 & ~n20909 ;
  assign n31856 = n31855 ^ n31690 ^ 1'b0 ;
  assign n31858 = n31857 ^ n31856 ^ n26900 ;
  assign n31859 = n6778 ^ x93 ^ 1'b0 ;
  assign n31860 = ~n7487 & n31859 ;
  assign n31861 = n31860 ^ n17982 ^ n3994 ;
  assign n31862 = n4352 | n31861 ;
  assign n31863 = n2943 | n31862 ;
  assign n31864 = n31863 ^ n11121 ^ 1'b0 ;
  assign n31867 = n15120 ^ n8739 ^ 1'b0 ;
  assign n31868 = ~n4465 & n31867 ;
  assign n31865 = n10645 ^ n8267 ^ 1'b0 ;
  assign n31866 = x203 & n31865 ;
  assign n31869 = n31868 ^ n31866 ^ n27386 ;
  assign n31870 = n31076 ^ n29378 ^ 1'b0 ;
  assign n31871 = n23003 | n31870 ;
  assign n31872 = n31871 ^ n30281 ^ 1'b0 ;
  assign n31873 = n31869 & n31872 ;
  assign n31874 = ( n11669 & ~n31864 ) | ( n11669 & n31873 ) | ( ~n31864 & n31873 ) ;
  assign n31875 = n12940 ^ n4363 ^ 1'b0 ;
  assign n31876 = n11760 & ~n31875 ;
  assign n31877 = x205 | n7520 ;
  assign n31878 = ( n1245 & ~n1266 ) | ( n1245 & n6784 ) | ( ~n1266 & n6784 ) ;
  assign n31879 = n4114 & n5042 ;
  assign n31880 = n31879 ^ n15805 ^ 1'b0 ;
  assign n31881 = n20183 | n31880 ;
  assign n31882 = n3256 | n20585 ;
  assign n31883 = n10504 ^ n1059 ^ 1'b0 ;
  assign n31884 = ( ~n31881 & n31882 ) | ( ~n31881 & n31883 ) | ( n31882 & n31883 ) ;
  assign n31885 = ( n330 & ~n2833 ) | ( n330 & n3258 ) | ( ~n2833 & n3258 ) ;
  assign n31886 = ( ~n8730 & n8878 ) | ( ~n8730 & n27621 ) | ( n8878 & n27621 ) ;
  assign n31887 = x218 & ~n26888 ;
  assign n31888 = ~n20484 & n31887 ;
  assign n31889 = n31888 ^ n5383 ^ 1'b0 ;
  assign n31890 = ~n31886 & n31889 ;
  assign n31891 = n14435 ^ n8179 ^ 1'b0 ;
  assign n31892 = n11339 ^ n5422 ^ 1'b0 ;
  assign n31893 = n10945 & n31892 ;
  assign n31894 = n28161 ^ n15457 ^ n5015 ;
  assign n31895 = ( n17282 & n31893 ) | ( n17282 & ~n31894 ) | ( n31893 & ~n31894 ) ;
  assign n31896 = n3072 | n9032 ;
  assign n31897 = n9411 ^ n9160 ^ 1'b0 ;
  assign n31898 = n6706 ^ n5556 ^ 1'b0 ;
  assign n31899 = ~n19674 & n31898 ;
  assign n31900 = n18814 & n31899 ;
  assign n31901 = n31897 & n31900 ;
  assign n31902 = n29941 ^ n17987 ^ n8084 ;
  assign n31903 = ( ~n3837 & n15896 ) | ( ~n3837 & n27168 ) | ( n15896 & n27168 ) ;
  assign n31904 = n16823 ^ n8282 ^ 1'b0 ;
  assign n31905 = ( n14669 & ~n23803 ) | ( n14669 & n31904 ) | ( ~n23803 & n31904 ) ;
  assign n31906 = n31905 ^ n11751 ^ n1353 ;
  assign n31907 = ( n15172 & n29807 ) | ( n15172 & ~n31906 ) | ( n29807 & ~n31906 ) ;
  assign n31908 = n23063 ^ n20845 ^ 1'b0 ;
  assign n31909 = n28173 & ~n31908 ;
  assign n31910 = n31909 ^ n17330 ^ 1'b0 ;
  assign n31911 = n31910 ^ n23558 ^ 1'b0 ;
  assign n31912 = n10396 | n31911 ;
  assign n31913 = n8936 & ~n31912 ;
  assign n31914 = ~n9468 & n12742 ;
  assign n31915 = n468 | n2793 ;
  assign n31916 = n31915 ^ n2718 ^ 1'b0 ;
  assign n31917 = n30707 ^ n28804 ^ 1'b0 ;
  assign n31918 = n30464 | n31917 ;
  assign n31919 = ( n4656 & ~n31916 ) | ( n4656 & n31918 ) | ( ~n31916 & n31918 ) ;
  assign n31920 = n31919 ^ n2798 ^ 1'b0 ;
  assign n31921 = n25809 ^ n17615 ^ 1'b0 ;
  assign n31922 = n31920 & ~n31921 ;
  assign n31925 = n12575 & ~n14208 ;
  assign n31926 = n12654 & n31925 ;
  assign n31923 = ( n9640 & ~n12263 ) | ( n9640 & n18421 ) | ( ~n12263 & n18421 ) ;
  assign n31924 = ~n9013 & n31923 ;
  assign n31927 = n31926 ^ n31924 ^ n7028 ;
  assign n31928 = ( n4054 & n8114 ) | ( n4054 & ~n10271 ) | ( n8114 & ~n10271 ) ;
  assign n31929 = n26917 ^ n4139 ^ 1'b0 ;
  assign n31930 = n2798 & n6225 ;
  assign n31931 = n31930 ^ n1393 ^ 1'b0 ;
  assign n31932 = n16679 ^ n9043 ^ 1'b0 ;
  assign n31933 = n31932 ^ n26248 ^ 1'b0 ;
  assign n31934 = n31931 & ~n31933 ;
  assign n31935 = ( n9429 & n31929 ) | ( n9429 & ~n31934 ) | ( n31929 & ~n31934 ) ;
  assign n31936 = n9644 & ~n17290 ;
  assign n31937 = n31936 ^ n16620 ^ 1'b0 ;
  assign n31938 = n20400 & n20952 ;
  assign n31939 = n31938 ^ n26018 ^ 1'b0 ;
  assign n31940 = n27160 ^ n11129 ^ 1'b0 ;
  assign n31941 = ~n18951 & n31940 ;
  assign n31942 = n31941 ^ n19815 ^ n9579 ;
  assign n31943 = n3670 & ~n10559 ;
  assign n31944 = ( ~n2194 & n11995 ) | ( ~n2194 & n31943 ) | ( n11995 & n31943 ) ;
  assign n31945 = n31055 ^ n26724 ^ n17035 ;
  assign n31946 = n1390 | n27037 ;
  assign n31947 = n15506 | n31946 ;
  assign n31948 = n31947 ^ n946 ^ 1'b0 ;
  assign n31949 = n31948 ^ n13686 ^ n1265 ;
  assign n31950 = n31949 ^ n21576 ^ n3375 ;
  assign n31951 = n2059 & n31950 ;
  assign n31952 = ~n11868 & n31951 ;
  assign n31953 = n31952 ^ n14691 ^ 1'b0 ;
  assign n31954 = n1791 | n31953 ;
  assign n31955 = n28305 ^ n20301 ^ 1'b0 ;
  assign n31956 = n14701 | n31955 ;
  assign n31957 = n21363 & ~n31956 ;
  assign n31958 = n20636 & n31957 ;
  assign n31959 = ~n15845 & n25957 ;
  assign n31960 = n23103 & n31959 ;
  assign n31963 = x210 & ~n6025 ;
  assign n31961 = ~n7083 & n29195 ;
  assign n31962 = n5360 & n31961 ;
  assign n31964 = n31963 ^ n31962 ^ 1'b0 ;
  assign n31965 = ~n16303 & n31964 ;
  assign n31966 = ~n12744 & n24889 ;
  assign n31967 = n4706 | n31966 ;
  assign n31968 = n13101 ^ n12296 ^ n1476 ;
  assign n31969 = ~n7135 & n7494 ;
  assign n31970 = n31969 ^ n5942 ^ 1'b0 ;
  assign n31971 = n17513 | n31970 ;
  assign n31972 = n4427 & ~n31971 ;
  assign n31973 = n1092 | n1986 ;
  assign n31974 = n31973 ^ n9613 ^ 1'b0 ;
  assign n31975 = ( n10542 & n31786 ) | ( n10542 & n31974 ) | ( n31786 & n31974 ) ;
  assign n31976 = ( ~n20196 & n31972 ) | ( ~n20196 & n31975 ) | ( n31972 & n31975 ) ;
  assign n31977 = ( n4264 & n15272 ) | ( n4264 & ~n16744 ) | ( n15272 & ~n16744 ) ;
  assign n31978 = n29778 & ~n31412 ;
  assign n31979 = x40 & n31978 ;
  assign n31980 = n12715 ^ n4759 ^ n4517 ;
  assign n31981 = ( n3091 & n24270 ) | ( n3091 & n31980 ) | ( n24270 & n31980 ) ;
  assign n31982 = n3735 & n11262 ;
  assign n31983 = n905 | n4658 ;
  assign n31984 = n3417 & ~n31983 ;
  assign n31985 = n14164 | n31984 ;
  assign n31986 = n31982 & ~n31985 ;
  assign n31987 = n13897 ^ n9170 ^ 1'b0 ;
  assign n31988 = n6331 & ~n31987 ;
  assign n31989 = n20979 & n31988 ;
  assign n31990 = ( ~n1502 & n6475 ) | ( ~n1502 & n23589 ) | ( n6475 & n23589 ) ;
  assign n31991 = n9096 & ~n31990 ;
  assign n31992 = n31991 ^ n31905 ^ n355 ;
  assign n31993 = ( n18210 & ~n19884 ) | ( n18210 & n31992 ) | ( ~n19884 & n31992 ) ;
  assign n31994 = n18387 ^ n9821 ^ n3572 ;
  assign n31995 = ( n2213 & ~n13574 ) | ( n2213 & n31994 ) | ( ~n13574 & n31994 ) ;
  assign n31996 = n977 | n9451 ;
  assign n31997 = n30040 | n31996 ;
  assign n31998 = n9552 | n31997 ;
  assign n31999 = n7067 & ~n16665 ;
  assign n32000 = n25505 ^ n7122 ^ 1'b0 ;
  assign n32001 = ~n11603 & n32000 ;
  assign n32002 = ( ~n1784 & n6874 ) | ( ~n1784 & n25454 ) | ( n6874 & n25454 ) ;
  assign n32003 = n14128 & n32002 ;
  assign n32004 = n32003 ^ n683 ^ 1'b0 ;
  assign n32005 = ( n5787 & n11722 ) | ( n5787 & ~n17828 ) | ( n11722 & ~n17828 ) ;
  assign n32006 = ( n8355 & ~n15054 ) | ( n8355 & n32005 ) | ( ~n15054 & n32005 ) ;
  assign n32007 = n32006 ^ n26338 ^ n16228 ;
  assign n32008 = ~n22855 & n32007 ;
  assign n32010 = ~n9629 & n21479 ;
  assign n32009 = n12277 ^ n12063 ^ x25 ;
  assign n32011 = n32010 ^ n32009 ^ 1'b0 ;
  assign n32012 = n23854 & ~n30460 ;
  assign n32013 = n10261 & ~n25108 ;
  assign n32014 = n7293 & n32013 ;
  assign n32015 = n29860 & n32014 ;
  assign n32016 = ( n6131 & n7689 ) | ( n6131 & n32015 ) | ( n7689 & n32015 ) ;
  assign n32017 = n1454 & n24769 ;
  assign n32018 = n9002 | n14601 ;
  assign n32019 = n32018 ^ n11350 ^ 1'b0 ;
  assign n32020 = n5978 & ~n8528 ;
  assign n32021 = n30366 & n32020 ;
  assign n32022 = x247 & n1801 ;
  assign n32023 = n32022 ^ n11892 ^ 1'b0 ;
  assign n32024 = ( n5853 & n10978 ) | ( n5853 & ~n32023 ) | ( n10978 & ~n32023 ) ;
  assign n32025 = x246 & n32024 ;
  assign n32026 = n32025 ^ n13316 ^ 1'b0 ;
  assign n32027 = n26404 ^ n12562 ^ 1'b0 ;
  assign n32028 = ~n29768 & n32027 ;
  assign n32029 = n12255 & n32028 ;
  assign n32032 = ( ~n4430 & n4944 ) | ( ~n4430 & n13991 ) | ( n4944 & n13991 ) ;
  assign n32030 = n10300 ^ n2684 ^ n1502 ;
  assign n32031 = n2949 | n32030 ;
  assign n32033 = n32032 ^ n32031 ^ 1'b0 ;
  assign n32034 = n32033 ^ n28134 ^ 1'b0 ;
  assign n32035 = n11850 | n32034 ;
  assign n32036 = ~n3589 & n12508 ;
  assign n32037 = ~x56 & n32036 ;
  assign n32038 = n4769 & n24473 ;
  assign n32039 = n2146 & n32038 ;
  assign n32044 = n28081 ^ n10756 ^ n7296 ;
  assign n32040 = n10334 ^ n8130 ^ 1'b0 ;
  assign n32041 = n6081 & n32040 ;
  assign n32042 = n19551 & n32041 ;
  assign n32043 = n32042 ^ n9374 ^ 1'b0 ;
  assign n32045 = n32044 ^ n32043 ^ n28810 ;
  assign n32046 = n32045 ^ n23469 ^ n17037 ;
  assign n32047 = ( n7270 & n17087 ) | ( n7270 & ~n28930 ) | ( n17087 & ~n28930 ) ;
  assign n32048 = n32047 ^ n15659 ^ n2376 ;
  assign n32051 = n8655 ^ n7819 ^ 1'b0 ;
  assign n32049 = n12222 | n23200 ;
  assign n32050 = n13354 | n32049 ;
  assign n32052 = n32051 ^ n32050 ^ n24859 ;
  assign n32053 = n18224 ^ n10079 ^ n8574 ;
  assign n32054 = x222 & n19709 ;
  assign n32055 = n28238 & n32054 ;
  assign n32056 = n1876 | n32055 ;
  assign n32057 = n6117 & n19363 ;
  assign n32058 = n448 & n32057 ;
  assign n32059 = n25371 ^ n1597 ^ 1'b0 ;
  assign n32060 = n22918 ^ n19621 ^ 1'b0 ;
  assign n32061 = ~n471 & n32060 ;
  assign n32062 = n12627 | n14648 ;
  assign n32063 = n10677 ^ n9917 ^ n6240 ;
  assign n32064 = n25783 & n32063 ;
  assign n32068 = n1521 & n2186 ;
  assign n32065 = n30080 ^ n2968 ^ 1'b0 ;
  assign n32066 = n15443 & n32065 ;
  assign n32067 = n5500 & ~n32066 ;
  assign n32069 = n32068 ^ n32067 ^ n15523 ;
  assign n32070 = n5238 | n9543 ;
  assign n32071 = n4540 & n5679 ;
  assign n32072 = n12805 & n32071 ;
  assign n32073 = ( n30788 & ~n32070 ) | ( n30788 & n32072 ) | ( ~n32070 & n32072 ) ;
  assign n32074 = n28171 ^ n17097 ^ 1'b0 ;
  assign n32075 = n21549 | n32074 ;
  assign n32076 = n13071 & ~n32075 ;
  assign n32077 = n25412 & n29476 ;
  assign n32079 = n11443 ^ n9030 ^ 1'b0 ;
  assign n32078 = n16730 ^ n11534 ^ n6721 ;
  assign n32080 = n32079 ^ n32078 ^ 1'b0 ;
  assign n32081 = n32080 ^ n4432 ^ 1'b0 ;
  assign n32082 = n6994 | n14371 ;
  assign n32083 = n32082 ^ n6146 ^ 1'b0 ;
  assign n32084 = n32083 ^ n3190 ^ 1'b0 ;
  assign n32085 = n10172 | n32084 ;
  assign n32086 = n32085 ^ n25261 ^ 1'b0 ;
  assign n32087 = n13873 ^ x160 ^ 1'b0 ;
  assign n32088 = n7630 ^ n7060 ^ n471 ;
  assign n32089 = n13996 ^ n4806 ^ x164 ;
  assign n32092 = n27631 ^ n14906 ^ n5037 ;
  assign n32090 = ( n5078 & n6291 ) | ( n5078 & ~n24690 ) | ( n6291 & ~n24690 ) ;
  assign n32091 = n17726 & n32090 ;
  assign n32093 = n32092 ^ n32091 ^ 1'b0 ;
  assign n32094 = ( ~n3831 & n32089 ) | ( ~n3831 & n32093 ) | ( n32089 & n32093 ) ;
  assign n32095 = n13055 ^ n11498 ^ n6907 ;
  assign n32098 = n16410 ^ n10996 ^ 1'b0 ;
  assign n32097 = n1251 & ~n16968 ;
  assign n32099 = n32098 ^ n32097 ^ 1'b0 ;
  assign n32096 = ~n17513 & n18753 ;
  assign n32100 = n32099 ^ n32096 ^ 1'b0 ;
  assign n32101 = n23527 ^ n11776 ^ 1'b0 ;
  assign n32102 = n706 | n32101 ;
  assign n32103 = n27627 ^ n15109 ^ n2191 ;
  assign n32104 = ( x0 & n16883 ) | ( x0 & n29819 ) | ( n16883 & n29819 ) ;
  assign n32112 = n4068 | n4163 ;
  assign n32106 = ( n2894 & ~n7696 ) | ( n2894 & n10699 ) | ( ~n7696 & n10699 ) ;
  assign n32105 = ~n2347 & n3783 ;
  assign n32107 = n32106 ^ n32105 ^ 1'b0 ;
  assign n32108 = n17168 & ~n32107 ;
  assign n32109 = n11082 ^ n2407 ^ 1'b0 ;
  assign n32110 = n32108 & n32109 ;
  assign n32111 = ~n9646 & n32110 ;
  assign n32113 = n32112 ^ n32111 ^ 1'b0 ;
  assign n32114 = n32104 & n32113 ;
  assign n32115 = ~n1850 & n9759 ;
  assign n32116 = n23329 & n31309 ;
  assign n32117 = n32115 & n32116 ;
  assign n32118 = n32117 ^ n20609 ^ 1'b0 ;
  assign n32119 = n8369 ^ n8098 ^ 1'b0 ;
  assign n32120 = n4832 & ~n32119 ;
  assign n32121 = ( n5849 & n8813 ) | ( n5849 & n32120 ) | ( n8813 & n32120 ) ;
  assign n32122 = n32121 ^ n3580 ^ 1'b0 ;
  assign n32123 = n18517 & ~n32122 ;
  assign n32124 = n32123 ^ n979 ^ 1'b0 ;
  assign n32125 = n32124 ^ n31771 ^ n15049 ;
  assign n32126 = x10 & ~n15220 ;
  assign n32127 = n26568 ^ n19423 ^ 1'b0 ;
  assign n32128 = n32126 & n32127 ;
  assign n32131 = n2723 & n4379 ;
  assign n32132 = ~n5862 & n32131 ;
  assign n32133 = n14543 & n32132 ;
  assign n32129 = ( ~n1300 & n21489 ) | ( ~n1300 & n22314 ) | ( n21489 & n22314 ) ;
  assign n32130 = ~n29985 & n32129 ;
  assign n32134 = n32133 ^ n32130 ^ 1'b0 ;
  assign n32135 = n32128 & ~n32134 ;
  assign n32136 = n16842 & ~n22958 ;
  assign n32137 = n9901 & n19862 ;
  assign n32138 = n32137 ^ n968 ^ 1'b0 ;
  assign n32139 = n32138 ^ n4471 ^ x214 ;
  assign n32140 = n28981 ^ n15534 ^ n2694 ;
  assign n32141 = ~n9779 & n15118 ;
  assign n32142 = n432 & n32141 ;
  assign n32143 = n32142 ^ n6426 ^ n4005 ;
  assign n32144 = n32143 ^ n16691 ^ 1'b0 ;
  assign n32145 = n27245 & ~n32144 ;
  assign n32146 = n27594 & n29575 ;
  assign n32147 = ~n29249 & n32146 ;
  assign n32148 = ( n6369 & n6505 ) | ( n6369 & n8677 ) | ( n6505 & n8677 ) ;
  assign n32149 = n13443 ^ n6002 ^ 1'b0 ;
  assign n32150 = n32148 & ~n32149 ;
  assign n32151 = n32150 ^ n22645 ^ 1'b0 ;
  assign n32152 = n29157 | n32151 ;
  assign n32153 = ( n366 & n5722 ) | ( n366 & n29832 ) | ( n5722 & n29832 ) ;
  assign n32154 = n3360 | n14624 ;
  assign n32155 = n32154 ^ n30130 ^ 1'b0 ;
  assign n32156 = n13188 & n32155 ;
  assign n32157 = ~n13706 & n32156 ;
  assign n32158 = ( n16204 & n32153 ) | ( n16204 & ~n32157 ) | ( n32153 & ~n32157 ) ;
  assign n32159 = ~n8622 & n14745 ;
  assign n32160 = ( n1583 & n29583 ) | ( n1583 & ~n32159 ) | ( n29583 & ~n32159 ) ;
  assign n32161 = n10507 | n18589 ;
  assign n32162 = n28612 & ~n32161 ;
  assign n32163 = ~n7055 & n14278 ;
  assign n32164 = n32162 & n32163 ;
  assign n32165 = n32164 ^ n14908 ^ 1'b0 ;
  assign n32166 = n11802 ^ n4287 ^ n4061 ;
  assign n32167 = n18582 ^ n2793 ^ 1'b0 ;
  assign n32168 = n4023 & n22937 ;
  assign n32169 = ~n32167 & n32168 ;
  assign n32170 = n2231 & ~n19220 ;
  assign n32171 = n32170 ^ n30420 ^ 1'b0 ;
  assign n32183 = n24505 ^ n5473 ^ n4717 ;
  assign n32180 = n18199 ^ n2071 ^ n547 ;
  assign n32181 = n21162 & n32180 ;
  assign n32182 = n32181 ^ n17198 ^ 1'b0 ;
  assign n32172 = n6111 ^ n3984 ^ 1'b0 ;
  assign n32173 = n26019 | n32172 ;
  assign n32174 = n15693 | n32173 ;
  assign n32175 = n32174 ^ n19708 ^ 1'b0 ;
  assign n32177 = ( n2945 & n10585 ) | ( n2945 & n15593 ) | ( n10585 & n15593 ) ;
  assign n32176 = n18205 ^ n10887 ^ 1'b0 ;
  assign n32178 = n32177 ^ n32176 ^ 1'b0 ;
  assign n32179 = n32175 & n32178 ;
  assign n32184 = n32183 ^ n32182 ^ n32179 ;
  assign n32185 = ( ~n17489 & n24651 ) | ( ~n17489 & n29686 ) | ( n24651 & n29686 ) ;
  assign n32186 = ~n17364 & n19255 ;
  assign n32187 = n32186 ^ n16955 ^ 1'b0 ;
  assign n32188 = ( ~n3435 & n32185 ) | ( ~n3435 & n32187 ) | ( n32185 & n32187 ) ;
  assign n32189 = n17933 ^ n12086 ^ 1'b0 ;
  assign n32190 = n1764 & ~n30217 ;
  assign n32191 = n32190 ^ n25446 ^ 1'b0 ;
  assign n32192 = ~n32189 & n32191 ;
  assign n32193 = n6488 & ~n15304 ;
  assign n32196 = n7826 | n8430 ;
  assign n32197 = n32196 ^ n3068 ^ 1'b0 ;
  assign n32194 = n1437 & ~n5324 ;
  assign n32195 = n32194 ^ n22864 ^ 1'b0 ;
  assign n32198 = n32197 ^ n32195 ^ 1'b0 ;
  assign n32199 = ( n6425 & ~n12713 ) | ( n6425 & n28473 ) | ( ~n12713 & n28473 ) ;
  assign n32200 = ( n17245 & n24597 ) | ( n17245 & n32199 ) | ( n24597 & n32199 ) ;
  assign n32201 = n2391 & ~n9088 ;
  assign n32202 = n32201 ^ n4323 ^ 1'b0 ;
  assign n32203 = n13957 ^ n3668 ^ 1'b0 ;
  assign n32204 = ~n2050 & n32203 ;
  assign n32205 = n28014 ^ n13277 ^ n4499 ;
  assign n32206 = ( n12317 & n13340 ) | ( n12317 & ~n23929 ) | ( n13340 & ~n23929 ) ;
  assign n32207 = n32206 ^ n10002 ^ 1'b0 ;
  assign n32208 = n17125 ^ n13289 ^ 1'b0 ;
  assign n32209 = n32208 ^ n10780 ^ 1'b0 ;
  assign n32212 = ( ~n1858 & n9094 ) | ( ~n1858 & n26687 ) | ( n9094 & n26687 ) ;
  assign n32210 = n15787 & ~n17048 ;
  assign n32211 = n32210 ^ n25847 ^ 1'b0 ;
  assign n32213 = n32212 ^ n32211 ^ 1'b0 ;
  assign n32214 = ~n32209 & n32213 ;
  assign n32215 = n31779 ^ n17683 ^ 1'b0 ;
  assign n32216 = ~n14438 & n19190 ;
  assign n32217 = ~n21633 & n32216 ;
  assign n32218 = n2669 | n15842 ;
  assign n32219 = n5233 & ~n32218 ;
  assign n32220 = ( ~n16929 & n19877 ) | ( ~n16929 & n32219 ) | ( n19877 & n32219 ) ;
  assign n32221 = n32220 ^ n23310 ^ n23075 ;
  assign n32222 = n22903 ^ n20490 ^ n2398 ;
  assign n32223 = n29334 ^ n7392 ^ 1'b0 ;
  assign n32224 = n32223 ^ n3509 ^ 1'b0 ;
  assign n32225 = x170 & ~n3031 ;
  assign n32226 = ( n1617 & n6272 ) | ( n1617 & n22394 ) | ( n6272 & n22394 ) ;
  assign n32227 = n32225 & ~n32226 ;
  assign n32228 = n32227 ^ n26145 ^ 1'b0 ;
  assign n32229 = n2074 & n9364 ;
  assign n32230 = n12334 | n32229 ;
  assign n32231 = n32230 ^ n21138 ^ 1'b0 ;
  assign n32232 = ~n2730 & n32231 ;
  assign n32233 = ( n13066 & n32228 ) | ( n13066 & n32232 ) | ( n32228 & n32232 ) ;
  assign n32234 = ( ~n22744 & n23536 ) | ( ~n22744 & n28331 ) | ( n23536 & n28331 ) ;
  assign n32236 = n15826 ^ n574 ^ 1'b0 ;
  assign n32237 = ~n11641 & n32236 ;
  assign n32238 = n4208 & n10731 ;
  assign n32239 = n6191 & n32238 ;
  assign n32240 = ~n32237 & n32239 ;
  assign n32241 = n13729 & ~n32240 ;
  assign n32242 = ~n16363 & n32241 ;
  assign n32235 = ( ~n2523 & n16551 ) | ( ~n2523 & n24895 ) | ( n16551 & n24895 ) ;
  assign n32243 = n32242 ^ n32235 ^ n15926 ;
  assign n32244 = ~n12399 & n32243 ;
  assign n32245 = n9088 | n24425 ;
  assign n32246 = n17027 ^ n6536 ^ 1'b0 ;
  assign n32247 = n32245 & n32246 ;
  assign n32248 = n4728 & n17890 ;
  assign n32249 = n5309 | n19587 ;
  assign n32250 = n3401 & ~n8437 ;
  assign n32251 = n12521 & n32250 ;
  assign n32252 = n32249 & n32251 ;
  assign n32256 = n15254 & n17321 ;
  assign n32253 = n3845 ^ n3705 ^ 1'b0 ;
  assign n32254 = n13252 | n32253 ;
  assign n32255 = n32254 ^ n14439 ^ n9364 ;
  assign n32257 = n32256 ^ n32255 ^ n31577 ;
  assign n32258 = n22590 ^ n4224 ^ 1'b0 ;
  assign n32261 = n11826 ^ n11140 ^ 1'b0 ;
  assign n32262 = n31685 ^ n5639 ^ 1'b0 ;
  assign n32263 = n32261 & ~n32262 ;
  assign n32259 = n10976 ^ n459 ^ 1'b0 ;
  assign n32260 = n26631 & ~n32259 ;
  assign n32264 = n32263 ^ n32260 ^ n13317 ;
  assign n32265 = ( n10185 & ~n13616 ) | ( n10185 & n16598 ) | ( ~n13616 & n16598 ) ;
  assign n32266 = n832 | n6549 ;
  assign n32267 = n8653 ^ n2500 ^ 1'b0 ;
  assign n32268 = n27513 ^ n372 ^ 1'b0 ;
  assign n32269 = n32267 | n32268 ;
  assign n32270 = n1705 & ~n32269 ;
  assign n32271 = n32270 ^ n15510 ^ 1'b0 ;
  assign n32272 = n18108 ^ n10820 ^ 1'b0 ;
  assign n32273 = n32272 ^ n4306 ^ 1'b0 ;
  assign n32277 = x150 & n15269 ;
  assign n32274 = n8091 ^ n2637 ^ 1'b0 ;
  assign n32275 = n12007 & ~n32274 ;
  assign n32276 = n20782 & ~n32275 ;
  assign n32278 = n32277 ^ n32276 ^ 1'b0 ;
  assign n32279 = n12999 & n19132 ;
  assign n32280 = ~n28264 & n32279 ;
  assign n32281 = n4965 & n28104 ;
  assign n32282 = n12343 ^ n4488 ^ 1'b0 ;
  assign n32283 = n9575 | n32282 ;
  assign n32284 = n18658 & ~n32283 ;
  assign n32285 = n32284 ^ n29664 ^ n8127 ;
  assign n32286 = n21429 ^ n11678 ^ x182 ;
  assign n32287 = n3874 & ~n8688 ;
  assign n32288 = x72 & ~n32287 ;
  assign n32289 = ~n15799 & n32288 ;
  assign n32290 = n23989 ^ n13156 ^ 1'b0 ;
  assign n32291 = ~n2440 & n32290 ;
  assign n32292 = n13964 ^ n462 ^ 1'b0 ;
  assign n32293 = ~n14529 & n32292 ;
  assign n32294 = n32293 ^ n24627 ^ n8394 ;
  assign n32295 = ( n7670 & n7947 ) | ( n7670 & ~n12814 ) | ( n7947 & ~n12814 ) ;
  assign n32296 = n17822 ^ n8747 ^ 1'b0 ;
  assign n32297 = n31555 | n32296 ;
  assign n32298 = n13218 ^ n1919 ^ 1'b0 ;
  assign n32299 = n6936 & n32298 ;
  assign n32300 = n1675 & n32299 ;
  assign n32301 = n32300 ^ n26543 ^ 1'b0 ;
  assign n32304 = ~n4177 & n5694 ;
  assign n32305 = n32304 ^ n8059 ^ 1'b0 ;
  assign n32306 = n8139 & ~n19450 ;
  assign n32307 = n32305 & ~n32306 ;
  assign n32308 = n9818 & n32307 ;
  assign n32309 = n30278 ^ n16834 ^ 1'b0 ;
  assign n32310 = ( ~n28148 & n32308 ) | ( ~n28148 & n32309 ) | ( n32308 & n32309 ) ;
  assign n32302 = ~n3197 & n3311 ;
  assign n32303 = ~n13334 & n32302 ;
  assign n32311 = n32310 ^ n32303 ^ 1'b0 ;
  assign n32312 = n8630 & ~n11025 ;
  assign n32313 = n28615 & n32312 ;
  assign n32314 = n24416 ^ n21868 ^ n7976 ;
  assign n32315 = n8647 | n27253 ;
  assign n32316 = n15632 ^ n2994 ^ 1'b0 ;
  assign n32317 = ( n11948 & ~n16738 ) | ( n11948 & n32316 ) | ( ~n16738 & n32316 ) ;
  assign n32318 = ~n802 & n6258 ;
  assign n32319 = n3366 & n32318 ;
  assign n32320 = n27440 & n29154 ;
  assign n32321 = ( ~n28462 & n32319 ) | ( ~n28462 & n32320 ) | ( n32319 & n32320 ) ;
  assign n32322 = n25437 ^ n6809 ^ 1'b0 ;
  assign n32323 = ~n19614 & n32322 ;
  assign n32324 = ~n2634 & n12562 ;
  assign n32325 = n32324 ^ n10981 ^ 1'b0 ;
  assign n32326 = ~n12531 & n32325 ;
  assign n32327 = x115 & ~n32326 ;
  assign n32328 = n12551 & ~n24075 ;
  assign n32329 = n22847 ^ n13000 ^ 1'b0 ;
  assign n32330 = n12043 & n32329 ;
  assign n32331 = n13102 & n32330 ;
  assign n32333 = ~n15063 & n22129 ;
  assign n32332 = n2628 | n28296 ;
  assign n32334 = n32333 ^ n32332 ^ 1'b0 ;
  assign n32335 = n20809 ^ n18899 ^ n2573 ;
  assign n32336 = n32335 ^ n28846 ^ n12488 ;
  assign n32337 = n14097 ^ n12694 ^ n9189 ;
  assign n32338 = ~n24244 & n32337 ;
  assign n32339 = n32336 & n32338 ;
  assign n32340 = n24765 ^ n21549 ^ 1'b0 ;
  assign n32341 = n11364 ^ n1735 ^ 1'b0 ;
  assign n32342 = ( n13456 & ~n28795 ) | ( n13456 & n32341 ) | ( ~n28795 & n32341 ) ;
  assign n32343 = n2265 | n9804 ;
  assign n32344 = ~n11694 & n32343 ;
  assign n32345 = n32344 ^ n14073 ^ 1'b0 ;
  assign n32346 = ( n4105 & n17828 ) | ( n4105 & ~n28118 ) | ( n17828 & ~n28118 ) ;
  assign n32347 = n13107 & ~n32346 ;
  assign n32348 = ~n23522 & n28316 ;
  assign n32349 = n10521 & n32348 ;
  assign n32350 = ~n13480 & n14688 ;
  assign n32351 = n32350 ^ n22388 ^ 1'b0 ;
  assign n32352 = ~n5892 & n32351 ;
  assign n32353 = ( n20831 & ~n21778 ) | ( n20831 & n30084 ) | ( ~n21778 & n30084 ) ;
  assign n32356 = n1923 | n4223 ;
  assign n32357 = n1923 & ~n32356 ;
  assign n32358 = n5074 & n32357 ;
  assign n32354 = ( ~n4575 & n14487 ) | ( ~n4575 & n17499 ) | ( n14487 & n17499 ) ;
  assign n32355 = ( n12111 & n22439 ) | ( n12111 & n32354 ) | ( n22439 & n32354 ) ;
  assign n32359 = n32358 ^ n32355 ^ n4871 ;
  assign n32360 = n31963 ^ n10179 ^ 1'b0 ;
  assign n32361 = n32359 & ~n32360 ;
  assign n32362 = n25463 ^ n21333 ^ 1'b0 ;
  assign n32363 = ~n376 & n807 ;
  assign n32364 = x129 & ~n7395 ;
  assign n32365 = n14430 ^ n7673 ^ 1'b0 ;
  assign n32366 = n7174 & ~n32365 ;
  assign n32367 = n32366 ^ n15552 ^ 1'b0 ;
  assign n32368 = n32367 ^ n12223 ^ n11699 ;
  assign n32369 = n32368 ^ n4662 ^ n3770 ;
  assign n32370 = n5565 | n12705 ;
  assign n32371 = x31 & ~n32370 ;
  assign n32372 = ( n4533 & n27214 ) | ( n4533 & n32371 ) | ( n27214 & n32371 ) ;
  assign n32374 = n11308 & ~n21419 ;
  assign n32375 = n11453 & n32374 ;
  assign n32373 = n17589 & n28440 ;
  assign n32376 = n32375 ^ n32373 ^ 1'b0 ;
  assign n32377 = ~n2492 & n11545 ;
  assign n32378 = n32377 ^ n28954 ^ 1'b0 ;
  assign n32379 = n16287 & n22390 ;
  assign n32380 = n32379 ^ x85 ^ 1'b0 ;
  assign n32381 = ~n4237 & n20372 ;
  assign n32382 = n32381 ^ n26757 ^ 1'b0 ;
  assign n32383 = n7424 ^ n3516 ^ 1'b0 ;
  assign n32385 = n345 & ~n2533 ;
  assign n32386 = n2533 & n32385 ;
  assign n32387 = n2989 & ~n32386 ;
  assign n32388 = ~n2989 & n32387 ;
  assign n32389 = n1278 | n1864 ;
  assign n32390 = n1864 & ~n32389 ;
  assign n32391 = n32390 ^ n614 ^ 1'b0 ;
  assign n32392 = ( n18673 & n32388 ) | ( n18673 & n32391 ) | ( n32388 & n32391 ) ;
  assign n32384 = ~n11832 & n13963 ;
  assign n32393 = n32392 ^ n32384 ^ n23676 ;
  assign n32394 = n29627 ^ n19266 ^ 1'b0 ;
  assign n32395 = n25909 ^ n5745 ^ 1'b0 ;
  assign n32396 = ~n9817 & n10066 ;
  assign n32400 = ( n16655 & n20855 ) | ( n16655 & n28513 ) | ( n20855 & n28513 ) ;
  assign n32397 = n12684 ^ n7411 ^ n787 ;
  assign n32398 = ~n22263 & n32397 ;
  assign n32399 = ~n23552 & n32398 ;
  assign n32401 = n32400 ^ n32399 ^ 1'b0 ;
  assign n32402 = n11757 & n14955 ;
  assign n32403 = n17611 | n27456 ;
  assign n32410 = n4844 | n9766 ;
  assign n32411 = n32410 ^ n6335 ^ 1'b0 ;
  assign n32412 = ( ~n11657 & n20436 ) | ( ~n11657 & n32411 ) | ( n20436 & n32411 ) ;
  assign n32405 = ( n1690 & n20824 ) | ( n1690 & n26008 ) | ( n20824 & n26008 ) ;
  assign n32406 = n2408 & ~n32405 ;
  assign n32407 = ~n10069 & n32406 ;
  assign n32408 = n32407 ^ n26929 ^ 1'b0 ;
  assign n32404 = n27649 ^ n8670 ^ 1'b0 ;
  assign n32409 = n32408 ^ n32404 ^ n736 ;
  assign n32413 = n32412 ^ n32409 ^ 1'b0 ;
  assign n32414 = n32403 & n32413 ;
  assign n32415 = ( n1260 & ~n12522 ) | ( n1260 & n22220 ) | ( ~n12522 & n22220 ) ;
  assign n32416 = n32415 ^ n3781 ^ n2723 ;
  assign n32417 = n6244 ^ n6132 ^ x25 ;
  assign n32418 = n32417 ^ n30365 ^ n6645 ;
  assign n32419 = n17751 | n27937 ;
  assign n32420 = n32419 ^ n22006 ^ 1'b0 ;
  assign n32421 = n32420 ^ n31010 ^ n22389 ;
  assign n32422 = n10851 ^ n632 ^ 1'b0 ;
  assign n32423 = n14369 ^ n13054 ^ 1'b0 ;
  assign n32424 = n9622 & n32423 ;
  assign n32425 = n32424 ^ n5507 ^ 1'b0 ;
  assign n32426 = n7222 & ~n17977 ;
  assign n32427 = ~n32425 & n32426 ;
  assign n32428 = ~n26626 & n30523 ;
  assign n32429 = n9994 ^ n4965 ^ 1'b0 ;
  assign n32430 = ~n8020 & n32429 ;
  assign n32431 = n12047 & ~n25243 ;
  assign n32432 = n32431 ^ n21629 ^ 1'b0 ;
  assign n32433 = n15710 & ~n31036 ;
  assign n32434 = n32432 & n32433 ;
  assign n32435 = n32434 ^ n1137 ^ 1'b0 ;
  assign n32436 = ~n6891 & n32435 ;
  assign n32437 = n26241 ^ n11095 ^ 1'b0 ;
  assign n32438 = ( n2497 & n14065 ) | ( n2497 & n14240 ) | ( n14065 & n14240 ) ;
  assign n32439 = n8574 & ~n32438 ;
  assign n32440 = n32439 ^ n2289 ^ 1'b0 ;
  assign n32441 = ( ~n19584 & n30072 ) | ( ~n19584 & n32440 ) | ( n30072 & n32440 ) ;
  assign n32442 = n21738 ^ n692 ^ 1'b0 ;
  assign n32443 = n10426 ^ n636 ^ 1'b0 ;
  assign n32444 = n14473 & ~n18409 ;
  assign n32447 = n1938 & n2291 ;
  assign n32448 = n32447 ^ n21803 ^ 1'b0 ;
  assign n32445 = n17101 ^ n13567 ^ 1'b0 ;
  assign n32446 = n2718 | n32445 ;
  assign n32449 = n32448 ^ n32446 ^ n16412 ;
  assign n32450 = n32449 ^ n4542 ^ 1'b0 ;
  assign n32451 = n24990 & ~n32450 ;
  assign n32453 = ~n7043 & n8337 ;
  assign n32454 = n7600 & n32453 ;
  assign n32455 = n32454 ^ n1647 ^ 1'b0 ;
  assign n32456 = n32455 ^ n15835 ^ 1'b0 ;
  assign n32452 = n8425 | n16222 ;
  assign n32457 = n32456 ^ n32452 ^ 1'b0 ;
  assign n32458 = n18097 & n21219 ;
  assign n32459 = n32458 ^ n23329 ^ 1'b0 ;
  assign n32460 = n31708 | n32459 ;
  assign n32461 = n6332 & n11237 ;
  assign n32462 = n8132 & n32461 ;
  assign n32463 = n32462 ^ n27993 ^ 1'b0 ;
  assign n32464 = n32460 | n32463 ;
  assign n32465 = n14448 & ~n15063 ;
  assign n32466 = n32465 ^ n7170 ^ 1'b0 ;
  assign n32467 = n12494 ^ n7759 ^ n4946 ;
  assign n32468 = n17141 & ~n32467 ;
  assign n32469 = n32468 ^ n9605 ^ 1'b0 ;
  assign n32471 = n8292 | n12308 ;
  assign n32470 = n6130 & n8713 ;
  assign n32472 = n32471 ^ n32470 ^ 1'b0 ;
  assign n32473 = ( n1888 & n32469 ) | ( n1888 & ~n32472 ) | ( n32469 & ~n32472 ) ;
  assign n32474 = n18336 & n32473 ;
  assign n32475 = n32466 & n32474 ;
  assign n32476 = n5455 | n6382 ;
  assign n32477 = ( n1745 & ~n10753 ) | ( n1745 & n32476 ) | ( ~n10753 & n32476 ) ;
  assign n32478 = ~n8052 & n19646 ;
  assign n32479 = n32478 ^ n27023 ^ n11565 ;
  assign n32480 = n27181 ^ n5268 ^ 1'b0 ;
  assign n32481 = n13848 | n32480 ;
  assign n32482 = n24171 ^ n19173 ^ 1'b0 ;
  assign n32483 = n15764 ^ n13535 ^ n2422 ;
  assign n32484 = n32483 ^ n17720 ^ 1'b0 ;
  assign n32485 = ( n6634 & n10389 ) | ( n6634 & n17330 ) | ( n10389 & n17330 ) ;
  assign n32486 = n13194 ^ n7867 ^ n1040 ;
  assign n32487 = n32486 ^ n29087 ^ n19653 ;
  assign n32488 = n23234 ^ n17751 ^ n3548 ;
  assign n32489 = n4123 ^ n1506 ^ 1'b0 ;
  assign n32490 = n6423 & ~n32489 ;
  assign n32491 = n32490 ^ n7930 ^ n2135 ;
  assign n32492 = n18861 ^ n13375 ^ n10281 ;
  assign n32493 = ~n21041 & n23733 ;
  assign n32494 = n32492 & n32493 ;
  assign n32502 = n29170 ^ n16675 ^ 1'b0 ;
  assign n32501 = n17643 ^ n4840 ^ 1'b0 ;
  assign n32499 = n11120 & n12726 ;
  assign n32500 = n32499 ^ n13096 ^ n6238 ;
  assign n32503 = n32502 ^ n32501 ^ n32500 ;
  assign n32495 = n3495 & ~n17513 ;
  assign n32496 = n32495 ^ n21580 ^ 1'b0 ;
  assign n32497 = n1977 | n32341 ;
  assign n32498 = n32496 & ~n32497 ;
  assign n32504 = n32503 ^ n32498 ^ 1'b0 ;
  assign n32505 = n13800 ^ n3617 ^ n1491 ;
  assign n32506 = n32505 ^ n14471 ^ 1'b0 ;
  assign n32507 = ~n4779 & n32506 ;
  assign n32508 = ~n5451 & n32507 ;
  assign n32509 = n31014 ^ n3175 ^ 1'b0 ;
  assign n32510 = ~n11937 & n32509 ;
  assign n32511 = ( ~n2638 & n7210 ) | ( ~n2638 & n25378 ) | ( n7210 & n25378 ) ;
  assign n32512 = ~n7153 & n28535 ;
  assign n32513 = ( n1470 & n3787 ) | ( n1470 & ~n5728 ) | ( n3787 & ~n5728 ) ;
  assign n32514 = ( n4447 & ~n26853 ) | ( n4447 & n32513 ) | ( ~n26853 & n32513 ) ;
  assign n32515 = n32514 ^ n23952 ^ n10367 ;
  assign n32516 = ( n3286 & ~n21846 ) | ( n3286 & n22688 ) | ( ~n21846 & n22688 ) ;
  assign n32517 = n32516 ^ n22926 ^ 1'b0 ;
  assign n32518 = n32517 ^ n30700 ^ n23268 ;
  assign n32519 = n3170 | n4464 ;
  assign n32520 = ~n6438 & n31655 ;
  assign n32521 = ~x146 & n32520 ;
  assign n32522 = n4244 | n11234 ;
  assign n32523 = n32522 ^ n8424 ^ 1'b0 ;
  assign n32529 = n2528 & ~n7095 ;
  assign n32527 = n1118 ^ n790 ^ 1'b0 ;
  assign n32526 = n17097 & ~n17742 ;
  assign n32528 = n32527 ^ n32526 ^ 1'b0 ;
  assign n32524 = n23184 | n27877 ;
  assign n32525 = n30384 | n32524 ;
  assign n32530 = n32529 ^ n32528 ^ n32525 ;
  assign n32531 = n3481 | n25178 ;
  assign n32532 = n28870 & ~n32531 ;
  assign n32533 = n12738 & n13989 ;
  assign n32534 = ~n1687 & n11579 ;
  assign n32535 = n25951 & n32534 ;
  assign n32536 = n15797 ^ n5797 ^ n2515 ;
  assign n32537 = n27778 & n32536 ;
  assign n32538 = n10875 & ~n24564 ;
  assign n32539 = n8955 & n32538 ;
  assign n32540 = ( ~n594 & n22767 ) | ( ~n594 & n32539 ) | ( n22767 & n32539 ) ;
  assign n32541 = n4942 ^ n2705 ^ 1'b0 ;
  assign n32542 = n2637 & ~n27486 ;
  assign n32543 = n32542 ^ n3798 ^ x1 ;
  assign n32544 = ( n1067 & n4444 ) | ( n1067 & n17649 ) | ( n4444 & n17649 ) ;
  assign n32545 = n26334 ^ n7755 ^ 1'b0 ;
  assign n32546 = n32544 & n32545 ;
  assign n32547 = n15075 & n32546 ;
  assign n32548 = n5425 & n32547 ;
  assign n32549 = n32548 ^ n9561 ^ n9510 ;
  assign n32550 = n1688 | n3672 ;
  assign n32551 = x203 | n32550 ;
  assign n32552 = n32551 ^ n23850 ^ n10017 ;
  assign n32553 = n10994 & ~n32552 ;
  assign n32554 = ( n2646 & ~n10461 ) | ( n2646 & n32553 ) | ( ~n10461 & n32553 ) ;
  assign n32555 = n17614 & n27112 ;
  assign n32556 = n13716 ^ n5533 ^ 1'b0 ;
  assign n32557 = n32556 ^ n31589 ^ 1'b0 ;
  assign n32558 = n25574 & ~n27651 ;
  assign n32559 = ~n12193 & n32558 ;
  assign n32560 = n5825 & n32559 ;
  assign n32561 = n29410 ^ n20585 ^ n3340 ;
  assign n32562 = ( n6455 & n10472 ) | ( n6455 & ~n10802 ) | ( n10472 & ~n10802 ) ;
  assign n32563 = n23459 | n32562 ;
  assign n32564 = ( n7136 & n10130 ) | ( n7136 & ~n20754 ) | ( n10130 & ~n20754 ) ;
  assign n32565 = n18604 ^ n7717 ^ 1'b0 ;
  assign n32566 = n14594 | n32565 ;
  assign n32567 = x108 & ~n13420 ;
  assign n32568 = n12718 ^ n9607 ^ n6589 ;
  assign n32569 = n24995 & ~n32568 ;
  assign n32570 = ~n32567 & n32569 ;
  assign n32571 = n574 & ~n905 ;
  assign n32572 = n32571 ^ n870 ^ 1'b0 ;
  assign n32573 = n13527 ^ n9137 ^ 1'b0 ;
  assign n32574 = ~n1093 & n32573 ;
  assign n32575 = n32574 ^ n19154 ^ 1'b0 ;
  assign n32576 = n8543 ^ n3169 ^ 1'b0 ;
  assign n32577 = n2758 & n22389 ;
  assign n32578 = n32577 ^ n4976 ^ 1'b0 ;
  assign n32579 = ( n2002 & ~n16651 ) | ( n2002 & n32578 ) | ( ~n16651 & n32578 ) ;
  assign n32580 = n32579 ^ n4720 ^ 1'b0 ;
  assign n32581 = n6784 & n16508 ;
  assign n32582 = n10398 & n32581 ;
  assign n32583 = x237 & n9314 ;
  assign n32584 = n32583 ^ n10216 ^ 1'b0 ;
  assign n32585 = n30367 & ~n32584 ;
  assign n32586 = n11013 | n32585 ;
  assign n32587 = n32586 ^ n4893 ^ 1'b0 ;
  assign n32588 = ~n1417 & n10534 ;
  assign n32589 = n32588 ^ n2241 ^ 1'b0 ;
  assign n32590 = ( n23249 & n26911 ) | ( n23249 & ~n32589 ) | ( n26911 & ~n32589 ) ;
  assign n32591 = ( n6610 & ~n6697 ) | ( n6610 & n11513 ) | ( ~n6697 & n11513 ) ;
  assign n32592 = n12841 & ~n21251 ;
  assign n32593 = ~n4073 & n32592 ;
  assign n32594 = ( n3067 & ~n4924 ) | ( n3067 & n32593 ) | ( ~n4924 & n32593 ) ;
  assign n32595 = n25992 | n32594 ;
  assign n32596 = n32591 & ~n32595 ;
  assign n32597 = n18664 & ~n32596 ;
  assign n32598 = ~n32590 & n32597 ;
  assign n32599 = n18301 & ~n19879 ;
  assign n32600 = n32599 ^ n27027 ^ n3830 ;
  assign n32601 = ( ~n4160 & n28320 ) | ( ~n4160 & n32600 ) | ( n28320 & n32600 ) ;
  assign n32602 = ( n12562 & ~n14492 ) | ( n12562 & n19293 ) | ( ~n14492 & n19293 ) ;
  assign n32603 = n14263 ^ n4389 ^ 1'b0 ;
  assign n32604 = n30464 | n32603 ;
  assign n32605 = n3109 & n14029 ;
  assign n32606 = n32605 ^ n21183 ^ 1'b0 ;
  assign n32607 = n32606 ^ n3720 ^ 1'b0 ;
  assign n32608 = n13987 & n32607 ;
  assign n32610 = n19628 ^ n6304 ^ 1'b0 ;
  assign n32611 = ~n5673 & n32610 ;
  assign n32609 = n3516 ^ n2719 ^ 1'b0 ;
  assign n32612 = n32611 ^ n32609 ^ n25442 ;
  assign n32613 = n11039 | n18840 ;
  assign n32614 = ( n11365 & n16348 ) | ( n11365 & n32613 ) | ( n16348 & n32613 ) ;
  assign n32615 = n20685 & ~n32614 ;
  assign n32616 = n17500 ^ n4384 ^ 1'b0 ;
  assign n32617 = n21062 ^ n9798 ^ 1'b0 ;
  assign n32618 = n4067 & ~n32617 ;
  assign n32619 = ( n19573 & n32616 ) | ( n19573 & n32618 ) | ( n32616 & n32618 ) ;
  assign n32620 = n30082 ^ n9008 ^ 1'b0 ;
  assign n32621 = n14173 ^ n8839 ^ 1'b0 ;
  assign n32622 = ~n3032 & n32621 ;
  assign n32623 = n16999 | n18642 ;
  assign n32624 = n2748 & ~n32623 ;
  assign n32626 = n5112 | n11616 ;
  assign n32627 = n10288 & ~n32626 ;
  assign n32625 = ~n802 & n1859 ;
  assign n32628 = n32627 ^ n32625 ^ 1'b0 ;
  assign n32629 = x168 & n1186 ;
  assign n32630 = n6216 ^ n466 ^ 1'b0 ;
  assign n32631 = n20001 | n32630 ;
  assign n32632 = ( n1556 & n11914 ) | ( n1556 & ~n32631 ) | ( n11914 & ~n32631 ) ;
  assign n32633 = n26192 ^ n8538 ^ 1'b0 ;
  assign n32634 = ( ~n32629 & n32632 ) | ( ~n32629 & n32633 ) | ( n32632 & n32633 ) ;
  assign n32635 = ( ~n1093 & n11037 ) | ( ~n1093 & n13449 ) | ( n11037 & n13449 ) ;
  assign n32636 = x122 & ~n6512 ;
  assign n32637 = n29436 & n32636 ;
  assign n32638 = ~n32635 & n32637 ;
  assign n32639 = n32638 ^ n9556 ^ n4342 ;
  assign n32640 = n17870 ^ n12401 ^ n10235 ;
  assign n32641 = ( ~n8405 & n17739 ) | ( ~n8405 & n23614 ) | ( n17739 & n23614 ) ;
  assign n32642 = ( n8814 & n12236 ) | ( n8814 & n18705 ) | ( n12236 & n18705 ) ;
  assign n32643 = n26934 ^ n9738 ^ n3160 ;
  assign n32644 = n32643 ^ n15507 ^ n5970 ;
  assign n32645 = n32642 & ~n32644 ;
  assign n32646 = n32645 ^ n10318 ^ 1'b0 ;
  assign n32647 = n404 & ~n30450 ;
  assign n32648 = n32647 ^ n17796 ^ 1'b0 ;
  assign n32649 = n18573 ^ n2619 ^ 1'b0 ;
  assign n32650 = n18366 & n21798 ;
  assign n32651 = n32650 ^ n26937 ^ 1'b0 ;
  assign n32652 = n2989 | n32651 ;
  assign n32653 = ( n14996 & n25689 ) | ( n14996 & n32652 ) | ( n25689 & n32652 ) ;
  assign n32654 = n6917 & n12813 ;
  assign n32655 = n5741 & n19116 ;
  assign n32656 = n32655 ^ n20366 ^ 1'b0 ;
  assign n32657 = n32654 & n32656 ;
  assign n32658 = n22481 ^ n21242 ^ 1'b0 ;
  assign n32659 = ( n284 & n809 ) | ( n284 & ~n2698 ) | ( n809 & ~n2698 ) ;
  assign n32660 = n13144 | n22353 ;
  assign n32661 = n19314 ^ n8222 ^ n1007 ;
  assign n32662 = ( ~n3500 & n13156 ) | ( ~n3500 & n21502 ) | ( n13156 & n21502 ) ;
  assign n32663 = n32662 ^ n1383 ^ 1'b0 ;
  assign n32664 = n16356 & n32663 ;
  assign n32665 = n16508 ^ n6096 ^ n616 ;
  assign n32666 = n18148 | n32665 ;
  assign n32667 = n32664 & n32666 ;
  assign n32668 = n9762 & n14769 ;
  assign n32669 = n4550 & n32668 ;
  assign n32670 = n32669 ^ n6667 ^ n4692 ;
  assign n32671 = n19171 ^ n6087 ^ 1'b0 ;
  assign n32672 = ~n13042 & n22970 ;
  assign n32673 = n3381 & n32672 ;
  assign n32674 = ~n15274 & n32673 ;
  assign n32675 = n21635 ^ n10715 ^ 1'b0 ;
  assign n32676 = n27510 ^ n8842 ^ n1482 ;
  assign n32677 = n32676 ^ n31621 ^ n20222 ;
  assign n32678 = n4585 ^ n757 ^ 1'b0 ;
  assign n32679 = ~n19069 & n32678 ;
  assign n32680 = n32679 ^ n23137 ^ 1'b0 ;
  assign n32681 = n32680 ^ n28340 ^ n25063 ;
  assign n32682 = n28704 ^ n19938 ^ n4637 ;
  assign n32683 = n32682 ^ n32591 ^ n10755 ;
  assign n32684 = n23093 ^ n3701 ^ 1'b0 ;
  assign n32685 = n5368 & n6647 ;
  assign n32686 = n8154 & n13342 ;
  assign n32687 = n5983 & ~n11947 ;
  assign n32688 = n32687 ^ n13531 ^ 1'b0 ;
  assign n32689 = ~n10741 & n16128 ;
  assign n32690 = ~n32688 & n32689 ;
  assign n32691 = n8962 ^ n7409 ^ 1'b0 ;
  assign n32692 = n12648 & n32691 ;
  assign n32693 = ( n20763 & n32690 ) | ( n20763 & n32692 ) | ( n32690 & n32692 ) ;
  assign n32694 = n20777 ^ n19711 ^ n9767 ;
  assign n32695 = ( n1260 & ~n4704 ) | ( n1260 & n32694 ) | ( ~n4704 & n32694 ) ;
  assign n32696 = n18399 ^ n1108 ^ 1'b0 ;
  assign n32697 = n32696 ^ n22259 ^ 1'b0 ;
  assign n32698 = n4612 & ~n32697 ;
  assign n32699 = ~n10102 & n11413 ;
  assign n32700 = n23761 ^ n12823 ^ n6453 ;
  assign n32701 = ~n32699 & n32700 ;
  assign n32702 = n32701 ^ n26145 ^ 1'b0 ;
  assign n32703 = n26427 | n29264 ;
  assign n32704 = n32703 ^ n23803 ^ 1'b0 ;
  assign n32705 = n4136 & ~n31963 ;
  assign n32706 = n6365 & n14517 ;
  assign n32707 = n32705 & n32706 ;
  assign n32708 = ~n6411 & n29104 ;
  assign n32709 = n32708 ^ n32150 ^ 1'b0 ;
  assign n32710 = n27243 ^ n22470 ^ 1'b0 ;
  assign n32711 = n6301 ^ n4014 ^ 1'b0 ;
  assign n32712 = n6079 & ~n32711 ;
  assign n32713 = n30600 ^ n18836 ^ 1'b0 ;
  assign n32714 = n32712 & ~n32713 ;
  assign n32715 = ( ~n7579 & n24974 ) | ( ~n7579 & n32714 ) | ( n24974 & n32714 ) ;
  assign n32717 = n3422 & n7922 ;
  assign n32718 = ( ~n20355 & n25999 ) | ( ~n20355 & n32717 ) | ( n25999 & n32717 ) ;
  assign n32719 = ~n2388 & n7163 ;
  assign n32720 = n32719 ^ n19781 ^ 1'b0 ;
  assign n32721 = n32718 & n32720 ;
  assign n32716 = n24989 & ~n30925 ;
  assign n32722 = n32721 ^ n32716 ^ 1'b0 ;
  assign n32723 = n4553 & ~n6170 ;
  assign n32724 = n32723 ^ n15884 ^ n1390 ;
  assign n32725 = ~n19164 & n32724 ;
  assign n32730 = n12851 ^ n5050 ^ 1'b0 ;
  assign n32731 = n1196 & ~n32730 ;
  assign n32726 = n19507 | n29848 ;
  assign n32727 = n1208 | n32726 ;
  assign n32728 = ~n11428 & n32727 ;
  assign n32729 = ~n1911 & n32728 ;
  assign n32732 = n32731 ^ n32729 ^ n15142 ;
  assign n32733 = n26911 ^ n9564 ^ n6139 ;
  assign n32734 = ( n20637 & n32657 ) | ( n20637 & ~n32733 ) | ( n32657 & ~n32733 ) ;
  assign n32735 = n6520 & ~n19818 ;
  assign n32736 = n20032 ^ n13776 ^ n4598 ;
  assign n32737 = n13506 & n32736 ;
  assign n32738 = n8878 ^ n4287 ^ n4274 ;
  assign n32739 = n32738 ^ n6586 ^ n6033 ;
  assign n32740 = n19468 | n32739 ;
  assign n32741 = n17956 ^ n13382 ^ 1'b0 ;
  assign n32742 = n23512 & n32741 ;
  assign n32743 = n15153 ^ n11350 ^ 1'b0 ;
  assign n32744 = ( ~n6712 & n8110 ) | ( ~n6712 & n32743 ) | ( n8110 & n32743 ) ;
  assign n32745 = n7830 | n30868 ;
  assign n32746 = ( n5366 & n6762 ) | ( n5366 & n12682 ) | ( n6762 & n12682 ) ;
  assign n32747 = ( n32519 & n32745 ) | ( n32519 & ~n32746 ) | ( n32745 & ~n32746 ) ;
  assign n32749 = ~n5779 & n7285 ;
  assign n32750 = n32749 ^ n259 ^ 1'b0 ;
  assign n32748 = n21952 & ~n22868 ;
  assign n32751 = n32750 ^ n32748 ^ 1'b0 ;
  assign n32753 = n14452 ^ n13321 ^ n7257 ;
  assign n32752 = n2247 & ~n13042 ;
  assign n32754 = n32753 ^ n32752 ^ 1'b0 ;
  assign n32755 = n9816 & ~n32754 ;
  assign n32756 = n5078 ^ n812 ^ 1'b0 ;
  assign n32757 = ~n7709 & n32756 ;
  assign n32758 = n4124 & ~n6956 ;
  assign n32759 = n10926 & n32758 ;
  assign n32760 = ~n14890 & n32759 ;
  assign n32761 = n24355 ^ n6777 ^ 1'b0 ;
  assign n32762 = n12186 | n15005 ;
  assign n32763 = n32762 ^ n22456 ^ 1'b0 ;
  assign n32764 = ( n32760 & ~n32761 ) | ( n32760 & n32763 ) | ( ~n32761 & n32763 ) ;
  assign n32765 = n32764 ^ n2803 ^ n2544 ;
  assign n32766 = n16018 ^ n5529 ^ 1'b0 ;
  assign n32767 = ~n7415 & n13088 ;
  assign n32768 = ~n9360 & n32767 ;
  assign n32769 = n7192 ^ n5871 ^ 1'b0 ;
  assign n32770 = n12580 & ~n32769 ;
  assign n32771 = ~n6155 & n32770 ;
  assign n32772 = n32768 & n32771 ;
  assign n32773 = n11545 ^ n1971 ^ 1'b0 ;
  assign n32774 = ~n32772 & n32773 ;
  assign n32775 = ( n4552 & n5172 ) | ( n4552 & ~n12355 ) | ( n5172 & ~n12355 ) ;
  assign n32776 = ( n1945 & n31021 ) | ( n1945 & n32775 ) | ( n31021 & n32775 ) ;
  assign n32777 = ( n26980 & ~n32774 ) | ( n26980 & n32776 ) | ( ~n32774 & n32776 ) ;
  assign n32778 = n9203 ^ n1672 ^ 1'b0 ;
  assign n32780 = n13216 ^ n3846 ^ 1'b0 ;
  assign n32779 = n25207 ^ n23952 ^ n13203 ;
  assign n32781 = n32780 ^ n32779 ^ n23543 ;
  assign n32782 = n15455 ^ n2411 ^ 1'b0 ;
  assign n32783 = n32375 & ~n32782 ;
  assign n32784 = ( ~n5916 & n8201 ) | ( ~n5916 & n27640 ) | ( n8201 & n27640 ) ;
  assign n32785 = n29566 ^ n21571 ^ 1'b0 ;
  assign n32786 = ~n1396 & n32785 ;
  assign n32787 = n32786 ^ n32453 ^ 1'b0 ;
  assign n32788 = n3136 & n32787 ;
  assign n32790 = n1363 | n6931 ;
  assign n32791 = n1681 | n32790 ;
  assign n32789 = n9662 | n10694 ;
  assign n32792 = n32791 ^ n32789 ^ n4794 ;
  assign n32793 = n32792 ^ n30224 ^ n14207 ;
  assign n32794 = ( n8630 & n12672 ) | ( n8630 & n17948 ) | ( n12672 & n17948 ) ;
  assign n32795 = n31394 ^ n14197 ^ n5704 ;
  assign n32796 = n15120 ^ n3184 ^ n2247 ;
  assign n32797 = ~n20868 & n32796 ;
  assign n32798 = n32797 ^ n24697 ^ 1'b0 ;
  assign n32799 = n25096 ^ n10677 ^ n5133 ;
  assign n32800 = n17511 | n32799 ;
  assign n32801 = ~n11987 & n32800 ;
  assign n32802 = n12457 & n32801 ;
  assign n32803 = n10709 | n15115 ;
  assign n32804 = n23027 & ~n32803 ;
  assign n32805 = n10513 | n11794 ;
  assign n32806 = n19195 ^ n12927 ^ n11476 ;
  assign n32807 = n15297 & ~n32806 ;
  assign n32808 = ( ~n25882 & n32805 ) | ( ~n25882 & n32807 ) | ( n32805 & n32807 ) ;
  assign n32809 = n17794 ^ n7311 ^ 1'b0 ;
  assign n32810 = ~n13897 & n32809 ;
  assign n32811 = n853 & n11013 ;
  assign n32812 = n29965 ^ n14056 ^ 1'b0 ;
  assign n32813 = n21385 & n23249 ;
  assign n32814 = n32812 & n32813 ;
  assign n32815 = n18172 & ~n32814 ;
  assign n32816 = n32811 & n32815 ;
  assign n32817 = n32816 ^ n32558 ^ 1'b0 ;
  assign n32818 = ~n17544 & n17952 ;
  assign n32819 = n14815 ^ n476 ^ 1'b0 ;
  assign n32820 = n16844 & n32819 ;
  assign n32821 = n9561 & n32820 ;
  assign n32822 = n10072 ^ n7916 ^ n1799 ;
  assign n32823 = n32822 ^ n30994 ^ n11463 ;
  assign n32824 = ~n6691 & n32823 ;
  assign n32825 = ( n5177 & ~n20670 ) | ( n5177 & n23343 ) | ( ~n20670 & n23343 ) ;
  assign n32826 = ~n5817 & n8740 ;
  assign n32827 = ( n3085 & n3402 ) | ( n3085 & n32826 ) | ( n3402 & n32826 ) ;
  assign n32828 = n13236 ^ n10881 ^ n7136 ;
  assign n32830 = n7526 ^ n3131 ^ n1941 ;
  assign n32831 = n11103 | n32830 ;
  assign n32832 = n32831 ^ n9328 ^ 1'b0 ;
  assign n32829 = n32308 ^ n20046 ^ 1'b0 ;
  assign n32833 = n32832 ^ n32829 ^ n3885 ;
  assign n32834 = ( n881 & n12563 ) | ( n881 & ~n32833 ) | ( n12563 & ~n32833 ) ;
  assign n32835 = n15426 ^ n8536 ^ 1'b0 ;
  assign n32836 = n3643 & n32835 ;
  assign n32837 = ~n25262 & n32836 ;
  assign n32838 = n14498 & n32837 ;
  assign n32839 = n6330 ^ n3647 ^ 1'b0 ;
  assign n32840 = ( ~n7981 & n8545 ) | ( ~n7981 & n9137 ) | ( n8545 & n9137 ) ;
  assign n32841 = n32840 ^ n9457 ^ 1'b0 ;
  assign n32842 = n32839 & ~n32841 ;
  assign n32843 = n15949 ^ n14722 ^ n12411 ;
  assign n32844 = n30834 & ~n32843 ;
  assign n32845 = n32844 ^ n20441 ^ 1'b0 ;
  assign n32846 = n6720 & ~n11996 ;
  assign n32847 = n16611 & n32846 ;
  assign n32848 = n30943 ^ n29372 ^ 1'b0 ;
  assign n32849 = n32848 ^ n25349 ^ n7970 ;
  assign n32850 = n13594 & ~n28926 ;
  assign n32851 = n32850 ^ n15543 ^ n636 ;
  assign n32852 = n10371 ^ n8436 ^ 1'b0 ;
  assign n32853 = n28279 ^ n9531 ^ 1'b0 ;
  assign n32854 = n32853 ^ n20231 ^ 1'b0 ;
  assign n32855 = n7610 & n30870 ;
  assign n32856 = n32855 ^ n4007 ^ 1'b0 ;
  assign n32857 = n5965 ^ n568 ^ 1'b0 ;
  assign n32858 = n17060 | n32857 ;
  assign n32859 = n32858 ^ n11702 ^ 1'b0 ;
  assign n32860 = ~n8554 & n32859 ;
  assign n32861 = n32860 ^ n30050 ^ n7869 ;
  assign n32862 = n20346 ^ n18382 ^ 1'b0 ;
  assign n32863 = n12627 & ~n32862 ;
  assign n32864 = n32863 ^ n8175 ^ n1336 ;
  assign n32865 = ~n26907 & n30502 ;
  assign n32866 = n11954 | n32865 ;
  assign n32867 = ( n7920 & ~n12026 ) | ( n7920 & n32866 ) | ( ~n12026 & n32866 ) ;
  assign n32868 = n5953 & ~n23964 ;
  assign n32869 = ( n32864 & n32867 ) | ( n32864 & n32868 ) | ( n32867 & n32868 ) ;
  assign n32873 = ( x106 & n7304 ) | ( x106 & ~n8413 ) | ( n7304 & ~n8413 ) ;
  assign n32874 = n32873 ^ n17162 ^ 1'b0 ;
  assign n32875 = n10041 | n32874 ;
  assign n32870 = n17775 ^ n10645 ^ n6501 ;
  assign n32871 = ( n5424 & ~n28505 ) | ( n5424 & n32870 ) | ( ~n28505 & n32870 ) ;
  assign n32872 = ( n6672 & n6908 ) | ( n6672 & ~n32871 ) | ( n6908 & ~n32871 ) ;
  assign n32876 = n32875 ^ n32872 ^ 1'b0 ;
  assign n32881 = n12936 ^ n7865 ^ 1'b0 ;
  assign n32882 = n3361 | n32881 ;
  assign n32878 = n13012 ^ n3876 ^ 1'b0 ;
  assign n32879 = ~n5585 & n32878 ;
  assign n32877 = n8493 & n28027 ;
  assign n32880 = n32879 ^ n32877 ^ 1'b0 ;
  assign n32883 = n32882 ^ n32880 ^ n18134 ;
  assign n32884 = n10318 ^ n1328 ^ 1'b0 ;
  assign n32885 = ~n16831 & n32884 ;
  assign n32886 = n32885 ^ n9297 ^ 1'b0 ;
  assign n32887 = n24455 & n32886 ;
  assign n32888 = n32887 ^ n21680 ^ 1'b0 ;
  assign n32889 = ~n3459 & n5535 ;
  assign n32890 = n32889 ^ n15598 ^ 1'b0 ;
  assign n32895 = n12977 & ~n23485 ;
  assign n32896 = n5907 & n32895 ;
  assign n32891 = n18505 ^ n10161 ^ n6428 ;
  assign n32892 = n22082 ^ n4866 ^ 1'b0 ;
  assign n32893 = n10714 & n32892 ;
  assign n32894 = ~n32891 & n32893 ;
  assign n32897 = n32896 ^ n32894 ^ n18248 ;
  assign n32898 = ( n1649 & n10227 ) | ( n1649 & ~n20457 ) | ( n10227 & ~n20457 ) ;
  assign n32899 = ( n5844 & n13897 ) | ( n5844 & ~n25546 ) | ( n13897 & ~n25546 ) ;
  assign n32900 = ~n5240 & n11088 ;
  assign n32901 = n32900 ^ n20298 ^ 1'b0 ;
  assign n32902 = n22305 ^ n8056 ^ n2881 ;
  assign n32903 = n25163 | n32902 ;
  assign n32904 = n32903 ^ n20731 ^ 1'b0 ;
  assign n32905 = n749 & ~n31050 ;
  assign n32906 = n32905 ^ n9903 ^ 1'b0 ;
  assign n32908 = n13780 ^ n13491 ^ 1'b0 ;
  assign n32909 = n32908 ^ n25444 ^ 1'b0 ;
  assign n32910 = n25675 & n32909 ;
  assign n32907 = n18298 ^ n17284 ^ n9114 ;
  assign n32911 = n32910 ^ n32907 ^ n3227 ;
  assign n32912 = n27461 ^ n21051 ^ n12728 ;
  assign n32913 = n4291 & n12645 ;
  assign n32914 = ( n23547 & ~n30575 ) | ( n23547 & n32913 ) | ( ~n30575 & n32913 ) ;
  assign n32915 = ~n1265 & n3690 ;
  assign n32916 = ~n11384 & n32915 ;
  assign n32917 = n3321 ^ n2832 ^ 1'b0 ;
  assign n32918 = n1233 | n32917 ;
  assign n32919 = n9652 & ~n32918 ;
  assign n32920 = ~n10034 & n32919 ;
  assign n32921 = ~n12483 & n25574 ;
  assign n32922 = n32921 ^ n15486 ^ 1'b0 ;
  assign n32923 = ( n11260 & ~n13920 ) | ( n11260 & n32922 ) | ( ~n13920 & n32922 ) ;
  assign n32924 = n20371 ^ n6674 ^ 1'b0 ;
  assign n32925 = n32923 & n32924 ;
  assign n32926 = n7862 | n20270 ;
  assign n32927 = n32926 ^ n30313 ^ 1'b0 ;
  assign n32928 = n32927 ^ n19699 ^ n16668 ;
  assign n32933 = n11299 ^ n4037 ^ 1'b0 ;
  assign n32934 = n32933 ^ n21284 ^ 1'b0 ;
  assign n32935 = ( n7208 & ~n25808 ) | ( n7208 & n32934 ) | ( ~n25808 & n32934 ) ;
  assign n32929 = n480 & n10411 ;
  assign n32930 = ~n7173 & n32929 ;
  assign n32931 = n32930 ^ n27828 ^ n21728 ;
  assign n32932 = n32931 ^ n17904 ^ n6088 ;
  assign n32936 = n32935 ^ n32932 ^ n17592 ;
  assign n32937 = n21706 ^ n6197 ^ 1'b0 ;
  assign n32938 = ~n18571 & n32502 ;
  assign n32939 = n9879 & n32938 ;
  assign n32940 = n32939 ^ n30010 ^ n21085 ;
  assign n32941 = n10247 | n22575 ;
  assign n32942 = n32941 ^ n18373 ^ 1'b0 ;
  assign n32943 = n11325 | n18680 ;
  assign n32944 = n32943 ^ n14634 ^ 1'b0 ;
  assign n32945 = ~n1511 & n9884 ;
  assign n32946 = n32945 ^ n28373 ^ 1'b0 ;
  assign n32947 = n3811 & n32946 ;
  assign n32948 = n32947 ^ n1863 ^ 1'b0 ;
  assign n32949 = n32948 ^ n4852 ^ 1'b0 ;
  assign n32950 = n30883 & n32949 ;
  assign n32951 = n12254 ^ n6560 ^ 1'b0 ;
  assign n32952 = n32951 ^ n2324 ^ 1'b0 ;
  assign n32953 = ~n291 & n19409 ;
  assign n32954 = ( n15120 & n18889 ) | ( n15120 & n32953 ) | ( n18889 & n32953 ) ;
  assign n32955 = ( ~x11 & n11553 ) | ( ~x11 & n25980 ) | ( n11553 & n25980 ) ;
  assign n32956 = n13579 ^ n7963 ^ n5070 ;
  assign n32957 = ( ~n13428 & n32955 ) | ( ~n13428 & n32956 ) | ( n32955 & n32956 ) ;
  assign n32958 = n18069 & ~n22530 ;
  assign n32959 = n27753 & n32958 ;
  assign n32960 = n26220 ^ n19972 ^ n768 ;
  assign n32961 = n30786 & ~n32960 ;
  assign n32962 = ~n13393 & n32961 ;
  assign n32963 = n18148 ^ n11750 ^ n7622 ;
  assign n32964 = ( n5143 & ~n8614 ) | ( n5143 & n32963 ) | ( ~n8614 & n32963 ) ;
  assign n32965 = n15398 ^ n10052 ^ n2412 ;
  assign n32966 = n31314 ^ n22395 ^ n12788 ;
  assign n32967 = n32966 ^ n26283 ^ 1'b0 ;
  assign n32968 = ( n30265 & n32965 ) | ( n30265 & ~n32967 ) | ( n32965 & ~n32967 ) ;
  assign n32969 = n17314 ^ n7895 ^ 1'b0 ;
  assign n32970 = n26228 & n32969 ;
  assign n32971 = n325 & n12655 ;
  assign n32972 = n16065 | n29376 ;
  assign n32973 = n32971 & ~n32972 ;
  assign n32975 = ( n279 & n2545 ) | ( n279 & n15274 ) | ( n2545 & n15274 ) ;
  assign n32974 = n449 & ~n26470 ;
  assign n32976 = n32975 ^ n32974 ^ 1'b0 ;
  assign n32977 = ( ~n9001 & n14349 ) | ( ~n9001 & n32867 ) | ( n14349 & n32867 ) ;
  assign n32978 = n8616 | n14272 ;
  assign n32979 = n12880 & n32978 ;
  assign n32980 = n11865 ^ n598 ^ 1'b0 ;
  assign n32981 = ( n3817 & n5014 ) | ( n3817 & n32980 ) | ( n5014 & n32980 ) ;
  assign n32982 = n28214 ^ n25799 ^ n1311 ;
  assign n32983 = n9501 & ~n32982 ;
  assign n32984 = ~n14905 & n16780 ;
  assign n32985 = n32984 ^ n16479 ^ n3385 ;
  assign n32986 = n31021 | n32985 ;
  assign n32987 = n32986 ^ n30657 ^ 1'b0 ;
  assign n32988 = ~n14328 & n20674 ;
  assign n32989 = ~n32987 & n32988 ;
  assign n32990 = n21187 ^ n18847 ^ n5435 ;
  assign n32991 = ~n2527 & n25661 ;
  assign n32992 = n32990 & n32991 ;
  assign n32993 = n32992 ^ n11702 ^ 1'b0 ;
  assign n32994 = n17040 ^ n11681 ^ n1298 ;
  assign n32995 = n5601 & n32994 ;
  assign n32996 = n5799 & n32995 ;
  assign n32997 = n9458 & n11770 ;
  assign n32998 = ( n12688 & n14471 ) | ( n12688 & ~n32997 ) | ( n14471 & ~n32997 ) ;
  assign n32999 = n4390 | n14041 ;
  assign n33000 = n21119 ^ n16046 ^ 1'b0 ;
  assign n33001 = n9113 & n33000 ;
  assign n33002 = n28777 ^ n5435 ^ 1'b0 ;
  assign n33003 = ~n11541 & n21071 ;
  assign n33004 = n22884 ^ n19646 ^ 1'b0 ;
  assign n33005 = ~n17758 & n33004 ;
  assign n33006 = n21851 & ~n27561 ;
  assign n33007 = ( n3190 & n23695 ) | ( n3190 & ~n26455 ) | ( n23695 & ~n26455 ) ;
  assign n33008 = n5104 & ~n33007 ;
  assign n33009 = n6006 | n17999 ;
  assign n33010 = ~n4688 & n8726 ;
  assign n33011 = ~n5086 & n21406 ;
  assign n33012 = n18291 ^ n15164 ^ n6680 ;
  assign n33013 = ~n7643 & n9566 ;
  assign n33014 = n30003 & n33013 ;
  assign n33015 = n18833 ^ n17664 ^ n2886 ;
  assign n33016 = n10294 & ~n33015 ;
  assign n33017 = ( n18067 & ~n30976 ) | ( n18067 & n33016 ) | ( ~n30976 & n33016 ) ;
  assign n33018 = n33017 ^ n29226 ^ n15585 ;
  assign n33019 = ( n5607 & n7926 ) | ( n5607 & n10009 ) | ( n7926 & n10009 ) ;
  assign n33020 = ( ~n2904 & n21398 ) | ( ~n2904 & n33019 ) | ( n21398 & n33019 ) ;
  assign n33021 = ( n462 & n25001 ) | ( n462 & n27082 ) | ( n25001 & n27082 ) ;
  assign n33022 = n7903 ^ n5474 ^ 1'b0 ;
  assign n33023 = n1548 & ~n7086 ;
  assign n33024 = n33023 ^ n14555 ^ 1'b0 ;
  assign n33025 = n12357 & ~n33024 ;
  assign n33026 = n33025 ^ n542 ^ 1'b0 ;
  assign n33027 = n11565 | n31526 ;
  assign n33028 = n33027 ^ n575 ^ 1'b0 ;
  assign n33029 = n19255 ^ n10030 ^ 1'b0 ;
  assign n33030 = n11730 ^ n7327 ^ 1'b0 ;
  assign n33031 = n33029 & ~n33030 ;
  assign n33032 = n20569 ^ n4823 ^ 1'b0 ;
  assign n33033 = ~n13770 & n33032 ;
  assign n33034 = ~n17524 & n33033 ;
  assign n33035 = n33034 ^ n6345 ^ 1'b0 ;
  assign n33036 = n18046 & ~n29060 ;
  assign n33037 = ( n22120 & n24095 ) | ( n22120 & n33036 ) | ( n24095 & n33036 ) ;
  assign n33038 = n22082 ^ n19731 ^ 1'b0 ;
  assign n33039 = x49 | n18224 ;
  assign n33040 = n24201 & n33039 ;
  assign n33042 = n14370 & n14421 ;
  assign n33043 = n1858 & n33042 ;
  assign n33044 = n3813 & ~n33043 ;
  assign n33045 = ~n14838 & n33044 ;
  assign n33041 = n6051 & n30481 ;
  assign n33046 = n33045 ^ n33041 ^ 1'b0 ;
  assign n33047 = n17525 ^ n2847 ^ n1614 ;
  assign n33048 = n5500 & ~n22292 ;
  assign n33049 = n33047 & n33048 ;
  assign n33050 = n16600 ^ n8486 ^ 1'b0 ;
  assign n33051 = ~n33049 & n33050 ;
  assign n33052 = ( n24497 & n25780 ) | ( n24497 & ~n28781 ) | ( n25780 & ~n28781 ) ;
  assign n33053 = ~n10420 & n33052 ;
  assign n33054 = n28255 ^ n18000 ^ n2503 ;
  assign n33055 = n8092 & ~n24910 ;
  assign n33056 = ( ~n1878 & n1887 ) | ( ~n1878 & n16136 ) | ( n1887 & n16136 ) ;
  assign n33057 = n23103 ^ n5279 ^ 1'b0 ;
  assign n33058 = n33056 & n33057 ;
  assign n33059 = ~n1186 & n32562 ;
  assign n33064 = n2698 | n9910 ;
  assign n33060 = n10816 ^ n9365 ^ 1'b0 ;
  assign n33061 = n6025 & n33060 ;
  assign n33062 = n9433 ^ n7867 ^ n3322 ;
  assign n33063 = n33061 & ~n33062 ;
  assign n33065 = n33064 ^ n33063 ^ n23671 ;
  assign n33066 = n22923 ^ n22592 ^ n10504 ;
  assign n33069 = n6334 & ~n11578 ;
  assign n33070 = n16683 & n33069 ;
  assign n33067 = ( n9927 & n17501 ) | ( n9927 & n32112 ) | ( n17501 & n32112 ) ;
  assign n33068 = ~n11134 & n33067 ;
  assign n33071 = n33070 ^ n33068 ^ 1'b0 ;
  assign n33073 = n4941 & n9936 ;
  assign n33074 = n2843 & n33073 ;
  assign n33075 = ( n5310 & n10129 ) | ( n5310 & n33074 ) | ( n10129 & n33074 ) ;
  assign n33072 = n17444 ^ n14561 ^ n6174 ;
  assign n33076 = n33075 ^ n33072 ^ 1'b0 ;
  assign n33077 = n13553 | n33076 ;
  assign n33078 = n7073 | n14075 ;
  assign n33079 = n12766 & ~n33078 ;
  assign n33080 = n16911 & n33079 ;
  assign n33081 = n12829 & ~n33080 ;
  assign n33082 = n27232 ^ n22717 ^ 1'b0 ;
  assign n33083 = n18657 ^ n9472 ^ n4442 ;
  assign n33084 = n33083 ^ n17147 ^ n2582 ;
  assign n33085 = n8438 ^ n2372 ^ 1'b0 ;
  assign n33086 = ~n355 & n8336 ;
  assign n33087 = n33086 ^ n11847 ^ 1'b0 ;
  assign n33088 = n26268 & n33087 ;
  assign n33089 = ( n7070 & n25541 ) | ( n7070 & ~n28813 ) | ( n25541 & ~n28813 ) ;
  assign n33090 = n33089 ^ n25408 ^ 1'b0 ;
  assign n33091 = ~n8952 & n18185 ;
  assign n33092 = n9478 & ~n30982 ;
  assign n33093 = n18245 & n33092 ;
  assign n33094 = n10042 & ~n33093 ;
  assign n33095 = n8763 & ~n31833 ;
  assign n33096 = n2103 & n14685 ;
  assign n33097 = n33096 ^ n19665 ^ n18657 ;
  assign n33098 = n8568 ^ n2338 ^ n1108 ;
  assign n33099 = ( x208 & n3565 ) | ( x208 & ~n33098 ) | ( n3565 & ~n33098 ) ;
  assign n33100 = n2110 & ~n10531 ;
  assign n33101 = n27204 | n33100 ;
  assign n33102 = n7740 & ~n33101 ;
  assign n33103 = ( n6149 & ~n15283 ) | ( n6149 & n23152 ) | ( ~n15283 & n23152 ) ;
  assign n33104 = ~n2215 & n5795 ;
  assign n33105 = ~n33103 & n33104 ;
  assign n33106 = ( n6554 & n17573 ) | ( n6554 & ~n17799 ) | ( n17573 & ~n17799 ) ;
  assign n33107 = n13538 ^ n7850 ^ 1'b0 ;
  assign n33108 = n26081 ^ n20881 ^ 1'b0 ;
  assign n33109 = n21661 & ~n33108 ;
  assign n33110 = ~n1685 & n10432 ;
  assign n33111 = n2960 & n33110 ;
  assign n33112 = ~n1538 & n20483 ;
  assign n33113 = ~x169 & n33112 ;
  assign n33114 = ~n4965 & n8985 ;
  assign n33115 = n16882 ^ n13308 ^ 1'b0 ;
  assign n33116 = n33115 ^ n2125 ^ 1'b0 ;
  assign n33117 = n9552 & ~n33116 ;
  assign n33118 = n19225 ^ n15688 ^ 1'b0 ;
  assign n33119 = ( n33114 & n33117 ) | ( n33114 & n33118 ) | ( n33117 & n33118 ) ;
  assign n33120 = n17753 ^ n7367 ^ 1'b0 ;
  assign n33121 = n3646 & n33120 ;
  assign n33122 = n33121 ^ n1357 ^ 1'b0 ;
  assign n33123 = n14274 & ~n33122 ;
  assign n33124 = n4688 ^ n1470 ^ 1'b0 ;
  assign n33125 = ~n3309 & n33124 ;
  assign n33126 = n2194 & n33125 ;
  assign n33127 = n33126 ^ x1 ^ 1'b0 ;
  assign n33128 = n33127 ^ n12103 ^ n3249 ;
  assign n33129 = ( n24750 & n33123 ) | ( n24750 & ~n33128 ) | ( n33123 & ~n33128 ) ;
  assign n33130 = n10078 ^ n9855 ^ n3172 ;
  assign n33131 = n6503 ^ n4603 ^ 1'b0 ;
  assign n33132 = n33130 | n33131 ;
  assign n33133 = n26900 ^ n6996 ^ 1'b0 ;
  assign n33134 = n33132 | n33133 ;
  assign n33135 = n33134 ^ n17754 ^ n6598 ;
  assign n33138 = n7935 ^ n2764 ^ 1'b0 ;
  assign n33139 = n1179 & n33138 ;
  assign n33140 = n33139 ^ n9557 ^ n2041 ;
  assign n33136 = n11458 & n14076 ;
  assign n33137 = n33136 ^ n19750 ^ 1'b0 ;
  assign n33141 = n33140 ^ n33137 ^ n26441 ;
  assign n33142 = n3513 | n14300 ;
  assign n33143 = n19223 & ~n33142 ;
  assign n33144 = n8447 ^ n6866 ^ 1'b0 ;
  assign n33145 = n17080 ^ n1705 ^ 1'b0 ;
  assign n33146 = n22238 & n33145 ;
  assign n33147 = n2892 & n5387 ;
  assign n33148 = n1630 & n33147 ;
  assign n33149 = ( n3462 & n19116 ) | ( n3462 & ~n33148 ) | ( n19116 & ~n33148 ) ;
  assign n33150 = n11955 & ~n18811 ;
  assign n33151 = ~n25342 & n33150 ;
  assign n33152 = n22559 ^ n20991 ^ n11536 ;
  assign n33153 = ~n18829 & n33152 ;
  assign n33154 = n16885 & n22801 ;
  assign n33155 = n13375 | n17734 ;
  assign n33156 = n33155 ^ n16294 ^ 1'b0 ;
  assign n33157 = n9005 | n11275 ;
  assign n33158 = n18672 & ~n33157 ;
  assign n33159 = ( n31563 & ~n33156 ) | ( n31563 & n33158 ) | ( ~n33156 & n33158 ) ;
  assign n33160 = ( n1240 & n2238 ) | ( n1240 & ~n4284 ) | ( n2238 & ~n4284 ) ;
  assign n33161 = n33160 ^ n6409 ^ 1'b0 ;
  assign n33162 = ~n9855 & n12407 ;
  assign n33163 = n20490 ^ n8306 ^ n914 ;
  assign n33164 = n33163 ^ n31126 ^ n11363 ;
  assign n33165 = n33164 ^ n3878 ^ n3172 ;
  assign n33166 = ( n2916 & n16540 ) | ( n2916 & n22416 ) | ( n16540 & n22416 ) ;
  assign n33167 = n10773 & n27882 ;
  assign n33168 = ~n14207 & n33167 ;
  assign n33169 = ~n33166 & n33168 ;
  assign n33170 = n459 & n18210 ;
  assign n33171 = n33170 ^ n8628 ^ 1'b0 ;
  assign n33172 = n33171 ^ n31361 ^ n1057 ;
  assign n33173 = n14251 ^ n1393 ^ 1'b0 ;
  assign n33174 = n33172 | n33173 ;
  assign n33175 = ~n3366 & n19819 ;
  assign n33176 = n33175 ^ n25143 ^ 1'b0 ;
  assign n33177 = x129 & ~n2260 ;
  assign n33178 = n6094 ^ n1061 ^ 1'b0 ;
  assign n33179 = n7218 & n32080 ;
  assign n33180 = ~n643 & n33179 ;
  assign n33181 = ( n262 & n5566 ) | ( n262 & ~n23313 ) | ( n5566 & ~n23313 ) ;
  assign n33182 = n2171 & ~n33181 ;
  assign n33183 = n33182 ^ n25744 ^ 1'b0 ;
  assign n33184 = n11449 | n33183 ;
  assign n33185 = n1535 & ~n33184 ;
  assign n33186 = n14805 | n33185 ;
  assign n33187 = n25419 | n33186 ;
  assign n33188 = ~n2169 & n14752 ;
  assign n33189 = n9772 & n33188 ;
  assign n33190 = n455 | n33189 ;
  assign n33191 = n17751 ^ n13070 ^ n1868 ;
  assign n33192 = n12120 & n21329 ;
  assign n33198 = n14368 ^ n1118 ^ 1'b0 ;
  assign n33199 = n10376 & ~n33198 ;
  assign n33196 = ( ~n289 & n1178 ) | ( ~n289 & n22343 ) | ( n1178 & n22343 ) ;
  assign n33194 = ~n4789 & n6859 ;
  assign n33195 = n33194 ^ n3568 ^ 1'b0 ;
  assign n33197 = n33196 ^ n33195 ^ 1'b0 ;
  assign n33193 = n13214 ^ n7552 ^ n2393 ;
  assign n33200 = n33199 ^ n33197 ^ n33193 ;
  assign n33201 = n21194 ^ n15231 ^ 1'b0 ;
  assign n33202 = ~n26110 & n33201 ;
  assign n33203 = n33202 ^ n7408 ^ 1'b0 ;
  assign n33204 = n17143 ^ n4224 ^ 1'b0 ;
  assign n33205 = n22782 | n33204 ;
  assign n33206 = n3392 | n33205 ;
  assign n33207 = n33203 & ~n33206 ;
  assign n33209 = n32326 ^ n5850 ^ n5288 ;
  assign n33208 = ~n1793 & n29454 ;
  assign n33210 = n33209 ^ n33208 ^ 1'b0 ;
  assign n33211 = ~n6840 & n13277 ;
  assign n33212 = n33211 ^ n21683 ^ 1'b0 ;
  assign n33213 = ~n13886 & n14606 ;
  assign n33214 = n33213 ^ n2654 ^ 1'b0 ;
  assign n33215 = ( ~n4312 & n28963 ) | ( ~n4312 & n33214 ) | ( n28963 & n33214 ) ;
  assign n33220 = n12806 & ~n20988 ;
  assign n33221 = ~n1091 & n33220 ;
  assign n33216 = ~n6528 & n9855 ;
  assign n33217 = x66 & n33216 ;
  assign n33218 = n33217 ^ n31824 ^ n22256 ;
  assign n33219 = n8298 & n33218 ;
  assign n33222 = n33221 ^ n33219 ^ 1'b0 ;
  assign n33223 = ( n2255 & ~n7619 ) | ( n2255 & n14463 ) | ( ~n7619 & n14463 ) ;
  assign n33224 = n33223 ^ n27293 ^ n6955 ;
  assign n33225 = n33224 ^ n8712 ^ n8075 ;
  assign n33226 = ( n13892 & n19895 ) | ( n13892 & ~n33225 ) | ( n19895 & ~n33225 ) ;
  assign n33227 = n6659 ^ n1873 ^ 1'b0 ;
  assign n33228 = ( n1252 & n2328 ) | ( n1252 & ~n3062 ) | ( n2328 & ~n3062 ) ;
  assign n33229 = n1030 | n33228 ;
  assign n33230 = n33229 ^ n7581 ^ 1'b0 ;
  assign n33231 = n15920 ^ n14935 ^ 1'b0 ;
  assign n33232 = n33231 ^ n23474 ^ n5470 ;
  assign n33233 = n33232 ^ n19785 ^ 1'b0 ;
  assign n33234 = n33230 & ~n33233 ;
  assign n33236 = n26143 ^ n9512 ^ 1'b0 ;
  assign n33237 = n28768 | n33236 ;
  assign n33235 = ( x4 & ~n14439 ) | ( x4 & n26430 ) | ( ~n14439 & n26430 ) ;
  assign n33238 = n33237 ^ n33235 ^ n21984 ;
  assign n33239 = n26578 & ~n27453 ;
  assign n33240 = ( ~n1763 & n11077 ) | ( ~n1763 & n33239 ) | ( n11077 & n33239 ) ;
  assign n33241 = n21728 ^ x69 ^ 1'b0 ;
  assign n33242 = n32211 ^ n4016 ^ 1'b0 ;
  assign n33243 = n33241 | n33242 ;
  assign n33244 = n33243 ^ n31251 ^ 1'b0 ;
  assign n33245 = n1750 & n23709 ;
  assign n33246 = n11564 | n33245 ;
  assign n33247 = ( ~n6710 & n22012 ) | ( ~n6710 & n33246 ) | ( n22012 & n33246 ) ;
  assign n33248 = n9532 | n14207 ;
  assign n33249 = n15523 & ~n33248 ;
  assign n33250 = ~n468 & n5020 ;
  assign n33251 = n33249 & n33250 ;
  assign n33252 = n764 & n19956 ;
  assign n33253 = n19034 ^ n17763 ^ 1'b0 ;
  assign n33254 = n23458 & ~n33253 ;
  assign n33255 = n27334 & n32164 ;
  assign n33256 = n18676 ^ n4040 ^ 1'b0 ;
  assign n33257 = x93 & ~n33256 ;
  assign n33258 = ~n20031 & n33257 ;
  assign n33259 = n12018 & ~n32681 ;
  assign n33260 = n33259 ^ n32946 ^ 1'b0 ;
  assign n33261 = ( ~x110 & n1179 ) | ( ~x110 & n15855 ) | ( n1179 & n15855 ) ;
  assign n33262 = ~n28897 & n33261 ;
  assign n33263 = ~n14858 & n33262 ;
  assign n33264 = n26251 ^ n9500 ^ 1'b0 ;
  assign n33265 = n22816 ^ n14524 ^ 1'b0 ;
  assign n33266 = n5369 & n33265 ;
  assign n33267 = ( n1052 & n18144 ) | ( n1052 & n21923 ) | ( n18144 & n21923 ) ;
  assign n33268 = n32753 & ~n33267 ;
  assign n33269 = ~n14529 & n33268 ;
  assign n33270 = n9547 ^ n1372 ^ 1'b0 ;
  assign n33271 = ~n16256 & n33270 ;
  assign n33272 = n33271 ^ n15334 ^ 1'b0 ;
  assign n33273 = ~n15708 & n20262 ;
  assign n33274 = n33272 & n33273 ;
  assign n33275 = ( ~n1661 & n6179 ) | ( ~n1661 & n32438 ) | ( n6179 & n32438 ) ;
  assign n33276 = ( n16204 & ~n26648 ) | ( n16204 & n28187 ) | ( ~n26648 & n28187 ) ;
  assign n33277 = n20663 ^ x180 ^ 1'b0 ;
  assign n33278 = n33088 ^ n17585 ^ 1'b0 ;
  assign n33279 = n11049 & ~n33278 ;
  assign n33280 = n33279 ^ n32934 ^ 1'b0 ;
  assign n33281 = n6132 & ~n18666 ;
  assign n33282 = n16716 & n33281 ;
  assign n33283 = n26764 ^ n23519 ^ n14632 ;
  assign n33284 = n29848 ^ n24707 ^ n19507 ;
  assign n33285 = n33284 ^ n1713 ^ 1'b0 ;
  assign n33286 = n21755 ^ n1650 ^ 1'b0 ;
  assign n33287 = n3369 | n6703 ;
  assign n33288 = ~n27365 & n32490 ;
  assign n33289 = ~n4307 & n33288 ;
  assign n33290 = ~n7327 & n14141 ;
  assign n33291 = n25422 | n33290 ;
  assign n33292 = n10440 & n11671 ;
  assign n33293 = ( n19602 & n22053 ) | ( n19602 & n25402 ) | ( n22053 & n25402 ) ;
  assign n33294 = ( n31508 & n33292 ) | ( n31508 & ~n33293 ) | ( n33292 & ~n33293 ) ;
  assign n33295 = n5817 | n7759 ;
  assign n33298 = n10580 ^ n5640 ^ 1'b0 ;
  assign n33296 = n8297 & ~n9317 ;
  assign n33297 = ~n17411 & n33296 ;
  assign n33299 = n33298 ^ n33297 ^ 1'b0 ;
  assign n33300 = n33299 ^ n11139 ^ 1'b0 ;
  assign n33303 = n15308 ^ n2677 ^ 1'b0 ;
  assign n33304 = n24027 ^ n16144 ^ 1'b0 ;
  assign n33305 = n12487 & ~n33304 ;
  assign n33306 = n33305 ^ n20210 ^ 1'b0 ;
  assign n33307 = n33303 | n33306 ;
  assign n33301 = n2403 | n25867 ;
  assign n33302 = n502 & ~n33301 ;
  assign n33308 = n33307 ^ n33302 ^ 1'b0 ;
  assign n33309 = n11515 | n33308 ;
  assign n33310 = n12963 ^ n2343 ^ 1'b0 ;
  assign n33311 = ~n19718 & n33310 ;
  assign n33312 = n19078 ^ n6689 ^ 1'b0 ;
  assign n33313 = ~n13166 & n20605 ;
  assign n33314 = ~n27625 & n33313 ;
  assign n33315 = ~n33312 & n33314 ;
  assign n33316 = n8180 & n19508 ;
  assign n33317 = n33316 ^ n21011 ^ n7366 ;
  assign n33318 = ~n5235 & n15862 ;
  assign n33319 = ( n25637 & ~n29348 ) | ( n25637 & n33318 ) | ( ~n29348 & n33318 ) ;
  assign n33320 = n33319 ^ n21343 ^ n6872 ;
  assign n33321 = n13500 & ~n18550 ;
  assign n33322 = ~n7510 & n23664 ;
  assign n33323 = n2647 & ~n11978 ;
  assign n33324 = ~n15661 & n33323 ;
  assign n33327 = n13910 ^ n4046 ^ n2470 ;
  assign n33325 = n6793 ^ n3151 ^ 1'b0 ;
  assign n33326 = n17982 & ~n33325 ;
  assign n33328 = n33327 ^ n33326 ^ n2376 ;
  assign n33329 = n33328 ^ n26472 ^ 1'b0 ;
  assign n33330 = n16333 ^ n11340 ^ 1'b0 ;
  assign n33331 = ~n17994 & n33330 ;
  assign n33332 = n33331 ^ n26755 ^ n1320 ;
  assign n33333 = n29557 ^ n2406 ^ 1'b0 ;
  assign n33334 = n32721 ^ n14624 ^ n12207 ;
  assign n33335 = n6502 & ~n17456 ;
  assign n33336 = n33335 ^ n27935 ^ n3314 ;
  assign n33337 = n14723 ^ n4405 ^ 1'b0 ;
  assign n33338 = n29030 & n33337 ;
  assign n33342 = n12192 ^ n6337 ^ 1'b0 ;
  assign n33343 = n25783 & n33342 ;
  assign n33344 = ( ~n8930 & n15438 ) | ( ~n8930 & n33343 ) | ( n15438 & n33343 ) ;
  assign n33339 = n13958 ^ n11638 ^ 1'b0 ;
  assign n33340 = n5384 & ~n33339 ;
  assign n33341 = n31622 & n33340 ;
  assign n33345 = n33344 ^ n33341 ^ 1'b0 ;
  assign n33346 = n12912 ^ n6380 ^ n3607 ;
  assign n33347 = n11289 & n33346 ;
  assign n33348 = ~n9060 & n33347 ;
  assign n33349 = n13030 & ~n33348 ;
  assign n33350 = n11144 ^ n5399 ^ 1'b0 ;
  assign n33351 = n29334 | n33350 ;
  assign n33352 = n666 & ~n33351 ;
  assign n33353 = ~n27893 & n33352 ;
  assign n33355 = n22026 ^ n18206 ^ 1'b0 ;
  assign n33356 = ~n31186 & n33355 ;
  assign n33354 = n8332 & ~n31608 ;
  assign n33357 = n33356 ^ n33354 ^ n5639 ;
  assign n33358 = ~n4917 & n11481 ;
  assign n33359 = n12682 & n33358 ;
  assign n33360 = n5349 ^ n3389 ^ n2103 ;
  assign n33361 = n27832 ^ n17787 ^ n15084 ;
  assign n33362 = ( ~n33359 & n33360 ) | ( ~n33359 & n33361 ) | ( n33360 & n33361 ) ;
  assign n33363 = n5209 ^ n3690 ^ 1'b0 ;
  assign n33364 = n14249 | n33363 ;
  assign n33365 = ~n1217 & n9018 ;
  assign n33366 = n20179 ^ n5199 ^ 1'b0 ;
  assign n33367 = n4034 & ~n33366 ;
  assign n33368 = ( ~n33364 & n33365 ) | ( ~n33364 & n33367 ) | ( n33365 & n33367 ) ;
  assign n33369 = x151 & n6912 ;
  assign n33370 = n33369 ^ n22932 ^ 1'b0 ;
  assign n33371 = n3475 & ~n33370 ;
  assign n33372 = n33371 ^ n2954 ^ 1'b0 ;
  assign n33373 = n33372 ^ n11086 ^ 1'b0 ;
  assign n33374 = n6322 & n11647 ;
  assign n33375 = n33374 ^ n7886 ^ 1'b0 ;
  assign n33376 = n10783 ^ n515 ^ 1'b0 ;
  assign n33377 = n33375 & n33376 ;
  assign n33378 = ( ~n938 & n5506 ) | ( ~n938 & n33377 ) | ( n5506 & n33377 ) ;
  assign n33379 = ( n23354 & n25473 ) | ( n23354 & ~n33378 ) | ( n25473 & ~n33378 ) ;
  assign n33380 = n1730 | n8635 ;
  assign n33381 = ~n20498 & n33380 ;
  assign n33382 = n33381 ^ n20579 ^ 1'b0 ;
  assign n33383 = n33382 ^ n15283 ^ 1'b0 ;
  assign n33384 = x153 & ~n33383 ;
  assign n33385 = n11153 | n31816 ;
  assign n33386 = ~n883 & n25284 ;
  assign n33387 = n25084 & n33386 ;
  assign n33389 = ( n10359 & n11200 ) | ( n10359 & ~n11641 ) | ( n11200 & ~n11641 ) ;
  assign n33388 = ( n15042 & n24807 ) | ( n15042 & ~n31504 ) | ( n24807 & ~n31504 ) ;
  assign n33390 = n33389 ^ n33388 ^ 1'b0 ;
  assign n33391 = ~n12614 & n33390 ;
  assign n33392 = n9944 & n33391 ;
  assign n33393 = n22491 ^ n12000 ^ n4083 ;
  assign n33394 = n32948 ^ n19951 ^ n8154 ;
  assign n33395 = ~n14038 & n17113 ;
  assign n33396 = n7500 & n33395 ;
  assign n33397 = n10703 ^ n7983 ^ 1'b0 ;
  assign n33398 = ~n1709 & n33397 ;
  assign n33399 = n33398 ^ n6442 ^ 1'b0 ;
  assign n33400 = ~n8124 & n33399 ;
  assign n33401 = ~n13658 & n29591 ;
  assign n33402 = n33401 ^ n8386 ^ 1'b0 ;
  assign n33403 = n30668 ^ n2871 ^ 1'b0 ;
  assign n33404 = n6374 & n33403 ;
  assign n33405 = ~n32503 & n33404 ;
  assign n33406 = n27029 & ~n33405 ;
  assign n33407 = n21962 & n33406 ;
  assign n33408 = n31205 ^ n29864 ^ n13850 ;
  assign n33409 = n33408 ^ n12113 ^ n2982 ;
  assign n33410 = n3792 & n7724 ;
  assign n33411 = n10396 & n33410 ;
  assign n33412 = n30834 ^ n9052 ^ 1'b0 ;
  assign n33413 = n27547 ^ n24451 ^ n9217 ;
  assign n33414 = n31912 ^ n16345 ^ 1'b0 ;
  assign n33415 = ~n24968 & n26478 ;
  assign n33416 = n33414 & n33415 ;
  assign n33417 = n17901 & n32037 ;
  assign n33418 = n5369 ^ n5019 ^ 1'b0 ;
  assign n33419 = n14945 & n33418 ;
  assign n33420 = n21757 & ~n32483 ;
  assign n33421 = ( n23493 & n33419 ) | ( n23493 & ~n33420 ) | ( n33419 & ~n33420 ) ;
  assign n33422 = ( n6695 & ~n17083 ) | ( n6695 & n26300 ) | ( ~n17083 & n26300 ) ;
  assign n33423 = ( n1582 & n8052 ) | ( n1582 & ~n9486 ) | ( n8052 & ~n9486 ) ;
  assign n33424 = n28244 ^ n5242 ^ 1'b0 ;
  assign n33425 = n15409 | n33424 ;
  assign n33426 = n33423 & ~n33425 ;
  assign n33427 = n3390 & n33426 ;
  assign n33428 = n33427 ^ n1673 ^ 1'b0 ;
  assign n33429 = n3810 & n33428 ;
  assign n33430 = n26768 ^ n6606 ^ 1'b0 ;
  assign n33431 = n25774 & n33430 ;
  assign n33432 = ~n14998 & n31420 ;
  assign n33433 = n3900 ^ n776 ^ 1'b0 ;
  assign n33434 = n30326 ^ n1018 ^ 1'b0 ;
  assign n33435 = n33434 ^ n18750 ^ 1'b0 ;
  assign n33436 = n2397 & ~n12291 ;
  assign n33437 = n32927 | n33436 ;
  assign n33438 = n21639 | n31325 ;
  assign n33439 = n29510 ^ n20525 ^ n13578 ;
  assign n33440 = n28315 ^ n2527 ^ 1'b0 ;
  assign n33441 = n3392 & n33440 ;
  assign n33442 = ( ~n840 & n6854 ) | ( ~n840 & n20710 ) | ( n6854 & n20710 ) ;
  assign n33443 = n33442 ^ n7700 ^ n7471 ;
  assign n33444 = ~n7939 & n16111 ;
  assign n33445 = n33444 ^ n2033 ^ 1'b0 ;
  assign n33446 = n33443 & ~n33445 ;
  assign n33447 = n20380 & ~n31974 ;
  assign n33448 = n33447 ^ n23110 ^ 1'b0 ;
  assign n33449 = n33446 | n33448 ;
  assign n33450 = n24742 ^ n6156 ^ 1'b0 ;
  assign n33451 = n23016 | n33450 ;
  assign n33452 = n7490 ^ n4051 ^ n521 ;
  assign n33453 = n3262 & n14899 ;
  assign n33454 = n10476 & n33453 ;
  assign n33455 = n33454 ^ n14791 ^ 1'b0 ;
  assign n33456 = n33452 | n33455 ;
  assign n33457 = ( n9980 & ~n12414 ) | ( n9980 & n33456 ) | ( ~n12414 & n33456 ) ;
  assign n33458 = n24602 & ~n31743 ;
  assign n33459 = n4274 ^ n1624 ^ 1'b0 ;
  assign n33460 = x134 & n33459 ;
  assign n33461 = ( n6423 & ~n9647 ) | ( n6423 & n15305 ) | ( ~n9647 & n15305 ) ;
  assign n33462 = ~n18419 & n25027 ;
  assign n33463 = ~n33461 & n33462 ;
  assign n33464 = ( n20605 & n33460 ) | ( n20605 & n33463 ) | ( n33460 & n33463 ) ;
  assign n33465 = n10631 ^ n4439 ^ n2931 ;
  assign n33467 = n4139 ^ n3646 ^ 1'b0 ;
  assign n33468 = n29449 & n33467 ;
  assign n33466 = n7178 | n8781 ;
  assign n33469 = n33468 ^ n33466 ^ 1'b0 ;
  assign n33470 = ( n6912 & n19570 ) | ( n6912 & n33469 ) | ( n19570 & n33469 ) ;
  assign n33471 = n12417 ^ n7101 ^ 1'b0 ;
  assign n33472 = ~n16322 & n33471 ;
  assign n33473 = n1983 | n8156 ;
  assign n33474 = n33473 ^ n495 ^ 1'b0 ;
  assign n33475 = n27021 | n33474 ;
  assign n33476 = n1664 | n33475 ;
  assign n33477 = ~n9989 & n16483 ;
  assign n33478 = ~n33476 & n33477 ;
  assign n33479 = ( n33470 & n33472 ) | ( n33470 & n33478 ) | ( n33472 & n33478 ) ;
  assign n33480 = n11496 | n33479 ;
  assign n33481 = n33480 ^ n17876 ^ 1'b0 ;
  assign n33482 = n17465 ^ n5092 ^ 1'b0 ;
  assign n33483 = n699 | n11800 ;
  assign n33484 = n33483 ^ n10631 ^ 1'b0 ;
  assign n33485 = n18311 & ~n33484 ;
  assign n33486 = ~n2231 & n7027 ;
  assign n33487 = ( n18573 & n23784 ) | ( n18573 & n33486 ) | ( n23784 & n33486 ) ;
  assign n33488 = n33487 ^ n8241 ^ 1'b0 ;
  assign n33489 = n33485 & ~n33488 ;
  assign n33490 = n23684 ^ n20158 ^ n4870 ;
  assign n33491 = n33490 ^ n28010 ^ 1'b0 ;
  assign n33493 = n14539 & n18361 ;
  assign n33492 = n5898 & ~n11250 ;
  assign n33494 = n33493 ^ n33492 ^ n13255 ;
  assign n33495 = ( n2317 & n5517 ) | ( n2317 & n17359 ) | ( n5517 & n17359 ) ;
  assign n33496 = n33495 ^ n29237 ^ 1'b0 ;
  assign n33497 = ~x44 & n25737 ;
  assign n33498 = n4098 ^ n2808 ^ 1'b0 ;
  assign n33499 = n6176 | n33498 ;
  assign n33500 = n6246 & ~n23142 ;
  assign n33501 = n33500 ^ n32811 ^ 1'b0 ;
  assign n33502 = n4873 & ~n5104 ;
  assign n33503 = n8191 & n21241 ;
  assign n33504 = ~n33502 & n33503 ;
  assign n33505 = n23419 ^ n15085 ^ n2845 ;
  assign n33506 = ( n5264 & n31544 ) | ( n5264 & ~n33505 ) | ( n31544 & ~n33505 ) ;
  assign n33507 = n33506 ^ n25815 ^ n19066 ;
  assign n33508 = n932 | n6681 ;
  assign n33509 = n33508 ^ n14105 ^ 1'b0 ;
  assign n33510 = n33509 ^ n16208 ^ n6120 ;
  assign n33511 = ( n4564 & ~n7125 ) | ( n4564 & n19818 ) | ( ~n7125 & n19818 ) ;
  assign n33512 = ( n15244 & n19829 ) | ( n15244 & n33511 ) | ( n19829 & n33511 ) ;
  assign n33513 = ~n2536 & n5090 ;
  assign n33514 = n29654 ^ x25 ^ 1'b0 ;
  assign n33515 = ( ~n18467 & n33513 ) | ( ~n18467 & n33514 ) | ( n33513 & n33514 ) ;
  assign n33516 = ~n5639 & n7094 ;
  assign n33517 = n33516 ^ n23488 ^ n13758 ;
  assign n33518 = n3512 & ~n14573 ;
  assign n33519 = n20548 ^ n6996 ^ 1'b0 ;
  assign n33520 = n33519 ^ n32553 ^ n17894 ;
  assign n33521 = n13028 ^ n4279 ^ 1'b0 ;
  assign n33522 = n2291 & n25618 ;
  assign n33523 = ~n666 & n27199 ;
  assign n33524 = n15597 ^ n3720 ^ 1'b0 ;
  assign n33525 = n20236 & n33524 ;
  assign n33526 = ( n10502 & n17682 ) | ( n10502 & n33525 ) | ( n17682 & n33525 ) ;
  assign n33527 = ( ~n7500 & n8400 ) | ( ~n7500 & n26528 ) | ( n8400 & n26528 ) ;
  assign n33528 = ( n11371 & n33526 ) | ( n11371 & ~n33527 ) | ( n33526 & ~n33527 ) ;
  assign n33529 = ( n12675 & n18484 ) | ( n12675 & ~n33501 ) | ( n18484 & ~n33501 ) ;
  assign n33530 = ( n5894 & n30026 ) | ( n5894 & ~n31434 ) | ( n30026 & ~n31434 ) ;
  assign n33531 = n33530 ^ n12008 ^ 1'b0 ;
  assign n33532 = ~n14592 & n33531 ;
  assign n33533 = n24850 ^ n1149 ^ 1'b0 ;
  assign n33534 = n30808 | n33533 ;
  assign n33535 = n31205 | n33534 ;
  assign n33536 = n21816 | n31174 ;
  assign n33539 = n6406 ^ n2994 ^ 1'b0 ;
  assign n33537 = n2724 & ~n2838 ;
  assign n33538 = ~n11143 & n33537 ;
  assign n33540 = n33539 ^ n33538 ^ n5741 ;
  assign n33541 = x93 & n2948 ;
  assign n33542 = n11632 ^ n5082 ^ 1'b0 ;
  assign n33543 = n33542 ^ n6328 ^ 1'b0 ;
  assign n33544 = n10127 & ~n33543 ;
  assign n33545 = n33544 ^ n6563 ^ 1'b0 ;
  assign n33546 = ~n33541 & n33545 ;
  assign n33547 = n3525 & ~n33546 ;
  assign n33548 = n33547 ^ n24430 ^ 1'b0 ;
  assign n33549 = n16058 & ~n33548 ;
  assign n33550 = n28150 ^ n4241 ^ 1'b0 ;
  assign n33551 = n28300 ^ n3383 ^ 1'b0 ;
  assign n33552 = n8442 | n8881 ;
  assign n33553 = n33552 ^ n29374 ^ 1'b0 ;
  assign n33554 = n25074 ^ n4156 ^ 1'b0 ;
  assign n33555 = ~n3330 & n33554 ;
  assign n33556 = n17237 ^ n11536 ^ n6063 ;
  assign n33557 = ( n3222 & n30420 ) | ( n3222 & n33513 ) | ( n30420 & n33513 ) ;
  assign n33558 = ( ~n6889 & n7581 ) | ( ~n6889 & n10053 ) | ( n7581 & n10053 ) ;
  assign n33559 = ~n8108 & n17876 ;
  assign n33560 = ~n33558 & n33559 ;
  assign n33561 = n6101 ^ n3021 ^ n2160 ;
  assign n33562 = n4823 | n33561 ;
  assign n33563 = n10376 | n33562 ;
  assign n33564 = n33563 ^ n7408 ^ 1'b0 ;
  assign n33565 = n10599 | n33564 ;
  assign n33566 = n24377 ^ n1134 ^ 1'b0 ;
  assign n33567 = n33566 ^ n25986 ^ 1'b0 ;
  assign n33568 = n26289 ^ n8953 ^ 1'b0 ;
  assign n33569 = n18786 & ~n33568 ;
  assign n33570 = n33569 ^ n31437 ^ x78 ;
  assign n33571 = x159 & ~n8758 ;
  assign n33573 = n5193 & ~n13491 ;
  assign n33574 = n33573 ^ n10111 ^ 1'b0 ;
  assign n33575 = n6865 & n33574 ;
  assign n33576 = n6244 & n33575 ;
  assign n33572 = n4826 & ~n27210 ;
  assign n33577 = n33576 ^ n33572 ^ n26501 ;
  assign n33578 = n6706 & n33577 ;
  assign n33579 = n13456 | n33578 ;
  assign n33580 = n5499 & n26911 ;
  assign n33581 = n23156 & ~n25191 ;
  assign n33582 = n25323 ^ n2040 ^ 1'b0 ;
  assign n33583 = n11693 | n33582 ;
  assign n33584 = x105 & ~n31708 ;
  assign n33585 = n33584 ^ n4963 ^ n2686 ;
  assign n33586 = ( n276 & n2649 ) | ( n276 & n3568 ) | ( n2649 & n3568 ) ;
  assign n33587 = ~n12682 & n33586 ;
  assign n33588 = n4979 & n33587 ;
  assign n33589 = n33588 ^ n17917 ^ n9320 ;
  assign n33590 = n18764 | n33589 ;
  assign n33591 = n13143 ^ n6281 ^ 1'b0 ;
  assign n33592 = n16417 ^ n10354 ^ 1'b0 ;
  assign n33593 = n33591 & ~n33592 ;
  assign n33594 = ~n23419 & n33593 ;
  assign n33595 = n33594 ^ n15906 ^ n12285 ;
  assign n33597 = n22366 & ~n28164 ;
  assign n33596 = n12031 & n28467 ;
  assign n33598 = n33597 ^ n33596 ^ 1'b0 ;
  assign n33599 = ~n11102 & n12881 ;
  assign n33600 = n33598 & n33599 ;
  assign n33601 = n2677 & n10113 ;
  assign n33602 = n16754 ^ n2062 ^ 1'b0 ;
  assign n33603 = n33601 & ~n33602 ;
  assign n33604 = ~n13674 & n30647 ;
  assign n33605 = n33604 ^ n9294 ^ 1'b0 ;
  assign n33606 = ( n11147 & n19218 ) | ( n11147 & ~n33605 ) | ( n19218 & ~n33605 ) ;
  assign n33607 = ( n666 & n33603 ) | ( n666 & n33606 ) | ( n33603 & n33606 ) ;
  assign n33608 = n15807 & ~n19775 ;
  assign n33609 = ~n33607 & n33608 ;
  assign n33610 = n30204 ^ n18588 ^ 1'b0 ;
  assign n33611 = ~n9359 & n28817 ;
  assign n33615 = n25130 ^ n5844 ^ n4868 ;
  assign n33612 = n3995 & ~n7898 ;
  assign n33613 = ~n32956 & n33612 ;
  assign n33614 = n24707 & n33613 ;
  assign n33616 = n33615 ^ n33614 ^ n30346 ;
  assign n33617 = ( n4113 & ~n9562 ) | ( n4113 & n30118 ) | ( ~n9562 & n30118 ) ;
  assign n33618 = n25060 ^ n14594 ^ 1'b0 ;
  assign n33619 = n24027 ^ n7904 ^ n5767 ;
  assign n33620 = n10605 & n24744 ;
  assign n33621 = n4589 & n33620 ;
  assign n33622 = n14627 & ~n17509 ;
  assign n33623 = ~n14052 & n33622 ;
  assign n33624 = n5919 | n33623 ;
  assign n33625 = n2718 & ~n33624 ;
  assign n33626 = n33327 ^ n25923 ^ 1'b0 ;
  assign n33627 = n19496 | n33626 ;
  assign n33628 = n15302 ^ n10900 ^ n7669 ;
  assign n33629 = n33628 ^ n23617 ^ n15846 ;
  assign n33630 = n33629 ^ n24814 ^ n8946 ;
  assign n33631 = ~n4615 & n7655 ;
  assign n33632 = ( n6428 & n23790 ) | ( n6428 & ~n25352 ) | ( n23790 & ~n25352 ) ;
  assign n33633 = n15794 ^ n10863 ^ 1'b0 ;
  assign n33634 = ( n284 & ~n1662 ) | ( n284 & n11043 ) | ( ~n1662 & n11043 ) ;
  assign n33635 = ( n640 & ~n12694 ) | ( n640 & n16631 ) | ( ~n12694 & n16631 ) ;
  assign n33636 = n33634 | n33635 ;
  assign n33637 = n33636 ^ n6404 ^ 1'b0 ;
  assign n33638 = ( n7185 & n33633 ) | ( n7185 & n33637 ) | ( n33633 & n33637 ) ;
  assign n33639 = n26614 & ~n33638 ;
  assign n33640 = ~n33632 & n33639 ;
  assign n33641 = n13464 ^ n4432 ^ n4171 ;
  assign n33642 = n12775 ^ n6299 ^ 1'b0 ;
  assign n33643 = n8208 & n33642 ;
  assign n33644 = n33643 ^ n6321 ^ 1'b0 ;
  assign n33645 = n33644 ^ n26781 ^ n18345 ;
  assign n33646 = n33641 | n33645 ;
  assign n33648 = n6285 | n8517 ;
  assign n33647 = ( ~n8705 & n9831 ) | ( ~n8705 & n15727 ) | ( n9831 & n15727 ) ;
  assign n33649 = n33648 ^ n33647 ^ 1'b0 ;
  assign n33650 = n20459 | n33649 ;
  assign n33651 = n405 & ~n12921 ;
  assign n33652 = n33650 & n33651 ;
  assign n33653 = n1776 | n33652 ;
  assign n33654 = n33653 ^ n17756 ^ 1'b0 ;
  assign n33656 = n12098 ^ n1689 ^ 1'b0 ;
  assign n33655 = n11864 ^ n4581 ^ n1604 ;
  assign n33657 = n33656 ^ n33655 ^ n9013 ;
  assign n33658 = ( ~n3995 & n11292 ) | ( ~n3995 & n12899 ) | ( n11292 & n12899 ) ;
  assign n33659 = n33658 ^ n13929 ^ n409 ;
  assign n33660 = n33659 ^ n11371 ^ 1'b0 ;
  assign n33661 = ( n5167 & n11737 ) | ( n5167 & n26956 ) | ( n11737 & n26956 ) ;
  assign n33662 = n10796 | n18565 ;
  assign n33663 = n3634 | n33662 ;
  assign n33664 = n33663 ^ n5935 ^ 1'b0 ;
  assign n33665 = n33661 & n33664 ;
  assign n33666 = n11607 & ~n17870 ;
  assign n33670 = n11173 ^ n7755 ^ n6070 ;
  assign n33667 = ~n1128 & n10588 ;
  assign n33668 = ~n8292 & n33667 ;
  assign n33669 = n28733 | n33668 ;
  assign n33671 = n33670 ^ n33669 ^ 1'b0 ;
  assign n33672 = n19911 ^ n19689 ^ 1'b0 ;
  assign n33673 = n4371 | n33672 ;
  assign n33674 = n6632 & ~n15317 ;
  assign n33675 = n19228 ^ n18673 ^ 1'b0 ;
  assign n33676 = ~n32459 & n33675 ;
  assign n33677 = n33676 ^ n24115 ^ 1'b0 ;
  assign n33678 = ~n33674 & n33677 ;
  assign n33679 = n19256 & n32417 ;
  assign n33680 = n33679 ^ n29580 ^ 1'b0 ;
  assign n33681 = n2276 & ~n33680 ;
  assign n33682 = n22595 & ~n24312 ;
  assign n33683 = n19084 & n33682 ;
  assign n33684 = n33683 ^ n22652 ^ 1'b0 ;
  assign n33685 = ( n6546 & n24749 ) | ( n6546 & n33684 ) | ( n24749 & n33684 ) ;
  assign n33686 = n2760 | n8103 ;
  assign n33687 = n33686 ^ n4520 ^ 1'b0 ;
  assign n33688 = ( n10595 & n26762 ) | ( n10595 & n33687 ) | ( n26762 & n33687 ) ;
  assign n33689 = n21167 & ~n33688 ;
  assign n33690 = n3780 & ~n33689 ;
  assign n33691 = ( n6648 & n13757 ) | ( n6648 & n18734 ) | ( n13757 & n18734 ) ;
  assign n33692 = n29237 ^ n5424 ^ n1470 ;
  assign n33693 = n33692 ^ n11126 ^ 1'b0 ;
  assign n33694 = n11002 | n16023 ;
  assign n33695 = n33694 ^ n30310 ^ 1'b0 ;
  assign n33696 = ~n31883 & n33695 ;
  assign n33697 = n33696 ^ n32830 ^ 1'b0 ;
  assign n33698 = n2127 & n28304 ;
  assign n33699 = n7491 & n33698 ;
  assign n33700 = n7511 & n12338 ;
  assign n33701 = ~n6369 & n33700 ;
  assign n33702 = n33701 ^ n11340 ^ 1'b0 ;
  assign n33703 = n24128 | n33702 ;
  assign n33704 = n33703 ^ n24309 ^ 1'b0 ;
  assign n33705 = ( n4825 & n5154 ) | ( n4825 & ~n20747 ) | ( n5154 & ~n20747 ) ;
  assign n33706 = n33705 ^ n13176 ^ 1'b0 ;
  assign n33707 = n33704 & n33706 ;
  assign n33708 = n17082 & n20832 ;
  assign n33709 = ~n17982 & n33708 ;
  assign n33712 = ( ~x96 & n25939 ) | ( ~x96 & n26522 ) | ( n25939 & n26522 ) ;
  assign n33713 = ( n9005 & ~n19431 ) | ( n9005 & n33712 ) | ( ~n19431 & n33712 ) ;
  assign n33710 = n26868 ^ n21017 ^ 1'b0 ;
  assign n33711 = ( n1877 & n24560 ) | ( n1877 & ~n33710 ) | ( n24560 & ~n33710 ) ;
  assign n33714 = n33713 ^ n33711 ^ n17697 ;
  assign n33715 = n25306 & n25571 ;
  assign n33716 = ~n4516 & n33715 ;
  assign n33717 = ( x109 & n4083 ) | ( x109 & n25944 ) | ( n4083 & n25944 ) ;
  assign n33718 = ~n4455 & n32968 ;
  assign n33719 = ~n33717 & n33718 ;
  assign n33720 = n12390 & ~n33719 ;
  assign n33721 = n33720 ^ n32556 ^ 1'b0 ;
  assign n33722 = n26305 ^ n12160 ^ n7375 ;
  assign n33724 = n7986 ^ n5507 ^ 1'b0 ;
  assign n33723 = n33134 ^ n32132 ^ 1'b0 ;
  assign n33725 = n33724 ^ n33723 ^ n25491 ;
  assign n33726 = ( n10815 & n12601 ) | ( n10815 & n17497 ) | ( n12601 & n17497 ) ;
  assign n33727 = ( n14901 & ~n33127 ) | ( n14901 & n33726 ) | ( ~n33127 & n33726 ) ;
  assign n33728 = n12682 ^ n11628 ^ 1'b0 ;
  assign n33729 = n10294 & ~n33728 ;
  assign n33730 = n29454 ^ n9766 ^ n9710 ;
  assign n33731 = n33730 ^ n20802 ^ n6848 ;
  assign n33732 = ( n3668 & ~n10212 ) | ( n3668 & n19803 ) | ( ~n10212 & n19803 ) ;
  assign n33733 = ( n11058 & n27883 ) | ( n11058 & n33732 ) | ( n27883 & n33732 ) ;
  assign n33734 = ( n8767 & ~n11084 ) | ( n8767 & n13755 ) | ( ~n11084 & n13755 ) ;
  assign n33735 = n33734 ^ n414 ^ 1'b0 ;
  assign n33736 = n33735 ^ n12146 ^ n6545 ;
  assign n33737 = n21547 ^ n11795 ^ 1'b0 ;
  assign n33738 = n5763 & n28695 ;
  assign n33739 = n20780 & n33738 ;
  assign n33740 = n30833 ^ n1740 ^ 1'b0 ;
  assign n33741 = n33740 ^ n18699 ^ n7159 ;
  assign n33742 = ~n4005 & n13579 ;
  assign n33743 = n33742 ^ n25904 ^ 1'b0 ;
  assign n33744 = n33743 ^ n15147 ^ n14239 ;
  assign n33745 = n19945 ^ n9976 ^ 1'b0 ;
  assign n33746 = ( n1127 & n21435 ) | ( n1127 & ~n21906 ) | ( n21435 & ~n21906 ) ;
  assign n33747 = ( n21930 & n33745 ) | ( n21930 & ~n33746 ) | ( n33745 & ~n33746 ) ;
  assign n33749 = ~x0 & n7549 ;
  assign n33750 = n10801 & n33749 ;
  assign n33748 = n3888 & n25067 ;
  assign n33751 = n33750 ^ n33748 ^ 1'b0 ;
  assign n33752 = ~n14221 & n27469 ;
  assign n33753 = ~n6252 & n33752 ;
  assign n33754 = n33753 ^ n3096 ^ 1'b0 ;
  assign n33755 = ( n10523 & n17193 ) | ( n10523 & ~n33754 ) | ( n17193 & ~n33754 ) ;
  assign n33757 = n16416 ^ n15575 ^ n4242 ;
  assign n33756 = n10630 ^ n663 ^ 1'b0 ;
  assign n33758 = n33757 ^ n33756 ^ n12796 ;
  assign n33759 = ( ~n2492 & n3945 ) | ( ~n2492 & n25171 ) | ( n3945 & n25171 ) ;
  assign n33760 = ( n10623 & n18985 ) | ( n10623 & ~n25399 ) | ( n18985 & ~n25399 ) ;
  assign n33761 = n17782 & n33760 ;
  assign n33762 = ~n7759 & n7917 ;
  assign n33763 = n33762 ^ n28606 ^ 1'b0 ;
  assign n33764 = n32873 ^ n19511 ^ n7252 ;
  assign n33765 = ( ~n18089 & n33763 ) | ( ~n18089 & n33764 ) | ( n33763 & n33764 ) ;
  assign n33766 = n30895 ^ n25968 ^ n2488 ;
  assign n33767 = ( n1001 & n4672 ) | ( n1001 & ~n11460 ) | ( n4672 & ~n11460 ) ;
  assign n33768 = n7688 | n33767 ;
  assign n33769 = n33768 ^ n6042 ^ 1'b0 ;
  assign n33770 = n3844 ^ n2862 ^ 1'b0 ;
  assign n33771 = n13575 & n33770 ;
  assign n33772 = ( ~n33156 & n33225 ) | ( ~n33156 & n33771 ) | ( n33225 & n33771 ) ;
  assign n33773 = n15152 ^ n8174 ^ n2533 ;
  assign n33774 = n33773 ^ n19597 ^ 1'b0 ;
  assign n33775 = n20747 | n33774 ;
  assign n33776 = n33775 ^ n21454 ^ n7123 ;
  assign n33777 = n33776 ^ n24938 ^ 1'b0 ;
  assign n33778 = ~n11762 & n33777 ;
  assign n33779 = n33778 ^ n21305 ^ 1'b0 ;
  assign n33780 = n8254 & n14247 ;
  assign n33781 = n33780 ^ n15230 ^ 1'b0 ;
  assign n33782 = n21982 ^ n16162 ^ 1'b0 ;
  assign n33783 = n33781 & n33782 ;
  assign n33784 = x244 & ~n870 ;
  assign n33785 = n33784 ^ n23850 ^ 1'b0 ;
  assign n33786 = n13512 ^ n9559 ^ 1'b0 ;
  assign n33787 = ( n21406 & n23438 ) | ( n21406 & n33786 ) | ( n23438 & n33786 ) ;
  assign n33788 = n7331 & ~n8463 ;
  assign n33789 = n33659 ^ n10626 ^ 1'b0 ;
  assign n33790 = n26300 & ~n33789 ;
  assign n33791 = ( n7527 & n33788 ) | ( n7527 & n33790 ) | ( n33788 & n33790 ) ;
  assign n33792 = ~x214 & n14366 ;
  assign n33793 = n13480 | n33792 ;
  assign n33794 = n6967 & ~n33793 ;
  assign n33795 = x106 & n20362 ;
  assign n33796 = n27753 ^ n10872 ^ 1'b0 ;
  assign n33797 = n4711 & n33796 ;
  assign n33798 = n12113 ^ n4581 ^ n1886 ;
  assign n33799 = n17861 ^ n13125 ^ n4708 ;
  assign n33800 = n18240 | n25148 ;
  assign n33801 = n33799 & ~n33800 ;
  assign n33802 = n33798 | n33801 ;
  assign n33803 = ~n17633 & n33802 ;
  assign n33804 = ~n20444 & n33803 ;
  assign n33805 = n19453 ^ n904 ^ 1'b0 ;
  assign n33806 = n4686 & n33805 ;
  assign n33807 = n20742 ^ n12977 ^ n5445 ;
  assign n33808 = n33807 ^ n33447 ^ 1'b0 ;
  assign n33809 = n16387 ^ n4212 ^ 1'b0 ;
  assign n33812 = n13819 ^ n7597 ^ n4037 ;
  assign n33810 = n6440 & n9499 ;
  assign n33811 = n5171 & n33810 ;
  assign n33813 = n33812 ^ n33811 ^ n4675 ;
  assign n33814 = n18746 ^ n17632 ^ n11738 ;
  assign n33815 = ( n23674 & ~n29924 ) | ( n23674 & n33814 ) | ( ~n29924 & n33814 ) ;
  assign n33816 = n6770 & n23015 ;
  assign n33817 = n33816 ^ n21606 ^ n4251 ;
  assign n33818 = ~n9225 & n32258 ;
  assign n33819 = n11164 ^ n7424 ^ 1'b0 ;
  assign n33821 = n26024 ^ n14380 ^ 1'b0 ;
  assign n33822 = ( n15234 & ~n19707 ) | ( n15234 & n33821 ) | ( ~n19707 & n33821 ) ;
  assign n33820 = n5724 | n31159 ;
  assign n33823 = n33822 ^ n33820 ^ n13208 ;
  assign n33824 = ( ~n3311 & n6242 ) | ( ~n3311 & n20974 ) | ( n6242 & n20974 ) ;
  assign n33826 = n16918 & n23598 ;
  assign n33827 = n33826 ^ n10197 ^ 1'b0 ;
  assign n33825 = n2525 & n5746 ;
  assign n33828 = n33827 ^ n33825 ^ 1'b0 ;
  assign n33829 = ( ~n28235 & n33824 ) | ( ~n28235 & n33828 ) | ( n33824 & n33828 ) ;
  assign n33830 = n16471 ^ n14551 ^ n3704 ;
  assign n33831 = n1729 | n33830 ;
  assign n33832 = n28998 ^ n18008 ^ n1511 ;
  assign n33833 = ( ~n29661 & n33831 ) | ( ~n29661 & n33832 ) | ( n33831 & n33832 ) ;
  assign n33834 = ~n8976 & n28204 ;
  assign n33835 = n33834 ^ n32254 ^ 1'b0 ;
  assign n33836 = n10727 & ~n16063 ;
  assign n33837 = ~n33835 & n33836 ;
  assign n33838 = n19722 & ~n33837 ;
  assign n33839 = ( n7926 & n23709 ) | ( n7926 & n25043 ) | ( n23709 & n25043 ) ;
  assign n33840 = ( n19827 & n26818 ) | ( n19827 & ~n33839 ) | ( n26818 & ~n33839 ) ;
  assign n33841 = ( n24247 & ~n31532 ) | ( n24247 & n33840 ) | ( ~n31532 & n33840 ) ;
  assign n33842 = ~n3546 & n12826 ;
  assign n33844 = n31571 ^ n8952 ^ 1'b0 ;
  assign n33843 = n12872 & ~n33193 ;
  assign n33845 = n33844 ^ n33843 ^ 1'b0 ;
  assign n33846 = n16985 ^ n7326 ^ n3782 ;
  assign n33848 = ~n386 & n12976 ;
  assign n33849 = ~n3581 & n33848 ;
  assign n33850 = n27766 | n33849 ;
  assign n33847 = n27783 & n30728 ;
  assign n33851 = n33850 ^ n33847 ^ n19642 ;
  assign n33852 = ( n7241 & n13315 ) | ( n7241 & ~n15879 ) | ( n13315 & ~n15879 ) ;
  assign n33853 = n22631 & ~n22958 ;
  assign n33854 = n5439 ^ n4995 ^ 1'b0 ;
  assign n33855 = n33853 | n33854 ;
  assign n33856 = n348 & n1743 ;
  assign n33857 = n33856 ^ n31539 ^ 1'b0 ;
  assign n33858 = n33857 ^ n21160 ^ 1'b0 ;
  assign n33859 = n5173 ^ n1445 ^ 1'b0 ;
  assign n33860 = ( ~n1363 & n11483 ) | ( ~n1363 & n14130 ) | ( n11483 & n14130 ) ;
  assign n33861 = n33860 ^ n3932 ^ 1'b0 ;
  assign n33862 = ~n13600 & n33861 ;
  assign n33863 = ~n33859 & n33862 ;
  assign n33864 = n11501 ^ n1988 ^ 1'b0 ;
  assign n33865 = n33864 ^ n22847 ^ 1'b0 ;
  assign n33866 = n4302 ^ n1279 ^ 1'b0 ;
  assign n33867 = ( n26614 & n33865 ) | ( n26614 & ~n33866 ) | ( n33865 & ~n33866 ) ;
  assign n33868 = n19420 ^ n6557 ^ 1'b0 ;
  assign n33869 = n4765 & ~n10793 ;
  assign n33870 = n262 & n33869 ;
  assign n33871 = n14783 | n18585 ;
  assign n33872 = n12063 & ~n33871 ;
  assign n33873 = n33872 ^ n12819 ^ n8018 ;
  assign n33874 = ( n18680 & n19290 ) | ( n18680 & n31277 ) | ( n19290 & n31277 ) ;
  assign n33875 = ( n12687 & n33873 ) | ( n12687 & ~n33874 ) | ( n33873 & ~n33874 ) ;
  assign n33876 = ( ~n3205 & n32180 ) | ( ~n3205 & n33875 ) | ( n32180 & n33875 ) ;
  assign n33877 = n1697 | n13869 ;
  assign n33878 = n33877 ^ n13578 ^ n12722 ;
  assign n33879 = n22690 & n23286 ;
  assign n33880 = n33879 ^ n1698 ^ 1'b0 ;
  assign n33881 = ( ~n8022 & n23664 ) | ( ~n8022 & n33880 ) | ( n23664 & n33880 ) ;
  assign n33882 = ( n4242 & ~n9769 ) | ( n4242 & n24762 ) | ( ~n9769 & n24762 ) ;
  assign n33883 = ( x248 & ~n27487 ) | ( x248 & n30948 ) | ( ~n27487 & n30948 ) ;
  assign n33885 = n28316 ^ n15170 ^ n690 ;
  assign n33884 = ~n19492 & n27089 ;
  assign n33886 = n33885 ^ n33884 ^ 1'b0 ;
  assign n33887 = n27574 ^ n12289 ^ 1'b0 ;
  assign n33888 = n4027 ^ x73 ^ 1'b0 ;
  assign n33889 = n807 | n22524 ;
  assign n33890 = ( n22531 & ~n33888 ) | ( n22531 & n33889 ) | ( ~n33888 & n33889 ) ;
  assign n33891 = n33578 ^ n16638 ^ 1'b0 ;
  assign n33892 = n31473 & n33891 ;
  assign n33893 = n6297 | n18472 ;
  assign n33894 = n2499 | n33893 ;
  assign n33897 = n31704 ^ n25135 ^ 1'b0 ;
  assign n33895 = ~n9306 & n15550 ;
  assign n33896 = n33895 ^ n10004 ^ 1'b0 ;
  assign n33898 = n33897 ^ n33896 ^ n22184 ;
  assign n33899 = n33894 & ~n33898 ;
  assign n33900 = n33899 ^ n8390 ^ 1'b0 ;
  assign n33901 = ( n5710 & n11138 ) | ( n5710 & ~n30575 ) | ( n11138 & ~n30575 ) ;
  assign n33902 = n33901 ^ n2247 ^ 1'b0 ;
  assign n33903 = ~n20867 & n33902 ;
  assign n33904 = n9430 & n14288 ;
  assign n33905 = n30815 & n33904 ;
  assign n33906 = n8453 | n27976 ;
  assign n33907 = n32499 | n33906 ;
  assign n33908 = ( n29415 & n33409 ) | ( n29415 & n33907 ) | ( n33409 & n33907 ) ;
  assign n33909 = n14283 | n28660 ;
  assign n33910 = n9521 | n33909 ;
  assign n33911 = ( ~n3930 & n9481 ) | ( ~n3930 & n33910 ) | ( n9481 & n33910 ) ;
  assign n33912 = n15301 ^ n8382 ^ 1'b0 ;
  assign n33914 = ~n381 & n10149 ;
  assign n33915 = n6640 & ~n33914 ;
  assign n33913 = n9566 ^ n8743 ^ n8740 ;
  assign n33916 = n33915 ^ n33913 ^ n16078 ;
  assign n33923 = n18085 & n21949 ;
  assign n33924 = n33923 ^ n20842 ^ 1'b0 ;
  assign n33917 = n3068 ^ n1654 ^ 1'b0 ;
  assign n33918 = n4129 | n33917 ;
  assign n33919 = n19258 ^ n13229 ^ n9184 ;
  assign n33920 = n33919 ^ n11583 ^ 1'b0 ;
  assign n33921 = n11659 & n33920 ;
  assign n33922 = ~n33918 & n33921 ;
  assign n33925 = n33924 ^ n33922 ^ 1'b0 ;
  assign n33926 = n27452 ^ n24424 ^ 1'b0 ;
  assign n33927 = n22658 ^ n14723 ^ n5554 ;
  assign n33928 = n33927 ^ n868 ^ 1'b0 ;
  assign n33929 = ( n389 & ~n5990 ) | ( n389 & n14644 ) | ( ~n5990 & n14644 ) ;
  assign n33930 = n16230 & n33929 ;
  assign n33935 = n15731 ^ n8231 ^ 1'b0 ;
  assign n33936 = n5070 & n17257 ;
  assign n33937 = ~n5122 & n33936 ;
  assign n33938 = ( n3254 & ~n16924 ) | ( n3254 & n33937 ) | ( ~n16924 & n33937 ) ;
  assign n33939 = n33935 & ~n33938 ;
  assign n33940 = n33939 ^ n22332 ^ n15196 ;
  assign n33934 = n22807 ^ n3062 ^ 1'b0 ;
  assign n33931 = n10263 & ~n14966 ;
  assign n33932 = ~n5390 & n33931 ;
  assign n33933 = n2400 & n33932 ;
  assign n33941 = n33940 ^ n33934 ^ n33933 ;
  assign n33944 = n23598 & n25225 ;
  assign n33945 = n33944 ^ n26470 ^ n5322 ;
  assign n33942 = x127 | n28536 ;
  assign n33943 = ~n8776 & n33942 ;
  assign n33946 = n33945 ^ n33943 ^ 1'b0 ;
  assign n33947 = n15734 ^ n7990 ^ 1'b0 ;
  assign n33948 = n23440 | n31151 ;
  assign n33949 = n23145 & ~n33948 ;
  assign n33950 = ~n2094 & n33030 ;
  assign n33951 = n10257 | n25293 ;
  assign n33952 = n12064 | n33951 ;
  assign n33953 = n21236 ^ n2041 ^ 1'b0 ;
  assign n33954 = n32994 & n33953 ;
  assign n33955 = n5424 & ~n33954 ;
  assign n33956 = n25658 ^ n21051 ^ n15600 ;
  assign n33958 = n8613 & n26450 ;
  assign n33957 = n4698 & n33442 ;
  assign n33959 = n33958 ^ n33957 ^ 1'b0 ;
  assign n33960 = n488 & ~n21753 ;
  assign n33961 = n33960 ^ n13027 ^ 1'b0 ;
  assign n33962 = n11288 | n16538 ;
  assign n33963 = n18365 | n33944 ;
  assign n33964 = n24716 & ~n33963 ;
  assign n33965 = n3170 ^ n1122 ^ 1'b0 ;
  assign n33966 = n3320 & n33965 ;
  assign n33967 = ( n22324 & n29527 ) | ( n22324 & n33966 ) | ( n29527 & n33966 ) ;
  assign n33968 = ( ~n2220 & n7771 ) | ( ~n2220 & n33967 ) | ( n7771 & n33967 ) ;
  assign n33972 = ( n4748 & n9240 ) | ( n4748 & n29738 ) | ( n9240 & n29738 ) ;
  assign n33973 = ( n11434 & n11863 ) | ( n11434 & n33972 ) | ( n11863 & n33972 ) ;
  assign n33969 = ~n8263 & n20617 ;
  assign n33970 = ~n5679 & n33969 ;
  assign n33971 = ( n21087 & n24434 ) | ( n21087 & n33970 ) | ( n24434 & n33970 ) ;
  assign n33974 = n33973 ^ n33971 ^ n29589 ;
  assign n33975 = n6323 | n10247 ;
  assign n33976 = n33975 ^ n32496 ^ n15291 ;
  assign n33977 = n29939 ^ n20256 ^ 1'b0 ;
  assign n33978 = n29173 ^ n19920 ^ 1'b0 ;
  assign n33979 = ~n15985 & n33978 ;
  assign n33980 = n20355 ^ n16154 ^ 1'b0 ;
  assign n33981 = n4671 ^ n3905 ^ 1'b0 ;
  assign n33982 = n12035 ^ n8600 ^ 1'b0 ;
  assign n33983 = n8389 & n33982 ;
  assign n33984 = n14321 ^ n2633 ^ 1'b0 ;
  assign n33985 = x202 & ~n33984 ;
  assign n33986 = n3177 | n12779 ;
  assign n33987 = n33985 | n33986 ;
  assign n33988 = ~n885 & n1384 ;
  assign n33989 = n1229 & ~n33988 ;
  assign n33990 = n1052 & n20294 ;
  assign n33991 = ~n33989 & n33990 ;
  assign n33992 = n4871 & ~n12750 ;
  assign n33993 = n23498 | n33992 ;
  assign n33994 = n8043 | n33993 ;
  assign n33996 = n17571 ^ n13023 ^ 1'b0 ;
  assign n33997 = ~n26122 & n33996 ;
  assign n33995 = n23279 ^ n15330 ^ n4555 ;
  assign n33998 = n33997 ^ n33995 ^ 1'b0 ;
  assign n33999 = ( n12222 & n33994 ) | ( n12222 & ~n33998 ) | ( n33994 & ~n33998 ) ;
  assign n34000 = n18587 ^ n17683 ^ 1'b0 ;
  assign n34001 = n4065 & ~n34000 ;
  assign n34002 = ~n16049 & n34001 ;
  assign n34003 = n34002 ^ n29672 ^ n11987 ;
  assign n34004 = n21671 ^ n18173 ^ n17196 ;
  assign n34007 = ( x121 & ~n14936 ) | ( x121 & n14945 ) | ( ~n14936 & n14945 ) ;
  assign n34005 = n18688 ^ n7203 ^ n7163 ;
  assign n34006 = n2515 & ~n34005 ;
  assign n34008 = n34007 ^ n34006 ^ n1171 ;
  assign n34009 = n19291 ^ n1236 ^ 1'b0 ;
  assign n34010 = n26813 | n34009 ;
  assign n34011 = n25481 | n34010 ;
  assign n34012 = n6712 & ~n34011 ;
  assign n34014 = ( ~n4095 & n27130 ) | ( ~n4095 & n32611 ) | ( n27130 & n32611 ) ;
  assign n34013 = n5357 & ~n23967 ;
  assign n34015 = n34014 ^ n34013 ^ n6219 ;
  assign n34016 = n7703 | n32712 ;
  assign n34017 = n3986 & ~n4288 ;
  assign n34018 = ~n8992 & n34017 ;
  assign n34019 = n34018 ^ n16530 ^ n9275 ;
  assign n34020 = n16252 | n34019 ;
  assign n34023 = ( n7017 & ~n9809 ) | ( n7017 & n14026 ) | ( ~n9809 & n14026 ) ;
  assign n34022 = ( n9892 & n16438 ) | ( n9892 & ~n16755 ) | ( n16438 & ~n16755 ) ;
  assign n34021 = n25589 ^ n19314 ^ n7228 ;
  assign n34024 = n34023 ^ n34022 ^ n34021 ;
  assign n34025 = ( n7787 & n9161 ) | ( n7787 & ~n25167 ) | ( n9161 & ~n25167 ) ;
  assign n34026 = n17209 & ~n25242 ;
  assign n34027 = n34026 ^ n22519 ^ 1'b0 ;
  assign n34028 = n10724 | n34027 ;
  assign n34029 = ( ~n12703 & n23170 ) | ( ~n12703 & n34028 ) | ( n23170 & n34028 ) ;
  assign n34030 = n17212 & n34029 ;
  assign n34031 = ~n11549 & n34030 ;
  assign n34032 = ( n12101 & n34025 ) | ( n12101 & ~n34031 ) | ( n34025 & ~n34031 ) ;
  assign n34033 = ( n4498 & n17667 ) | ( n4498 & n23906 ) | ( n17667 & n23906 ) ;
  assign n34034 = n5474 & n26248 ;
  assign n34035 = n34033 & n34034 ;
  assign n34036 = n3861 | n8886 ;
  assign n34037 = n22013 & ~n34036 ;
  assign n34038 = n903 & ~n34037 ;
  assign n34039 = n21122 & n34038 ;
  assign n34040 = n18457 ^ n12941 ^ n2178 ;
  assign n34041 = n34040 ^ n17962 ^ n12946 ;
  assign n34042 = n3641 & n34041 ;
  assign n34043 = n19078 ^ n17533 ^ 1'b0 ;
  assign n34044 = n13319 & n34043 ;
  assign n34045 = n28777 ^ n12621 ^ 1'b0 ;
  assign n34046 = ( ~n8304 & n29494 ) | ( ~n8304 & n29833 ) | ( n29494 & n29833 ) ;
  assign n34047 = n9048 ^ x161 ^ 1'b0 ;
  assign n34048 = n22629 & ~n34047 ;
  assign n34049 = n34048 ^ n3273 ^ 1'b0 ;
  assign n34050 = n3870 & ~n8440 ;
  assign n34051 = n5656 & n34050 ;
  assign n34052 = n34051 ^ n13870 ^ n11707 ;
  assign n34053 = n27817 ^ n3070 ^ 1'b0 ;
  assign n34054 = n11053 & n34053 ;
  assign n34055 = n16716 & ~n33417 ;
  assign n34056 = n3652 & n4450 ;
  assign n34057 = ~n2450 & n34056 ;
  assign n34058 = n31195 | n33801 ;
  assign n34059 = n7324 | n34058 ;
  assign n34060 = n30927 & n34059 ;
  assign n34061 = n12614 ^ n11768 ^ 1'b0 ;
  assign n34062 = ( n5322 & n6017 ) | ( n5322 & n30559 ) | ( n6017 & n30559 ) ;
  assign n34063 = ~n4177 & n25345 ;
  assign n34064 = ( ~n457 & n2363 ) | ( ~n457 & n16449 ) | ( n2363 & n16449 ) ;
  assign n34065 = n34064 ^ n24201 ^ n1346 ;
  assign n34066 = ( n7285 & n17977 ) | ( n7285 & n34065 ) | ( n17977 & n34065 ) ;
  assign n34067 = ~n6506 & n28861 ;
  assign n34068 = n34067 ^ n15448 ^ 1'b0 ;
  assign n34069 = ( ~n5268 & n15621 ) | ( ~n5268 & n30791 ) | ( n15621 & n30791 ) ;
  assign n34070 = n16854 ^ n905 ^ 1'b0 ;
  assign n34071 = n34070 ^ n13183 ^ x73 ;
  assign n34072 = n34071 ^ n13713 ^ 1'b0 ;
  assign n34073 = n34069 & n34072 ;
  assign n34074 = ( x67 & n1162 ) | ( x67 & ~n19699 ) | ( n1162 & ~n19699 ) ;
  assign n34075 = n32061 & ~n34074 ;
  assign n34081 = ( ~n7904 & n11066 ) | ( ~n7904 & n12077 ) | ( n11066 & n12077 ) ;
  assign n34080 = ~n284 & n7702 ;
  assign n34076 = n7392 | n8453 ;
  assign n34077 = n34076 ^ n9463 ^ 1'b0 ;
  assign n34078 = ( n9025 & n9250 ) | ( n9025 & n34077 ) | ( n9250 & n34077 ) ;
  assign n34079 = ( ~n7331 & n32068 ) | ( ~n7331 & n34078 ) | ( n32068 & n34078 ) ;
  assign n34082 = n34081 ^ n34080 ^ n34079 ;
  assign n34083 = n23456 & n24129 ;
  assign n34084 = n5589 | n7228 ;
  assign n34085 = n8660 & ~n34084 ;
  assign n34086 = ( n11650 & n12237 ) | ( n11650 & n24469 ) | ( n12237 & n24469 ) ;
  assign n34087 = ~n34085 & n34086 ;
  assign n34088 = n15827 & n34087 ;
  assign n34089 = n34088 ^ n12953 ^ 1'b0 ;
  assign n34090 = ~n30758 & n34089 ;
  assign n34091 = n10780 ^ n4044 ^ 1'b0 ;
  assign n34092 = ~n2596 & n5823 ;
  assign n34093 = n23686 & n34092 ;
  assign n34094 = ~n5840 & n31099 ;
  assign n34095 = n9352 ^ n8506 ^ 1'b0 ;
  assign n34096 = n29237 & ~n34095 ;
  assign n34097 = n34094 & n34096 ;
  assign n34098 = ( n34091 & n34093 ) | ( n34091 & ~n34097 ) | ( n34093 & ~n34097 ) ;
  assign n34099 = ~n1276 & n20271 ;
  assign n34100 = ( n14496 & n17392 ) | ( n14496 & ~n33328 ) | ( n17392 & ~n33328 ) ;
  assign n34101 = ( ~n5091 & n9903 ) | ( ~n5091 & n17058 ) | ( n9903 & n17058 ) ;
  assign n34102 = n34101 ^ n1346 ^ 1'b0 ;
  assign n34103 = n15533 | n25605 ;
  assign n34104 = n34103 ^ n13770 ^ 1'b0 ;
  assign n34105 = n9488 & n29792 ;
  assign n34106 = n3515 & n34105 ;
  assign n34107 = n34106 ^ n1845 ^ 1'b0 ;
  assign n34108 = n6996 ^ n1645 ^ 1'b0 ;
  assign n34109 = n34108 ^ n9976 ^ 1'b0 ;
  assign n34110 = ~n3521 & n34109 ;
  assign n34111 = n11147 | n20551 ;
  assign n34112 = n34111 ^ n20475 ^ n11401 ;
  assign n34113 = ( n2689 & n31276 ) | ( n2689 & n34112 ) | ( n31276 & n34112 ) ;
  assign n34117 = ~n4537 & n15029 ;
  assign n34118 = n3960 & n34117 ;
  assign n34114 = n13028 ^ n10990 ^ 1'b0 ;
  assign n34115 = n11461 & ~n34114 ;
  assign n34116 = n15199 & n34115 ;
  assign n34119 = n34118 ^ n34116 ^ n9096 ;
  assign n34120 = n5235 | n30915 ;
  assign n34121 = ( ~n6990 & n16356 ) | ( ~n6990 & n19255 ) | ( n16356 & n19255 ) ;
  assign n34122 = n34121 ^ n14584 ^ 1'b0 ;
  assign n34123 = n19199 ^ n724 ^ 1'b0 ;
  assign n34124 = n4983 | n12524 ;
  assign n34125 = n32727 | n34124 ;
  assign n34126 = ~n5217 & n34125 ;
  assign n34127 = ~n12351 & n34126 ;
  assign n34133 = ( x35 & n18783 ) | ( x35 & ~n20831 ) | ( n18783 & ~n20831 ) ;
  assign n34128 = ~n751 & n5775 ;
  assign n34129 = n34128 ^ n2529 ^ 1'b0 ;
  assign n34130 = n20236 & ~n34129 ;
  assign n34131 = ~n5457 & n34130 ;
  assign n34132 = ~n13480 & n34131 ;
  assign n34134 = n34133 ^ n34132 ^ 1'b0 ;
  assign n34135 = n2688 & n16789 ;
  assign n34136 = n9628 | n34135 ;
  assign n34137 = n6476 ^ n1750 ^ 1'b0 ;
  assign n34138 = ( n5599 & n12708 ) | ( n5599 & ~n34137 ) | ( n12708 & ~n34137 ) ;
  assign n34139 = n8608 & ~n14808 ;
  assign n34140 = ( n14080 & ~n30543 ) | ( n14080 & n34139 ) | ( ~n30543 & n34139 ) ;
  assign n34141 = n30253 ^ n13720 ^ 1'b0 ;
  assign n34142 = n20168 ^ n19297 ^ 1'b0 ;
  assign n34143 = ( ~n4229 & n5133 ) | ( ~n4229 & n28164 ) | ( n5133 & n28164 ) ;
  assign n34144 = ( n17442 & ~n31014 ) | ( n17442 & n34143 ) | ( ~n31014 & n34143 ) ;
  assign n34145 = ~n2070 & n3964 ;
  assign n34146 = n34145 ^ n6949 ^ n6320 ;
  assign n34147 = ~n993 & n34146 ;
  assign n34148 = n28458 & n34147 ;
  assign n34149 = ( n8697 & ~n10233 ) | ( n8697 & n11342 ) | ( ~n10233 & n11342 ) ;
  assign n34150 = ~n11553 & n26621 ;
  assign n34151 = ~n34149 & n34150 ;
  assign n34152 = ~n4125 & n28426 ;
  assign n34153 = ( n2970 & n31832 ) | ( n2970 & ~n34071 ) | ( n31832 & ~n34071 ) ;
  assign n34154 = n16483 ^ n4045 ^ 1'b0 ;
  assign n34155 = n34153 | n34154 ;
  assign n34156 = n34155 ^ n13601 ^ 1'b0 ;
  assign n34157 = n28179 ^ n11795 ^ 1'b0 ;
  assign n34158 = n33578 ^ n29324 ^ n14047 ;
  assign n34159 = n25572 & ~n31665 ;
  assign n34161 = n18852 ^ n5784 ^ n2234 ;
  assign n34160 = n14892 | n23484 ;
  assign n34162 = n34161 ^ n34160 ^ 1'b0 ;
  assign n34163 = n34162 ^ n3031 ^ 1'b0 ;
  assign n34165 = ( n2159 & n2195 ) | ( n2159 & n11296 ) | ( n2195 & n11296 ) ;
  assign n34166 = ~n443 & n34165 ;
  assign n34167 = n34166 ^ n3063 ^ 1'b0 ;
  assign n34164 = n26119 ^ n25566 ^ n4165 ;
  assign n34168 = n34167 ^ n34164 ^ 1'b0 ;
  assign n34169 = n19296 | n34168 ;
  assign n34170 = n34169 ^ n18509 ^ 1'b0 ;
  assign n34171 = n31010 ^ n17444 ^ 1'b0 ;
  assign n34172 = n8792 | n10480 ;
  assign n34173 = n3852 | n21059 ;
  assign n34174 = ~n1057 & n19790 ;
  assign n34175 = n12950 ^ n12428 ^ n12417 ;
  assign n34176 = n34175 ^ n7490 ^ 1'b0 ;
  assign n34179 = n7487 | n16994 ;
  assign n34180 = n25249 | n34179 ;
  assign n34177 = n11834 ^ n6596 ^ 1'b0 ;
  assign n34178 = x73 & ~n34177 ;
  assign n34181 = n34180 ^ n34178 ^ n16673 ;
  assign n34182 = n22980 & ~n31539 ;
  assign n34183 = n34182 ^ n16630 ^ n15690 ;
  assign n34184 = ( n34176 & n34181 ) | ( n34176 & n34183 ) | ( n34181 & n34183 ) ;
  assign n34185 = n15835 ^ n4618 ^ 1'b0 ;
  assign n34186 = n7191 & n34185 ;
  assign n34187 = n23619 ^ n18780 ^ 1'b0 ;
  assign n34188 = n34187 ^ n25473 ^ 1'b0 ;
  assign n34192 = ( n12899 & n23564 ) | ( n12899 & ~n25617 ) | ( n23564 & ~n25617 ) ;
  assign n34189 = n6530 & ~n9535 ;
  assign n34190 = n34189 ^ n1068 ^ 1'b0 ;
  assign n34191 = ~n16470 & n34190 ;
  assign n34193 = n34192 ^ n34191 ^ 1'b0 ;
  assign n34194 = ~n10386 & n34193 ;
  assign n34195 = ~n11257 & n34194 ;
  assign n34196 = n27910 ^ n6344 ^ n2022 ;
  assign n34200 = n15290 | n23454 ;
  assign n34201 = n27982 | n34200 ;
  assign n34199 = n23319 & n26435 ;
  assign n34197 = n1496 & n15800 ;
  assign n34198 = n8926 & ~n34197 ;
  assign n34202 = n34201 ^ n34199 ^ n34198 ;
  assign n34203 = n17952 | n34104 ;
  assign n34204 = n21011 ^ n10457 ^ 1'b0 ;
  assign n34207 = ( n1852 & n2490 ) | ( n1852 & ~n11566 ) | ( n2490 & ~n11566 ) ;
  assign n34205 = n3607 ^ n2887 ^ 1'b0 ;
  assign n34206 = n24342 | n34205 ;
  assign n34208 = n34207 ^ n34206 ^ n15020 ;
  assign n34209 = x28 & ~n2494 ;
  assign n34210 = n34209 ^ n10934 ^ 1'b0 ;
  assign n34211 = n17132 | n34210 ;
  assign n34212 = n5281 ^ n3066 ^ 1'b0 ;
  assign n34213 = n19283 ^ n10514 ^ n7125 ;
  assign n34214 = n16530 & ~n29533 ;
  assign n34215 = ( n4741 & ~n34213 ) | ( n4741 & n34214 ) | ( ~n34213 & n34214 ) ;
  assign n34216 = n3298 & ~n26706 ;
  assign n34217 = n17465 ^ n7119 ^ 1'b0 ;
  assign n34218 = n15509 | n34217 ;
  assign n34219 = ( n14131 & ~n28113 ) | ( n14131 & n34218 ) | ( ~n28113 & n34218 ) ;
  assign n34221 = n4409 | n6073 ;
  assign n34222 = n3312 & ~n34221 ;
  assign n34223 = n34222 ^ n4983 ^ n3004 ;
  assign n34220 = n3433 ^ n1778 ^ 1'b0 ;
  assign n34224 = n34223 ^ n34220 ^ n2490 ;
  assign n34225 = n26004 & ~n34224 ;
  assign n34226 = n34219 & n34225 ;
  assign n34227 = n14230 | n34226 ;
  assign n34228 = n34216 & ~n34227 ;
  assign n34229 = n12748 ^ n2411 ^ 1'b0 ;
  assign n34230 = ( n13918 & n30278 ) | ( n13918 & n34229 ) | ( n30278 & n34229 ) ;
  assign n34231 = n3530 ^ n3120 ^ n1345 ;
  assign n34237 = x130 & n1250 ;
  assign n34238 = ~n1250 & n34237 ;
  assign n34239 = n34238 ^ n30166 ^ 1'b0 ;
  assign n34232 = ~n1726 & n5486 ;
  assign n34233 = n1726 & n34232 ;
  assign n34234 = n34233 ^ n12504 ^ 1'b0 ;
  assign n34235 = n10369 & ~n34234 ;
  assign n34236 = n34234 & n34235 ;
  assign n34240 = n34239 ^ n34236 ^ n496 ;
  assign n34241 = ( ~n9047 & n16722 ) | ( ~n9047 & n34240 ) | ( n16722 & n34240 ) ;
  assign n34242 = n25073 ^ n4093 ^ 1'b0 ;
  assign n34243 = n15430 | n34242 ;
  assign n34244 = n23230 & ~n34243 ;
  assign n34245 = n34241 & n34244 ;
  assign n34246 = n16650 ^ n2184 ^ 1'b0 ;
  assign n34247 = ~n34245 & n34246 ;
  assign n34248 = ( ~n1344 & n34231 ) | ( ~n1344 & n34247 ) | ( n34231 & n34247 ) ;
  assign n34249 = ~n843 & n20609 ;
  assign n34250 = n34249 ^ n1705 ^ 1'b0 ;
  assign n34251 = n3195 & n9491 ;
  assign n34252 = ( n26941 & n34250 ) | ( n26941 & n34251 ) | ( n34250 & n34251 ) ;
  assign n34253 = n30930 ^ n1475 ^ 1'b0 ;
  assign n34254 = n10386 & ~n34253 ;
  assign n34255 = n22483 & n34254 ;
  assign n34257 = n13075 ^ n5132 ^ 1'b0 ;
  assign n34256 = n3713 & ~n5974 ;
  assign n34258 = n34257 ^ n34256 ^ 1'b0 ;
  assign n34259 = n3996 | n5755 ;
  assign n34260 = n34259 ^ n8361 ^ 1'b0 ;
  assign n34261 = n34260 ^ n33490 ^ 1'b0 ;
  assign n34262 = n4067 & n30579 ;
  assign n34263 = n34262 ^ n4364 ^ 1'b0 ;
  assign n34264 = ( n1236 & n9082 ) | ( n1236 & ~n33831 ) | ( n9082 & ~n33831 ) ;
  assign n34265 = ( x218 & ~x242 ) | ( x218 & n6297 ) | ( ~x242 & n6297 ) ;
  assign n34266 = n1591 & ~n14188 ;
  assign n34267 = n34265 & n34266 ;
  assign n34269 = n8515 ^ n6044 ^ 1'b0 ;
  assign n34268 = n3581 & n25174 ;
  assign n34270 = n34269 ^ n34268 ^ 1'b0 ;
  assign n34271 = n12784 ^ n11559 ^ 1'b0 ;
  assign n34272 = n10913 | n34271 ;
  assign n34273 = n11809 & ~n34272 ;
  assign n34274 = n5981 & n34273 ;
  assign n34276 = n7165 ^ n989 ^ 1'b0 ;
  assign n34277 = n34276 ^ n20640 ^ 1'b0 ;
  assign n34278 = n16131 & n34277 ;
  assign n34275 = n16771 & ~n24012 ;
  assign n34279 = n34278 ^ n34275 ^ 1'b0 ;
  assign n34280 = ~n16806 & n19251 ;
  assign n34281 = n22560 ^ n14937 ^ n12925 ;
  assign n34282 = n5250 | n17719 ;
  assign n34283 = ( n3542 & n7668 ) | ( n3542 & n34282 ) | ( n7668 & n34282 ) ;
  assign n34284 = n34283 ^ n16608 ^ x210 ;
  assign n34285 = n14686 ^ n8918 ^ n1366 ;
  assign n34286 = n34285 ^ n27857 ^ 1'b0 ;
  assign n34290 = n8066 & n29129 ;
  assign n34291 = n9944 & n34290 ;
  assign n34292 = n7926 & ~n34291 ;
  assign n34293 = n10263 & ~n14218 ;
  assign n34294 = n34292 & n34293 ;
  assign n34287 = n825 | n28727 ;
  assign n34288 = n34287 ^ n10050 ^ 1'b0 ;
  assign n34289 = ( n1748 & n32078 ) | ( n1748 & ~n34288 ) | ( n32078 & ~n34288 ) ;
  assign n34295 = n34294 ^ n34289 ^ n9745 ;
  assign n34296 = n3994 & n22956 ;
  assign n34297 = ~n34295 & n34296 ;
  assign n34298 = n31682 ^ n2114 ^ 1'b0 ;
  assign n34299 = n3172 ^ n1632 ^ 1'b0 ;
  assign n34300 = n6575 ^ n6103 ^ 1'b0 ;
  assign n34301 = n13418 | n34300 ;
  assign n34302 = n26472 ^ n12069 ^ x88 ;
  assign n34303 = ( n434 & n34301 ) | ( n434 & n34302 ) | ( n34301 & n34302 ) ;
  assign n34308 = n15798 ^ n12005 ^ 1'b0 ;
  assign n34309 = ~n1020 & n34308 ;
  assign n34306 = ( n857 & ~n13622 ) | ( n857 & n16928 ) | ( ~n13622 & n16928 ) ;
  assign n34304 = n28756 ^ n9016 ^ 1'b0 ;
  assign n34305 = n23904 | n34304 ;
  assign n34307 = n34306 ^ n34305 ^ n1090 ;
  assign n34310 = n34309 ^ n34307 ^ n11048 ;
  assign n34311 = n12573 ^ n12465 ^ 1'b0 ;
  assign n34312 = n19718 ^ n17662 ^ 1'b0 ;
  assign n34313 = n7491 | n8352 ;
  assign n34314 = n441 & ~n34313 ;
  assign n34315 = ~n15041 & n20015 ;
  assign n34316 = n30815 & n34315 ;
  assign n34317 = ( n18261 & ~n34314 ) | ( n18261 & n34316 ) | ( ~n34314 & n34316 ) ;
  assign n34318 = n7173 ^ n6486 ^ 1'b0 ;
  assign n34319 = ( n10422 & ~n11821 ) | ( n10422 & n34318 ) | ( ~n11821 & n34318 ) ;
  assign n34320 = n6793 ^ n6270 ^ n2766 ;
  assign n34321 = n34320 ^ n6548 ^ 1'b0 ;
  assign n34322 = n14255 & ~n34321 ;
  assign n34323 = n1455 & n34322 ;
  assign n34324 = n28467 ^ n13761 ^ n1028 ;
  assign n34325 = ~n11249 & n34324 ;
  assign n34326 = n34325 ^ n6372 ^ 1'b0 ;
  assign n34327 = n17734 ^ n9825 ^ 1'b0 ;
  assign n34328 = n34327 ^ n6070 ^ 1'b0 ;
  assign n34329 = n6188 ^ n2191 ^ n2024 ;
  assign n34330 = n34329 ^ n28929 ^ 1'b0 ;
  assign n34332 = n2276 & n3422 ;
  assign n34333 = n34332 ^ n2746 ^ 1'b0 ;
  assign n34331 = ~n3669 & n10872 ;
  assign n34334 = n34333 ^ n34331 ^ 1'b0 ;
  assign n34335 = n34334 ^ n4429 ^ 1'b0 ;
  assign n34336 = n10233 & n34335 ;
  assign n34337 = n31434 ^ n16979 ^ n11599 ;
  assign n34338 = n6843 & n14086 ;
  assign n34339 = n16554 & n34338 ;
  assign n34340 = ~n1186 & n8070 ;
  assign n34341 = n34339 & n34340 ;
  assign n34342 = n3309 | n34341 ;
  assign n34343 = ( n1205 & ~n9965 ) | ( n1205 & n34342 ) | ( ~n9965 & n34342 ) ;
  assign n34344 = n25070 | n34343 ;
  assign n34345 = n27208 ^ n9851 ^ n5357 ;
  assign n34346 = n9851 & n14611 ;
  assign n34347 = n34346 ^ n9512 ^ 1'b0 ;
  assign n34350 = n16777 ^ n4323 ^ 1'b0 ;
  assign n34351 = n34350 ^ n24448 ^ n19820 ;
  assign n34348 = n14114 ^ n8813 ^ n6277 ;
  assign n34349 = n34348 ^ n4436 ^ n1209 ;
  assign n34352 = n34351 ^ n34349 ^ n14155 ;
  assign n34353 = n32918 ^ n8368 ^ 1'b0 ;
  assign n34359 = n19278 ^ n483 ^ 1'b0 ;
  assign n34354 = ~n2157 & n11438 ;
  assign n34355 = n34354 ^ n355 ^ 1'b0 ;
  assign n34356 = n34355 ^ n7810 ^ n2766 ;
  assign n34357 = n19769 & ~n26034 ;
  assign n34358 = n34356 & n34357 ;
  assign n34360 = n34359 ^ n34358 ^ n21743 ;
  assign n34361 = ( n8625 & n14312 ) | ( n8625 & ~n20617 ) | ( n14312 & ~n20617 ) ;
  assign n34362 = n34361 ^ n13942 ^ n9585 ;
  assign n34363 = n27051 ^ n8409 ^ 1'b0 ;
  assign n34364 = n21888 & n34363 ;
  assign n34365 = n9364 & ~n10290 ;
  assign n34366 = ( n14269 & n18285 ) | ( n14269 & ~n34365 ) | ( n18285 & ~n34365 ) ;
  assign n34367 = ( n34362 & n34364 ) | ( n34362 & ~n34366 ) | ( n34364 & ~n34366 ) ;
  assign n34368 = ~n24865 & n34367 ;
  assign n34369 = n4653 & ~n23588 ;
  assign n34370 = n29858 ^ n7884 ^ n1769 ;
  assign n34371 = ~n27481 & n34370 ;
  assign n34372 = ~n32274 & n34371 ;
  assign n34373 = n21350 ^ n2834 ^ 1'b0 ;
  assign n34374 = ~n34372 & n34373 ;
  assign n34375 = n33724 ^ n30998 ^ 1'b0 ;
  assign n34376 = n812 & n29358 ;
  assign n34377 = n34376 ^ n33792 ^ x120 ;
  assign n34378 = ( x250 & n16454 ) | ( x250 & ~n32467 ) | ( n16454 & ~n32467 ) ;
  assign n34379 = n3659 & n15156 ;
  assign n34380 = n34379 ^ n6629 ^ 1'b0 ;
  assign n34381 = n34380 ^ n10738 ^ 1'b0 ;
  assign n34382 = x170 & n34381 ;
  assign n34383 = ~n24594 & n34382 ;
  assign n34384 = n22264 | n27222 ;
  assign n34385 = n3512 & ~n34384 ;
  assign n34386 = n17474 | n32494 ;
  assign n34387 = n29840 & ~n34386 ;
  assign n34388 = n26939 ^ n5678 ^ 1'b0 ;
  assign n34392 = n5065 | n19414 ;
  assign n34389 = n2663 & ~n28187 ;
  assign n34390 = n34389 ^ n14210 ^ 1'b0 ;
  assign n34391 = n18359 & ~n34390 ;
  assign n34393 = n34392 ^ n34391 ^ n11545 ;
  assign n34395 = ( ~n1504 & n15307 ) | ( ~n1504 & n21629 ) | ( n15307 & n21629 ) ;
  assign n34396 = n6586 & n34395 ;
  assign n34397 = n34396 ^ n2778 ^ 1'b0 ;
  assign n34394 = n27094 ^ n23327 ^ 1'b0 ;
  assign n34398 = n34397 ^ n34394 ^ n1508 ;
  assign n34399 = ( ~n4462 & n29070 ) | ( ~n4462 & n34398 ) | ( n29070 & n34398 ) ;
  assign n34400 = n22042 ^ n11401 ^ 1'b0 ;
  assign n34401 = ( n27996 & ~n28384 ) | ( n27996 & n34400 ) | ( ~n28384 & n34400 ) ;
  assign n34402 = n8038 & ~n8533 ;
  assign n34403 = n12199 & ~n34402 ;
  assign n34404 = n10630 ^ n5057 ^ 1'b0 ;
  assign n34405 = n18443 | n34404 ;
  assign n34406 = n12083 ^ x10 ^ 1'b0 ;
  assign n34408 = n15080 ^ n14385 ^ 1'b0 ;
  assign n34409 = n25695 & n34408 ;
  assign n34407 = n12866 & ~n20836 ;
  assign n34410 = n34409 ^ n34407 ^ 1'b0 ;
  assign n34411 = ( n6077 & n34406 ) | ( n6077 & ~n34410 ) | ( n34406 & ~n34410 ) ;
  assign n34412 = n33454 ^ n13684 ^ 1'b0 ;
  assign n34413 = n34412 ^ n12032 ^ n10603 ;
  assign n34414 = n34413 ^ n3553 ^ 1'b0 ;
  assign n34415 = n19687 & n31588 ;
  assign n34416 = ~n4132 & n29013 ;
  assign n34417 = n34416 ^ n24441 ^ 1'b0 ;
  assign n34418 = n30137 ^ n6224 ^ 1'b0 ;
  assign n34419 = n3917 & ~n17710 ;
  assign n34420 = n34419 ^ n24109 ^ 1'b0 ;
  assign n34421 = ( ~x92 & n952 ) | ( ~x92 & n23103 ) | ( n952 & n23103 ) ;
  assign n34422 = n32694 ^ n14345 ^ x83 ;
  assign n34423 = n492 & ~n34422 ;
  assign n34424 = ~n16201 & n34423 ;
  assign n34425 = n34421 | n34424 ;
  assign n34426 = n1512 & n18741 ;
  assign n34427 = n34425 & n34426 ;
  assign n34428 = ~n6073 & n6745 ;
  assign n34429 = n5360 & n34428 ;
  assign n34430 = n32160 ^ n17987 ^ n11669 ;
  assign n34431 = n30143 ^ n1623 ^ 1'b0 ;
  assign n34432 = n8154 & n34431 ;
  assign n34433 = n4653 ^ n287 ^ 1'b0 ;
  assign n34434 = n6595 & ~n34433 ;
  assign n34435 = n11196 | n34434 ;
  assign n34436 = n4506 ^ n2896 ^ 1'b0 ;
  assign n34437 = n13105 & ~n34436 ;
  assign n34438 = n34437 ^ n2638 ^ 1'b0 ;
  assign n34439 = ~n34435 & n34438 ;
  assign n34440 = n34439 ^ n5974 ^ 1'b0 ;
  assign n34441 = ( n30998 & n34432 ) | ( n30998 & ~n34440 ) | ( n34432 & ~n34440 ) ;
  assign n34445 = ~n6675 & n11565 ;
  assign n34446 = n7937 & n34445 ;
  assign n34447 = n34446 ^ n17119 ^ 1'b0 ;
  assign n34448 = n24560 & ~n34447 ;
  assign n34442 = n7927 & ~n30287 ;
  assign n34443 = n34442 ^ n31254 ^ 1'b0 ;
  assign n34444 = n15038 | n34443 ;
  assign n34449 = n34448 ^ n34444 ^ 1'b0 ;
  assign n34450 = n19144 & n32121 ;
  assign n34451 = n4620 & ~n29304 ;
  assign n34452 = ~n7017 & n34451 ;
  assign n34453 = ( n6028 & n14802 ) | ( n6028 & n16345 ) | ( n14802 & n16345 ) ;
  assign n34454 = ( ~n15965 & n34452 ) | ( ~n15965 & n34453 ) | ( n34452 & n34453 ) ;
  assign n34455 = n7738 & n14584 ;
  assign n34456 = n9365 & n34455 ;
  assign n34457 = ( n3952 & ~n26610 ) | ( n3952 & n34456 ) | ( ~n26610 & n34456 ) ;
  assign n34458 = n15598 & ~n34457 ;
  assign n34459 = n26736 & n34458 ;
  assign n34460 = n7482 ^ n2461 ^ 1'b0 ;
  assign n34464 = n2051 | n2290 ;
  assign n34465 = n10342 & ~n34464 ;
  assign n34461 = ~n24941 & n33137 ;
  assign n34462 = n34461 ^ n11035 ^ 1'b0 ;
  assign n34463 = n23074 & n34462 ;
  assign n34466 = n34465 ^ n34463 ^ 1'b0 ;
  assign n34467 = ( n9601 & n24408 ) | ( n9601 & n24497 ) | ( n24408 & n24497 ) ;
  assign n34468 = n2184 & n21660 ;
  assign n34469 = n34467 & n34468 ;
  assign n34470 = n33629 & n34469 ;
  assign n34471 = n18481 ^ n12283 ^ 1'b0 ;
  assign n34472 = ~n22518 & n34471 ;
  assign n34473 = n31085 ^ n10156 ^ 1'b0 ;
  assign n34474 = n19525 & ~n34473 ;
  assign n34475 = n8716 ^ n3534 ^ 1'b0 ;
  assign n34476 = ~n34474 & n34475 ;
  assign n34477 = ~n28264 & n34476 ;
  assign n34478 = n9327 | n34477 ;
  assign n34479 = n4124 | n34478 ;
  assign n34480 = n724 | n3817 ;
  assign n34481 = n34480 ^ n10712 ^ n6941 ;
  assign n34482 = ~n6478 & n15632 ;
  assign n34485 = n3860 | n14573 ;
  assign n34483 = n10275 ^ n5635 ^ n2254 ;
  assign n34484 = ~n25968 & n34483 ;
  assign n34486 = n34485 ^ n34484 ^ n8747 ;
  assign n34487 = ( n11923 & n31748 ) | ( n11923 & ~n34486 ) | ( n31748 & ~n34486 ) ;
  assign n34488 = n392 & n25615 ;
  assign n34489 = n34488 ^ n18337 ^ 1'b0 ;
  assign n34490 = x187 & n2968 ;
  assign n34491 = n23644 ^ n11327 ^ n3697 ;
  assign n34492 = n11912 & ~n34491 ;
  assign n34493 = n34490 & n34492 ;
  assign n34494 = n1357 | n15573 ;
  assign n34495 = n34493 & ~n34494 ;
  assign n34496 = n1258 | n3772 ;
  assign n34497 = n13007 | n34496 ;
  assign n34498 = n21179 & ~n27802 ;
  assign n34499 = n34498 ^ n15436 ^ 1'b0 ;
  assign n34500 = ~n22855 & n34499 ;
  assign n34501 = ( n6831 & n12266 ) | ( n6831 & n13420 ) | ( n12266 & n13420 ) ;
  assign n34502 = n18543 & ~n34501 ;
  assign n34503 = n1088 | n34502 ;
  assign n34504 = n17403 ^ n15653 ^ 1'b0 ;
  assign n34505 = n28775 & ~n34504 ;
  assign n34506 = n10307 ^ n9025 ^ 1'b0 ;
  assign n34507 = n24154 & ~n34506 ;
  assign n34510 = n10527 ^ n4958 ^ 1'b0 ;
  assign n34509 = n1314 | n3840 ;
  assign n34511 = n34510 ^ n34509 ^ 1'b0 ;
  assign n34508 = n3353 & n3541 ;
  assign n34512 = n34511 ^ n34508 ^ n21285 ;
  assign n34513 = n34512 ^ n6766 ^ n5729 ;
  assign n34514 = n18229 & n31879 ;
  assign n34515 = n9623 & ~n29840 ;
  assign n34516 = n34515 ^ n15264 ^ 1'b0 ;
  assign n34517 = n14991 ^ n1491 ^ 1'b0 ;
  assign n34518 = n34516 & ~n34517 ;
  assign n34519 = n21744 & n27253 ;
  assign n34520 = n4790 & ~n34519 ;
  assign n34521 = n20475 ^ n8188 ^ 1'b0 ;
  assign n34522 = n34521 ^ n27684 ^ n16496 ;
  assign n34523 = n23132 & n34522 ;
  assign n34524 = n13085 ^ n6878 ^ 1'b0 ;
  assign n34525 = n34524 ^ n20534 ^ n6220 ;
  assign n34526 = n21350 & ~n30381 ;
  assign n34527 = ( n14636 & ~n34525 ) | ( n14636 & n34526 ) | ( ~n34525 & n34526 ) ;
  assign n34532 = n11339 ^ n8052 ^ n5492 ;
  assign n34533 = n8455 ^ n2349 ^ 1'b0 ;
  assign n34534 = n6194 | n34533 ;
  assign n34535 = n34532 & ~n34534 ;
  assign n34529 = n17768 & ~n22167 ;
  assign n34530 = n16236 & n34529 ;
  assign n34528 = n4710 | n17319 ;
  assign n34531 = n34530 ^ n34528 ^ 1'b0 ;
  assign n34536 = n34535 ^ n34531 ^ 1'b0 ;
  assign n34537 = n17048 ^ n11122 ^ n1145 ;
  assign n34538 = n1385 & ~n4028 ;
  assign n34539 = n34537 & n34538 ;
  assign n34540 = n13422 | n20886 ;
  assign n34541 = n317 | n34540 ;
  assign n34542 = n5263 | n32438 ;
  assign n34543 = n766 | n34542 ;
  assign n34544 = n15340 ^ n6838 ^ 1'b0 ;
  assign n34545 = n34544 ^ n1133 ^ 1'b0 ;
  assign n34546 = ( n6809 & ~n15895 ) | ( n6809 & n29143 ) | ( ~n15895 & n29143 ) ;
  assign n34547 = n21053 ^ n11342 ^ 1'b0 ;
  assign n34548 = n21637 & ~n33844 ;
  assign n34549 = n15621 & ~n24519 ;
  assign n34550 = n34549 ^ n27202 ^ 1'b0 ;
  assign n34551 = n4318 & ~n18112 ;
  assign n34552 = ~n1408 & n34551 ;
  assign n34553 = n34552 ^ n23920 ^ 1'b0 ;
  assign n34554 = n34553 ^ n11433 ^ 1'b0 ;
  assign n34555 = n25609 & n34554 ;
  assign n34556 = n8701 ^ n1853 ^ 1'b0 ;
  assign n34557 = n34556 ^ n10195 ^ n4047 ;
  assign n34558 = ~n1616 & n34557 ;
  assign n34559 = n34558 ^ n5506 ^ 1'b0 ;
  assign n34560 = n14074 & n23536 ;
  assign n34561 = ( ~n15380 & n34559 ) | ( ~n15380 & n34560 ) | ( n34559 & n34560 ) ;
  assign n34562 = n4404 ^ n1468 ^ 1'b0 ;
  assign n34563 = n23551 ^ n9481 ^ n7753 ;
  assign n34564 = n8436 & n19429 ;
  assign n34565 = ~n29416 & n34564 ;
  assign n34566 = ~n2498 & n17057 ;
  assign n34567 = n6229 | n10406 ;
  assign n34568 = n17092 & ~n34567 ;
  assign n34569 = n34566 | n34568 ;
  assign n34570 = ~n12873 & n20831 ;
  assign n34571 = n13294 ^ n3887 ^ 1'b0 ;
  assign n34572 = ( n25114 & n26136 ) | ( n25114 & n34571 ) | ( n26136 & n34571 ) ;
  assign n34573 = n6275 & ~n12422 ;
  assign n34574 = ~n13164 & n33130 ;
  assign n34575 = ( n18040 & ~n21168 ) | ( n18040 & n34574 ) | ( ~n21168 & n34574 ) ;
  assign n34576 = n26199 & n34575 ;
  assign n34577 = n34576 ^ n26467 ^ 1'b0 ;
  assign n34578 = n3324 ^ n1554 ^ 1'b0 ;
  assign n34579 = n14443 | n34578 ;
  assign n34580 = ~n9302 & n34579 ;
  assign n34581 = ~n23267 & n34580 ;
  assign n34582 = n15333 & n33509 ;
  assign n34583 = n34582 ^ n11683 ^ 1'b0 ;
  assign n34584 = ( n1290 & n10714 ) | ( n1290 & n26772 ) | ( n10714 & n26772 ) ;
  assign n34585 = n34584 ^ n33588 ^ n19030 ;
  assign n34586 = ( ~n1099 & n2638 ) | ( ~n1099 & n4060 ) | ( n2638 & n4060 ) ;
  assign n34587 = ( ~n23563 & n32672 ) | ( ~n23563 & n34586 ) | ( n32672 & n34586 ) ;
  assign n34588 = n34587 ^ n20586 ^ n17000 ;
  assign n34589 = n14198 ^ n4429 ^ 1'b0 ;
  assign n34590 = n34589 ^ n21448 ^ 1'b0 ;
  assign n34591 = ~n18916 & n34590 ;
  assign n34592 = n14592 ^ n3858 ^ 1'b0 ;
  assign n34593 = n19336 & ~n34592 ;
  assign n34594 = n1497 & ~n3668 ;
  assign n34595 = n24853 & n34594 ;
  assign n34596 = n4540 & ~n34595 ;
  assign n34597 = n34596 ^ n28275 ^ 1'b0 ;
  assign n34598 = n7402 & n14551 ;
  assign n34599 = n34598 ^ n14617 ^ 1'b0 ;
  assign n34600 = n19009 & n31539 ;
  assign n34601 = n34600 ^ n17970 ^ 1'b0 ;
  assign n34602 = n34599 | n34601 ;
  assign n34603 = ~n12133 & n26089 ;
  assign n34604 = n6043 | n14569 ;
  assign n34605 = n34604 ^ n13899 ^ 1'b0 ;
  assign n34606 = n29514 & ~n34605 ;
  assign n34607 = ~n13932 & n20271 ;
  assign n34608 = n9592 & ~n12003 ;
  assign n34609 = n34608 ^ n1922 ^ 1'b0 ;
  assign n34610 = n11971 ^ n1388 ^ 1'b0 ;
  assign n34611 = n15869 | n34610 ;
  assign n34612 = n26817 | n34611 ;
  assign n34619 = n22847 ^ n15270 ^ n14038 ;
  assign n34620 = n34619 ^ n27130 ^ n13764 ;
  assign n34613 = n14277 ^ n757 ^ 1'b0 ;
  assign n34614 = n1336 & ~n34613 ;
  assign n34615 = ~n4053 & n34614 ;
  assign n34616 = n34615 ^ n7182 ^ 1'b0 ;
  assign n34617 = ~n18356 & n34616 ;
  assign n34618 = ~n13797 & n34617 ;
  assign n34621 = n34620 ^ n34618 ^ 1'b0 ;
  assign n34622 = n34612 & n34621 ;
  assign n34624 = ~n4882 & n10340 ;
  assign n34625 = n15221 & n24417 ;
  assign n34626 = n18394 ^ n9015 ^ 1'b0 ;
  assign n34627 = n4117 | n34626 ;
  assign n34628 = ( n34624 & n34625 ) | ( n34624 & n34627 ) | ( n34625 & n34627 ) ;
  assign n34623 = ~n19054 & n33685 ;
  assign n34629 = n34628 ^ n34623 ^ 1'b0 ;
  assign n34630 = n21688 ^ n17858 ^ 1'b0 ;
  assign n34631 = x143 & ~n34630 ;
  assign n34633 = n7878 ^ n5532 ^ n4819 ;
  assign n34634 = n34633 ^ n7399 ^ 1'b0 ;
  assign n34635 = n21589 | n34634 ;
  assign n34632 = n7626 & ~n13526 ;
  assign n34636 = n34635 ^ n34632 ^ 1'b0 ;
  assign n34637 = n21983 ^ n7966 ^ n420 ;
  assign n34638 = n34637 ^ n23922 ^ n7174 ;
  assign n34639 = n32089 ^ n7831 ^ 1'b0 ;
  assign n34642 = n12814 ^ n2746 ^ 1'b0 ;
  assign n34641 = ~n3341 & n7134 ;
  assign n34643 = n34642 ^ n34641 ^ 1'b0 ;
  assign n34640 = ~n13953 & n19133 ;
  assign n34644 = n34643 ^ n34640 ^ 1'b0 ;
  assign n34645 = n15513 ^ n10834 ^ n7215 ;
  assign n34646 = ( n14086 & ~n15981 ) | ( n14086 & n34645 ) | ( ~n15981 & n34645 ) ;
  assign n34647 = n21385 ^ n12971 ^ n1472 ;
  assign n34648 = n25859 & n34647 ;
  assign n34649 = n34646 & n34648 ;
  assign n34650 = n26646 ^ n13163 ^ 1'b0 ;
  assign n34651 = n16058 & ~n34650 ;
  assign n34652 = n12465 | n23653 ;
  assign n34653 = n25550 | n34652 ;
  assign n34654 = n9387 & ~n34653 ;
  assign n34655 = n34654 ^ n29190 ^ 1'b0 ;
  assign n34656 = n12193 ^ n1438 ^ 1'b0 ;
  assign n34657 = n30173 ^ x12 ^ 1'b0 ;
  assign n34658 = n20063 ^ n8717 ^ 1'b0 ;
  assign n34659 = n17244 ^ n15057 ^ 1'b0 ;
  assign n34660 = n29000 | n34659 ;
  assign n34661 = n7522 | n34660 ;
  assign n34662 = n19708 ^ n706 ^ 1'b0 ;
  assign n34663 = n5288 ^ n2867 ^ 1'b0 ;
  assign n34664 = n16274 | n34663 ;
  assign n34665 = n27168 ^ n16036 ^ n11411 ;
  assign n34666 = n6393 | n15698 ;
  assign n34667 = ( ~n8913 & n17088 ) | ( ~n8913 & n34666 ) | ( n17088 & n34666 ) ;
  assign n34668 = n3646 ^ n3283 ^ 1'b0 ;
  assign n34669 = n8823 & ~n10862 ;
  assign n34670 = n7844 & n34669 ;
  assign n34671 = n34670 ^ n13462 ^ 1'b0 ;
  assign n34672 = n25652 & n32028 ;
  assign n34673 = n29708 ^ n13295 ^ 1'b0 ;
  assign n34674 = n24403 & n34673 ;
  assign n34675 = n8568 & ~n11373 ;
  assign n34676 = n34675 ^ n11087 ^ 1'b0 ;
  assign n34677 = n34676 ^ n15744 ^ n11999 ;
  assign n34678 = n34677 ^ n10840 ^ 1'b0 ;
  assign n34679 = n12573 & n22948 ;
  assign n34680 = n34679 ^ n21780 ^ n17708 ;
  assign n34681 = ~n10692 & n34144 ;
  assign n34682 = n34681 ^ n5671 ^ 1'b0 ;
  assign n34683 = n3810 | n26605 ;
  assign n34684 = ~n4875 & n34683 ;
  assign n34690 = n4860 & ~n13749 ;
  assign n34687 = n27622 ^ n7422 ^ 1'b0 ;
  assign n34688 = ~n11524 & n26654 ;
  assign n34689 = n34687 | n34688 ;
  assign n34691 = n34690 ^ n34689 ^ 1'b0 ;
  assign n34685 = n33137 ^ n5109 ^ n4656 ;
  assign n34686 = ( ~n4766 & n32473 ) | ( ~n4766 & n34685 ) | ( n32473 & n34685 ) ;
  assign n34692 = n34691 ^ n34686 ^ 1'b0 ;
  assign n34693 = n1800 | n10481 ;
  assign n34694 = n34693 ^ n31276 ^ 1'b0 ;
  assign n34695 = ~n3365 & n34694 ;
  assign n34696 = n13832 & n31823 ;
  assign n34697 = ~n16313 & n34696 ;
  assign n34698 = n10544 & ~n11873 ;
  assign n34699 = n34698 ^ n33405 ^ 1'b0 ;
  assign n34700 = n3257 & ~n16585 ;
  assign n34702 = n7480 & ~n18492 ;
  assign n34701 = n2052 & ~n3924 ;
  assign n34703 = n34702 ^ n34701 ^ 1'b0 ;
  assign n34704 = ( ~n18318 & n34700 ) | ( ~n18318 & n34703 ) | ( n34700 & n34703 ) ;
  assign n34705 = ( ~n7527 & n11356 ) | ( ~n7527 & n21494 ) | ( n11356 & n21494 ) ;
  assign n34706 = n8986 & ~n34705 ;
  assign n34707 = n34706 ^ n22164 ^ n12611 ;
  assign n34708 = n24192 ^ n22853 ^ n20400 ;
  assign n34709 = n10815 & n15999 ;
  assign n34710 = n34709 ^ n9914 ^ 1'b0 ;
  assign n34711 = n18832 ^ n10080 ^ 1'b0 ;
  assign n34712 = n15843 & n34711 ;
  assign n34713 = n34710 | n34712 ;
  assign n34714 = n34713 ^ n31256 ^ n22452 ;
  assign n34715 = n431 & n15514 ;
  assign n34716 = n23182 ^ n17103 ^ n15915 ;
  assign n34717 = n33939 ^ n33045 ^ n23419 ;
  assign n34718 = n10956 ^ n7846 ^ n4619 ;
  assign n34719 = n30203 ^ n26736 ^ n17782 ;
  assign n34720 = n6553 & ~n34719 ;
  assign n34721 = n34720 ^ n5676 ^ 1'b0 ;
  assign n34722 = n22527 ^ n5984 ^ 1'b0 ;
  assign n34723 = n13632 ^ x106 ^ 1'b0 ;
  assign n34724 = n26180 ^ n7108 ^ 1'b0 ;
  assign n34725 = n34723 | n34724 ;
  assign n34726 = n1342 | n12240 ;
  assign n34727 = n9779 & ~n34726 ;
  assign n34728 = n14664 ^ n7704 ^ 1'b0 ;
  assign n34729 = ~n1022 & n34728 ;
  assign n34730 = ( n2889 & ~n19148 ) | ( n2889 & n34729 ) | ( ~n19148 & n34729 ) ;
  assign n34731 = ~n12498 & n13994 ;
  assign n34732 = n1217 & n34731 ;
  assign n34733 = n843 ^ n730 ^ 1'b0 ;
  assign n34734 = ( n9126 & ~n34732 ) | ( n9126 & n34733 ) | ( ~n34732 & n34733 ) ;
  assign n34735 = ( n33156 & ~n34730 ) | ( n33156 & n34734 ) | ( ~n34730 & n34734 ) ;
  assign n34736 = n15896 | n32415 ;
  assign n34737 = n25352 | n34736 ;
  assign n34738 = n9901 & n31249 ;
  assign n34739 = ~n15203 & n34738 ;
  assign n34740 = n32151 | n32212 ;
  assign n34741 = n1214 & n5941 ;
  assign n34742 = ~n32057 & n34741 ;
  assign n34743 = n33717 & ~n34742 ;
  assign n34744 = n24712 & n34743 ;
  assign n34745 = ( ~n15624 & n21950 ) | ( ~n15624 & n34744 ) | ( n21950 & n34744 ) ;
  assign n34746 = n20193 ^ n3837 ^ n1543 ;
  assign n34750 = n18404 ^ n11327 ^ n10282 ;
  assign n34751 = n34750 ^ n24502 ^ 1'b0 ;
  assign n34747 = n2924 | n6332 ;
  assign n34748 = n34747 ^ n6865 ^ n4044 ;
  assign n34749 = n3381 & ~n34748 ;
  assign n34752 = n34751 ^ n34749 ^ 1'b0 ;
  assign n34753 = n7698 & ~n17866 ;
  assign n34754 = n17969 ^ n13911 ^ 1'b0 ;
  assign n34755 = ~n34753 & n34754 ;
  assign n34760 = n21152 ^ n8455 ^ 1'b0 ;
  assign n34758 = n16383 ^ n1449 ^ 1'b0 ;
  assign n34759 = n23971 | n34758 ;
  assign n34756 = ( ~n5637 & n19522 ) | ( ~n5637 & n22397 ) | ( n19522 & n22397 ) ;
  assign n34757 = n34756 ^ n27430 ^ 1'b0 ;
  assign n34761 = n34760 ^ n34759 ^ n34757 ;
  assign n34763 = n14482 & n24997 ;
  assign n34764 = n34763 ^ n8889 ^ 1'b0 ;
  assign n34762 = ( ~n2321 & n6582 ) | ( ~n2321 & n11946 ) | ( n6582 & n11946 ) ;
  assign n34765 = n34764 ^ n34762 ^ 1'b0 ;
  assign n34766 = ( ~n885 & n4588 ) | ( ~n885 & n10034 ) | ( n4588 & n10034 ) ;
  assign n34767 = n34766 ^ n13480 ^ 1'b0 ;
  assign n34768 = n23087 ^ n1150 ^ 1'b0 ;
  assign n34769 = n21216 & n34768 ;
  assign n34770 = n4134 | n16732 ;
  assign n34771 = n15919 ^ n13541 ^ 1'b0 ;
  assign n34772 = n34771 ^ n15101 ^ n9760 ;
  assign n34773 = n26753 ^ n12738 ^ 1'b0 ;
  assign n34774 = n8377 | n34773 ;
  assign n34775 = n21344 & ~n34774 ;
  assign n34776 = n24611 ^ n18337 ^ n16994 ;
  assign n34777 = n25235 ^ n6800 ^ n2726 ;
  assign n34778 = n34777 ^ n22567 ^ n19825 ;
  assign n34779 = n34778 ^ n27208 ^ 1'b0 ;
  assign n34780 = n34779 ^ n16426 ^ 1'b0 ;
  assign n34781 = n12993 & ~n34780 ;
  assign n34782 = n11266 ^ n668 ^ x253 ;
  assign n34783 = n11959 & n34782 ;
  assign n34784 = n34783 ^ n1317 ^ 1'b0 ;
  assign n34785 = n7339 & ~n18382 ;
  assign n34786 = n28016 ^ n25112 ^ 1'b0 ;
  assign n34787 = ( ~n3780 & n9096 ) | ( ~n3780 & n24408 ) | ( n9096 & n24408 ) ;
  assign n34790 = n27281 ^ n7673 ^ x49 ;
  assign n34791 = n9312 & ~n34790 ;
  assign n34788 = n11666 ^ n4816 ^ 1'b0 ;
  assign n34789 = n34788 ^ n25835 ^ n11553 ;
  assign n34792 = n34791 ^ n34789 ^ n26272 ;
  assign n34793 = n2180 | n7833 ;
  assign n34794 = n34793 ^ n31139 ^ n29018 ;
  assign n34795 = n10884 ^ x147 ^ 1'b0 ;
  assign n34796 = n34794 | n34795 ;
  assign n34797 = n7642 ^ n3699 ^ 1'b0 ;
  assign n34798 = n34797 ^ n29758 ^ 1'b0 ;
  assign n34799 = ~n3191 & n29429 ;
  assign n34800 = n18823 ^ n18203 ^ n1542 ;
  assign n34801 = n9626 ^ n2189 ^ n1118 ;
  assign n34802 = ( n9098 & n10943 ) | ( n9098 & n31856 ) | ( n10943 & n31856 ) ;
  assign n34803 = n16997 ^ n8865 ^ 1'b0 ;
  assign n34804 = ~n976 & n34803 ;
  assign n34805 = n12465 | n31515 ;
  assign n34806 = n30787 ^ n14896 ^ 1'b0 ;
  assign n34807 = ~n19881 & n34806 ;
  assign n34808 = ( n1674 & ~n10863 ) | ( n1674 & n17858 ) | ( ~n10863 & n17858 ) ;
  assign n34809 = ( ~n10476 & n27764 ) | ( ~n10476 & n34808 ) | ( n27764 & n34808 ) ;
  assign n34810 = n10430 ^ n7490 ^ n2040 ;
  assign n34811 = ( n2335 & n25117 ) | ( n2335 & n34810 ) | ( n25117 & n34810 ) ;
  assign n34812 = n34811 ^ n24589 ^ n24494 ;
  assign n34814 = n16419 & ~n17744 ;
  assign n34815 = ~x198 & n34814 ;
  assign n34816 = n34815 ^ n5763 ^ 1'b0 ;
  assign n34813 = n17660 & ~n31296 ;
  assign n34817 = n34816 ^ n34813 ^ 1'b0 ;
  assign n34818 = ( ~n8151 & n31183 ) | ( ~n8151 & n31667 ) | ( n31183 & n31667 ) ;
  assign n34819 = ~n34817 & n34818 ;
  assign n34820 = n34812 & n34819 ;
  assign n34821 = n8345 | n34820 ;
  assign n34822 = n12578 ^ n10987 ^ 1'b0 ;
  assign n34823 = n24157 ^ n23444 ^ n17561 ;
  assign n34824 = n2026 | n14679 ;
  assign n34825 = n21010 ^ n946 ^ 1'b0 ;
  assign n34826 = n34824 & ~n34825 ;
  assign n34827 = n34826 ^ n29419 ^ 1'b0 ;
  assign n34828 = n1743 & n29696 ;
  assign n34829 = n34828 ^ n17102 ^ n7413 ;
  assign n34830 = ~n27212 & n34829 ;
  assign n34831 = n1315 & ~n1864 ;
  assign n34832 = ~n12903 & n18361 ;
  assign n34833 = ~n34831 & n34832 ;
  assign n34834 = n34833 ^ n29212 ^ 1'b0 ;
  assign n34835 = ~n25160 & n34834 ;
  assign n34836 = n15230 ^ n7641 ^ n6140 ;
  assign n34843 = n3550 & ~n5239 ;
  assign n34844 = n27066 & n34843 ;
  assign n34837 = n17446 ^ n2553 ^ 1'b0 ;
  assign n34838 = n8719 | n34837 ;
  assign n34839 = ( n9150 & n18823 ) | ( n9150 & ~n34838 ) | ( n18823 & ~n34838 ) ;
  assign n34840 = n34839 ^ n5565 ^ 1'b0 ;
  assign n34841 = n5547 & n34840 ;
  assign n34842 = n34841 ^ n12139 ^ n7173 ;
  assign n34845 = n34844 ^ n34842 ^ 1'b0 ;
  assign n34846 = n16049 & ~n33615 ;
  assign n34847 = ~n14027 & n34846 ;
  assign n34848 = n34845 & ~n34847 ;
  assign n34849 = n336 & ~n14892 ;
  assign n34850 = n34849 ^ n6940 ^ n1542 ;
  assign n34851 = ~n14804 & n23115 ;
  assign n34852 = n28233 & ~n34851 ;
  assign n34853 = n34852 ^ n6852 ^ 1'b0 ;
  assign n34854 = n34850 & ~n34853 ;
  assign n34855 = ( n4088 & ~n16268 ) | ( n4088 & n34854 ) | ( ~n16268 & n34854 ) ;
  assign n34856 = n27590 ^ n2391 ^ 1'b0 ;
  assign n34857 = n20814 | n27900 ;
  assign n34858 = n4757 | n30289 ;
  assign n34859 = n34858 ^ n20526 ^ 1'b0 ;
  assign n34860 = n32130 | n34859 ;
  assign n34861 = n26302 ^ n9865 ^ 1'b0 ;
  assign n34862 = n34861 ^ n21894 ^ 1'b0 ;
  assign n34863 = n29761 & n34862 ;
  assign n34864 = ~n23923 & n34863 ;
  assign n34865 = n10334 & n34864 ;
  assign n34867 = ( n14368 & n22181 ) | ( n14368 & n34764 ) | ( n22181 & n34764 ) ;
  assign n34868 = n34867 ^ n29563 ^ n301 ;
  assign n34866 = n20389 ^ n9743 ^ n9396 ;
  assign n34869 = n34868 ^ n34866 ^ 1'b0 ;
  assign n34870 = n1881 ^ n1494 ^ 1'b0 ;
  assign n34871 = n936 & ~n34870 ;
  assign n34872 = n34871 ^ n34600 ^ 1'b0 ;
  assign n34873 = ( n4268 & n14316 ) | ( n4268 & ~n24377 ) | ( n14316 & ~n24377 ) ;
  assign n34874 = ~n8490 & n34873 ;
  assign n34875 = n8635 & n34874 ;
  assign n34876 = n34875 ^ n9058 ^ n443 ;
  assign n34877 = ~n27641 & n34876 ;
  assign n34879 = n24890 | n27908 ;
  assign n34880 = n5440 & ~n34879 ;
  assign n34878 = n15691 ^ n9735 ^ 1'b0 ;
  assign n34881 = n34880 ^ n34878 ^ n9531 ;
  assign n34882 = n1091 & ~n25565 ;
  assign n34883 = n14600 & n34882 ;
  assign n34884 = n16496 | n34883 ;
  assign n34885 = ~n829 & n24301 ;
  assign n34886 = n11738 & ~n23247 ;
  assign n34887 = n27649 ^ n13401 ^ n12460 ;
  assign n34888 = n34886 | n34887 ;
  assign n34889 = x78 & ~n2314 ;
  assign n34890 = n34889 ^ n23528 ^ 1'b0 ;
  assign n34891 = n15631 | n34890 ;
  assign n34892 = n7185 ^ n4165 ^ n3830 ;
  assign n34893 = n34892 ^ n11341 ^ n5276 ;
  assign n34894 = n7918 ^ n4697 ^ 1'b0 ;
  assign n34895 = n2683 & n34894 ;
  assign n34896 = ( ~n6693 & n17685 ) | ( ~n6693 & n34895 ) | ( n17685 & n34895 ) ;
  assign n34897 = n15832 ^ n10556 ^ 1'b0 ;
  assign n34898 = n6123 ^ n3902 ^ 1'b0 ;
  assign n34899 = n34897 | n34898 ;
  assign n34903 = n19160 ^ n18691 ^ 1'b0 ;
  assign n34904 = ~n15985 & n34903 ;
  assign n34900 = n23484 ^ n11945 ^ n6229 ;
  assign n34901 = n34900 ^ n25301 ^ 1'b0 ;
  assign n34902 = n15274 & n34901 ;
  assign n34905 = n34904 ^ n34902 ^ n1924 ;
  assign n34906 = n25536 ^ n15280 ^ 1'b0 ;
  assign n34907 = n1007 & ~n18823 ;
  assign n34908 = n18218 & n34907 ;
  assign n34909 = n4694 | n9517 ;
  assign n34910 = n5239 & ~n34909 ;
  assign n34911 = ( n1208 & ~n5970 ) | ( n1208 & n34910 ) | ( ~n5970 & n34910 ) ;
  assign n34912 = ( ~n21621 & n34908 ) | ( ~n21621 & n34911 ) | ( n34908 & n34911 ) ;
  assign n34913 = n34380 | n34912 ;
  assign n34914 = n33865 | n34913 ;
  assign n34915 = n11669 & n34914 ;
  assign n34916 = n34915 ^ n4242 ^ 1'b0 ;
  assign n34917 = n25872 ^ n7302 ^ 1'b0 ;
  assign n34918 = n863 | n34917 ;
  assign n34919 = n27303 ^ n15333 ^ 1'b0 ;
  assign n34920 = ~n15844 & n34919 ;
  assign n34921 = ( n18778 & ~n21319 ) | ( n18778 & n21403 ) | ( ~n21319 & n21403 ) ;
  assign n34922 = n34921 ^ n14613 ^ n12143 ;
  assign n34923 = n435 & ~n8431 ;
  assign n34924 = ( ~n4877 & n27628 ) | ( ~n4877 & n34923 ) | ( n27628 & n34923 ) ;
  assign n34925 = n2743 | n10958 ;
  assign n34926 = n25507 & n34925 ;
  assign n34927 = n34926 ^ n26998 ^ n11475 ;
  assign n34928 = n20438 ^ n13337 ^ 1'b0 ;
  assign n34929 = n33127 | n34928 ;
  assign n34930 = n355 & n4360 ;
  assign n34931 = n7374 & n34930 ;
  assign n34932 = n26639 ^ n6967 ^ 1'b0 ;
  assign n34933 = ~n34931 & n34932 ;
  assign n34934 = n32990 ^ n9080 ^ 1'b0 ;
  assign n34939 = n29824 | n34276 ;
  assign n34940 = n9102 | n34939 ;
  assign n34935 = n16106 ^ n545 ^ 1'b0 ;
  assign n34936 = n9486 | n34935 ;
  assign n34937 = n34936 ^ n5250 ^ 1'b0 ;
  assign n34938 = n31608 | n34937 ;
  assign n34941 = n34940 ^ n34938 ^ n23216 ;
  assign n34942 = n22305 & ~n26008 ;
  assign n34943 = n28618 & n34942 ;
  assign n34944 = ~n17661 & n34943 ;
  assign n34945 = n34944 ^ n34365 ^ 1'b0 ;
  assign n34946 = n3941 & ~n21633 ;
  assign n34947 = n34946 ^ n6630 ^ n5892 ;
  assign n34948 = n16203 ^ n13151 ^ n6714 ;
  assign n34949 = n20970 | n34948 ;
  assign n34950 = n34949 ^ n20373 ^ 1'b0 ;
  assign n34951 = n25941 & n34950 ;
  assign n34952 = ~n18403 & n23630 ;
  assign n34953 = ~n6570 & n34952 ;
  assign n34954 = ( n2123 & n6743 ) | ( n2123 & n19827 ) | ( n6743 & n19827 ) ;
  assign n34955 = n27877 ^ n3459 ^ n1763 ;
  assign n34956 = n23024 ^ n10199 ^ n3174 ;
  assign n34957 = n14561 ^ n1933 ^ 1'b0 ;
  assign n34958 = n20458 ^ n18616 ^ 1'b0 ;
  assign n34959 = ~n34957 & n34958 ;
  assign n34960 = n2693 & ~n10107 ;
  assign n34961 = ~n2008 & n34960 ;
  assign n34962 = n34961 ^ n5169 ^ n671 ;
  assign n34963 = n15675 ^ n10729 ^ n3000 ;
  assign n34964 = ( n10042 & n12867 ) | ( n10042 & n19805 ) | ( n12867 & n19805 ) ;
  assign n34966 = n26980 ^ n24089 ^ 1'b0 ;
  assign n34967 = n22465 & n34966 ;
  assign n34965 = n21192 | n33303 ;
  assign n34968 = n34967 ^ n34965 ^ 1'b0 ;
  assign n34970 = n23527 & n27226 ;
  assign n34971 = n1350 & n34970 ;
  assign n34972 = x55 & ~n28840 ;
  assign n34973 = n34971 & n34972 ;
  assign n34969 = ~n8809 & n17157 ;
  assign n34974 = n34973 ^ n34969 ^ 1'b0 ;
  assign n34975 = ( ~n8282 & n12280 ) | ( ~n8282 & n27232 ) | ( n12280 & n27232 ) ;
  assign n34976 = n12048 | n13276 ;
  assign n34977 = n34976 ^ n25016 ^ 1'b0 ;
  assign n34978 = ( n4530 & ~n8210 ) | ( n4530 & n34977 ) | ( ~n8210 & n34977 ) ;
  assign n34979 = n12422 & n12620 ;
  assign n34980 = n13824 & n34979 ;
  assign n34981 = n19457 ^ n8634 ^ 1'b0 ;
  assign n34982 = n7134 ^ n987 ^ 1'b0 ;
  assign n34983 = ~n34981 & n34982 ;
  assign n34984 = ( n5057 & n34980 ) | ( n5057 & n34983 ) | ( n34980 & n34983 ) ;
  assign n34985 = ~n4823 & n5285 ;
  assign n34986 = n2142 & n34985 ;
  assign n34989 = n8011 & ~n11590 ;
  assign n34990 = ~x52 & n34989 ;
  assign n34991 = ( ~n2846 & n29348 ) | ( ~n2846 & n34990 ) | ( n29348 & n34990 ) ;
  assign n34987 = n8540 | n23210 ;
  assign n34988 = n34987 ^ n20286 ^ 1'b0 ;
  assign n34992 = n34991 ^ n34988 ^ 1'b0 ;
  assign n34993 = n34986 | n34992 ;
  assign n34994 = n34993 ^ n22325 ^ n12216 ;
  assign n34995 = n18659 & n34994 ;
  assign n34996 = n3106 & ~n14060 ;
  assign n34997 = n34995 & n34996 ;
  assign n34998 = n30352 & n32987 ;
  assign n34999 = n34998 ^ n17096 ^ 1'b0 ;
  assign n35000 = n30143 ^ n11816 ^ n4708 ;
  assign n35004 = n2354 ^ n526 ^ 1'b0 ;
  assign n35005 = n1858 | n35004 ;
  assign n35006 = n35005 ^ n19695 ^ n10146 ;
  assign n35003 = n20046 & n20601 ;
  assign n35007 = n35006 ^ n35003 ^ 1'b0 ;
  assign n35001 = n9745 & n31359 ;
  assign n35002 = n35001 ^ n14634 ^ n4632 ;
  assign n35008 = n35007 ^ n35002 ^ n14740 ;
  assign n35009 = n35008 ^ n7673 ^ n3772 ;
  assign n35010 = n35000 | n35009 ;
  assign n35011 = n11447 & ~n25143 ;
  assign n35012 = ( ~n3093 & n19259 ) | ( ~n3093 & n35011 ) | ( n19259 & n35011 ) ;
  assign n35013 = n9078 | n23178 ;
  assign n35014 = n35013 ^ n1984 ^ 1'b0 ;
  assign n35015 = ( n17751 & ~n34301 ) | ( n17751 & n35014 ) | ( ~n34301 & n35014 ) ;
  assign n35016 = n10924 & n35015 ;
  assign n35017 = n22643 | n26079 ;
  assign n35018 = n35017 ^ n17850 ^ 1'b0 ;
  assign n35019 = ~n5274 & n31866 ;
  assign n35020 = n35019 ^ n8950 ^ 1'b0 ;
  assign n35021 = n23457 & n35020 ;
  assign n35022 = ~n2215 & n35021 ;
  assign n35023 = n35022 ^ n3923 ^ 1'b0 ;
  assign n35024 = ~n17685 & n22401 ;
  assign n35026 = n25284 ^ n23305 ^ 1'b0 ;
  assign n35027 = n4819 & ~n35026 ;
  assign n35028 = n35027 ^ n12140 ^ n7431 ;
  assign n35029 = ( n14540 & n25844 ) | ( n14540 & ~n35028 ) | ( n25844 & ~n35028 ) ;
  assign n35025 = n4291 & ~n13073 ;
  assign n35030 = n35029 ^ n35025 ^ n20178 ;
  assign n35031 = n18248 ^ n10111 ^ 1'b0 ;
  assign n35032 = ( ~n3122 & n8483 ) | ( ~n3122 & n16514 ) | ( n8483 & n16514 ) ;
  assign n35033 = n13921 & ~n30455 ;
  assign n35034 = n6879 & n35033 ;
  assign n35035 = n4368 & n6427 ;
  assign n35036 = n35035 ^ n18351 ^ 1'b0 ;
  assign n35037 = ~n17834 & n20096 ;
  assign n35038 = n29064 & n35037 ;
  assign n35039 = n15731 | n35038 ;
  assign n35040 = n18664 ^ n18364 ^ n1320 ;
  assign n35041 = n22063 ^ n13317 ^ 1'b0 ;
  assign n35042 = n35041 ^ n33312 ^ n16427 ;
  assign n35043 = n1352 & n18911 ;
  assign n35044 = n5162 & n35043 ;
  assign n35045 = n35044 ^ n18247 ^ n14667 ;
  assign n35046 = x169 & n26193 ;
  assign n35047 = n8959 | n14436 ;
  assign n35048 = n35047 ^ n21335 ^ 1'b0 ;
  assign n35049 = n11843 & ~n35048 ;
  assign n35050 = n35049 ^ n4499 ^ 1'b0 ;
  assign n35051 = n2783 | n35050 ;
  assign n35052 = n17592 & ~n24750 ;
  assign n35053 = n29403 ^ n10316 ^ n4622 ;
  assign n35054 = n28611 ^ n4730 ^ 1'b0 ;
  assign n35055 = n7402 & n35054 ;
  assign n35056 = ( n18171 & n35053 ) | ( n18171 & ~n35055 ) | ( n35053 & ~n35055 ) ;
  assign n35057 = n35056 ^ n5836 ^ 1'b0 ;
  assign n35058 = ~n3069 & n22325 ;
  assign n35059 = ~n14075 & n35058 ;
  assign n35060 = ( ~n9351 & n9478 ) | ( ~n9351 & n35059 ) | ( n9478 & n35059 ) ;
  assign n35061 = n35060 ^ n32574 ^ n28196 ;
  assign n35062 = n26467 ^ n23146 ^ 1'b0 ;
  assign n35063 = ( ~n2024 & n3306 ) | ( ~n2024 & n35062 ) | ( n3306 & n35062 ) ;
  assign n35064 = n1551 | n28827 ;
  assign n35065 = n8226 | n35064 ;
  assign n35066 = n10898 & n20331 ;
  assign n35067 = n35066 ^ n20551 ^ 1'b0 ;
  assign n35068 = ~n25927 & n35067 ;
  assign n35069 = n23569 ^ n13715 ^ x241 ;
  assign n35070 = n35069 ^ n27899 ^ n23267 ;
  assign n35071 = n18144 & ~n35070 ;
  assign n35072 = ( ~n10904 & n15333 ) | ( ~n10904 & n16177 ) | ( n15333 & n16177 ) ;
  assign n35073 = n27463 | n35072 ;
  assign n35074 = n35073 ^ n19077 ^ 1'b0 ;
  assign n35075 = n31061 & ~n35074 ;
  assign n35076 = n16028 & n18249 ;
  assign n35077 = ~n11185 & n35076 ;
  assign n35078 = n35077 ^ n8427 ^ 1'b0 ;
  assign n35082 = n8475 ^ n4847 ^ 1'b0 ;
  assign n35083 = n9919 & n35082 ;
  assign n35079 = n30851 ^ n27554 ^ n2113 ;
  assign n35080 = ( n827 & ~n8726 ) | ( n827 & n35079 ) | ( ~n8726 & n35079 ) ;
  assign n35081 = n35080 ^ n867 ^ 1'b0 ;
  assign n35084 = n35083 ^ n35081 ^ n12821 ;
  assign n35085 = ( n15522 & ~n23166 ) | ( n15522 & n27912 ) | ( ~n23166 & n27912 ) ;
  assign n35086 = n3897 ^ n1491 ^ 1'b0 ;
  assign n35087 = ( n6874 & n10919 ) | ( n6874 & ~n10936 ) | ( n10919 & ~n10936 ) ;
  assign n35088 = ~n1936 & n18133 ;
  assign n35089 = ~n12803 & n35088 ;
  assign n35090 = n8787 & n18650 ;
  assign n35091 = n35089 & n35090 ;
  assign n35095 = n3307 | n13101 ;
  assign n35093 = n9411 ^ n7569 ^ 1'b0 ;
  assign n35094 = n13385 & ~n35093 ;
  assign n35096 = n35095 ^ n35094 ^ n19112 ;
  assign n35092 = n14988 ^ n1720 ^ 1'b0 ;
  assign n35097 = n35096 ^ n35092 ^ n8075 ;
  assign n35098 = n35097 ^ n32176 ^ 1'b0 ;
  assign n35099 = ~n11517 & n20104 ;
  assign n35100 = n15919 ^ n883 ^ 1'b0 ;
  assign n35101 = ~n35099 & n35100 ;
  assign n35102 = n10116 & n35101 ;
  assign n35103 = n12928 & ~n24184 ;
  assign n35104 = n35103 ^ n29204 ^ n15448 ;
  assign n35105 = n17876 | n21532 ;
  assign n35106 = n2140 & ~n35105 ;
  assign n35107 = n35106 ^ n9872 ^ 1'b0 ;
  assign n35108 = n27568 ^ n15244 ^ 1'b0 ;
  assign n35109 = n29414 ^ n14684 ^ 1'b0 ;
  assign n35110 = n35108 | n35109 ;
  assign n35111 = n26793 ^ n19569 ^ n9311 ;
  assign n35112 = n4147 & n10312 ;
  assign n35113 = n22021 ^ n7962 ^ n1277 ;
  assign n35114 = n35113 ^ n5399 ^ 1'b0 ;
  assign n35115 = ( n15654 & n22724 ) | ( n15654 & ~n35114 ) | ( n22724 & ~n35114 ) ;
  assign n35116 = ( n19712 & n35112 ) | ( n19712 & n35115 ) | ( n35112 & n35115 ) ;
  assign n35117 = ~n1562 & n8992 ;
  assign n35118 = n35117 ^ n841 ^ 1'b0 ;
  assign n35119 = n639 | n763 ;
  assign n35120 = n35118 & ~n35119 ;
  assign n35123 = ( n7566 & n12011 ) | ( n7566 & ~n24192 ) | ( n12011 & ~n24192 ) ;
  assign n35124 = n22310 & n35123 ;
  assign n35121 = n10903 & n14859 ;
  assign n35122 = n35121 ^ n27879 ^ n21416 ;
  assign n35125 = n35124 ^ n35122 ^ 1'b0 ;
  assign n35126 = ~n20395 & n35125 ;
  assign n35128 = n20486 ^ n11240 ^ 1'b0 ;
  assign n35129 = ~n20493 & n35128 ;
  assign n35127 = n4591 | n14937 ;
  assign n35130 = n35129 ^ n35127 ^ 1'b0 ;
  assign n35131 = n30040 | n34002 ;
  assign n35132 = n1517 | n9396 ;
  assign n35133 = n35132 ^ n12117 ^ 1'b0 ;
  assign n35134 = n6352 ^ n429 ^ 1'b0 ;
  assign n35135 = ~n35133 & n35134 ;
  assign n35136 = n35135 ^ n6100 ^ 1'b0 ;
  assign n35137 = ~n14805 & n30133 ;
  assign n35138 = ~n29648 & n35137 ;
  assign n35139 = n35138 ^ n5100 ^ 1'b0 ;
  assign n35140 = n3004 & n11295 ;
  assign n35141 = n35140 ^ n27276 ^ n16369 ;
  assign n35142 = ~n3883 & n35141 ;
  assign n35143 = n35142 ^ n1678 ^ 1'b0 ;
  assign n35144 = ~n35139 & n35143 ;
  assign n35145 = n613 & ~n27240 ;
  assign n35146 = n24361 & n35145 ;
  assign n35151 = n33575 ^ n11746 ^ n3278 ;
  assign n35147 = ( n2760 & ~n18327 ) | ( n2760 & n18484 ) | ( ~n18327 & n18484 ) ;
  assign n35148 = n18926 ^ n11913 ^ 1'b0 ;
  assign n35149 = n35147 & ~n35148 ;
  assign n35150 = n6553 & n35149 ;
  assign n35152 = n35151 ^ n35150 ^ 1'b0 ;
  assign n35153 = n1629 & n35152 ;
  assign n35154 = ( ~n444 & n5458 ) | ( ~n444 & n5669 ) | ( n5458 & n5669 ) ;
  assign n35156 = n25613 ^ n13942 ^ n5445 ;
  assign n35157 = n22325 ^ n20711 ^ 1'b0 ;
  assign n35158 = n35156 & ~n35157 ;
  assign n35159 = n35158 ^ n14859 ^ 1'b0 ;
  assign n35160 = ~n11437 & n35159 ;
  assign n35155 = n14321 & ~n34825 ;
  assign n35161 = n35160 ^ n35155 ^ 1'b0 ;
  assign n35162 = n35161 ^ n29167 ^ n12718 ;
  assign n35163 = n35162 ^ n11993 ^ 1'b0 ;
  assign n35164 = n35154 | n35163 ;
  assign n35165 = n33775 ^ n28865 ^ 1'b0 ;
  assign n35166 = n21932 ^ n10513 ^ 1'b0 ;
  assign n35167 = n11857 | n15397 ;
  assign n35168 = n35167 ^ n9267 ^ 1'b0 ;
  assign n35169 = n18052 & n35168 ;
  assign n35170 = ( n9182 & n13175 ) | ( n9182 & ~n29782 ) | ( n13175 & ~n29782 ) ;
  assign n35172 = n831 & ~n4427 ;
  assign n35173 = n35172 ^ n4053 ^ 1'b0 ;
  assign n35171 = n17046 & n32377 ;
  assign n35174 = n35173 ^ n35171 ^ 1'b0 ;
  assign n35175 = n27424 ^ n2475 ^ n1367 ;
  assign n35176 = n25093 & ~n35175 ;
  assign n35177 = n35174 & n35176 ;
  assign n35178 = n7969 & ~n16021 ;
  assign n35179 = n35178 ^ n3327 ^ 1'b0 ;
  assign n35181 = n6398 ^ n1824 ^ n388 ;
  assign n35180 = n13021 ^ n11356 ^ n6417 ;
  assign n35182 = n35181 ^ n35180 ^ n20855 ;
  assign n35183 = n16818 | n35182 ;
  assign n35184 = n35183 ^ n4973 ^ 1'b0 ;
  assign n35185 = n30455 ^ n12522 ^ 1'b0 ;
  assign n35186 = ( ~n9874 & n16340 ) | ( ~n9874 & n35185 ) | ( n16340 & n35185 ) ;
  assign n35187 = n24095 ^ n5676 ^ 1'b0 ;
  assign n35188 = ~n16741 & n35187 ;
  assign n35189 = n27433 ^ n23067 ^ n10806 ;
  assign n35190 = n20120 & ~n35189 ;
  assign n35191 = n35190 ^ n3410 ^ 1'b0 ;
  assign n35192 = n31504 ^ n24038 ^ 1'b0 ;
  assign n35193 = n22865 ^ n20545 ^ 1'b0 ;
  assign n35194 = n33680 ^ n2645 ^ n1729 ;
  assign n35196 = x122 & n29396 ;
  assign n35197 = ~n335 & n35196 ;
  assign n35195 = ~n7617 & n30074 ;
  assign n35198 = n35197 ^ n35195 ^ 1'b0 ;
  assign n35199 = n9026 & n18404 ;
  assign n35200 = n35199 ^ n12311 ^ 1'b0 ;
  assign n35201 = ~n19415 & n35200 ;
  assign n35202 = n1062 & n28464 ;
  assign n35203 = n35202 ^ n24983 ^ 1'b0 ;
  assign n35204 = ( ~n2623 & n14789 ) | ( ~n2623 & n25879 ) | ( n14789 & n25879 ) ;
  assign n35205 = n15282 ^ n11178 ^ 1'b0 ;
  assign n35206 = n35204 | n35205 ;
  assign n35207 = n25323 ^ n8486 ^ n5075 ;
  assign n35208 = ~n1889 & n7709 ;
  assign n35209 = n8580 & ~n30982 ;
  assign n35210 = ~n1522 & n35209 ;
  assign n35211 = ~n18981 & n35210 ;
  assign n35212 = n13643 & n19209 ;
  assign n35213 = n7794 | n10605 ;
  assign n35214 = ~n702 & n35213 ;
  assign n35215 = n11879 & n33563 ;
  assign n35216 = n7729 & ~n35215 ;
  assign n35217 = n35214 & n35216 ;
  assign n35218 = n30807 ^ n27673 ^ n19731 ;
  assign n35219 = n17148 ^ n6679 ^ 1'b0 ;
  assign n35220 = n35218 | n35219 ;
  assign n35224 = n13376 | n13571 ;
  assign n35221 = n7994 & ~n22259 ;
  assign n35222 = n35221 ^ n24145 ^ 1'b0 ;
  assign n35223 = n14578 & n35222 ;
  assign n35225 = n35224 ^ n35223 ^ 1'b0 ;
  assign n35226 = n31960 & n35225 ;
  assign n35227 = n12957 | n30878 ;
  assign n35228 = ( n7079 & ~n34332 ) | ( n7079 & n35227 ) | ( ~n34332 & n35227 ) ;
  assign n35229 = n29278 ^ n20465 ^ 1'b0 ;
  assign n35230 = n35229 ^ n14138 ^ 1'b0 ;
  assign n35232 = ( n6425 & n7342 ) | ( n6425 & ~n12570 ) | ( n7342 & ~n12570 ) ;
  assign n35231 = n1600 & ~n11127 ;
  assign n35233 = n35232 ^ n35231 ^ n20266 ;
  assign n35236 = n32930 ^ n13748 ^ 1'b0 ;
  assign n35237 = n16942 & n35236 ;
  assign n35234 = n6369 & ~n8227 ;
  assign n35235 = n10136 | n35234 ;
  assign n35238 = n35237 ^ n35235 ^ 1'b0 ;
  assign n35239 = n21074 ^ n10399 ^ 1'b0 ;
  assign n35240 = n15542 ^ n10799 ^ 1'b0 ;
  assign n35241 = n35240 ^ n14251 ^ n1593 ;
  assign n35242 = ( n5328 & n12299 ) | ( n5328 & n26736 ) | ( n12299 & n26736 ) ;
  assign n35243 = n9659 | n35242 ;
  assign n35244 = n14725 | n35243 ;
  assign n35245 = n28347 | n35244 ;
  assign n35246 = n3148 | n15202 ;
  assign n35247 = n35246 ^ n32272 ^ 1'b0 ;
  assign n35248 = ~n9887 & n35247 ;
  assign n35249 = ( n8960 & n18327 ) | ( n8960 & ~n35248 ) | ( n18327 & ~n35248 ) ;
  assign n35250 = ~n17334 & n35249 ;
  assign n35251 = n5392 & n35250 ;
  assign n35252 = ( ~n1327 & n7510 ) | ( ~n1327 & n8442 ) | ( n7510 & n8442 ) ;
  assign n35253 = n5372 & ~n35252 ;
  assign n35254 = n35253 ^ n25249 ^ 1'b0 ;
  assign n35255 = n10846 ^ n3366 ^ 1'b0 ;
  assign n35256 = ( n6520 & ~n35254 ) | ( n6520 & n35255 ) | ( ~n35254 & n35255 ) ;
  assign n35257 = n33501 | n35256 ;
  assign n35258 = n26883 ^ n9449 ^ 1'b0 ;
  assign n35259 = ~n11950 & n35258 ;
  assign n35260 = n16338 ^ n10373 ^ 1'b0 ;
  assign n35261 = ~n21780 & n35260 ;
  assign n35262 = n35261 ^ n16004 ^ 1'b0 ;
  assign n35263 = n24377 ^ n22631 ^ 1'b0 ;
  assign n35264 = n8559 ^ n3498 ^ 1'b0 ;
  assign n35265 = n35264 ^ n7544 ^ 1'b0 ;
  assign n35266 = n10454 & n31271 ;
  assign n35267 = n2934 & n35266 ;
  assign n35268 = n35267 ^ n29498 ^ 1'b0 ;
  assign n35269 = n35265 & n35268 ;
  assign n35270 = n12103 | n17817 ;
  assign n35271 = n35270 ^ n1164 ^ 1'b0 ;
  assign n35272 = n26038 ^ n21736 ^ 1'b0 ;
  assign n35273 = ~n32486 & n35272 ;
  assign n35276 = ~n18671 & n23812 ;
  assign n35277 = n35276 ^ n6739 ^ 1'b0 ;
  assign n35274 = ~n15152 & n27622 ;
  assign n35275 = n23637 & ~n35274 ;
  assign n35278 = n35277 ^ n35275 ^ 1'b0 ;
  assign n35281 = n12960 ^ n4359 ^ 1'b0 ;
  assign n35282 = n4601 & ~n35281 ;
  assign n35279 = n1469 | n7682 ;
  assign n35280 = n35279 ^ n5250 ^ 1'b0 ;
  assign n35283 = n35282 ^ n35280 ^ 1'b0 ;
  assign n35284 = n6981 & ~n35283 ;
  assign n35285 = n10672 | n27379 ;
  assign n35286 = n16115 & ~n35285 ;
  assign n35287 = n14313 ^ n11469 ^ n8970 ;
  assign n35288 = ( n1292 & ~n1650 ) | ( n1292 & n8519 ) | ( ~n1650 & n8519 ) ;
  assign n35289 = n35288 ^ n29612 ^ n6326 ;
  assign n35290 = ( n2042 & n5336 ) | ( n2042 & n6311 ) | ( n5336 & n6311 ) ;
  assign n35291 = ~n17282 & n35290 ;
  assign n35292 = n35291 ^ n23313 ^ 1'b0 ;
  assign n35293 = n35292 ^ n4924 ^ x234 ;
  assign n35294 = n1081 & ~n9981 ;
  assign n35295 = ( n21268 & ~n32517 ) | ( n21268 & n35294 ) | ( ~n32517 & n35294 ) ;
  assign n35296 = ( ~x57 & x77 ) | ( ~x57 & n4835 ) | ( x77 & n4835 ) ;
  assign n35297 = ( n1656 & n2425 ) | ( n1656 & n25613 ) | ( n2425 & n25613 ) ;
  assign n35298 = ( n15706 & n16534 ) | ( n15706 & n35297 ) | ( n16534 & n35297 ) ;
  assign n35299 = n6306 ^ n702 ^ 1'b0 ;
  assign n35300 = n35299 ^ n12783 ^ 1'b0 ;
  assign n35301 = n35298 & ~n35300 ;
  assign n35302 = n35301 ^ n31152 ^ n25444 ;
  assign n35303 = ~n777 & n35302 ;
  assign n35304 = n35303 ^ n10827 ^ n8752 ;
  assign n35305 = n35304 ^ n26369 ^ 1'b0 ;
  assign n35306 = n22468 & n29224 ;
  assign n35307 = n35306 ^ n3225 ^ 1'b0 ;
  assign n35308 = n35307 ^ n4384 ^ 1'b0 ;
  assign n35309 = n955 & n35308 ;
  assign n35310 = n30239 | n35309 ;
  assign n35311 = n8921 ^ n5212 ^ n1408 ;
  assign n35312 = n21375 & ~n35311 ;
  assign n35313 = n35312 ^ n3658 ^ 1'b0 ;
  assign n35314 = n34677 & n35313 ;
  assign n35315 = n24450 ^ n20542 ^ n13963 ;
  assign n35316 = n17662 & n26076 ;
  assign n35317 = n35316 ^ n13423 ^ n9545 ;
  assign n35318 = n9002 & ~n35317 ;
  assign n35319 = n25238 ^ n20970 ^ 1'b0 ;
  assign n35320 = ( n4542 & ~n7505 ) | ( n4542 & n31904 ) | ( ~n7505 & n31904 ) ;
  assign n35321 = n16549 & ~n25645 ;
  assign n35322 = n2474 & n5652 ;
  assign n35323 = ~n9976 & n10534 ;
  assign n35324 = n35322 & n35323 ;
  assign n35325 = n27302 ^ n2662 ^ 1'b0 ;
  assign n35326 = n3502 | n35325 ;
  assign n35327 = n30657 ^ n5722 ^ 1'b0 ;
  assign n35328 = n34910 ^ n5451 ^ 1'b0 ;
  assign n35329 = n35327 | n35328 ;
  assign n35330 = n35329 ^ n10772 ^ 1'b0 ;
  assign n35331 = n19545 ^ n16563 ^ 1'b0 ;
  assign n35332 = n11909 & n28492 ;
  assign n35333 = ( n15390 & n18710 ) | ( n15390 & ~n35332 ) | ( n18710 & ~n35332 ) ;
  assign n35334 = ( n2697 & n8008 ) | ( n2697 & n8187 ) | ( n8008 & n8187 ) ;
  assign n35335 = n24631 & ~n35334 ;
  assign n35336 = n24233 ^ n15568 ^ 1'b0 ;
  assign n35337 = n18181 ^ n7579 ^ 1'b0 ;
  assign n35338 = ~n10715 & n17500 ;
  assign n35339 = ( n4991 & n20377 ) | ( n4991 & ~n35338 ) | ( n20377 & ~n35338 ) ;
  assign n35340 = n17970 ^ n7490 ^ 1'b0 ;
  assign n35341 = n5892 ^ n1159 ^ 1'b0 ;
  assign n35342 = n1101 & n35341 ;
  assign n35343 = ( n7745 & ~n17502 ) | ( n7745 & n35342 ) | ( ~n17502 & n35342 ) ;
  assign n35344 = ~n15956 & n35343 ;
  assign n35345 = n35344 ^ n2011 ^ 1'b0 ;
  assign n35346 = n18363 ^ n4437 ^ n3322 ;
  assign n35347 = ( n10650 & ~n32417 ) | ( n10650 & n35346 ) | ( ~n32417 & n35346 ) ;
  assign n35348 = n24148 & ~n29436 ;
  assign n35349 = n35347 & n35348 ;
  assign n35350 = n16336 | n18407 ;
  assign n35351 = ( ~n3088 & n7274 ) | ( ~n3088 & n32306 ) | ( n7274 & n32306 ) ;
  assign n35353 = ~n830 & n5949 ;
  assign n35354 = n31111 & ~n35353 ;
  assign n35355 = n1474 & n35354 ;
  assign n35352 = ( ~n393 & n1616 ) | ( ~n393 & n25658 ) | ( n1616 & n25658 ) ;
  assign n35356 = n35355 ^ n35352 ^ n8198 ;
  assign n35357 = n12313 ^ n659 ^ 1'b0 ;
  assign n35358 = n2330 & n13327 ;
  assign n35359 = n16201 & n35358 ;
  assign n35360 = n35359 ^ n8786 ^ 1'b0 ;
  assign n35361 = ( n5683 & n10265 ) | ( n5683 & ~n13283 ) | ( n10265 & ~n13283 ) ;
  assign n35362 = n31505 & n35361 ;
  assign n35363 = ~n18549 & n35362 ;
  assign n35367 = ~n8146 & n19615 ;
  assign n35368 = ~n2740 & n35367 ;
  assign n35364 = n2328 & ~n5759 ;
  assign n35365 = n35364 ^ n15910 ^ 1'b0 ;
  assign n35366 = ~n18513 & n35365 ;
  assign n35369 = n35368 ^ n35366 ^ n32418 ;
  assign n35370 = ( n780 & n2686 ) | ( n780 & n4449 ) | ( n2686 & n4449 ) ;
  assign n35371 = n12571 ^ n4478 ^ 1'b0 ;
  assign n35372 = ~n8702 & n32171 ;
  assign n35373 = n13334 ^ n4827 ^ n979 ;
  assign n35374 = ( ~n3920 & n13941 ) | ( ~n3920 & n35373 ) | ( n13941 & n35373 ) ;
  assign n35375 = n24351 & ~n35374 ;
  assign n35376 = n35375 ^ n13879 ^ 1'b0 ;
  assign n35377 = n4440 | n34688 ;
  assign n35378 = n35376 | n35377 ;
  assign n35379 = n1434 | n34805 ;
  assign n35380 = n20227 ^ n16934 ^ n12752 ;
  assign n35381 = ( ~n28336 & n32757 ) | ( ~n28336 & n35380 ) | ( n32757 & n35380 ) ;
  assign n35382 = n8178 | n10002 ;
  assign n35383 = n6005 | n35382 ;
  assign n35384 = n7770 ^ n471 ^ 1'b0 ;
  assign n35385 = n35384 ^ n31525 ^ 1'b0 ;
  assign n35386 = n25686 | n35385 ;
  assign n35387 = ~n11685 & n31286 ;
  assign n35388 = n13725 | n35387 ;
  assign n35389 = n22343 & ~n35388 ;
  assign n35390 = n30468 ^ n17095 ^ n3736 ;
  assign n35391 = n35280 ^ n17851 ^ n17327 ;
  assign n35392 = n6942 ^ n450 ^ 1'b0 ;
  assign n35393 = n18717 & n35392 ;
  assign n35394 = ~n12570 & n35393 ;
  assign n35395 = n5481 & n35394 ;
  assign n35396 = n10334 | n13698 ;
  assign n35397 = ~n35395 & n35396 ;
  assign n35398 = n11229 & ~n13857 ;
  assign n35399 = n26123 & n35398 ;
  assign n35400 = n2191 & ~n7744 ;
  assign n35401 = n35400 ^ n25401 ^ 1'b0 ;
  assign n35403 = ( n9150 & ~n17573 ) | ( n9150 & n17799 ) | ( ~n17573 & n17799 ) ;
  assign n35402 = n14579 & ~n27018 ;
  assign n35404 = n35403 ^ n35402 ^ 1'b0 ;
  assign n35405 = n22485 & n27993 ;
  assign n35406 = n33775 ^ n30305 ^ 1'b0 ;
  assign n35407 = n11747 & n35406 ;
  assign n35408 = n35405 & n35407 ;
  assign n35409 = n13646 | n16993 ;
  assign n35410 = n35409 ^ n2201 ^ 1'b0 ;
  assign n35411 = n35410 ^ n25404 ^ n6617 ;
  assign n35412 = n8099 ^ n2825 ^ 1'b0 ;
  assign n35413 = n13367 | n16914 ;
  assign n35414 = n35413 ^ n9757 ^ 1'b0 ;
  assign n35415 = ( n4398 & n23484 ) | ( n4398 & ~n35414 ) | ( n23484 & ~n35414 ) ;
  assign n35416 = n26902 & ~n35415 ;
  assign n35417 = n13966 & n34749 ;
  assign n35418 = n35417 ^ n30124 ^ 1'b0 ;
  assign n35419 = n20339 ^ n12726 ^ 1'b0 ;
  assign n35420 = n10128 & n35419 ;
  assign n35421 = n7668 ^ n5529 ^ 1'b0 ;
  assign n35422 = n35420 & n35421 ;
  assign n35423 = n20204 ^ n14311 ^ n12201 ;
  assign n35426 = n30714 ^ n659 ^ 1'b0 ;
  assign n35424 = n7475 | n11475 ;
  assign n35425 = n18284 & ~n35424 ;
  assign n35427 = n35426 ^ n35425 ^ n2119 ;
  assign n35428 = ~n5042 & n14336 ;
  assign n35429 = ~n14336 & n35428 ;
  assign n35430 = n3478 & ~n35429 ;
  assign n35431 = ( n9779 & ~n18490 ) | ( n9779 & n35430 ) | ( ~n18490 & n35430 ) ;
  assign n35432 = n831 & ~n12168 ;
  assign n35433 = n26852 ^ n9615 ^ n6254 ;
  assign n35434 = n35432 | n35433 ;
  assign n35439 = ( n15290 & n15950 ) | ( n15290 & ~n19453 ) | ( n15950 & ~n19453 ) ;
  assign n35438 = n5173 & ~n8939 ;
  assign n35440 = n35439 ^ n35438 ^ n8062 ;
  assign n35441 = ( n6994 & ~n17850 ) | ( n6994 & n35440 ) | ( ~n17850 & n35440 ) ;
  assign n35435 = n10195 & ~n12201 ;
  assign n35436 = n35435 ^ n31361 ^ 1'b0 ;
  assign n35437 = n12888 & n35436 ;
  assign n35442 = n35441 ^ n35437 ^ 1'b0 ;
  assign n35443 = n1984 & ~n12308 ;
  assign n35444 = n35443 ^ n27863 ^ 1'b0 ;
  assign n35445 = n28757 ^ n25392 ^ n25229 ;
  assign n35446 = n35444 & n35445 ;
  assign n35447 = ~n22917 & n29589 ;
  assign n35448 = ( ~n4457 & n26871 ) | ( ~n4457 & n35447 ) | ( n26871 & n35447 ) ;
  assign n35449 = ( ~n10650 & n16694 ) | ( ~n10650 & n35448 ) | ( n16694 & n35448 ) ;
  assign n35450 = ( n650 & n16906 ) | ( n650 & ~n28067 ) | ( n16906 & ~n28067 ) ;
  assign n35451 = n35450 ^ n6013 ^ 1'b0 ;
  assign n35452 = n9211 & n35451 ;
  assign n35453 = ~n1158 & n21206 ;
  assign n35454 = n35453 ^ n3095 ^ 1'b0 ;
  assign n35455 = ~n11071 & n31424 ;
  assign n35456 = n35455 ^ n9010 ^ 1'b0 ;
  assign n35457 = n4102 & n26335 ;
  assign n35461 = n5624 ^ n1950 ^ 1'b0 ;
  assign n35460 = ( ~n5100 & n5222 ) | ( ~n5100 & n7703 ) | ( n5222 & n7703 ) ;
  assign n35458 = n3823 & ~n9808 ;
  assign n35459 = ~n19090 & n35458 ;
  assign n35462 = n35461 ^ n35460 ^ n35459 ;
  assign n35463 = ~n13518 & n21171 ;
  assign n35464 = n12757 ^ n6413 ^ 1'b0 ;
  assign n35465 = n30700 ^ n14492 ^ n8626 ;
  assign n35466 = n16818 | n35465 ;
  assign n35467 = n9130 & ~n35466 ;
  assign n35468 = n29773 ^ n15180 ^ 1'b0 ;
  assign n35469 = n698 | n35468 ;
  assign n35470 = ( n19505 & n23059 ) | ( n19505 & ~n25453 ) | ( n23059 & ~n25453 ) ;
  assign n35471 = n35470 ^ n18717 ^ n2980 ;
  assign n35472 = n8619 ^ n8337 ^ 1'b0 ;
  assign n35473 = ( n26308 & n30650 ) | ( n26308 & n35472 ) | ( n30650 & n35472 ) ;
  assign n35474 = n15477 ^ n10827 ^ n2665 ;
  assign n35475 = n35474 ^ n28452 ^ n23460 ;
  assign n35476 = n35475 ^ n16759 ^ 1'b0 ;
  assign n35477 = ( n20290 & ~n20977 ) | ( n20290 & n35476 ) | ( ~n20977 & n35476 ) ;
  assign n35478 = n12940 ^ n12023 ^ 1'b0 ;
  assign n35479 = n20015 & ~n31242 ;
  assign n35480 = n9124 | n10546 ;
  assign n35481 = n33193 ^ n31864 ^ n11453 ;
  assign n35482 = n32032 ^ n22900 ^ 1'b0 ;
  assign n35483 = n5049 & ~n35482 ;
  assign n35484 = n35483 ^ n700 ^ 1'b0 ;
  assign n35485 = ( n1566 & n9976 ) | ( n1566 & n22116 ) | ( n9976 & n22116 ) ;
  assign n35486 = ( n24985 & n28611 ) | ( n24985 & n35485 ) | ( n28611 & n35485 ) ;
  assign n35488 = n7710 & n11032 ;
  assign n35489 = n11279 & n35488 ;
  assign n35490 = n35489 ^ n9570 ^ n8760 ;
  assign n35487 = n15675 & n26940 ;
  assign n35491 = n35490 ^ n35487 ^ 1'b0 ;
  assign n35492 = n4062 ^ n1685 ^ 1'b0 ;
  assign n35493 = ( n16063 & n31793 ) | ( n16063 & ~n35492 ) | ( n31793 & ~n35492 ) ;
  assign n35494 = n12492 & ~n35493 ;
  assign n35495 = n15569 ^ n4279 ^ 1'b0 ;
  assign n35496 = ~n11498 & n35495 ;
  assign n35497 = n35496 ^ n21379 ^ 1'b0 ;
  assign n35498 = n35497 ^ n6866 ^ n2746 ;
  assign n35499 = n11718 ^ n6909 ^ n1660 ;
  assign n35503 = ( n3330 & ~n4028 ) | ( n3330 & n20592 ) | ( ~n4028 & n20592 ) ;
  assign n35500 = n3921 & n11760 ;
  assign n35501 = ~n4318 & n35500 ;
  assign n35502 = n20887 | n35501 ;
  assign n35504 = n35503 ^ n35502 ^ 1'b0 ;
  assign n35505 = ( ~n6417 & n18570 ) | ( ~n6417 & n35504 ) | ( n18570 & n35504 ) ;
  assign n35506 = ( n16352 & n29914 ) | ( n16352 & ~n35505 ) | ( n29914 & ~n35505 ) ;
  assign n35507 = n33989 ^ n32812 ^ n9458 ;
  assign n35508 = n6540 & n8985 ;
  assign n35509 = ~n8985 & n35508 ;
  assign n35510 = n17427 | n35509 ;
  assign n35511 = n17427 & ~n35510 ;
  assign n35512 = n35158 & ~n35511 ;
  assign n35513 = n35507 & n35512 ;
  assign n35514 = n12910 | n35513 ;
  assign n35515 = n35514 ^ n6598 ^ 1'b0 ;
  assign n35516 = n27051 & ~n35158 ;
  assign n35517 = n35447 ^ n14097 ^ 1'b0 ;
  assign n35518 = n7472 & ~n23034 ;
  assign n35519 = n444 & ~n31923 ;
  assign n35520 = n24396 & n35519 ;
  assign n35521 = ( n24291 & n27947 ) | ( n24291 & n35520 ) | ( n27947 & n35520 ) ;
  assign n35522 = n22301 ^ n4560 ^ 1'b0 ;
  assign n35523 = n2997 & ~n35522 ;
  assign n35526 = n12415 | n16584 ;
  assign n35527 = n35526 ^ n681 ^ 1'b0 ;
  assign n35524 = n14808 | n32717 ;
  assign n35525 = n35524 ^ n13040 ^ 1'b0 ;
  assign n35528 = n35527 ^ n35525 ^ n19290 ;
  assign n35529 = ( n4003 & n35523 ) | ( n4003 & ~n35528 ) | ( n35523 & ~n35528 ) ;
  assign n35530 = ( n19391 & ~n35521 ) | ( n19391 & n35529 ) | ( ~n35521 & n35529 ) ;
  assign n35531 = ( n8427 & n17924 ) | ( n8427 & ~n23704 ) | ( n17924 & ~n23704 ) ;
  assign n35532 = ( n4066 & n12024 ) | ( n4066 & ~n35531 ) | ( n12024 & ~n35531 ) ;
  assign n35533 = ( ~n3611 & n4240 ) | ( ~n3611 & n15212 ) | ( n4240 & n15212 ) ;
  assign n35534 = n35533 ^ n7969 ^ n7505 ;
  assign n35535 = n2177 | n35534 ;
  assign n35536 = n35532 & n35535 ;
  assign n35537 = n13459 & n35536 ;
  assign n35538 = n35537 ^ n17169 ^ n14628 ;
  assign n35541 = ( n4934 & ~n21152 ) | ( n4934 & n33771 ) | ( ~n21152 & n33771 ) ;
  assign n35542 = n8032 & n22896 ;
  assign n35543 = ~n35541 & n35542 ;
  assign n35539 = n6367 ^ n673 ^ 1'b0 ;
  assign n35540 = n5816 | n35539 ;
  assign n35544 = n35543 ^ n35540 ^ 1'b0 ;
  assign n35546 = n24155 ^ n8032 ^ n887 ;
  assign n35545 = n22564 & ~n29111 ;
  assign n35547 = n35546 ^ n35545 ^ 1'b0 ;
  assign n35548 = n17322 ^ n12313 ^ 1'b0 ;
  assign n35552 = n17023 ^ n17010 ^ n4466 ;
  assign n35549 = n19579 ^ n8625 ^ n2547 ;
  assign n35550 = n35549 ^ n20349 ^ 1'b0 ;
  assign n35551 = ~n18833 & n35550 ;
  assign n35553 = n35552 ^ n35551 ^ 1'b0 ;
  assign n35554 = n35548 | n35553 ;
  assign n35555 = n23796 ^ n13927 ^ 1'b0 ;
  assign n35556 = n35555 ^ n4823 ^ 1'b0 ;
  assign n35557 = n15788 & ~n35556 ;
  assign n35558 = n1900 & n8477 ;
  assign n35559 = n17305 ^ n12912 ^ n6646 ;
  assign n35560 = n3867 | n6683 ;
  assign n35561 = n35560 ^ n24662 ^ n15942 ;
  assign n35562 = n14304 ^ n5146 ^ 1'b0 ;
  assign n35563 = n35562 ^ n24986 ^ n22422 ;
  assign n35565 = n4751 ^ n2730 ^ n1522 ;
  assign n35564 = n10746 & ~n11260 ;
  assign n35566 = n35565 ^ n35564 ^ 1'b0 ;
  assign n35567 = ( n4404 & n7770 ) | ( n4404 & n9760 ) | ( n7770 & n9760 ) ;
  assign n35568 = n35567 ^ n21894 ^ 1'b0 ;
  assign n35569 = n7103 | n25435 ;
  assign n35570 = n35568 | n35569 ;
  assign n35571 = n9586 | n10943 ;
  assign n35572 = n17818 & ~n35571 ;
  assign n35573 = n35572 ^ n1997 ^ 1'b0 ;
  assign n35574 = n9648 & n35573 ;
  assign n35575 = n27745 ^ n24868 ^ n2943 ;
  assign n35576 = ( n613 & n1156 ) | ( n613 & ~n35575 ) | ( n1156 & ~n35575 ) ;
  assign n35577 = n22871 ^ n21317 ^ 1'b0 ;
  assign n35578 = n35577 ^ n19393 ^ n15273 ;
  assign n35579 = n34986 ^ n27600 ^ n3764 ;
  assign n35580 = n3627 & n8392 ;
  assign n35581 = n15258 & n35580 ;
  assign n35582 = ( n4256 & ~n12820 ) | ( n4256 & n35581 ) | ( ~n12820 & n35581 ) ;
  assign n35583 = n34114 ^ n4119 ^ 1'b0 ;
  assign n35584 = n35582 | n35583 ;
  assign n35585 = n7001 | n19378 ;
  assign n35586 = n35585 ^ n10090 ^ 1'b0 ;
  assign n35587 = n6460 & n35586 ;
  assign n35588 = n23920 ^ n19504 ^ n7003 ;
  assign n35589 = ~n19923 & n35588 ;
  assign n35590 = n35589 ^ n4810 ^ 1'b0 ;
  assign n35591 = ( n21833 & n29409 ) | ( n21833 & ~n31373 ) | ( n29409 & ~n31373 ) ;
  assign n35594 = n6843 ^ n2615 ^ n976 ;
  assign n35595 = ( ~n7410 & n26719 ) | ( ~n7410 & n35594 ) | ( n26719 & n35594 ) ;
  assign n35592 = n1108 & n27877 ;
  assign n35593 = ~n13713 & n35592 ;
  assign n35596 = n35595 ^ n35593 ^ 1'b0 ;
  assign n35597 = n21119 ^ n8632 ^ 1'b0 ;
  assign n35598 = ~n9069 & n35597 ;
  assign n35599 = ~n28087 & n35598 ;
  assign n35600 = x201 & ~n30486 ;
  assign n35601 = n3488 & n35600 ;
  assign n35602 = n13943 ^ n4986 ^ 1'b0 ;
  assign n35603 = n767 | n7642 ;
  assign n35604 = n1823 | n35603 ;
  assign n35605 = n35604 ^ n17148 ^ 1'b0 ;
  assign n35606 = n13536 | n35605 ;
  assign n35607 = n13207 ^ n5470 ^ 1'b0 ;
  assign n35608 = n35607 ^ n14471 ^ n4635 ;
  assign n35609 = n35608 ^ n23021 ^ n9220 ;
  assign n35610 = n20352 | n33443 ;
  assign n35611 = n5681 ^ n1263 ^ 1'b0 ;
  assign n35612 = n8161 & ~n35611 ;
  assign n35613 = n13650 ^ n2600 ^ 1'b0 ;
  assign n35614 = ~n18764 & n35613 ;
  assign n35616 = n6191 & ~n15372 ;
  assign n35617 = n22590 & n35616 ;
  assign n35615 = n20064 | n33573 ;
  assign n35618 = n35617 ^ n35615 ^ 1'b0 ;
  assign n35619 = n35614 & n35618 ;
  assign n35620 = n1266 & n15511 ;
  assign n35621 = n3509 & n35620 ;
  assign n35622 = n6169 & ~n10398 ;
  assign n35623 = n27000 ^ n17332 ^ n17218 ;
  assign n35624 = n3169 & n8896 ;
  assign n35625 = ~n9855 & n35624 ;
  assign n35626 = n24907 & ~n35625 ;
  assign n35627 = n14613 ^ n13042 ^ n2500 ;
  assign n35628 = n35627 ^ n7766 ^ n2821 ;
  assign n35629 = ( n15809 & n28941 ) | ( n15809 & ~n32432 ) | ( n28941 & ~n32432 ) ;
  assign n35630 = n14354 ^ n13021 ^ n3475 ;
  assign n35631 = n35630 ^ n20072 ^ 1'b0 ;
  assign n35632 = n9641 & n35631 ;
  assign n35633 = n3206 & n35632 ;
  assign n35634 = n35633 ^ n22846 ^ 1'b0 ;
  assign n35635 = n21642 ^ n3264 ^ n1445 ;
  assign n35636 = n5038 | n13578 ;
  assign n35637 = n35636 ^ n21321 ^ 1'b0 ;
  assign n35638 = n35635 | n35637 ;
  assign n35639 = n10813 | n23170 ;
  assign n35640 = ( n693 & n1281 ) | ( n693 & n14805 ) | ( n1281 & n14805 ) ;
  assign n35641 = n35640 ^ n35070 ^ n22167 ;
  assign n35642 = n6530 | n12540 ;
  assign n35643 = n35642 ^ n14247 ^ 1'b0 ;
  assign n35644 = n35643 ^ n11874 ^ n10542 ;
  assign n35645 = n18295 ^ n5324 ^ 1'b0 ;
  assign n35646 = n4066 | n16675 ;
  assign n35647 = ( n14694 & ~n19989 ) | ( n14694 & n35646 ) | ( ~n19989 & n35646 ) ;
  assign n35648 = n28775 ^ n13027 ^ n7213 ;
  assign n35649 = ( n10584 & n28800 ) | ( n10584 & n35648 ) | ( n28800 & n35648 ) ;
  assign n35650 = ( n12093 & ~n29389 ) | ( n12093 & n35649 ) | ( ~n29389 & n35649 ) ;
  assign n35651 = n12309 ^ n3507 ^ n868 ;
  assign n35652 = n2215 | n35651 ;
  assign n35653 = ~n15643 & n35652 ;
  assign n35654 = n13864 & n15457 ;
  assign n35655 = n35654 ^ n4465 ^ 1'b0 ;
  assign n35656 = n16788 ^ n2417 ^ 1'b0 ;
  assign n35657 = n21950 & n35656 ;
  assign n35658 = n35657 ^ n4868 ^ 1'b0 ;
  assign n35659 = n22012 | n35658 ;
  assign n35660 = n35659 ^ n7639 ^ 1'b0 ;
  assign n35661 = n16461 ^ n1775 ^ 1'b0 ;
  assign n35662 = ~n8588 & n35661 ;
  assign n35663 = n22343 ^ n1681 ^ 1'b0 ;
  assign n35664 = n2086 & ~n35663 ;
  assign n35665 = n35664 ^ n24182 ^ 1'b0 ;
  assign n35666 = n35662 & ~n35665 ;
  assign n35667 = ~n21753 & n24791 ;
  assign n35668 = ~n2476 & n2798 ;
  assign n35669 = ~n2798 & n35668 ;
  assign n35670 = n22631 & ~n35669 ;
  assign n35671 = n5035 & ~n6190 ;
  assign n35672 = ~n5035 & n35671 ;
  assign n35673 = n1672 & ~n4242 ;
  assign n35674 = n35672 & n35673 ;
  assign n35675 = n11498 | n35674 ;
  assign n35676 = n8183 ^ n4566 ^ 1'b0 ;
  assign n35677 = ~n35675 & n35676 ;
  assign n35678 = ~n35670 & n35677 ;
  assign n35679 = n35678 ^ n28685 ^ 1'b0 ;
  assign n35680 = n11913 ^ n11357 ^ n9258 ;
  assign n35684 = ( n18670 & n23783 ) | ( n18670 & ~n24487 ) | ( n23783 & ~n24487 ) ;
  assign n35681 = x202 & n4653 ;
  assign n35682 = n35681 ^ n9111 ^ 1'b0 ;
  assign n35683 = n16334 & n35682 ;
  assign n35685 = n35684 ^ n35683 ^ 1'b0 ;
  assign n35686 = n5538 ^ n4714 ^ 1'b0 ;
  assign n35687 = ~n13573 & n35686 ;
  assign n35688 = ~n3440 & n35687 ;
  assign n35689 = n35688 ^ n18317 ^ 1'b0 ;
  assign n35690 = n28970 ^ n18668 ^ 1'b0 ;
  assign n35691 = n9966 & n35690 ;
  assign n35692 = ( x146 & n11407 ) | ( x146 & ~n35691 ) | ( n11407 & ~n35691 ) ;
  assign n35693 = n3384 | n35692 ;
  assign n35694 = n35693 ^ n29921 ^ n2781 ;
  assign n35695 = n8078 & n35694 ;
  assign n35696 = n35689 & n35695 ;
  assign n35698 = n5066 & ~n6599 ;
  assign n35697 = n2748 | n11356 ;
  assign n35699 = n35698 ^ n35697 ^ 1'b0 ;
  assign n35700 = n5014 ^ n3061 ^ 1'b0 ;
  assign n35701 = n28481 ^ n18143 ^ n14016 ;
  assign n35702 = n23567 & n35701 ;
  assign n35703 = n35702 ^ n19953 ^ 1'b0 ;
  assign n35704 = x121 & n1133 ;
  assign n35705 = ~n1824 & n35704 ;
  assign n35706 = ( n305 & n3772 ) | ( n305 & ~n5980 ) | ( n3772 & ~n5980 ) ;
  assign n35707 = n2999 & ~n8358 ;
  assign n35708 = ~n35706 & n35707 ;
  assign n35709 = ( n33291 & n35705 ) | ( n33291 & ~n35708 ) | ( n35705 & ~n35708 ) ;
  assign n35712 = n19624 ^ n10621 ^ 1'b0 ;
  assign n35713 = ~n15947 & n35712 ;
  assign n35710 = ~n4144 & n28087 ;
  assign n35711 = n24538 & n35710 ;
  assign n35714 = n35713 ^ n35711 ^ n12485 ;
  assign n35716 = n33196 ^ n3060 ^ 1'b0 ;
  assign n35717 = n8298 & ~n35716 ;
  assign n35718 = ( n18265 & n19858 ) | ( n18265 & n35717 ) | ( n19858 & n35717 ) ;
  assign n35715 = n29931 ^ n19386 ^ 1'b0 ;
  assign n35719 = n35718 ^ n35715 ^ 1'b0 ;
  assign n35720 = n8296 ^ n3156 ^ 1'b0 ;
  assign n35721 = ~n29197 & n35720 ;
  assign n35722 = n24396 ^ n21029 ^ n17980 ;
  assign n35724 = n8662 | n17671 ;
  assign n35725 = ~n10125 & n35724 ;
  assign n35726 = n35725 ^ n9046 ^ 1'b0 ;
  assign n35723 = n13720 & ~n29060 ;
  assign n35727 = n35726 ^ n35723 ^ 1'b0 ;
  assign n35728 = ~n8156 & n35727 ;
  assign n35729 = n35728 ^ n7296 ^ 1'b0 ;
  assign n35730 = n20374 ^ n6048 ^ n3275 ;
  assign n35731 = ( n4332 & n7724 ) | ( n4332 & ~n28287 ) | ( n7724 & ~n28287 ) ;
  assign n35732 = ~n10591 & n35731 ;
  assign n35733 = n35732 ^ n28941 ^ 1'b0 ;
  assign n35734 = x45 & n12931 ;
  assign n35735 = ~n11826 & n35734 ;
  assign n35736 = n25683 ^ n10406 ^ 1'b0 ;
  assign n35737 = n26417 & ~n35736 ;
  assign n35740 = n8706 & n9644 ;
  assign n35738 = n17657 | n24488 ;
  assign n35739 = n35738 ^ n27740 ^ n21855 ;
  assign n35741 = n35740 ^ n35739 ^ 1'b0 ;
  assign n35748 = n9365 & n18037 ;
  assign n35749 = n35748 ^ n20516 ^ n1754 ;
  assign n35742 = n11940 ^ n7178 ^ 1'b0 ;
  assign n35743 = n13946 & n35742 ;
  assign n35744 = n14542 & n21011 ;
  assign n35745 = ~n5895 & n35744 ;
  assign n35746 = n35743 & ~n35745 ;
  assign n35747 = n35746 ^ n15058 ^ 1'b0 ;
  assign n35750 = n35749 ^ n35747 ^ n3177 ;
  assign n35751 = n24033 ^ n9908 ^ n5787 ;
  assign n35752 = ( n26708 & n31403 ) | ( n26708 & n35751 ) | ( n31403 & n35751 ) ;
  assign n35753 = n35752 ^ n9416 ^ 1'b0 ;
  assign n35754 = n25316 ^ n12013 ^ n2377 ;
  assign n35755 = ( ~n12996 & n20860 ) | ( ~n12996 & n35754 ) | ( n20860 & n35754 ) ;
  assign n35756 = n5430 & ~n14956 ;
  assign n35757 = n15828 & n35756 ;
  assign n35758 = n9450 | n22514 ;
  assign n35759 = n35758 ^ n22034 ^ 1'b0 ;
  assign n35760 = n35292 ^ n32197 ^ n16608 ;
  assign n35761 = n19688 ^ n14047 ^ n974 ;
  assign n35762 = ( n8758 & n22647 ) | ( n8758 & n33361 ) | ( n22647 & n33361 ) ;
  assign n35763 = ( n1192 & n12027 ) | ( n1192 & ~n14457 ) | ( n12027 & ~n14457 ) ;
  assign n35764 = n12707 | n35763 ;
  assign n35765 = n1537 | n26153 ;
  assign n35766 = n12767 & ~n23660 ;
  assign n35767 = ~n16681 & n35766 ;
  assign n35768 = n19084 | n25805 ;
  assign n35769 = n35768 ^ n18314 ^ 1'b0 ;
  assign n35770 = x63 & n9312 ;
  assign n35771 = n35770 ^ n8134 ^ 1'b0 ;
  assign n35772 = n812 | n35771 ;
  assign n35773 = n26693 | n35772 ;
  assign n35774 = ( n2338 & n25441 ) | ( n2338 & ~n35773 ) | ( n25441 & ~n35773 ) ;
  assign n35775 = ( n9236 & ~n30081 ) | ( n9236 & n31291 ) | ( ~n30081 & n31291 ) ;
  assign n35776 = n30749 | n35775 ;
  assign n35777 = ( n5589 & n12741 ) | ( n5589 & ~n16234 ) | ( n12741 & ~n16234 ) ;
  assign n35778 = n7196 | n12910 ;
  assign n35779 = n35778 ^ n22471 ^ n11368 ;
  assign n35780 = ( n24859 & n34226 ) | ( n24859 & n35779 ) | ( n34226 & n35779 ) ;
  assign n35781 = ( ~n35739 & n35777 ) | ( ~n35739 & n35780 ) | ( n35777 & n35780 ) ;
  assign n35782 = n19743 & n35471 ;
  assign n35783 = n30723 ^ n21898 ^ n2839 ;
  assign n35784 = n7058 | n35783 ;
  assign n35785 = n3759 ^ n3238 ^ 1'b0 ;
  assign n35786 = n9595 & n35785 ;
  assign n35787 = n35786 ^ n13335 ^ 1'b0 ;
  assign n35788 = n1989 & ~n35787 ;
  assign n35789 = n698 | n11050 ;
  assign n35790 = n35788 | n35789 ;
  assign n35791 = ( n3317 & ~n8265 ) | ( n3317 & n28936 ) | ( ~n8265 & n28936 ) ;
  assign n35792 = n33687 ^ n31295 ^ n2743 ;
  assign n35793 = ( n1934 & ~n2628 ) | ( n1934 & n32796 ) | ( ~n2628 & n32796 ) ;
  assign n35794 = ( ~n1125 & n1627 ) | ( ~n1125 & n2324 ) | ( n1627 & n2324 ) ;
  assign n35795 = n9397 | n35794 ;
  assign n35796 = n25637 ^ n10045 ^ n8605 ;
  assign n35797 = n27295 & ~n35796 ;
  assign n35798 = n35797 ^ n16895 ^ 1'b0 ;
  assign n35799 = n2287 & ~n22186 ;
  assign n35800 = n35799 ^ n31152 ^ 1'b0 ;
  assign n35801 = n8330 & n31320 ;
  assign n35802 = ( n1666 & n35800 ) | ( n1666 & n35801 ) | ( n35800 & n35801 ) ;
  assign n35803 = n34729 ^ n19198 ^ n5177 ;
  assign n35804 = ( n4471 & n16489 ) | ( n4471 & n17970 ) | ( n16489 & n17970 ) ;
  assign n35805 = n13324 & n14992 ;
  assign n35806 = n35805 ^ n10410 ^ 1'b0 ;
  assign n35807 = n7665 & n34014 ;
  assign n35808 = n20814 & n35807 ;
  assign n35809 = n8411 & n14207 ;
  assign n35810 = ( n21278 & ~n25487 ) | ( n21278 & n31577 ) | ( ~n25487 & n31577 ) ;
  assign n35811 = ( n804 & n35809 ) | ( n804 & ~n35810 ) | ( n35809 & ~n35810 ) ;
  assign n35812 = n20453 ^ n8033 ^ 1'b0 ;
  assign n35813 = n21583 & n35812 ;
  assign n35814 = ( x220 & n30778 ) | ( x220 & ~n35813 ) | ( n30778 & ~n35813 ) ;
  assign n35816 = ~n4061 & n15588 ;
  assign n35815 = ( n2149 & n2851 ) | ( n2149 & n20476 ) | ( n2851 & n20476 ) ;
  assign n35817 = n35816 ^ n35815 ^ 1'b0 ;
  assign n35818 = ( n6367 & n15044 ) | ( n6367 & n31541 ) | ( n15044 & n31541 ) ;
  assign n35819 = n18527 | n29580 ;
  assign n35820 = n35819 ^ n3697 ^ 1'b0 ;
  assign n35821 = n9894 | n35820 ;
  assign n35822 = n17463 & ~n35821 ;
  assign n35823 = n35822 ^ n12580 ^ 1'b0 ;
  assign n35824 = n3769 ^ n2777 ^ 1'b0 ;
  assign n35825 = n1093 & n35824 ;
  assign n35826 = n22977 | n33570 ;
  assign n35827 = n35826 ^ n31904 ^ 1'b0 ;
  assign n35828 = n8315 | n8676 ;
  assign n35829 = n380 & n3466 ;
  assign n35830 = ( n16751 & n30845 ) | ( n16751 & n35829 ) | ( n30845 & n35829 ) ;
  assign n35831 = n35830 ^ n6092 ^ n5091 ;
  assign n35832 = n35831 ^ n23363 ^ 1'b0 ;
  assign n35833 = ( ~n880 & n15057 ) | ( ~n880 & n15571 ) | ( n15057 & n15571 ) ;
  assign n35834 = ( n12180 & ~n31401 ) | ( n12180 & n35833 ) | ( ~n31401 & n35833 ) ;
  assign n35835 = n9875 | n12538 ;
  assign n35836 = n1494 & ~n35835 ;
  assign n35837 = n553 & ~n35836 ;
  assign n35838 = n25690 ^ n6414 ^ 1'b0 ;
  assign n35839 = ( n13356 & n35837 ) | ( n13356 & n35838 ) | ( n35837 & n35838 ) ;
  assign n35840 = n30689 ^ n14341 ^ 1'b0 ;
  assign n35841 = n18127 & n25833 ;
  assign n35842 = n4045 & n35841 ;
  assign n35843 = n35842 ^ n9635 ^ 1'b0 ;
  assign n35844 = n13205 & n35843 ;
  assign n35845 = n17256 & ~n21838 ;
  assign n35846 = n19303 ^ n15116 ^ 1'b0 ;
  assign n35847 = n1374 | n35846 ;
  assign n35848 = n35847 ^ n16721 ^ 1'b0 ;
  assign n35849 = n1345 | n26119 ;
  assign n35850 = n9009 | n35849 ;
  assign n35851 = n35850 ^ n5791 ^ n2653 ;
  assign n35852 = n14849 ^ n6853 ^ n704 ;
  assign n35853 = n15595 ^ n1870 ^ 1'b0 ;
  assign n35857 = n10481 | n18680 ;
  assign n35858 = n35857 ^ n16964 ^ 1'b0 ;
  assign n35854 = n21236 & ~n30102 ;
  assign n35855 = n35854 ^ n7206 ^ 1'b0 ;
  assign n35856 = n15486 & ~n35855 ;
  assign n35859 = n35858 ^ n35856 ^ 1'b0 ;
  assign n35860 = ( n20780 & ~n35853 ) | ( n20780 & n35859 ) | ( ~n35853 & n35859 ) ;
  assign n35864 = n26911 ^ n24089 ^ n7817 ;
  assign n35865 = n24547 ^ n21333 ^ 1'b0 ;
  assign n35866 = ~n35864 & n35865 ;
  assign n35861 = n4388 & ~n7808 ;
  assign n35862 = n35861 ^ x158 ^ 1'b0 ;
  assign n35863 = n24505 & ~n35862 ;
  assign n35867 = n35866 ^ n35863 ^ 1'b0 ;
  assign n35868 = ( n605 & ~n5716 ) | ( n605 & n7927 ) | ( ~n5716 & n7927 ) ;
  assign n35869 = n35868 ^ n15919 ^ n3765 ;
  assign n35870 = ( n2557 & n5116 ) | ( n2557 & ~n35869 ) | ( n5116 & ~n35869 ) ;
  assign n35871 = n9756 | n35870 ;
  assign n35872 = n20336 ^ n18292 ^ n16743 ;
  assign n35873 = n17134 | n24716 ;
  assign n35876 = n32721 ^ n12350 ^ 1'b0 ;
  assign n35877 = n4072 & n35876 ;
  assign n35874 = n10494 | n10952 ;
  assign n35875 = n35874 ^ n16656 ^ 1'b0 ;
  assign n35878 = n35877 ^ n35875 ^ 1'b0 ;
  assign n35879 = n6379 ^ n1457 ^ 1'b0 ;
  assign n35880 = n4232 | n17933 ;
  assign n35881 = n35880 ^ n7781 ^ 1'b0 ;
  assign n35882 = n12477 ^ n5315 ^ 1'b0 ;
  assign n35883 = n35881 & ~n35882 ;
  assign n35884 = n35883 ^ n27181 ^ n21810 ;
  assign n35885 = ~n16526 & n20433 ;
  assign n35886 = ( n27063 & n28770 ) | ( n27063 & ~n35885 ) | ( n28770 & ~n35885 ) ;
  assign n35887 = ( ~n1312 & n7473 ) | ( ~n1312 & n20042 ) | ( n7473 & n20042 ) ;
  assign n35888 = ~n11814 & n11945 ;
  assign n35889 = n35888 ^ n19297 ^ n11850 ;
  assign n35890 = n3512 | n15720 ;
  assign n35891 = n12713 & ~n20816 ;
  assign n35894 = n8227 & n24992 ;
  assign n35892 = ( n593 & ~n7363 ) | ( n593 & n26323 ) | ( ~n7363 & n26323 ) ;
  assign n35893 = n10060 & ~n35892 ;
  assign n35895 = n35894 ^ n35893 ^ 1'b0 ;
  assign n35896 = ( n3996 & ~n4866 ) | ( n3996 & n8279 ) | ( ~n4866 & n8279 ) ;
  assign n35897 = n871 & n17461 ;
  assign n35898 = ~n4318 & n35897 ;
  assign n35899 = n35898 ^ n6430 ^ 1'b0 ;
  assign n35900 = n11493 & ~n35899 ;
  assign n35901 = n15308 & ~n26732 ;
  assign n35902 = ~n35900 & n35901 ;
  assign n35903 = n35902 ^ n6763 ^ 1'b0 ;
  assign n35904 = n35896 & n35903 ;
  assign n35905 = n35904 ^ n6722 ^ n6311 ;
  assign n35906 = n23458 ^ n8605 ^ 1'b0 ;
  assign n35907 = ( ~n5816 & n16977 ) | ( ~n5816 & n26736 ) | ( n16977 & n26736 ) ;
  assign n35908 = ( n22807 & ~n34365 ) | ( n22807 & n35907 ) | ( ~n34365 & n35907 ) ;
  assign n35909 = ( n10835 & n35906 ) | ( n10835 & ~n35908 ) | ( n35906 & ~n35908 ) ;
  assign n35910 = n23163 ^ n19649 ^ 1'b0 ;
  assign n35912 = n27673 ^ n1775 ^ 1'b0 ;
  assign n35913 = n13043 | n35912 ;
  assign n35914 = n35913 ^ n18776 ^ n8403 ;
  assign n35911 = ~n609 & n30481 ;
  assign n35915 = n35914 ^ n35911 ^ 1'b0 ;
  assign n35916 = n10133 | n22310 ;
  assign n35917 = n29595 & n35916 ;
  assign n35918 = ~n2284 & n35917 ;
  assign n35919 = ( n10325 & n21823 ) | ( n10325 & n26183 ) | ( n21823 & n26183 ) ;
  assign n35920 = ( n5185 & n8393 ) | ( n5185 & ~n24555 ) | ( n8393 & ~n24555 ) ;
  assign n35921 = n27333 & n35920 ;
  assign n35922 = n35921 ^ n20164 ^ 1'b0 ;
  assign n35923 = n35922 ^ n4566 ^ 1'b0 ;
  assign n35924 = n35919 & n35923 ;
  assign n35925 = ~n5092 & n14062 ;
  assign n35926 = ~n423 & n33973 ;
  assign n35927 = n24894 ^ n13468 ^ 1'b0 ;
  assign n35928 = ( n5105 & ~n34730 ) | ( n5105 & n35927 ) | ( ~n34730 & n35927 ) ;
  assign n35929 = ( ~n12026 & n22117 ) | ( ~n12026 & n35928 ) | ( n22117 & n35928 ) ;
  assign n35930 = ~n1776 & n25251 ;
  assign n35931 = n35930 ^ n20595 ^ 1'b0 ;
  assign n35932 = n35931 ^ n5474 ^ n428 ;
  assign n35940 = n14870 ^ n11490 ^ n2013 ;
  assign n35935 = ( x50 & ~n3034 ) | ( x50 & n15912 ) | ( ~n3034 & n15912 ) ;
  assign n35936 = n35935 ^ n31161 ^ n767 ;
  assign n35937 = n16858 & n35936 ;
  assign n35938 = n2536 & n35937 ;
  assign n35939 = n6960 | n35938 ;
  assign n35941 = n35940 ^ n35939 ^ 1'b0 ;
  assign n35933 = n13131 ^ n2867 ^ 1'b0 ;
  assign n35934 = n5947 & n35933 ;
  assign n35942 = n35941 ^ n35934 ^ n34049 ;
  assign n35943 = n3791 & n8691 ;
  assign n35944 = ~n15462 & n35943 ;
  assign n35945 = ( n18217 & n18889 ) | ( n18217 & n35944 ) | ( n18889 & n35944 ) ;
  assign n35946 = ( n25882 & n28589 ) | ( n25882 & n35945 ) | ( n28589 & n35945 ) ;
  assign n35947 = n35946 ^ n13401 ^ 1'b0 ;
  assign n35948 = n10370 ^ n750 ^ 1'b0 ;
  assign n35949 = ( ~n2406 & n22094 ) | ( ~n2406 & n35948 ) | ( n22094 & n35948 ) ;
  assign n35950 = ~n10478 & n35949 ;
  assign n35951 = n35950 ^ n27457 ^ 1'b0 ;
  assign n35952 = n15994 & n28778 ;
  assign n35953 = ( n6021 & n17566 ) | ( n6021 & n31519 ) | ( n17566 & n31519 ) ;
  assign n35954 = n10307 & ~n21231 ;
  assign n35955 = n23946 ^ n11594 ^ n2076 ;
  assign n35956 = ~n35954 & n35955 ;
  assign n35957 = ( n18530 & n18847 ) | ( n18530 & ~n23129 ) | ( n18847 & ~n23129 ) ;
  assign n35958 = n16237 ^ n12478 ^ n3248 ;
  assign n35959 = n35958 ^ n13197 ^ 1'b0 ;
  assign n35960 = n16955 & n35959 ;
  assign n35961 = ~n35957 & n35960 ;
  assign n35962 = n11959 & n18447 ;
  assign n35963 = ( n15283 & n25460 ) | ( n15283 & n25689 ) | ( n25460 & n25689 ) ;
  assign n35964 = n8552 & n13364 ;
  assign n35965 = n35964 ^ n6216 ^ 1'b0 ;
  assign n35966 = n30010 ^ n26852 ^ n7163 ;
  assign n35967 = n33391 & ~n35966 ;
  assign n35968 = n35967 ^ n35154 ^ 1'b0 ;
  assign n35969 = ~n13670 & n22599 ;
  assign n35970 = ~n1585 & n35969 ;
  assign n35971 = n2400 & n4758 ;
  assign n35975 = ( n7679 & ~n20609 ) | ( n7679 & n27446 ) | ( ~n20609 & n27446 ) ;
  assign n35974 = n7767 ^ n6352 ^ n1827 ;
  assign n35972 = ( n9769 & n9777 ) | ( n9769 & ~n21464 ) | ( n9777 & ~n21464 ) ;
  assign n35973 = n35972 ^ n3247 ^ 1'b0 ;
  assign n35976 = n35975 ^ n35974 ^ n35973 ;
  assign n35977 = ~n25108 & n34070 ;
  assign n35978 = n29268 & n35977 ;
  assign n35982 = n1385 & n6881 ;
  assign n35981 = n30046 ^ n12337 ^ n10721 ;
  assign n35979 = x231 & n8549 ;
  assign n35980 = ( n6090 & n23045 ) | ( n6090 & ~n35979 ) | ( n23045 & ~n35979 ) ;
  assign n35983 = n35982 ^ n35981 ^ n35980 ;
  assign n35984 = n6433 ^ n2461 ^ 1'b0 ;
  assign n35985 = n668 & n17002 ;
  assign n35986 = n35985 ^ n17520 ^ 1'b0 ;
  assign n35987 = ~n1888 & n4152 ;
  assign n35988 = n20741 & n35987 ;
  assign n35994 = ~n4340 & n7470 ;
  assign n35990 = n13674 ^ n10966 ^ 1'b0 ;
  assign n35989 = n3571 | n22899 ;
  assign n35991 = n35990 ^ n35989 ^ 1'b0 ;
  assign n35992 = n10755 | n35991 ;
  assign n35993 = n10267 & ~n35992 ;
  assign n35995 = n35994 ^ n35993 ^ 1'b0 ;
  assign n35996 = n12439 ^ n5129 ^ 1'b0 ;
  assign n35997 = n32468 ^ n8651 ^ 1'b0 ;
  assign n35998 = n30143 & n35997 ;
  assign n35999 = n7968 | n34997 ;
  assign n36000 = n35999 ^ n7674 ^ 1'b0 ;
  assign n36001 = n7345 & n14530 ;
  assign n36002 = n36001 ^ n9562 ^ 1'b0 ;
  assign n36003 = n10144 | n27561 ;
  assign n36004 = n34320 | n36003 ;
  assign n36005 = n23486 & ~n32320 ;
  assign n36006 = n15319 ^ n12317 ^ n5445 ;
  assign n36007 = n22322 & n36006 ;
  assign n36008 = ( n22767 & n24186 ) | ( n22767 & n36007 ) | ( n24186 & n36007 ) ;
  assign n36010 = n11295 & n13363 ;
  assign n36009 = n32183 ^ n3663 ^ 1'b0 ;
  assign n36011 = n36010 ^ n36009 ^ n7158 ;
  assign n36012 = n27236 ^ n17517 ^ n7914 ;
  assign n36013 = n33246 & ~n36012 ;
  assign n36014 = n36013 ^ n17009 ^ 1'b0 ;
  assign n36015 = n13166 ^ n564 ^ 1'b0 ;
  assign n36016 = n7373 & n36015 ;
  assign n36017 = n8234 ^ n6858 ^ 1'b0 ;
  assign n36018 = n36016 & ~n36017 ;
  assign n36019 = n2430 & n13712 ;
  assign n36020 = n36019 ^ n26128 ^ 1'b0 ;
  assign n36021 = n32908 ^ n18302 ^ 1'b0 ;
  assign n36022 = ~n6856 & n8047 ;
  assign n36023 = ~n490 & n36022 ;
  assign n36024 = n7579 & ~n36023 ;
  assign n36025 = ~n36021 & n36024 ;
  assign n36026 = n36025 ^ n10759 ^ n9242 ;
  assign n36027 = n1278 | n36026 ;
  assign n36028 = n36027 ^ n31683 ^ 1'b0 ;
  assign n36029 = n28188 ^ n17673 ^ n14401 ;
  assign n36030 = ~n11289 & n15641 ;
  assign n36031 = n36029 | n36030 ;
  assign n36032 = n12454 & ~n12566 ;
  assign n36033 = ( n17148 & ~n26886 ) | ( n17148 & n36032 ) | ( ~n26886 & n36032 ) ;
  assign n36034 = n6267 & ~n31703 ;
  assign n36035 = n36034 ^ n13454 ^ 1'b0 ;
  assign n36036 = n295 & n36035 ;
  assign n36037 = ~n36033 & n36036 ;
  assign n36038 = n20602 | n36037 ;
  assign n36039 = n10903 ^ n7475 ^ n3763 ;
  assign n36040 = n7126 & n32655 ;
  assign n36041 = n7138 & n36040 ;
  assign n36042 = n36041 ^ n18651 ^ 1'b0 ;
  assign n36043 = n29713 ^ n19565 ^ n16826 ;
  assign n36044 = n36043 ^ n16751 ^ 1'b0 ;
  assign n36045 = ~n26368 & n29514 ;
  assign n36046 = ~n6895 & n36045 ;
  assign n36047 = n31966 ^ n27740 ^ 1'b0 ;
  assign n36048 = n30221 & n33875 ;
  assign n36049 = ~n2642 & n36048 ;
  assign n36050 = n30195 ^ n6856 ^ 1'b0 ;
  assign n36051 = ~n36049 & n36050 ;
  assign n36052 = ~n36047 & n36051 ;
  assign n36053 = ( n5063 & n18963 ) | ( n5063 & ~n29792 ) | ( n18963 & ~n29792 ) ;
  assign n36054 = n16333 ^ n9139 ^ n6211 ;
  assign n36055 = n19167 | n30664 ;
  assign n36056 = n19628 | n36055 ;
  assign n36057 = ~n26982 & n36056 ;
  assign n36058 = n36057 ^ n28740 ^ 1'b0 ;
  assign n36059 = ~n15991 & n17014 ;
  assign n36060 = n12274 ^ n7375 ^ 1'b0 ;
  assign n36061 = ~n36059 & n36060 ;
  assign n36062 = n36061 ^ n20060 ^ 1'b0 ;
  assign n36063 = n27015 | n36062 ;
  assign n36064 = n22162 ^ n22031 ^ 1'b0 ;
  assign n36065 = n5500 & n34165 ;
  assign n36066 = n36065 ^ n26289 ^ 1'b0 ;
  assign n36067 = n1252 & ~n36066 ;
  assign n36068 = ( n22726 & ~n29915 ) | ( n22726 & n36067 ) | ( ~n29915 & n36067 ) ;
  assign n36069 = n24120 ^ n10690 ^ 1'b0 ;
  assign n36070 = ~n8541 & n36069 ;
  assign n36071 = ( n15469 & n33030 ) | ( n15469 & n36070 ) | ( n33030 & n36070 ) ;
  assign n36072 = n36071 ^ n35005 ^ n9165 ;
  assign n36073 = n17524 ^ n14852 ^ n12125 ;
  assign n36074 = ~n2564 & n8368 ;
  assign n36075 = ~n1524 & n36074 ;
  assign n36076 = ~n7036 & n36075 ;
  assign n36077 = ( n21079 & ~n36073 ) | ( n21079 & n36076 ) | ( ~n36073 & n36076 ) ;
  assign n36081 = n7549 ^ n1757 ^ n787 ;
  assign n36079 = ( n7627 & n27799 ) | ( n7627 & ~n31496 ) | ( n27799 & ~n31496 ) ;
  assign n36078 = n2337 & ~n23932 ;
  assign n36080 = n36079 ^ n36078 ^ n1434 ;
  assign n36082 = n36081 ^ n36080 ^ 1'b0 ;
  assign n36083 = n36077 & n36082 ;
  assign n36084 = n36083 ^ n10843 ^ 1'b0 ;
  assign n36085 = ( ~n8307 & n23332 ) | ( ~n8307 & n29195 ) | ( n23332 & n29195 ) ;
  assign n36086 = n33976 ^ n24572 ^ 1'b0 ;
  assign n36087 = n36085 & ~n36086 ;
  assign n36088 = n27679 ^ n22943 ^ n18680 ;
  assign n36089 = n24793 ^ n18216 ^ 1'b0 ;
  assign n36090 = ~n16643 & n36089 ;
  assign n36091 = ( n15746 & n20042 ) | ( n15746 & ~n28334 ) | ( n20042 & ~n28334 ) ;
  assign n36092 = n15005 ^ n11893 ^ 1'b0 ;
  assign n36093 = n24890 ^ n13275 ^ n1022 ;
  assign n36094 = ( ~n1148 & n15566 ) | ( ~n1148 & n17134 ) | ( n15566 & n17134 ) ;
  assign n36095 = ~n4848 & n16927 ;
  assign n36096 = n6815 & n34229 ;
  assign n36097 = n36095 & n36096 ;
  assign n36098 = n36097 ^ n28601 ^ n8183 ;
  assign n36099 = ( x204 & ~n287 ) | ( x204 & n14074 ) | ( ~n287 & n14074 ) ;
  assign n36100 = n36099 ^ n16585 ^ 1'b0 ;
  assign n36101 = n2014 & ~n16330 ;
  assign n36102 = ( n13156 & n19206 ) | ( n13156 & n36101 ) | ( n19206 & n36101 ) ;
  assign n36103 = n2502 & ~n12093 ;
  assign n36104 = n36102 & n36103 ;
  assign n36105 = ~n24383 & n30704 ;
  assign n36106 = n19233 ^ n3018 ^ n2262 ;
  assign n36107 = n12123 | n34380 ;
  assign n36108 = n36107 ^ n16230 ^ 1'b0 ;
  assign n36109 = n36108 ^ n15734 ^ 1'b0 ;
  assign n36110 = n20315 ^ n18262 ^ 1'b0 ;
  assign n36111 = n25925 & n36110 ;
  assign n36112 = n2497 | n9969 ;
  assign n36113 = n21569 & ~n36112 ;
  assign n36114 = n22649 ^ n7708 ^ n7015 ;
  assign n36115 = n14375 ^ n6798 ^ 1'b0 ;
  assign n36116 = n14120 & ~n36115 ;
  assign n36117 = ~n36114 & n36116 ;
  assign n36118 = n36117 ^ n28847 ^ n8558 ;
  assign n36120 = n5716 & ~n29511 ;
  assign n36121 = n13027 & n36120 ;
  assign n36119 = ~n16731 & n34983 ;
  assign n36122 = n36121 ^ n36119 ^ n33937 ;
  assign n36123 = n14683 ^ n5310 ^ 1'b0 ;
  assign n36124 = ( ~n30374 & n34967 ) | ( ~n30374 & n36123 ) | ( n34967 & n36123 ) ;
  assign n36125 = n34359 ^ n7004 ^ n3566 ;
  assign n36126 = n19235 ^ n16410 ^ 1'b0 ;
  assign n36127 = ~n19265 & n36126 ;
  assign n36128 = n18393 & n19560 ;
  assign n36129 = ~n1576 & n36128 ;
  assign n36130 = ( n1068 & n8194 ) | ( n1068 & ~n17255 ) | ( n8194 & ~n17255 ) ;
  assign n36131 = n36130 ^ n14183 ^ 1'b0 ;
  assign n36132 = ~n21573 & n36131 ;
  assign n36133 = ~n9089 & n9500 ;
  assign n36134 = ~n10993 & n36133 ;
  assign n36135 = ~n11252 & n17527 ;
  assign n36136 = n36135 ^ n14061 ^ 1'b0 ;
  assign n36137 = n12493 & n25361 ;
  assign n36138 = n7343 & ~n27576 ;
  assign n36139 = x98 | n11687 ;
  assign n36140 = n36139 ^ n16481 ^ 1'b0 ;
  assign n36141 = n25459 & n36140 ;
  assign n36143 = n16960 | n20193 ;
  assign n36144 = n36143 ^ n29156 ^ 1'b0 ;
  assign n36142 = n11190 & ~n30122 ;
  assign n36145 = n36144 ^ n36142 ^ 1'b0 ;
  assign n36146 = n10017 ^ n8726 ^ 1'b0 ;
  assign n36147 = n36146 ^ n35993 ^ n13869 ;
  assign n36148 = ( n629 & n20689 ) | ( n629 & n22475 ) | ( n20689 & n22475 ) ;
  assign n36149 = n36148 ^ n28565 ^ n15784 ;
  assign n36150 = ( n17350 & n25516 ) | ( n17350 & ~n31972 ) | ( n25516 & ~n31972 ) ;
  assign n36151 = n4142 ^ n2476 ^ n700 ;
  assign n36152 = ( n19255 & n26556 ) | ( n19255 & ~n36151 ) | ( n26556 & ~n36151 ) ;
  assign n36153 = ~n7029 & n22631 ;
  assign n36154 = n36153 ^ n857 ^ 1'b0 ;
  assign n36156 = ~n4157 & n22891 ;
  assign n36155 = n3457 | n7058 ;
  assign n36157 = n36156 ^ n36155 ^ 1'b0 ;
  assign n36158 = n36157 ^ n34382 ^ 1'b0 ;
  assign n36159 = ( ~n8297 & n13578 ) | ( ~n8297 & n28247 ) | ( n13578 & n28247 ) ;
  assign n36160 = n36159 ^ n15550 ^ 1'b0 ;
  assign n36161 = n35617 ^ n34168 ^ n13208 ;
  assign n36162 = n4670 & n9666 ;
  assign n36163 = ~n7907 & n21489 ;
  assign n36164 = ( n1908 & ~n9351 ) | ( n1908 & n36163 ) | ( ~n9351 & n36163 ) ;
  assign n36165 = n14382 | n36164 ;
  assign n36166 = n13127 ^ n11948 ^ 1'b0 ;
  assign n36167 = n1908 & ~n36166 ;
  assign n36168 = n36167 ^ n10755 ^ 1'b0 ;
  assign n36169 = ( ~n11831 & n18230 ) | ( ~n11831 & n36168 ) | ( n18230 & n36168 ) ;
  assign n36170 = n36169 ^ n23917 ^ 1'b0 ;
  assign n36171 = ~n2944 & n23579 ;
  assign n36172 = n36171 ^ n10080 ^ 1'b0 ;
  assign n36173 = ( n9882 & n20886 ) | ( n9882 & ~n21139 ) | ( n20886 & ~n21139 ) ;
  assign n36174 = n3246 & ~n33769 ;
  assign n36175 = n36173 & n36174 ;
  assign n36176 = n10703 & ~n17929 ;
  assign n36177 = x27 & n19635 ;
  assign n36178 = ~n20874 & n36177 ;
  assign n36179 = ( n7688 & ~n36176 ) | ( n7688 & n36178 ) | ( ~n36176 & n36178 ) ;
  assign n36180 = n12660 | n22028 ;
  assign n36181 = n11266 & ~n36180 ;
  assign n36182 = n36181 ^ n22826 ^ x248 ;
  assign n36183 = n496 & n7918 ;
  assign n36185 = ( n1233 & n27622 ) | ( n1233 & ~n29431 ) | ( n27622 & ~n29431 ) ;
  assign n36184 = ( ~n8827 & n19931 ) | ( ~n8827 & n28082 ) | ( n19931 & n28082 ) ;
  assign n36186 = n36185 ^ n36184 ^ 1'b0 ;
  assign n36187 = n13662 & n15091 ;
  assign n36188 = n36187 ^ n34660 ^ 1'b0 ;
  assign n36189 = n17419 ^ n11431 ^ n6560 ;
  assign n36190 = n36189 ^ n10150 ^ 1'b0 ;
  assign n36191 = ~n7431 & n36190 ;
  assign n36196 = ~n3366 & n35264 ;
  assign n36197 = n8053 & n36196 ;
  assign n36198 = n36197 ^ n26680 ^ n16927 ;
  assign n36192 = ( ~n859 & n6558 ) | ( ~n859 & n6649 ) | ( n6558 & n6649 ) ;
  assign n36193 = n36192 ^ n1907 ^ 1'b0 ;
  assign n36194 = n28462 & n36193 ;
  assign n36195 = n36194 ^ n5725 ^ 1'b0 ;
  assign n36199 = n36198 ^ n36195 ^ 1'b0 ;
  assign n36201 = ( n3229 & n5541 ) | ( n3229 & ~n11120 ) | ( n5541 & ~n11120 ) ;
  assign n36200 = n6761 | n18821 ;
  assign n36202 = n36201 ^ n36200 ^ 1'b0 ;
  assign n36203 = ( ~x207 & n2812 ) | ( ~x207 & n23812 ) | ( n2812 & n23812 ) ;
  assign n36204 = n36203 ^ n27042 ^ n16732 ;
  assign n36205 = ( ~n9603 & n36202 ) | ( ~n9603 & n36204 ) | ( n36202 & n36204 ) ;
  assign n36206 = n36205 ^ n17272 ^ 1'b0 ;
  assign n36207 = n36206 ^ n31497 ^ n22203 ;
  assign n36212 = ( ~n4828 & n6999 ) | ( ~n4828 & n19053 ) | ( n6999 & n19053 ) ;
  assign n36210 = ( n3509 & n12356 ) | ( n3509 & n20125 ) | ( n12356 & n20125 ) ;
  assign n36208 = n22256 & n23875 ;
  assign n36209 = n36208 ^ n15052 ^ 1'b0 ;
  assign n36211 = n36210 ^ n36209 ^ n17779 ;
  assign n36213 = n36212 ^ n36211 ^ n35475 ;
  assign n36214 = n36076 ^ n34317 ^ 1'b0 ;
  assign n36215 = n393 | n1102 ;
  assign n36216 = n13220 & n27932 ;
  assign n36217 = n36215 & n36216 ;
  assign n36218 = n10679 ^ n2614 ^ 1'b0 ;
  assign n36219 = ~n10797 & n36218 ;
  assign n36220 = ( n5813 & n23118 ) | ( n5813 & n30780 ) | ( n23118 & n30780 ) ;
  assign n36221 = n36220 ^ n8541 ^ 1'b0 ;
  assign n36222 = n36219 & ~n36221 ;
  assign n36223 = n6339 ^ n2305 ^ 1'b0 ;
  assign n36224 = ( ~n12247 & n14275 ) | ( ~n12247 & n14558 ) | ( n14275 & n14558 ) ;
  assign n36225 = n27716 ^ n24802 ^ n19407 ;
  assign n36226 = ( n36223 & ~n36224 ) | ( n36223 & n36225 ) | ( ~n36224 & n36225 ) ;
  assign n36227 = ~n18967 & n21389 ;
  assign n36228 = n36227 ^ n8543 ^ 1'b0 ;
  assign n36229 = n6763 & ~n7952 ;
  assign n36230 = n11751 & ~n36229 ;
  assign n36231 = ~n22808 & n36230 ;
  assign n36232 = ~n9532 & n32033 ;
  assign n36233 = n33767 & n36232 ;
  assign n36235 = n4749 | n20145 ;
  assign n36234 = n14685 | n20948 ;
  assign n36236 = n36235 ^ n36234 ^ n3786 ;
  assign n36237 = ( n548 & n20546 ) | ( n548 & ~n21071 ) | ( n20546 & ~n21071 ) ;
  assign n36238 = n25528 & n35881 ;
  assign n36239 = n36238 ^ n15859 ^ 1'b0 ;
  assign n36240 = n36239 ^ n23695 ^ 1'b0 ;
  assign n36241 = n22016 & n36240 ;
  assign n36242 = ~n5457 & n9389 ;
  assign n36243 = ~n1563 & n36242 ;
  assign n36244 = ( n487 & n27052 ) | ( n487 & n36243 ) | ( n27052 & n36243 ) ;
  assign n36245 = n36244 ^ n22200 ^ 1'b0 ;
  assign n36246 = n17428 | n36245 ;
  assign n36247 = n18525 ^ n2815 ^ 1'b0 ;
  assign n36248 = n12152 & ~n36247 ;
  assign n36249 = n2642 | n31845 ;
  assign n36250 = n7204 & ~n35741 ;
  assign n36251 = ( n1178 & n2306 ) | ( n1178 & ~n33024 ) | ( n2306 & ~n33024 ) ;
  assign n36252 = n12096 ^ n9250 ^ 1'b0 ;
  assign n36255 = n669 ^ x106 ^ 1'b0 ;
  assign n36253 = ( n2701 & n18959 ) | ( n2701 & ~n20017 ) | ( n18959 & ~n20017 ) ;
  assign n36254 = n36253 ^ n8626 ^ 1'b0 ;
  assign n36256 = n36255 ^ n36254 ^ n21849 ;
  assign n36257 = n8067 & ~n35294 ;
  assign n36258 = x197 & ~n21677 ;
  assign n36259 = n36258 ^ n30591 ^ 1'b0 ;
  assign n36260 = ( n7713 & n11903 ) | ( n7713 & ~n15377 ) | ( n11903 & ~n15377 ) ;
  assign n36261 = n11814 & n36260 ;
  assign n36262 = n33511 & n36261 ;
  assign n36263 = ( n2918 & ~n5007 ) | ( n2918 & n14124 ) | ( ~n5007 & n14124 ) ;
  assign n36264 = n10128 & ~n28837 ;
  assign n36265 = n36263 & n36264 ;
  assign n36266 = n6835 ^ n5191 ^ 1'b0 ;
  assign n36267 = ( x112 & ~n12531 ) | ( x112 & n19304 ) | ( ~n12531 & n19304 ) ;
  assign n36268 = n36267 ^ n27568 ^ 1'b0 ;
  assign n36269 = ( n4830 & n7777 ) | ( n4830 & n36268 ) | ( n7777 & n36268 ) ;
  assign n36270 = n3565 ^ n2011 ^ n723 ;
  assign n36271 = ( n12718 & n20411 ) | ( n12718 & n27112 ) | ( n20411 & n27112 ) ;
  assign n36272 = ~n10056 & n19825 ;
  assign n36273 = ~n19314 & n36272 ;
  assign n36274 = n17075 | n23142 ;
  assign n36275 = n24428 & n36274 ;
  assign n36276 = n36275 ^ n2519 ^ 1'b0 ;
  assign n36277 = n21608 ^ n15068 ^ n4003 ;
  assign n36278 = n5827 & ~n15315 ;
  assign n36279 = ~n36277 & n36278 ;
  assign n36280 = ~n34820 & n36279 ;
  assign n36281 = n10418 & n16008 ;
  assign n36282 = ~n27485 & n36281 ;
  assign n36283 = n22134 ^ n14689 ^ n9089 ;
  assign n36284 = n23927 ^ n18323 ^ n4412 ;
  assign n36285 = ( n12195 & n22799 ) | ( n12195 & ~n36284 ) | ( n22799 & ~n36284 ) ;
  assign n36286 = n32745 ^ n22144 ^ 1'b0 ;
  assign n36287 = n13393 & ~n36286 ;
  assign n36288 = ( ~n12230 & n25293 ) | ( ~n12230 & n36287 ) | ( n25293 & n36287 ) ;
  assign n36289 = ~x27 & n8340 ;
  assign n36290 = ( n6331 & n13524 ) | ( n6331 & ~n34750 ) | ( n13524 & ~n34750 ) ;
  assign n36291 = n16814 ^ n4536 ^ 1'b0 ;
  assign n36292 = n36290 & n36291 ;
  assign n36293 = n18395 ^ n14583 ^ 1'b0 ;
  assign n36294 = n28532 & ~n36293 ;
  assign n36295 = n7406 & n24115 ;
  assign n36296 = n7903 ^ n6695 ^ 1'b0 ;
  assign n36297 = n36296 ^ n14336 ^ n9542 ;
  assign n36298 = n36297 ^ n33662 ^ 1'b0 ;
  assign n36299 = ~n7044 & n36298 ;
  assign n36300 = n18928 ^ n6526 ^ n3120 ;
  assign n36301 = ( n28286 & n30209 ) | ( n28286 & ~n36300 ) | ( n30209 & ~n36300 ) ;
  assign n36302 = ( ~n14634 & n20471 ) | ( ~n14634 & n36301 ) | ( n20471 & n36301 ) ;
  assign n36303 = n36302 ^ n5160 ^ 1'b0 ;
  assign n36304 = ~n18602 & n24415 ;
  assign n36305 = n36304 ^ n32546 ^ 1'b0 ;
  assign n36306 = n16143 ^ n10358 ^ n4906 ;
  assign n36307 = n7311 ^ n2410 ^ 1'b0 ;
  assign n36308 = ~n32772 & n36307 ;
  assign n36309 = n28057 ^ n11669 ^ x31 ;
  assign n36310 = n8251 | n19066 ;
  assign n36311 = n6819 | n14689 ;
  assign n36312 = n20486 | n22297 ;
  assign n36313 = n36312 ^ n19688 ^ 1'b0 ;
  assign n36314 = n36313 ^ n16947 ^ n3166 ;
  assign n36315 = n31768 & n36314 ;
  assign n36316 = n14065 | n33930 ;
  assign n36317 = n24589 | n36316 ;
  assign n36318 = n19278 ^ n11504 ^ 1'b0 ;
  assign n36319 = n13984 & ~n36318 ;
  assign n36320 = n23978 ^ n14174 ^ n6291 ;
  assign n36321 = n9467 | n33849 ;
  assign n36322 = n36320 | n36321 ;
  assign n36323 = n36322 ^ n34766 ^ n27623 ;
  assign n36324 = n8441 & ~n13795 ;
  assign n36325 = n35966 ^ n21944 ^ n13518 ;
  assign n36326 = n27984 ^ n4160 ^ 1'b0 ;
  assign n36327 = ( n4708 & n5369 ) | ( n4708 & n28676 ) | ( n5369 & n28676 ) ;
  assign n36328 = n36326 & ~n36327 ;
  assign n36329 = ( ~n19201 & n36325 ) | ( ~n19201 & n36328 ) | ( n36325 & n36328 ) ;
  assign n36330 = n10005 & ~n32753 ;
  assign n36331 = n23289 & n24219 ;
  assign n36332 = ~n36330 & n36331 ;
  assign n36333 = n10851 & n14156 ;
  assign n36334 = ~n19196 & n35407 ;
  assign n36335 = ( n1655 & ~n5122 ) | ( n1655 & n21888 ) | ( ~n5122 & n21888 ) ;
  assign n36336 = n2710 & n3738 ;
  assign n36337 = n36335 & n36336 ;
  assign n36338 = ( n9119 & ~n12089 ) | ( n9119 & n29664 ) | ( ~n12089 & n29664 ) ;
  assign n36339 = n830 & n36338 ;
  assign n36340 = n19569 ^ n18325 ^ 1'b0 ;
  assign n36341 = n8405 & ~n36340 ;
  assign n36342 = ( n9945 & n12376 ) | ( n9945 & ~n23042 ) | ( n12376 & ~n23042 ) ;
  assign n36347 = ~n1924 & n3601 ;
  assign n36344 = n6945 | n25669 ;
  assign n36345 = n36344 ^ n17731 ^ 1'b0 ;
  assign n36343 = n4077 & n17676 ;
  assign n36346 = n36345 ^ n36343 ^ n18931 ;
  assign n36348 = n36347 ^ n36346 ^ n316 ;
  assign n36349 = ( n29660 & n36342 ) | ( n29660 & ~n36348 ) | ( n36342 & ~n36348 ) ;
  assign n36350 = n6625 | n22181 ;
  assign n36351 = n36350 ^ n6567 ^ 1'b0 ;
  assign n36352 = n9908 | n24432 ;
  assign n36353 = n22270 | n36352 ;
  assign n36354 = n36353 ^ n18262 ^ n595 ;
  assign n36355 = n777 & ~n35328 ;
  assign n36356 = n7674 & ~n36355 ;
  assign n36357 = n36354 & n36356 ;
  assign n36358 = n16793 ^ n7751 ^ 1'b0 ;
  assign n36359 = n1855 ^ n1798 ^ 1'b0 ;
  assign n36360 = n24707 ^ n24040 ^ n7255 ;
  assign n36361 = n1337 | n36360 ;
  assign n36362 = n36361 ^ n18304 ^ 1'b0 ;
  assign n36363 = n36362 ^ n8163 ^ 1'b0 ;
  assign n36364 = n28206 | n36363 ;
  assign n36365 = ( n34948 & n36359 ) | ( n34948 & ~n36364 ) | ( n36359 & ~n36364 ) ;
  assign n36366 = ( x136 & ~n5381 ) | ( x136 & n11294 ) | ( ~n5381 & n11294 ) ;
  assign n36367 = ( ~n5221 & n19227 ) | ( ~n5221 & n36366 ) | ( n19227 & n36366 ) ;
  assign n36371 = n16561 ^ n7252 ^ 1'b0 ;
  assign n36368 = n15410 ^ n10907 ^ 1'b0 ;
  assign n36369 = n22602 ^ n15553 ^ 1'b0 ;
  assign n36370 = n36368 & ~n36369 ;
  assign n36372 = n36371 ^ n36370 ^ n23302 ;
  assign n36373 = n7634 ^ n5050 ^ 1'b0 ;
  assign n36374 = ~n14310 & n36373 ;
  assign n36375 = n2068 & n36374 ;
  assign n36376 = n31515 ^ n7454 ^ 1'b0 ;
  assign n36377 = n16481 & ~n36376 ;
  assign n36378 = n20805 ^ n3106 ^ 1'b0 ;
  assign n36379 = n30237 ^ n26721 ^ n2735 ;
  assign n36380 = n6820 | n25519 ;
  assign n36381 = n29249 & ~n31621 ;
  assign n36382 = n5466 & n36381 ;
  assign n36383 = ~n27590 & n36382 ;
  assign n36386 = n11230 & ~n13571 ;
  assign n36384 = n6983 & n22685 ;
  assign n36385 = n36384 ^ n5529 ^ 1'b0 ;
  assign n36387 = n36386 ^ n36385 ^ 1'b0 ;
  assign n36388 = n1095 | n16342 ;
  assign n36389 = ( n13798 & n30776 ) | ( n13798 & n36388 ) | ( n30776 & n36388 ) ;
  assign n36390 = n5970 & ~n15818 ;
  assign n36391 = n36390 ^ n5484 ^ 1'b0 ;
  assign n36392 = ( ~n6404 & n22584 ) | ( ~n6404 & n36391 ) | ( n22584 & n36391 ) ;
  assign n36393 = n36392 ^ n26464 ^ n24628 ;
  assign n36394 = n11062 | n15841 ;
  assign n36395 = n26270 ^ n25996 ^ n21158 ;
  assign n36396 = n13367 & ~n36395 ;
  assign n36397 = ~n9191 & n36396 ;
  assign n36398 = n32294 | n36397 ;
  assign n36399 = n26342 & ~n36398 ;
  assign n36400 = n21673 ^ n17561 ^ 1'b0 ;
  assign n36401 = n17703 & n36400 ;
  assign n36402 = n31932 ^ n8180 ^ 1'b0 ;
  assign n36403 = n36187 | n36402 ;
  assign n36405 = n23759 ^ n1720 ^ 1'b0 ;
  assign n36404 = n3796 & n24433 ;
  assign n36406 = n36405 ^ n36404 ^ 1'b0 ;
  assign n36407 = n7653 & n18159 ;
  assign n36408 = n7921 & n36407 ;
  assign n36409 = n13531 & ~n36408 ;
  assign n36413 = n1044 & ~n7440 ;
  assign n36414 = n36413 ^ n4308 ^ 1'b0 ;
  assign n36415 = n36414 ^ n14501 ^ 1'b0 ;
  assign n36416 = n36415 ^ n30717 ^ 1'b0 ;
  assign n36412 = n2467 & n14104 ;
  assign n36410 = ~n5773 & n16131 ;
  assign n36411 = n36410 ^ n18917 ^ n3070 ;
  assign n36417 = n36416 ^ n36412 ^ n36411 ;
  assign n36418 = ( n9673 & n16355 ) | ( n9673 & n26188 ) | ( n16355 & n26188 ) ;
  assign n36419 = n29348 ^ n18505 ^ 1'b0 ;
  assign n36420 = n8288 & ~n36419 ;
  assign n36421 = ~n900 & n36420 ;
  assign n36422 = n2853 & ~n7520 ;
  assign n36423 = ~n1888 & n36422 ;
  assign n36424 = n36423 ^ n13642 ^ 1'b0 ;
  assign n36428 = n9050 | n24054 ;
  assign n36429 = n36428 ^ n15170 ^ 1'b0 ;
  assign n36425 = n33730 ^ n21897 ^ n17695 ;
  assign n36426 = n13724 & n36425 ;
  assign n36427 = n36426 ^ n28519 ^ n11079 ;
  assign n36430 = n36429 ^ n36427 ^ n34314 ;
  assign n36431 = ( n23477 & ~n25549 ) | ( n23477 & n36430 ) | ( ~n25549 & n36430 ) ;
  assign n36432 = n32434 ^ n14548 ^ 1'b0 ;
  assign n36433 = n5196 | n7656 ;
  assign n36434 = n36433 ^ n5983 ^ 1'b0 ;
  assign n36435 = ( ~n1497 & n19235 ) | ( ~n1497 & n36434 ) | ( n19235 & n36434 ) ;
  assign n36436 = n36435 ^ n28338 ^ 1'b0 ;
  assign n36437 = n33221 ^ n19877 ^ n1320 ;
  assign n36438 = n10712 & n36437 ;
  assign n36442 = x94 & n27740 ;
  assign n36439 = ~n3701 & n26157 ;
  assign n36440 = n36439 ^ n14984 ^ 1'b0 ;
  assign n36441 = n12222 | n36440 ;
  assign n36443 = n36442 ^ n36441 ^ 1'b0 ;
  assign n36444 = n21248 & ~n26832 ;
  assign n36445 = n11296 & n36444 ;
  assign n36446 = n21974 ^ n7190 ^ 1'b0 ;
  assign n36447 = n20591 ^ n18230 ^ n17321 ;
  assign n36448 = ( x35 & n5383 ) | ( x35 & n6427 ) | ( n5383 & n6427 ) ;
  assign n36449 = ( n3437 & n23950 ) | ( n3437 & n36448 ) | ( n23950 & n36448 ) ;
  assign n36450 = ( n17290 & n36447 ) | ( n17290 & ~n36449 ) | ( n36447 & ~n36449 ) ;
  assign n36451 = n35123 ^ n3062 ^ n2764 ;
  assign n36452 = ~n9520 & n36451 ;
  assign n36453 = n6515 & ~n19640 ;
  assign n36454 = n2778 & n36453 ;
  assign n36455 = n36454 ^ n2542 ^ 1'b0 ;
  assign n36456 = n24814 ^ n7666 ^ n4129 ;
  assign n36457 = n12163 & n36456 ;
  assign n36458 = ( n19409 & n25374 ) | ( n19409 & n36457 ) | ( n25374 & n36457 ) ;
  assign n36459 = ( ~n10563 & n36455 ) | ( ~n10563 & n36458 ) | ( n36455 & n36458 ) ;
  assign n36460 = n14582 & n36411 ;
  assign n36461 = n36459 & n36460 ;
  assign n36462 = n4819 | n23106 ;
  assign n36463 = n36462 ^ n5100 ^ 1'b0 ;
  assign n36464 = n3022 & n15207 ;
  assign n36468 = n8412 & ~n13082 ;
  assign n36465 = n19465 & ~n24900 ;
  assign n36466 = n8727 & n36465 ;
  assign n36467 = ( n15641 & ~n21888 ) | ( n15641 & n36466 ) | ( ~n21888 & n36466 ) ;
  assign n36469 = n36468 ^ n36467 ^ 1'b0 ;
  assign n36470 = n36464 & ~n36469 ;
  assign n36471 = n6568 & n16442 ;
  assign n36472 = n36471 ^ n5593 ^ 1'b0 ;
  assign n36474 = n34485 ^ n14130 ^ 1'b0 ;
  assign n36475 = n5476 | n36474 ;
  assign n36473 = n13208 ^ n4032 ^ 1'b0 ;
  assign n36476 = n36475 ^ n36473 ^ 1'b0 ;
  assign n36477 = n1360 & n36476 ;
  assign n36478 = ~n6209 & n36477 ;
  assign n36479 = n13340 & n32420 ;
  assign n36480 = n36479 ^ n11019 ^ n10287 ;
  assign n36481 = n28243 ^ n26853 ^ 1'b0 ;
  assign n36482 = n10057 | n36481 ;
  assign n36483 = n36482 ^ n10389 ^ 1'b0 ;
  assign n36484 = n36483 ^ n19758 ^ n3264 ;
  assign n36485 = ( n1559 & ~n18338 ) | ( n1559 & n21622 ) | ( ~n18338 & n21622 ) ;
  assign n36486 = n29911 & ~n35855 ;
  assign n36487 = ~n36485 & n36486 ;
  assign n36488 = n36487 ^ n29366 ^ n10799 ;
  assign n36491 = ~n7561 & n18665 ;
  assign n36492 = n36491 ^ n3952 ^ 1'b0 ;
  assign n36489 = n19319 | n22980 ;
  assign n36490 = n36489 ^ n13035 ^ 1'b0 ;
  assign n36493 = n36492 ^ n36490 ^ 1'b0 ;
  assign n36494 = ~n26867 & n34336 ;
  assign n36495 = n36494 ^ n34730 ^ 1'b0 ;
  assign n36496 = n13450 ^ n8533 ^ 1'b0 ;
  assign n36497 = ~n15924 & n36496 ;
  assign n36498 = n21624 ^ n14802 ^ 1'b0 ;
  assign n36499 = n21835 | n36498 ;
  assign n36500 = ~n9444 & n29684 ;
  assign n36501 = ~n13435 & n36500 ;
  assign n36502 = ( ~n12649 & n30179 ) | ( ~n12649 & n36501 ) | ( n30179 & n36501 ) ;
  assign n36506 = n1348 & n5872 ;
  assign n36507 = n5166 & n36506 ;
  assign n36505 = n11561 | n13191 ;
  assign n36508 = n36507 ^ n36505 ^ 1'b0 ;
  assign n36503 = n19736 ^ n10759 ^ n2875 ;
  assign n36504 = ( ~n20436 & n21932 ) | ( ~n20436 & n36503 ) | ( n21932 & n36503 ) ;
  assign n36509 = n36508 ^ n36504 ^ n9637 ;
  assign n36510 = n33361 ^ n27193 ^ n1978 ;
  assign n36511 = ( n6868 & n19407 ) | ( n6868 & ~n27659 ) | ( n19407 & ~n27659 ) ;
  assign n36512 = n35386 ^ n22818 ^ 1'b0 ;
  assign n36513 = n36511 & ~n36512 ;
  assign n36514 = n11131 & n20076 ;
  assign n36515 = n25521 ^ n7542 ^ 1'b0 ;
  assign n36516 = n25971 | n36515 ;
  assign n36517 = ( n1435 & n20769 ) | ( n1435 & n36516 ) | ( n20769 & n36516 ) ;
  assign n36518 = ( n5359 & n28250 ) | ( n5359 & ~n36517 ) | ( n28250 & ~n36517 ) ;
  assign n36519 = n3029 | n23282 ;
  assign n36520 = n8851 & ~n36519 ;
  assign n36521 = n36520 ^ n8935 ^ n1537 ;
  assign n36522 = n15956 ^ n6173 ^ 1'b0 ;
  assign n36523 = n13624 ^ n6341 ^ 1'b0 ;
  assign n36524 = ~n36253 & n36523 ;
  assign n36525 = n36524 ^ n23425 ^ 1'b0 ;
  assign n36526 = n28608 ^ n12917 ^ n7388 ;
  assign n36527 = n36526 ^ n15805 ^ 1'b0 ;
  assign n36528 = n32496 & ~n36527 ;
  assign n36529 = n36528 ^ n31791 ^ 1'b0 ;
  assign n36530 = ~n32264 & n35515 ;
  assign n36531 = n36530 ^ n33942 ^ 1'b0 ;
  assign n36532 = ( ~n3079 & n3212 ) | ( ~n3079 & n35384 ) | ( n3212 & n35384 ) ;
  assign n36533 = ( n17375 & n32335 ) | ( n17375 & ~n36532 ) | ( n32335 & ~n36532 ) ;
  assign n36534 = n7834 & ~n28743 ;
  assign n36535 = ( ~n374 & n31796 ) | ( ~n374 & n36534 ) | ( n31796 & n36534 ) ;
  assign n36536 = ( n2571 & n36533 ) | ( n2571 & n36535 ) | ( n36533 & n36535 ) ;
  assign n36537 = n25780 ^ n16458 ^ 1'b0 ;
  assign n36538 = n14197 & ~n36537 ;
  assign n36539 = ~n6994 & n10694 ;
  assign n36540 = n36539 ^ n4351 ^ 1'b0 ;
  assign n36541 = n2363 & n36540 ;
  assign n36542 = n9782 ^ n3920 ^ 1'b0 ;
  assign n36543 = n33117 ^ n26764 ^ n14584 ;
  assign n36544 = n36543 ^ n27641 ^ 1'b0 ;
  assign n36545 = n11527 & n36544 ;
  assign n36546 = n15283 & n23743 ;
  assign n36547 = n36546 ^ n23640 ^ 1'b0 ;
  assign n36549 = ( ~n1030 & n9882 ) | ( ~n1030 & n10152 ) | ( n9882 & n10152 ) ;
  assign n36548 = n15399 & ~n19456 ;
  assign n36550 = n36549 ^ n36548 ^ 1'b0 ;
  assign n36551 = n36550 ^ n12784 ^ n11782 ;
  assign n36553 = n2477 & ~n23192 ;
  assign n36552 = n5917 & ~n34397 ;
  assign n36554 = n36553 ^ n36552 ^ 1'b0 ;
  assign n36555 = ~n7963 & n36554 ;
  assign n36556 = ~n36551 & n36555 ;
  assign n36557 = n10591 | n36556 ;
  assign n36558 = n36557 ^ n24035 ^ 1'b0 ;
  assign n36559 = n20164 ^ n9049 ^ 1'b0 ;
  assign n36560 = n36559 ^ n15473 ^ n5262 ;
  assign n36561 = n5476 & ~n12500 ;
  assign n36562 = ( n18017 & n24414 ) | ( n18017 & ~n30675 ) | ( n24414 & ~n30675 ) ;
  assign n36563 = n25821 ^ n10123 ^ 1'b0 ;
  assign n36564 = n36563 ^ n13668 ^ 1'b0 ;
  assign n36565 = n13074 ^ n2753 ^ 1'b0 ;
  assign n36566 = n24997 ^ x33 ^ 1'b0 ;
  assign n36567 = n36565 & n36566 ;
  assign n36568 = n30634 ^ n8802 ^ 1'b0 ;
  assign n36569 = n9030 & n36568 ;
  assign n36570 = n36569 ^ n28967 ^ n4333 ;
  assign n36571 = n25746 ^ n3975 ^ n2585 ;
  assign n36572 = n1385 | n5799 ;
  assign n36573 = ~n13987 & n36572 ;
  assign n36574 = n23991 ^ n20568 ^ 1'b0 ;
  assign n36575 = n36574 ^ n18451 ^ n10181 ;
  assign n36576 = n14155 ^ n1106 ^ 1'b0 ;
  assign n36577 = n2170 & n15379 ;
  assign n36578 = n7860 & ~n36577 ;
  assign n36579 = ~n3264 & n7227 ;
  assign n36580 = ~n7852 & n36579 ;
  assign n36581 = n9722 & ~n36580 ;
  assign n36582 = n36581 ^ n6380 ^ 1'b0 ;
  assign n36583 = n36582 ^ n26395 ^ 1'b0 ;
  assign n36584 = n11130 | n36583 ;
  assign n36585 = n14379 ^ n13382 ^ 1'b0 ;
  assign n36586 = n7643 | n36585 ;
  assign n36587 = n36586 ^ n6872 ^ 1'b0 ;
  assign n36588 = ~n8311 & n36587 ;
  assign n36589 = n36588 ^ n26160 ^ 1'b0 ;
  assign n36590 = n36285 | n36589 ;
  assign n36591 = n6240 & ~n36590 ;
  assign n36592 = ~n7754 & n20620 ;
  assign n36593 = n22840 & n36592 ;
  assign n36594 = n36593 ^ n25044 ^ n8281 ;
  assign n36595 = n22495 ^ n20104 ^ n5293 ;
  assign n36596 = ( x84 & n28243 ) | ( x84 & n36595 ) | ( n28243 & n36595 ) ;
  assign n36597 = n9647 | n27153 ;
  assign n36598 = n20012 & n29868 ;
  assign n36599 = n36598 ^ n3525 ^ 1'b0 ;
  assign n36600 = n32760 ^ n25347 ^ n21094 ;
  assign n36604 = n6523 ^ n5424 ^ n1171 ;
  assign n36605 = ( ~n417 & n14021 ) | ( ~n417 & n16994 ) | ( n14021 & n16994 ) ;
  assign n36606 = n18569 & ~n36605 ;
  assign n36607 = ~n36604 & n36606 ;
  assign n36601 = ( n2186 & n19027 ) | ( n2186 & ~n35403 ) | ( n19027 & ~n35403 ) ;
  assign n36602 = n33012 & ~n36601 ;
  assign n36603 = n17778 & n36602 ;
  assign n36608 = n36607 ^ n36603 ^ 1'b0 ;
  assign n36609 = n22160 ^ n17489 ^ 1'b0 ;
  assign n36610 = n20574 ^ n3711 ^ 1'b0 ;
  assign n36611 = n18734 | n36610 ;
  assign n36612 = n17308 | n18277 ;
  assign n36613 = n36612 ^ n5892 ^ 1'b0 ;
  assign n36614 = n18070 & ~n36613 ;
  assign n36615 = n13541 ^ n8073 ^ 1'b0 ;
  assign n36616 = ( ~n10988 & n11197 ) | ( ~n10988 & n22820 ) | ( n11197 & n22820 ) ;
  assign n36617 = n36616 ^ n35396 ^ 1'b0 ;
  assign n36618 = n36615 | n36617 ;
  assign n36619 = n17518 ^ n13032 ^ 1'b0 ;
  assign n36620 = n35316 ^ n29898 ^ n18764 ;
  assign n36621 = n36620 ^ n23081 ^ n3791 ;
  assign n36622 = n6893 ^ n1754 ^ 1'b0 ;
  assign n36623 = n9478 ^ n5599 ^ n2052 ;
  assign n36624 = n36623 ^ n24541 ^ 1'b0 ;
  assign n36625 = n36622 & ~n36624 ;
  assign n36626 = n8763 | n11285 ;
  assign n36627 = n36626 ^ n25850 ^ 1'b0 ;
  assign n36628 = n36625 & n36627 ;
  assign n36629 = ( n14581 & ~n25950 ) | ( n14581 & n36628 ) | ( ~n25950 & n36628 ) ;
  assign n36630 = ~n9475 & n24266 ;
  assign n36631 = n36630 ^ n20454 ^ n10694 ;
  assign n36632 = n15896 & n36631 ;
  assign n36633 = ( n33683 & n35960 ) | ( n33683 & n36632 ) | ( n35960 & n36632 ) ;
  assign n36634 = n21878 ^ n16441 ^ n1014 ;
  assign n36635 = ~n19414 & n24453 ;
  assign n36636 = n36634 & n36635 ;
  assign n36637 = ( n20315 & n25084 ) | ( n20315 & n29519 ) | ( n25084 & n29519 ) ;
  assign n36638 = n6602 ^ n4998 ^ 1'b0 ;
  assign n36639 = n36637 | n36638 ;
  assign n36642 = ( x148 & n5135 ) | ( x148 & n36414 ) | ( n5135 & n36414 ) ;
  assign n36643 = ( n5406 & n16685 ) | ( n5406 & ~n36642 ) | ( n16685 & ~n36642 ) ;
  assign n36640 = n605 & ~n34093 ;
  assign n36641 = n36640 ^ n24368 ^ 1'b0 ;
  assign n36644 = n36643 ^ n36641 ^ 1'b0 ;
  assign n36645 = ~n8124 & n23427 ;
  assign n36646 = n28734 ^ n12574 ^ 1'b0 ;
  assign n36647 = n11581 ^ n9637 ^ x93 ;
  assign n36648 = ( n1035 & n19172 ) | ( n1035 & ~n36647 ) | ( n19172 & ~n36647 ) ;
  assign n36649 = ( n1771 & n24391 ) | ( n1771 & ~n36648 ) | ( n24391 & ~n36648 ) ;
  assign n36650 = n12946 ^ n11591 ^ n11304 ;
  assign n36651 = n23865 ^ n14138 ^ n8151 ;
  assign n36652 = n5948 | n12830 ;
  assign n36653 = n36652 ^ n7125 ^ 1'b0 ;
  assign n36654 = ( n13755 & n36651 ) | ( n13755 & ~n36653 ) | ( n36651 & ~n36653 ) ;
  assign n36655 = ~n7638 & n16234 ;
  assign n36656 = ( n5460 & ~n16288 ) | ( n5460 & n29289 ) | ( ~n16288 & n29289 ) ;
  assign n36657 = n4168 & n36656 ;
  assign n36658 = ~n36227 & n36657 ;
  assign n36659 = ~n19972 & n30132 ;
  assign n36660 = n7830 & n36659 ;
  assign n36661 = ~n4124 & n8519 ;
  assign n36662 = n36661 ^ n21790 ^ n6466 ;
  assign n36663 = ~n18680 & n36662 ;
  assign n36664 = ( n2478 & ~n10017 ) | ( n2478 & n11112 ) | ( ~n10017 & n11112 ) ;
  assign n36665 = ( n770 & n12289 ) | ( n770 & n13780 ) | ( n12289 & n13780 ) ;
  assign n36666 = n937 ^ x96 ^ 1'b0 ;
  assign n36667 = n6511 & ~n36666 ;
  assign n36673 = n19992 ^ n19030 ^ 1'b0 ;
  assign n36674 = n10987 | n36673 ;
  assign n36668 = ~n6431 & n13452 ;
  assign n36669 = n36668 ^ n5802 ^ 1'b0 ;
  assign n36670 = ( n7367 & ~n11489 ) | ( n7367 & n36669 ) | ( ~n11489 & n36669 ) ;
  assign n36671 = n6866 ^ n5797 ^ 1'b0 ;
  assign n36672 = ~n36670 & n36671 ;
  assign n36675 = n36674 ^ n36672 ^ 1'b0 ;
  assign n36676 = n36667 & n36675 ;
  assign n36677 = n22504 ^ n11978 ^ n7377 ;
  assign n36680 = n12594 ^ n5500 ^ n3602 ;
  assign n36678 = n27250 ^ n12590 ^ n10919 ;
  assign n36679 = ~n13207 & n36678 ;
  assign n36681 = n36680 ^ n36679 ^ 1'b0 ;
  assign n36682 = n10178 & n12133 ;
  assign n36683 = ( n10122 & ~n11793 ) | ( n10122 & n36682 ) | ( ~n11793 & n36682 ) ;
  assign n36684 = ~n9226 & n36683 ;
  assign n36685 = n34125 ^ n15425 ^ 1'b0 ;
  assign n36686 = n10743 ^ n8978 ^ n6793 ;
  assign n36687 = ( ~n11667 & n21776 ) | ( ~n11667 & n23611 ) | ( n21776 & n23611 ) ;
  assign n36688 = n36687 ^ n1380 ^ 1'b0 ;
  assign n36689 = ( n32223 & ~n36686 ) | ( n32223 & n36688 ) | ( ~n36686 & n36688 ) ;
  assign n36690 = x135 & ~n8030 ;
  assign n36691 = n36690 ^ n21766 ^ 1'b0 ;
  assign n36692 = n16867 ^ n13459 ^ x9 ;
  assign n36693 = ( ~n7803 & n21101 ) | ( ~n7803 & n36692 ) | ( n21101 & n36692 ) ;
  assign n36694 = n21026 & ~n36693 ;
  assign n36695 = n7217 ^ n2410 ^ n1641 ;
  assign n36696 = n36695 ^ n4419 ^ 1'b0 ;
  assign n36697 = ~n8053 & n36696 ;
  assign n36698 = n36697 ^ n28387 ^ 1'b0 ;
  assign n36699 = n16193 & ~n36698 ;
  assign n36700 = n1764 | n6073 ;
  assign n36701 = ( n13480 & ~n20227 ) | ( n13480 & n24380 ) | ( ~n20227 & n24380 ) ;
  assign n36702 = n36701 ^ x200 ^ 1'b0 ;
  assign n36703 = n31181 & ~n36702 ;
  assign n36704 = ( n16555 & n36700 ) | ( n16555 & n36703 ) | ( n36700 & n36703 ) ;
  assign n36705 = n29856 ^ n7274 ^ 1'b0 ;
  assign n36706 = n36705 ^ n32961 ^ n23444 ;
  assign n36707 = n27870 & n31499 ;
  assign n36708 = n15190 ^ n7201 ^ 1'b0 ;
  assign n36709 = n24235 & n36708 ;
  assign n36710 = n23314 ^ n8249 ^ 1'b0 ;
  assign n36711 = n625 | n14636 ;
  assign n36712 = n36711 ^ n24472 ^ 1'b0 ;
  assign n36713 = n23271 & ~n25112 ;
  assign n36714 = n36713 ^ n3896 ^ 1'b0 ;
  assign n36715 = ( n7806 & ~n9752 ) | ( n7806 & n36714 ) | ( ~n9752 & n36714 ) ;
  assign n36716 = n27016 ^ n11378 ^ n703 ;
  assign n36717 = n24366 ^ n17517 ^ 1'b0 ;
  assign n36718 = n758 | n36717 ;
  assign n36719 = n36718 ^ n31037 ^ n13780 ;
  assign n36720 = n5641 | n24337 ;
  assign n36721 = n36229 ^ n24895 ^ n12107 ;
  assign n36722 = n36721 ^ n10432 ^ 1'b0 ;
  assign n36723 = ~n514 & n12653 ;
  assign n36724 = n36723 ^ n5370 ^ 1'b0 ;
  assign n36725 = n4959 | n9587 ;
  assign n36726 = n9904 ^ n8465 ^ 1'b0 ;
  assign n36727 = n34229 ^ n15156 ^ n7889 ;
  assign n36728 = n10053 ^ n8369 ^ n3076 ;
  assign n36729 = n36728 ^ n6851 ^ n2297 ;
  assign n36730 = n17723 ^ n3647 ^ 1'b0 ;
  assign n36731 = ( ~n20262 & n23587 ) | ( ~n20262 & n36730 ) | ( n23587 & n36730 ) ;
  assign n36732 = n18064 ^ n12450 ^ 1'b0 ;
  assign n36733 = ~n18720 & n36732 ;
  assign n36734 = n4945 ^ n3699 ^ 1'b0 ;
  assign n36735 = n3080 | n18243 ;
  assign n36736 = n36735 ^ n16486 ^ n9042 ;
  assign n36737 = n10631 & n36736 ;
  assign n36738 = n36734 & n36737 ;
  assign n36739 = n3189 & n16412 ;
  assign n36740 = n36739 ^ n5210 ^ 1'b0 ;
  assign n36741 = n36740 ^ n11556 ^ n7146 ;
  assign n36742 = n36741 ^ n20667 ^ n2890 ;
  assign n36743 = n13390 & n36742 ;
  assign n36744 = ~n2145 & n17488 ;
  assign n36745 = ( n2364 & n14785 ) | ( n2364 & ~n26025 ) | ( n14785 & ~n26025 ) ;
  assign n36746 = n11860 ^ n9840 ^ n7515 ;
  assign n36747 = ( n13467 & n34694 ) | ( n13467 & ~n36746 ) | ( n34694 & ~n36746 ) ;
  assign n36748 = n23558 & ~n31175 ;
  assign n36749 = n1374 | n26058 ;
  assign n36750 = n24989 ^ n14529 ^ 1'b0 ;
  assign n36751 = n20765 & ~n36750 ;
  assign n36752 = n6908 & n20609 ;
  assign n36753 = n18271 ^ n9154 ^ n6800 ;
  assign n36754 = n5420 ^ n4819 ^ 1'b0 ;
  assign n36755 = n36754 ^ n18377 ^ n9184 ;
  assign n36756 = ( n1522 & n36753 ) | ( n1522 & ~n36755 ) | ( n36753 & ~n36755 ) ;
  assign n36757 = ~n6620 & n12719 ;
  assign n36758 = n9808 & n36757 ;
  assign n36759 = n1629 & n36758 ;
  assign n36760 = n28280 ^ n11303 ^ 1'b0 ;
  assign n36761 = n2085 ^ n1906 ^ n1538 ;
  assign n36762 = n4150 & n36761 ;
  assign n36763 = n36760 & n36762 ;
  assign n36764 = n28868 ^ n28269 ^ 1'b0 ;
  assign n36765 = n31749 | n36764 ;
  assign n36767 = n14026 ^ n3247 ^ 1'b0 ;
  assign n36766 = ( n23700 & ~n26866 ) | ( n23700 & n29939 ) | ( ~n26866 & n29939 ) ;
  assign n36768 = n36767 ^ n36766 ^ 1'b0 ;
  assign n36769 = n36768 ^ n28520 ^ n15558 ;
  assign n36770 = ( n1070 & n3495 ) | ( n1070 & n33257 ) | ( n3495 & n33257 ) ;
  assign n36771 = ( ~n23354 & n32823 ) | ( ~n23354 & n36770 ) | ( n32823 & n36770 ) ;
  assign n36772 = ( n8808 & n26941 ) | ( n8808 & ~n28842 ) | ( n26941 & ~n28842 ) ;
  assign n36773 = n742 & n28182 ;
  assign n36774 = n1440 | n2793 ;
  assign n36775 = n9149 & ~n36774 ;
  assign n36776 = n3240 | n36775 ;
  assign n36777 = n5898 ^ n3736 ^ 1'b0 ;
  assign n36778 = n3568 & ~n10327 ;
  assign n36779 = ~n36777 & n36778 ;
  assign n36780 = n5356 ^ n3062 ^ 1'b0 ;
  assign n36781 = ~n2241 & n36780 ;
  assign n36782 = ~n15861 & n36781 ;
  assign n36783 = n36779 & n36782 ;
  assign n36784 = n11947 ^ n11177 ^ 1'b0 ;
  assign n36785 = n23268 ^ n1582 ^ 1'b0 ;
  assign n36786 = n36785 ^ n4975 ^ 1'b0 ;
  assign n36787 = ~n9139 & n36786 ;
  assign n36788 = ( n7676 & n36784 ) | ( n7676 & ~n36787 ) | ( n36784 & ~n36787 ) ;
  assign n36789 = n22395 ^ n10660 ^ 1'b0 ;
  assign n36790 = ( n10458 & n24963 ) | ( n10458 & ~n33767 ) | ( n24963 & ~n33767 ) ;
  assign n36791 = n16506 | n36790 ;
  assign n36792 = n36791 ^ n36582 ^ 1'b0 ;
  assign n36793 = n10029 ^ n3018 ^ n2705 ;
  assign n36794 = ( n3180 & n9659 ) | ( n3180 & ~n36793 ) | ( n9659 & ~n36793 ) ;
  assign n36795 = ~n30144 & n30409 ;
  assign n36802 = n4358 | n4682 ;
  assign n36796 = n7649 ^ n2110 ^ 1'b0 ;
  assign n36797 = ~n8709 & n36796 ;
  assign n36798 = n8393 & ~n11838 ;
  assign n36799 = ( n4801 & n36797 ) | ( n4801 & ~n36798 ) | ( n36797 & ~n36798 ) ;
  assign n36800 = n3598 | n36799 ;
  assign n36801 = n29297 | n36800 ;
  assign n36803 = n36802 ^ n36801 ^ 1'b0 ;
  assign n36804 = n13251 ^ n1675 ^ 1'b0 ;
  assign n36805 = n21637 ^ n18020 ^ 1'b0 ;
  assign n36806 = n5288 & n36805 ;
  assign n36807 = n36806 ^ n33064 ^ n11371 ;
  assign n36808 = n23104 | n31882 ;
  assign n36809 = ( n19848 & n29449 ) | ( n19848 & n36808 ) | ( n29449 & n36808 ) ;
  assign n36819 = ( n5229 & ~n16818 ) | ( n5229 & n25599 ) | ( ~n16818 & n25599 ) ;
  assign n36810 = ~n2862 & n11106 ;
  assign n36811 = n2871 & n36810 ;
  assign n36812 = ~n14361 & n33139 ;
  assign n36813 = n36811 & n36812 ;
  assign n36814 = n36813 ^ n2436 ^ 1'b0 ;
  assign n36815 = n7060 & n36814 ;
  assign n36816 = ~n13335 & n36815 ;
  assign n36817 = n19089 & n36816 ;
  assign n36818 = n25453 | n36817 ;
  assign n36820 = n36819 ^ n36818 ^ 1'b0 ;
  assign n36821 = ~n9857 & n27459 ;
  assign n36822 = ( n9997 & ~n31047 ) | ( n9997 & n36821 ) | ( ~n31047 & n36821 ) ;
  assign n36823 = n27965 & n36822 ;
  assign n36824 = n36823 ^ n16603 ^ 1'b0 ;
  assign n36825 = n16703 ^ n13645 ^ 1'b0 ;
  assign n36826 = n26019 | n36825 ;
  assign n36827 = n14018 & ~n36826 ;
  assign n36828 = n2314 | n2716 ;
  assign n36829 = n36827 & ~n36828 ;
  assign n36831 = n22060 ^ n18935 ^ 1'b0 ;
  assign n36830 = ~n13341 & n16749 ;
  assign n36832 = n36831 ^ n36830 ^ 1'b0 ;
  assign n36834 = n20528 ^ n8612 ^ 1'b0 ;
  assign n36835 = n33316 & n36834 ;
  assign n36833 = n7582 & ~n32704 ;
  assign n36836 = n36835 ^ n36833 ^ 1'b0 ;
  assign n36837 = ~n5532 & n19614 ;
  assign n36838 = n10641 & ~n36837 ;
  assign n36839 = n36838 ^ n5328 ^ 1'b0 ;
  assign n36840 = n17531 & n31155 ;
  assign n36841 = n36840 ^ n16359 ^ 1'b0 ;
  assign n36842 = ( ~n4047 & n5042 ) | ( ~n4047 & n9922 ) | ( n5042 & n9922 ) ;
  assign n36843 = n32343 ^ n8528 ^ 1'b0 ;
  assign n36844 = ( n2580 & n7480 ) | ( n2580 & n16970 ) | ( n7480 & n16970 ) ;
  assign n36845 = ( n25962 & ~n36843 ) | ( n25962 & n36844 ) | ( ~n36843 & n36844 ) ;
  assign n36846 = n1959 & ~n29576 ;
  assign n36847 = n36846 ^ n11773 ^ 1'b0 ;
  assign n36848 = ~n13811 & n27250 ;
  assign n36849 = n36848 ^ n12990 ^ 1'b0 ;
  assign n36850 = x154 & ~n13868 ;
  assign n36851 = n36850 ^ n1961 ^ 1'b0 ;
  assign n36852 = n36851 ^ n3401 ^ 1'b0 ;
  assign n36853 = ~n36849 & n36852 ;
  assign n36854 = n2925 ^ x222 ^ 1'b0 ;
  assign n36855 = ~n11687 & n36854 ;
  assign n36856 = n21624 & n36855 ;
  assign n36859 = ~n4137 & n8819 ;
  assign n36860 = ~n435 & n36859 ;
  assign n36861 = n36860 ^ n18304 ^ 1'b0 ;
  assign n36857 = n8253 & ~n19945 ;
  assign n36858 = n36857 ^ n11584 ^ 1'b0 ;
  assign n36862 = n36861 ^ n36858 ^ n3510 ;
  assign n36863 = ~n16549 & n20629 ;
  assign n36864 = n30358 ^ n10608 ^ n7836 ;
  assign n36865 = ~n3770 & n11398 ;
  assign n36866 = n7531 ^ n735 ^ 1'b0 ;
  assign n36867 = n36865 | n36866 ;
  assign n36868 = ( n7538 & ~n8063 ) | ( n7538 & n9634 ) | ( ~n8063 & n9634 ) ;
  assign n36869 = n36868 ^ n8581 ^ 1'b0 ;
  assign n36870 = ~n13676 & n36869 ;
  assign n36871 = ( n1283 & ~n16565 ) | ( n1283 & n28874 ) | ( ~n16565 & n28874 ) ;
  assign n36872 = n1208 & ~n36871 ;
  assign n36873 = n11188 & n36872 ;
  assign n36874 = ( n7503 & n23749 ) | ( n7503 & n24212 ) | ( n23749 & n24212 ) ;
  assign n36875 = n22677 ^ n9021 ^ 1'b0 ;
  assign n36876 = n17701 & ~n36875 ;
  assign n36877 = n2557 | n34878 ;
  assign n36878 = n36876 | n36877 ;
  assign n36879 = n36878 ^ n27633 ^ 1'b0 ;
  assign n36880 = ~n12891 & n14444 ;
  assign n36881 = n35396 & n36880 ;
  assign n36882 = n9127 | n28000 ;
  assign n36883 = n36882 ^ n4066 ^ 1'b0 ;
  assign n36884 = n23760 ^ n13443 ^ n9700 ;
  assign n36885 = n15305 ^ n8923 ^ n3548 ;
  assign n36886 = ( ~n1350 & n5369 ) | ( ~n1350 & n36885 ) | ( n5369 & n36885 ) ;
  assign n36887 = n36886 ^ n20259 ^ n7887 ;
  assign n36888 = ( n1538 & n14196 ) | ( n1538 & n36887 ) | ( n14196 & n36887 ) ;
  assign n36889 = n15657 ^ n1698 ^ n698 ;
  assign n36890 = n18106 ^ n5292 ^ 1'b0 ;
  assign n36891 = ( ~n35819 & n36889 ) | ( ~n35819 & n36890 ) | ( n36889 & n36890 ) ;
  assign n36892 = n3958 ^ n1953 ^ 1'b0 ;
  assign n36893 = n17771 ^ n13361 ^ n12917 ;
  assign n36894 = ( n18673 & n36892 ) | ( n18673 & n36893 ) | ( n36892 & n36893 ) ;
  assign n36895 = n36894 ^ n7770 ^ n5656 ;
  assign n36896 = n5150 ^ n2741 ^ 1'b0 ;
  assign n36897 = ~n3075 & n36896 ;
  assign n36898 = ( ~n19441 & n36895 ) | ( ~n19441 & n36897 ) | ( n36895 & n36897 ) ;
  assign n36899 = n4091 & n26020 ;
  assign n36900 = ~n8093 & n15570 ;
  assign n36901 = ( n13616 & n20269 ) | ( n13616 & n36900 ) | ( n20269 & n36900 ) ;
  assign n36902 = ( n4820 & ~n9134 ) | ( n4820 & n14944 ) | ( ~n9134 & n14944 ) ;
  assign n36904 = n1303 ^ n951 ^ 1'b0 ;
  assign n36905 = ~n10528 & n36904 ;
  assign n36903 = n5322 | n20859 ;
  assign n36906 = n36905 ^ n36903 ^ 1'b0 ;
  assign n36907 = n12030 & n36906 ;
  assign n36908 = n8657 | n13375 ;
  assign n36909 = n32568 & ~n36908 ;
  assign n36910 = n3973 & n8315 ;
  assign n36911 = n36910 ^ n16412 ^ 1'b0 ;
  assign n36912 = n7908 ^ n2599 ^ 1'b0 ;
  assign n36913 = n583 | n32834 ;
  assign n36914 = n6092 & ~n23184 ;
  assign n36915 = n36914 ^ n18318 ^ 1'b0 ;
  assign n36916 = ( n17828 & n21633 ) | ( n17828 & n36915 ) | ( n21633 & n36915 ) ;
  assign n36917 = n27570 ^ n24177 ^ n8250 ;
  assign n36918 = n5184 | n32501 ;
  assign n36919 = n36918 ^ n5912 ^ 1'b0 ;
  assign n36920 = ( n5013 & n32696 ) | ( n5013 & ~n36919 ) | ( n32696 & ~n36919 ) ;
  assign n36921 = n13121 | n26438 ;
  assign n36922 = n36921 ^ n27933 ^ 1'b0 ;
  assign n36923 = ~n36920 & n36922 ;
  assign n36924 = n17123 ^ n2390 ^ 1'b0 ;
  assign n36925 = n36923 & ~n36924 ;
  assign n36926 = n12299 ^ n10404 ^ n2649 ;
  assign n36927 = n36926 ^ n6444 ^ 1'b0 ;
  assign n36928 = n21020 ^ n17583 ^ n14983 ;
  assign n36929 = n36928 ^ n12598 ^ n3292 ;
  assign n36930 = ~n3395 & n6973 ;
  assign n36931 = ~n3309 & n12783 ;
  assign n36932 = n13817 | n36931 ;
  assign n36933 = n36932 ^ n16937 ^ 1'b0 ;
  assign n36934 = n20851 ^ n15730 ^ n5347 ;
  assign n36935 = ( n36930 & n36933 ) | ( n36930 & n36934 ) | ( n36933 & n36934 ) ;
  assign n36936 = ~n25288 & n36487 ;
  assign n36937 = n8250 & ~n15736 ;
  assign n36938 = ~n3319 & n36937 ;
  assign n36939 = n14239 ^ n10952 ^ 1'b0 ;
  assign n36940 = n26024 ^ n21903 ^ 1'b0 ;
  assign n36941 = n36939 & ~n36940 ;
  assign n36942 = n16046 ^ n9524 ^ 1'b0 ;
  assign n36943 = n21292 & ~n36942 ;
  assign n36944 = n907 & n36943 ;
  assign n36945 = n5785 & n12313 ;
  assign n36946 = n27146 ^ n21790 ^ n16255 ;
  assign n36947 = ( n6952 & n9980 ) | ( n6952 & ~n36946 ) | ( n9980 & ~n36946 ) ;
  assign n36948 = n5204 & n33705 ;
  assign n36951 = n3140 & ~n10579 ;
  assign n36952 = n36951 ^ n8543 ^ 1'b0 ;
  assign n36949 = n7458 & n17563 ;
  assign n36950 = n10547 & ~n36949 ;
  assign n36953 = n36952 ^ n36950 ^ 1'b0 ;
  assign n36954 = n25284 ^ n21917 ^ 1'b0 ;
  assign n36955 = ( n36948 & n36953 ) | ( n36948 & n36954 ) | ( n36953 & n36954 ) ;
  assign n36956 = n2985 & n13157 ;
  assign n36957 = ~n2064 & n36956 ;
  assign n36958 = n36957 ^ n35612 ^ 1'b0 ;
  assign n36959 = n34779 ^ n17682 ^ n6224 ;
  assign n36960 = n15875 & ~n36959 ;
  assign n36961 = n871 & n6209 ;
  assign n36962 = n4465 & n36961 ;
  assign n36963 = n36962 ^ n15386 ^ n6512 ;
  assign n36964 = n31969 ^ n6132 ^ 1'b0 ;
  assign n36965 = ( n2325 & ~n33710 ) | ( n2325 & n36964 ) | ( ~n33710 & n36964 ) ;
  assign n36966 = n20370 & ~n25355 ;
  assign n36967 = ~n4389 & n36966 ;
  assign n36968 = n16749 & n36967 ;
  assign n36969 = x230 & ~n10890 ;
  assign n36970 = n36969 ^ n36850 ^ n23105 ;
  assign n36971 = n12240 | n19263 ;
  assign n36972 = x151 | n36971 ;
  assign n36973 = n27243 & n36972 ;
  assign n36974 = ~n36970 & n36973 ;
  assign n36975 = n31235 & ~n36974 ;
  assign n36976 = n36975 ^ n9073 ^ 1'b0 ;
  assign n36977 = n27428 ^ n13416 ^ 1'b0 ;
  assign n36978 = n29052 & n36977 ;
  assign n36979 = ( n639 & n31585 ) | ( n639 & n36978 ) | ( n31585 & n36978 ) ;
  assign n36980 = n7508 | n27003 ;
  assign n36981 = n4062 & ~n36980 ;
  assign n36982 = n9972 | n13405 ;
  assign n36983 = n13340 & n36982 ;
  assign n36984 = ~n8825 & n36983 ;
  assign n36985 = n1219 & ~n6362 ;
  assign n36986 = n36985 ^ n26260 ^ 1'b0 ;
  assign n36987 = ( n6361 & n20018 ) | ( n6361 & n36934 ) | ( n20018 & n36934 ) ;
  assign n36988 = ( n7217 & ~n9218 ) | ( n7217 & n21185 ) | ( ~n9218 & n21185 ) ;
  assign n36989 = n7428 & n12713 ;
  assign n36990 = ~n36988 & n36989 ;
  assign n36992 = n9149 ^ n9038 ^ 1'b0 ;
  assign n36993 = n1783 & n36992 ;
  assign n36991 = n22535 ^ n984 ^ 1'b0 ;
  assign n36994 = n36993 ^ n36991 ^ n24227 ;
  assign n36995 = n12578 ^ n6563 ^ 1'b0 ;
  assign n36996 = ~n36994 & n36995 ;
  assign n36997 = ( n12615 & ~n14653 ) | ( n12615 & n36996 ) | ( ~n14653 & n36996 ) ;
  assign n36998 = n18836 & ~n35528 ;
  assign n36999 = n23605 ^ n16163 ^ 1'b0 ;
  assign n37000 = ~n28513 & n36999 ;
  assign n37001 = n5025 & n37000 ;
  assign n37003 = n16116 ^ n4509 ^ 1'b0 ;
  assign n37004 = n37003 ^ n23427 ^ n12798 ;
  assign n37002 = ~n2498 & n11739 ;
  assign n37005 = n37004 ^ n37002 ^ 1'b0 ;
  assign n37006 = n21042 & ~n37005 ;
  assign n37007 = n6568 & ~n29177 ;
  assign n37008 = n37007 ^ n23024 ^ 1'b0 ;
  assign n37009 = ( n17083 & ~n19547 ) | ( n17083 & n37008 ) | ( ~n19547 & n37008 ) ;
  assign n37010 = ( n3167 & n4629 ) | ( n3167 & ~n21921 ) | ( n4629 & ~n21921 ) ;
  assign n37011 = n6897 & ~n15969 ;
  assign n37012 = n37010 | n37011 ;
  assign n37013 = n37012 ^ n1810 ^ 1'b0 ;
  assign n37014 = n25829 ^ n22581 ^ 1'b0 ;
  assign n37015 = n28699 ^ n28307 ^ n400 ;
  assign n37016 = n11941 & ~n37015 ;
  assign n37017 = ~n3757 & n37016 ;
  assign n37018 = n2284 & n3206 ;
  assign n37019 = ( n2843 & n14712 ) | ( n2843 & ~n30122 ) | ( n14712 & ~n30122 ) ;
  assign n37020 = n21999 ^ n9359 ^ 1'b0 ;
  assign n37021 = n15590 & ~n37020 ;
  assign n37022 = n6060 & ~n7022 ;
  assign n37023 = n37022 ^ n18995 ^ 1'b0 ;
  assign n37024 = n29529 ^ n8383 ^ 1'b0 ;
  assign n37025 = n4974 | n37024 ;
  assign n37026 = n29431 | n37025 ;
  assign n37027 = n37023 | n37026 ;
  assign n37028 = n15266 & n15792 ;
  assign n37029 = n16208 & n37028 ;
  assign n37030 = n29835 ^ n19990 ^ 1'b0 ;
  assign n37031 = n37030 ^ n21621 ^ n17095 ;
  assign n37032 = ~n37029 & n37031 ;
  assign n37033 = n36741 & n37032 ;
  assign n37036 = n17753 ^ n2382 ^ 1'b0 ;
  assign n37037 = n20769 & n37036 ;
  assign n37034 = n10454 ^ n5697 ^ n4794 ;
  assign n37035 = n23565 & ~n37034 ;
  assign n37038 = n37037 ^ n37035 ^ n7617 ;
  assign n37039 = n24627 ^ n19539 ^ n18506 ;
  assign n37040 = ( n1757 & ~n37038 ) | ( n1757 & n37039 ) | ( ~n37038 & n37039 ) ;
  assign n37041 = n806 & ~n957 ;
  assign n37042 = ~n25941 & n37041 ;
  assign n37043 = n37042 ^ n4620 ^ 1'b0 ;
  assign n37044 = ( n1867 & n9279 ) | ( n1867 & n37043 ) | ( n9279 & n37043 ) ;
  assign n37045 = n7255 ^ n6931 ^ n1197 ;
  assign n37046 = n37045 ^ n10875 ^ n1192 ;
  assign n37047 = n257 & n37046 ;
  assign n37048 = n31502 & n37047 ;
  assign n37049 = ~n7192 & n37048 ;
  assign n37050 = n18651 | n26257 ;
  assign n37051 = ~n8088 & n37050 ;
  assign n37052 = ~n15296 & n17201 ;
  assign n37053 = n19623 & n37052 ;
  assign n37054 = n10934 | n16442 ;
  assign n37055 = n37054 ^ n35830 ^ 1'b0 ;
  assign n37056 = n37053 | n37055 ;
  assign n37057 = n15410 & n28906 ;
  assign n37058 = n19999 & n37057 ;
  assign n37059 = n33172 ^ n27487 ^ n22879 ;
  assign n37060 = n25841 ^ n18536 ^ n7081 ;
  assign n37061 = n37060 ^ n36761 ^ n2221 ;
  assign n37063 = n2606 & n3687 ;
  assign n37064 = ~n3687 & n37063 ;
  assign n37065 = n37064 ^ n6245 ^ 1'b0 ;
  assign n37066 = n37065 ^ n3549 ^ 1'b0 ;
  assign n37067 = n13579 & n37066 ;
  assign n37062 = n1635 & ~n4910 ;
  assign n37068 = n37067 ^ n37062 ^ 1'b0 ;
  assign n37070 = n434 & n35058 ;
  assign n37071 = n4134 & n37070 ;
  assign n37069 = n4819 & ~n10797 ;
  assign n37072 = n37071 ^ n37069 ^ 1'b0 ;
  assign n37075 = n3918 & n19107 ;
  assign n37074 = n28188 ^ n26693 ^ 1'b0 ;
  assign n37073 = n13563 & ~n20517 ;
  assign n37076 = n37075 ^ n37074 ^ n37073 ;
  assign n37077 = n26205 & ~n37076 ;
  assign n37078 = n37077 ^ n583 ^ 1'b0 ;
  assign n37079 = ~n5941 & n33542 ;
  assign n37080 = ( n11586 & n31881 ) | ( n11586 & n34566 ) | ( n31881 & n34566 ) ;
  assign n37081 = ( ~n28904 & n37079 ) | ( ~n28904 & n37080 ) | ( n37079 & n37080 ) ;
  assign n37083 = n23456 ^ n14858 ^ 1'b0 ;
  assign n37084 = n3502 | n37083 ;
  assign n37082 = ~x213 & n3107 ;
  assign n37085 = n37084 ^ n37082 ^ n9037 ;
  assign n37086 = n37085 ^ n5863 ^ 1'b0 ;
  assign n37087 = n28405 | n37086 ;
  assign n37088 = n37087 ^ n25592 ^ n18917 ;
  assign n37090 = n18289 & n22181 ;
  assign n37089 = n1366 & n13051 ;
  assign n37091 = n37090 ^ n37089 ^ n10018 ;
  assign n37092 = n37091 ^ n35249 ^ 1'b0 ;
  assign n37093 = n25858 & ~n37092 ;
  assign n37094 = n8120 & n22144 ;
  assign n37095 = n37094 ^ n3381 ^ 1'b0 ;
  assign n37096 = n6329 & ~n37095 ;
  assign n37097 = n29660 ^ n24056 ^ n17697 ;
  assign n37098 = ( ~n19571 & n29297 ) | ( ~n19571 & n37097 ) | ( n29297 & n37097 ) ;
  assign n37099 = x91 & n14364 ;
  assign n37100 = n37099 ^ n7593 ^ 1'b0 ;
  assign n37101 = n17508 | n37100 ;
  assign n37102 = n37101 ^ n5642 ^ 1'b0 ;
  assign n37103 = n21367 & n29582 ;
  assign n37104 = n37103 ^ n15927 ^ 1'b0 ;
  assign n37105 = ~n5242 & n16618 ;
  assign n37106 = n37105 ^ n20894 ^ 1'b0 ;
  assign n37107 = n37106 ^ n33713 ^ 1'b0 ;
  assign n37109 = n8955 & n24962 ;
  assign n37108 = n10760 ^ n3302 ^ n2403 ;
  assign n37110 = n37109 ^ n37108 ^ 1'b0 ;
  assign n37111 = n6555 ^ n5767 ^ 1'b0 ;
  assign n37112 = ~x3 & n16361 ;
  assign n37113 = n9456 & ~n37112 ;
  assign n37114 = ( n5913 & n37111 ) | ( n5913 & ~n37113 ) | ( n37111 & ~n37113 ) ;
  assign n37115 = n25501 ^ n2531 ^ x45 ;
  assign n37116 = ~n23106 & n25396 ;
  assign n37117 = ~n30579 & n37116 ;
  assign n37118 = n23106 ^ n20473 ^ n4081 ;
  assign n37119 = n1654 & n37118 ;
  assign n37120 = n5973 & n37119 ;
  assign n37121 = n16732 ^ n15258 ^ n7174 ;
  assign n37122 = n25771 | n26793 ;
  assign n37123 = n28443 & ~n37122 ;
  assign n37124 = n4535 | n37123 ;
  assign n37125 = n22457 | n37124 ;
  assign n37126 = ~n6527 & n37125 ;
  assign n37127 = ~n19973 & n37126 ;
  assign n37128 = n15839 & ~n18865 ;
  assign n37129 = n17517 & n37128 ;
  assign n37130 = ~n9949 & n19494 ;
  assign n37131 = ( ~n6169 & n19937 ) | ( ~n6169 & n37130 ) | ( n19937 & n37130 ) ;
  assign n37132 = n26457 ^ n17531 ^ 1'b0 ;
  assign n37133 = n2530 & ~n37132 ;
  assign n37134 = n10073 & ~n37133 ;
  assign n37135 = n23474 ^ n9416 ^ n944 ;
  assign n37136 = n20956 ^ n14492 ^ n2497 ;
  assign n37137 = n7323 ^ n6761 ^ n1011 ;
  assign n37138 = n37137 ^ n11459 ^ n8792 ;
  assign n37139 = n37138 ^ n6787 ^ n3334 ;
  assign n37140 = n11018 ^ n4134 ^ n262 ;
  assign n37141 = ( ~n6160 & n20077 ) | ( ~n6160 & n37140 ) | ( n20077 & n37140 ) ;
  assign n37142 = n37141 ^ n19901 ^ 1'b0 ;
  assign n37143 = n4315 | n37142 ;
  assign n37144 = ( n1004 & n6311 ) | ( n1004 & ~n10174 ) | ( n6311 & ~n10174 ) ;
  assign n37145 = n34599 ^ n20035 ^ n471 ;
  assign n37146 = n37144 & n37145 ;
  assign n37147 = n37146 ^ n36850 ^ 1'b0 ;
  assign n37148 = n18440 ^ n13812 ^ 1'b0 ;
  assign n37149 = ( n4112 & ~n10391 ) | ( n4112 & n12524 ) | ( ~n10391 & n12524 ) ;
  assign n37150 = n37149 ^ n33139 ^ n20339 ;
  assign n37151 = n12952 | n37150 ;
  assign n37152 = n31588 ^ n11638 ^ 1'b0 ;
  assign n37153 = n11169 & ~n37152 ;
  assign n37154 = n37153 ^ n3062 ^ n1220 ;
  assign n37158 = n30807 ^ n5167 ^ n3682 ;
  assign n37155 = n5438 & n6427 ;
  assign n37156 = n28693 ^ n23086 ^ n13866 ;
  assign n37157 = ~n37155 & n37156 ;
  assign n37159 = n37158 ^ n37157 ^ 1'b0 ;
  assign n37161 = ( x73 & ~n2680 ) | ( x73 & n24052 ) | ( ~n2680 & n24052 ) ;
  assign n37160 = ~n16271 & n36320 ;
  assign n37162 = n37161 ^ n37160 ^ 1'b0 ;
  assign n37163 = ~x206 & n3268 ;
  assign n37164 = x241 & ~n9849 ;
  assign n37165 = n37164 ^ n32272 ^ 1'b0 ;
  assign n37166 = n37165 ^ n2944 ^ 1'b0 ;
  assign n37167 = ~n1744 & n4790 ;
  assign n37168 = n24257 | n31950 ;
  assign n37169 = n37167 & ~n37168 ;
  assign n37170 = n13873 | n36755 ;
  assign n37171 = ( n9438 & ~n12387 ) | ( n9438 & n15221 ) | ( ~n12387 & n15221 ) ;
  assign n37172 = n1595 & ~n18978 ;
  assign n37173 = n12258 | n29548 ;
  assign n37174 = n37172 | n37173 ;
  assign n37175 = ~n20514 & n37174 ;
  assign n37176 = n37171 & n37175 ;
  assign n37177 = n2567 & n37176 ;
  assign n37178 = n4327 & ~n15953 ;
  assign n37179 = n37178 ^ n34717 ^ 1'b0 ;
  assign n37180 = n21913 & ~n35189 ;
  assign n37181 = n22133 & n37180 ;
  assign n37182 = n17463 ^ n14590 ^ 1'b0 ;
  assign n37183 = n1395 & n37182 ;
  assign n37184 = n27873 & n37183 ;
  assign n37185 = n3487 & n29225 ;
  assign n37186 = n37185 ^ n4638 ^ 1'b0 ;
  assign n37187 = ( n1109 & n30315 ) | ( n1109 & ~n37186 ) | ( n30315 & ~n37186 ) ;
  assign n37188 = n30645 ^ n12685 ^ n2712 ;
  assign n37189 = ( n10633 & n24226 ) | ( n10633 & ~n37188 ) | ( n24226 & ~n37188 ) ;
  assign n37194 = n1750 | n13145 ;
  assign n37195 = ( n6115 & n19847 ) | ( n6115 & ~n37194 ) | ( n19847 & ~n37194 ) ;
  assign n37190 = n26115 ^ n5030 ^ 1'b0 ;
  assign n37191 = n37190 ^ n9274 ^ 1'b0 ;
  assign n37192 = ~n14273 & n37191 ;
  assign n37193 = n3095 & ~n37192 ;
  assign n37196 = n37195 ^ n37193 ^ n23319 ;
  assign n37197 = n31871 ^ n14829 ^ 1'b0 ;
  assign n37198 = n23550 ^ n8056 ^ n3438 ;
  assign n37199 = n7500 & ~n28259 ;
  assign n37200 = n11248 ^ n1281 ^ 1'b0 ;
  assign n37201 = ~n16654 & n37200 ;
  assign n37202 = n16848 | n37201 ;
  assign n37203 = ~n8056 & n27229 ;
  assign n37204 = ~n3791 & n37203 ;
  assign n37205 = n9076 ^ n4446 ^ 1'b0 ;
  assign n37206 = n4833 & n32198 ;
  assign n37207 = n37206 ^ n18796 ^ 1'b0 ;
  assign n37208 = n8307 | n11230 ;
  assign n37209 = n37208 ^ n34797 ^ n20515 ;
  assign n37210 = n11587 ^ n2262 ^ 1'b0 ;
  assign n37211 = n3889 & n37210 ;
  assign n37212 = n37211 ^ n3951 ^ n462 ;
  assign n37213 = ~n6030 & n37212 ;
  assign n37218 = n12087 ^ n10509 ^ n9632 ;
  assign n37215 = n8930 & n14578 ;
  assign n37216 = ~x223 & n37215 ;
  assign n37214 = n13251 ^ n8203 ^ 1'b0 ;
  assign n37217 = n37216 ^ n37214 ^ n1837 ;
  assign n37219 = n37218 ^ n37217 ^ n14008 ;
  assign n37220 = n649 & ~n21927 ;
  assign n37221 = n37220 ^ n26834 ^ 1'b0 ;
  assign n37222 = n15932 & n26036 ;
  assign n37223 = n32211 & n37222 ;
  assign n37224 = ( n9087 & n16003 ) | ( n9087 & ~n16319 ) | ( n16003 & ~n16319 ) ;
  assign n37225 = n23573 & ~n37224 ;
  assign n37226 = ~n12400 & n37225 ;
  assign n37227 = n19290 ^ n7698 ^ n6862 ;
  assign n37228 = n17408 & ~n37227 ;
  assign n37229 = n37228 ^ n5741 ^ 1'b0 ;
  assign n37232 = n18387 ^ n10240 ^ 1'b0 ;
  assign n37230 = n26237 & ~n34074 ;
  assign n37231 = n37230 ^ n11962 ^ 1'b0 ;
  assign n37233 = n37232 ^ n37231 ^ n21396 ;
  assign n37234 = ( n7892 & n29138 ) | ( n7892 & ~n32043 ) | ( n29138 & ~n32043 ) ;
  assign n37235 = n4806 & ~n34062 ;
  assign n37236 = n25982 & n37235 ;
  assign n37237 = ~n13593 & n16120 ;
  assign n37238 = n37237 ^ n4773 ^ 1'b0 ;
  assign n37239 = n3035 & ~n37238 ;
  assign n37240 = n11693 & n37239 ;
  assign n37241 = n8167 | n8498 ;
  assign n37242 = n37241 ^ n12646 ^ 1'b0 ;
  assign n37243 = ~n1985 & n9321 ;
  assign n37244 = n17317 & n37243 ;
  assign n37246 = n27978 ^ n26123 ^ n12549 ;
  assign n37247 = ( n13714 & n30689 ) | ( n13714 & ~n37246 ) | ( n30689 & ~n37246 ) ;
  assign n37245 = n3559 & ~n37137 ;
  assign n37248 = n37247 ^ n37245 ^ 1'b0 ;
  assign n37249 = n11171 ^ n5107 ^ 1'b0 ;
  assign n37250 = ~n9756 & n37249 ;
  assign n37251 = n14945 & ~n31621 ;
  assign n37252 = ~n37250 & n37251 ;
  assign n37253 = n29563 & ~n37252 ;
  assign n37254 = n17347 ^ n11825 ^ n9766 ;
  assign n37255 = n6744 ^ n2168 ^ 1'b0 ;
  assign n37256 = n37255 ^ n12087 ^ 1'b0 ;
  assign n37257 = ~n10527 & n37256 ;
  assign n37258 = n7584 & n19465 ;
  assign n37259 = n6612 & n37258 ;
  assign n37260 = ( n584 & n5907 ) | ( n584 & ~n34192 ) | ( n5907 & ~n34192 ) ;
  assign n37261 = ( n1948 & n11230 ) | ( n1948 & n12556 ) | ( n11230 & n12556 ) ;
  assign n37262 = n23488 ^ n9839 ^ 1'b0 ;
  assign n37263 = x221 & ~n37262 ;
  assign n37264 = ~n25568 & n32476 ;
  assign n37265 = ~n1923 & n37264 ;
  assign n37266 = ~n2865 & n37265 ;
  assign n37267 = n5872 & ~n17924 ;
  assign n37268 = n37267 ^ n28225 ^ 1'b0 ;
  assign n37269 = n2028 | n3578 ;
  assign n37270 = n37269 ^ n28376 ^ 1'b0 ;
  assign n37271 = n13636 ^ n13101 ^ 1'b0 ;
  assign n37272 = n12249 & n37271 ;
  assign n37273 = n10039 & n37272 ;
  assign n37274 = ~n25061 & n27042 ;
  assign n37275 = n22008 & ~n29031 ;
  assign n37280 = ~n6423 & n6479 ;
  assign n37281 = n23137 & n37280 ;
  assign n37278 = n19858 ^ n2254 ^ 1'b0 ;
  assign n37279 = ~n19544 & n37278 ;
  assign n37276 = ( n2411 & n3945 ) | ( n2411 & n33344 ) | ( n3945 & n33344 ) ;
  assign n37277 = n37276 ^ n14396 ^ n4952 ;
  assign n37282 = n37281 ^ n37279 ^ n37277 ;
  assign n37283 = n15525 & n16888 ;
  assign n37284 = n25073 ^ n11597 ^ n8259 ;
  assign n37285 = n1866 & n37284 ;
  assign n37286 = n37285 ^ n18229 ^ 1'b0 ;
  assign n37287 = n31905 ^ n11099 ^ 1'b0 ;
  assign n37288 = n37286 | n37287 ;
  assign n37289 = n12993 ^ n10665 ^ 1'b0 ;
  assign n37290 = n10797 | n37289 ;
  assign n37291 = ( n4325 & n5362 ) | ( n4325 & ~n37290 ) | ( n5362 & ~n37290 ) ;
  assign n37292 = n31908 ^ n23486 ^ 1'b0 ;
  assign n37293 = n16616 ^ n8159 ^ 1'b0 ;
  assign n37294 = n5988 ^ x68 ^ 1'b0 ;
  assign n37295 = ~n15290 & n37294 ;
  assign n37296 = n6869 | n10942 ;
  assign n37297 = n37295 | n37296 ;
  assign n37298 = ~n26979 & n32720 ;
  assign n37299 = ~n12817 & n37298 ;
  assign n37302 = n14276 ^ n10650 ^ 1'b0 ;
  assign n37300 = ~n5169 & n8817 ;
  assign n37301 = n37300 ^ n32272 ^ n16922 ;
  assign n37303 = n37302 ^ n37301 ^ n5493 ;
  assign n37304 = n17203 ^ n756 ^ 1'b0 ;
  assign n37305 = n9217 & ~n37304 ;
  assign n37306 = n28238 ^ n19989 ^ n14741 ;
  assign n37307 = n35868 ^ n15418 ^ x231 ;
  assign n37308 = ( n37305 & ~n37306 ) | ( n37305 & n37307 ) | ( ~n37306 & n37307 ) ;
  assign n37309 = n2700 & n8497 ;
  assign n37310 = ( n3006 & ~n35726 ) | ( n3006 & n37309 ) | ( ~n35726 & n37309 ) ;
  assign n37311 = n32694 ^ n17510 ^ 1'b0 ;
  assign n37312 = ~n324 & n37311 ;
  assign n37313 = n37312 ^ n4866 ^ 1'b0 ;
  assign n37314 = n9064 & ~n37313 ;
  assign n37315 = n36415 ^ n4517 ^ 1'b0 ;
  assign n37316 = n37314 & n37315 ;
  assign n37317 = n3742 & ~n20041 ;
  assign n37318 = n37317 ^ n4043 ^ 1'b0 ;
  assign n37319 = n6740 & ~n37318 ;
  assign n37320 = n17560 & n37319 ;
  assign n37321 = ~n6660 & n7422 ;
  assign n37322 = n11937 & n37321 ;
  assign n37323 = n37322 ^ n4276 ^ 1'b0 ;
  assign n37324 = n37323 ^ n22564 ^ 1'b0 ;
  assign n37325 = n23087 ^ n19264 ^ 1'b0 ;
  assign n37326 = n30515 | n37325 ;
  assign n37329 = n11155 ^ n1888 ^ n1808 ;
  assign n37327 = n26182 ^ n18652 ^ n409 ;
  assign n37328 = n1204 & n37327 ;
  assign n37330 = n37329 ^ n37328 ^ 1'b0 ;
  assign n37331 = n977 | n7752 ;
  assign n37332 = n9054 & ~n37331 ;
  assign n37333 = n37332 ^ n33988 ^ n2333 ;
  assign n37334 = ~n7510 & n37333 ;
  assign n37335 = n37334 ^ n10267 ^ 1'b0 ;
  assign n37336 = ( ~n12314 & n22107 ) | ( ~n12314 & n32963 ) | ( n22107 & n32963 ) ;
  assign n37337 = n28961 ^ n14765 ^ n280 ;
  assign n37338 = n20298 ^ x5 ^ 1'b0 ;
  assign n37339 = x145 & n37338 ;
  assign n37340 = n37339 ^ n23738 ^ 1'b0 ;
  assign n37341 = n10645 ^ n8350 ^ n2217 ;
  assign n37342 = n20105 ^ n8805 ^ 1'b0 ;
  assign n37343 = n22113 & n37342 ;
  assign n37344 = n37343 ^ n20889 ^ 1'b0 ;
  assign n37345 = n12675 & n37344 ;
  assign n37346 = n37345 ^ n4808 ^ 1'b0 ;
  assign n37347 = n21994 ^ n961 ^ 1'b0 ;
  assign n37348 = n22674 ^ n4073 ^ 1'b0 ;
  assign n37349 = n9551 & n37348 ;
  assign n37350 = n4026 & n8430 ;
  assign n37351 = ~n7621 & n12269 ;
  assign n37352 = n14956 & n37351 ;
  assign n37353 = ( n22390 & n33241 ) | ( n22390 & n37352 ) | ( n33241 & n37352 ) ;
  assign n37354 = n24982 ^ n15771 ^ 1'b0 ;
  assign n37355 = ( n12773 & n33052 ) | ( n12773 & ~n37354 ) | ( n33052 & ~n37354 ) ;
  assign n37356 = n12147 ^ n11907 ^ n4564 ;
  assign n37357 = n1776 | n1851 ;
  assign n37358 = n17768 | n37357 ;
  assign n37359 = n37358 ^ n8382 ^ 1'b0 ;
  assign n37360 = n24868 ^ n11230 ^ 1'b0 ;
  assign n37361 = n15953 ^ n4812 ^ n968 ;
  assign n37362 = n15925 & ~n27141 ;
  assign n37363 = n37362 ^ n1199 ^ 1'b0 ;
  assign n37364 = ( ~n7843 & n37361 ) | ( ~n7843 & n37363 ) | ( n37361 & n37363 ) ;
  assign n37365 = n18245 | n32902 ;
  assign n37366 = n17505 ^ n16170 ^ n9578 ;
  assign n37367 = n31861 | n37366 ;
  assign n37368 = ~n3814 & n18783 ;
  assign n37369 = n37368 ^ n23809 ^ 1'b0 ;
  assign n37370 = n6825 & n7584 ;
  assign n37371 = n37370 ^ n19959 ^ n11806 ;
  assign n37372 = n37371 ^ n24275 ^ 1'b0 ;
  assign n37373 = ~n7581 & n15473 ;
  assign n37374 = n2531 & n37373 ;
  assign n37375 = n37374 ^ n28588 ^ n1309 ;
  assign n37376 = ( n8716 & ~n14047 ) | ( n8716 & n25444 ) | ( ~n14047 & n25444 ) ;
  assign n37377 = ( n7867 & n14139 ) | ( n7867 & n31504 ) | ( n14139 & n31504 ) ;
  assign n37378 = n31631 ^ n11174 ^ 1'b0 ;
  assign n37379 = n21049 ^ n3317 ^ 1'b0 ;
  assign n37380 = x202 & ~n37379 ;
  assign n37381 = n7238 & n37380 ;
  assign n37382 = n26760 ^ n13185 ^ n3712 ;
  assign n37383 = ( n1239 & n8930 ) | ( n1239 & n27618 ) | ( n8930 & n27618 ) ;
  assign n37384 = n3289 & n23784 ;
  assign n37385 = n15507 & ~n19854 ;
  assign n37386 = n37385 ^ n3362 ^ 1'b0 ;
  assign n37387 = n37386 ^ n31489 ^ n11022 ;
  assign n37388 = n37387 ^ n6950 ^ n5551 ;
  assign n37389 = n4501 ^ n627 ^ 1'b0 ;
  assign n37390 = ~n3520 & n37389 ;
  assign n37391 = n25587 & n37390 ;
  assign n37392 = n37391 ^ n33688 ^ 1'b0 ;
  assign n37393 = n1554 & ~n37392 ;
  assign n37394 = ~n8842 & n29217 ;
  assign n37395 = n2633 & n37394 ;
  assign n37396 = n10633 | n37395 ;
  assign n37397 = n28583 ^ n26007 ^ n23987 ;
  assign n37398 = n35462 ^ n11822 ^ n10706 ;
  assign n37399 = n22324 ^ n8942 ^ 1'b0 ;
  assign n37400 = ~n20331 & n37399 ;
  assign n37401 = n20947 & n21363 ;
  assign n37402 = n5533 & n37401 ;
  assign n37403 = n12404 ^ n6750 ^ 1'b0 ;
  assign n37405 = n3305 | n26288 ;
  assign n37406 = ( n7678 & ~n11914 ) | ( n7678 & n37405 ) | ( ~n11914 & n37405 ) ;
  assign n37407 = ( ~n5817 & n14749 ) | ( ~n5817 & n37406 ) | ( n14749 & n37406 ) ;
  assign n37404 = n7894 & ~n20349 ;
  assign n37408 = n37407 ^ n37404 ^ 1'b0 ;
  assign n37409 = n16766 & ~n32015 ;
  assign n37411 = ~n5169 & n11192 ;
  assign n37412 = ~n29625 & n37411 ;
  assign n37410 = n20169 | n20696 ;
  assign n37413 = n37412 ^ n37410 ^ 1'b0 ;
  assign n37414 = n16102 ^ n11319 ^ 1'b0 ;
  assign n37415 = n37414 ^ n25663 ^ 1'b0 ;
  assign n37416 = n20516 ^ n17230 ^ 1'b0 ;
  assign n37417 = n16626 ^ n15857 ^ n4057 ;
  assign n37418 = ( n15961 & n23375 ) | ( n15961 & n37417 ) | ( n23375 & n37417 ) ;
  assign n37419 = n16915 ^ n15950 ^ 1'b0 ;
  assign n37420 = n30724 & ~n37419 ;
  assign n37421 = n9671 & n23416 ;
  assign n37424 = n15657 ^ n7204 ^ 1'b0 ;
  assign n37422 = n12385 & ~n28526 ;
  assign n37423 = n32993 & ~n37422 ;
  assign n37425 = n37424 ^ n37423 ^ 1'b0 ;
  assign n37426 = ~x161 & n20855 ;
  assign n37427 = n37426 ^ n4169 ^ n3292 ;
  assign n37430 = n22683 ^ n10191 ^ n753 ;
  assign n37431 = ( n7424 & ~n9274 ) | ( n7424 & n37430 ) | ( ~n9274 & n37430 ) ;
  assign n37429 = n448 | n2769 ;
  assign n37432 = n37431 ^ n37429 ^ 1'b0 ;
  assign n37428 = n32291 & n33866 ;
  assign n37433 = n37432 ^ n37428 ^ 1'b0 ;
  assign n37434 = ( n22486 & n37427 ) | ( n22486 & n37433 ) | ( n37427 & n37433 ) ;
  assign n37435 = n25171 ^ n13768 ^ n12406 ;
  assign n37436 = n37435 ^ n32007 ^ 1'b0 ;
  assign n37437 = ( n4461 & n4842 ) | ( n4461 & ~n26693 ) | ( n4842 & ~n26693 ) ;
  assign n37438 = n7707 & ~n15630 ;
  assign n37439 = ~n12826 & n13745 ;
  assign n37440 = ~n8942 & n37439 ;
  assign n37443 = n33743 ^ n5162 ^ 1'b0 ;
  assign n37441 = ( n16466 & n29259 ) | ( n16466 & n30425 ) | ( n29259 & n30425 ) ;
  assign n37442 = n19424 & ~n37441 ;
  assign n37444 = n37443 ^ n37442 ^ 1'b0 ;
  assign n37445 = n23144 ^ n17934 ^ n9892 ;
  assign n37446 = ~n1352 & n12741 ;
  assign n37447 = n19573 & n37446 ;
  assign n37448 = n29671 ^ n22395 ^ 1'b0 ;
  assign n37449 = n2869 & n37448 ;
  assign n37450 = n23008 ^ n17648 ^ 1'b0 ;
  assign n37451 = n5716 & ~n9131 ;
  assign n37452 = n37451 ^ n2355 ^ 1'b0 ;
  assign n37453 = n12741 & ~n24091 ;
  assign n37454 = ~n5165 & n37453 ;
  assign n37455 = ( n3915 & n20556 ) | ( n3915 & n37454 ) | ( n20556 & n37454 ) ;
  assign n37456 = n37455 ^ n36326 ^ n5343 ;
  assign n37457 = n29053 ^ n940 ^ 1'b0 ;
  assign n37458 = ( n3874 & n25896 ) | ( n3874 & n37457 ) | ( n25896 & n37457 ) ;
  assign n37459 = n37458 ^ n6321 ^ 1'b0 ;
  assign n37460 = n5074 | n12940 ;
  assign n37461 = n25528 & ~n26000 ;
  assign n37462 = n25201 ^ x201 ^ 1'b0 ;
  assign n37463 = n1297 | n37462 ;
  assign n37464 = ( n908 & n10249 ) | ( n908 & n18636 ) | ( n10249 & n18636 ) ;
  assign n37465 = n23682 & ~n37464 ;
  assign n37466 = n37465 ^ n19849 ^ 1'b0 ;
  assign n37467 = n8128 | n37466 ;
  assign n37468 = n25195 ^ n21062 ^ 1'b0 ;
  assign n37469 = n2883 ^ n2571 ^ n883 ;
  assign n37470 = n37469 ^ n21314 ^ n14802 ;
  assign n37471 = n12434 ^ n5447 ^ n3290 ;
  assign n37473 = ( n1117 & ~n1821 ) | ( n1117 & n12042 ) | ( ~n1821 & n12042 ) ;
  assign n37472 = n25112 ^ n4214 ^ 1'b0 ;
  assign n37474 = n37473 ^ n37472 ^ n26173 ;
  assign n37475 = n37471 & n37474 ;
  assign n37476 = n6478 | n27302 ;
  assign n37477 = n37475 | n37476 ;
  assign n37478 = n8156 ^ n5222 ^ 1'b0 ;
  assign n37479 = n870 | n37478 ;
  assign n37480 = n5763 & n16183 ;
  assign n37481 = n36118 ^ n25930 ^ 1'b0 ;
  assign n37484 = n4595 & ~n14737 ;
  assign n37485 = ~n7386 & n37484 ;
  assign n37482 = n7136 & n24597 ;
  assign n37483 = n37482 ^ n14395 ^ 1'b0 ;
  assign n37486 = n37485 ^ n37483 ^ n1779 ;
  assign n37487 = n9113 ^ n5794 ^ 1'b0 ;
  assign n37488 = n37487 ^ n23042 ^ 1'b0 ;
  assign n37489 = n10037 & n37488 ;
  assign n37490 = n25882 & n37489 ;
  assign n37491 = n15258 | n25071 ;
  assign n37492 = n37491 ^ n13216 ^ 1'b0 ;
  assign n37493 = n37091 ^ n22181 ^ n3839 ;
  assign n37494 = n37493 ^ n23646 ^ 1'b0 ;
  assign n37495 = n37492 | n37494 ;
  assign n37496 = n35931 ^ n1042 ^ 1'b0 ;
  assign n37497 = ~n7204 & n37496 ;
  assign n37498 = ~n28330 & n37497 ;
  assign n37499 = ( n9084 & n11411 ) | ( n9084 & n29489 ) | ( n11411 & n29489 ) ;
  assign n37501 = ( n2884 & n3712 ) | ( n2884 & n13544 ) | ( n3712 & n13544 ) ;
  assign n37500 = n3120 & ~n13694 ;
  assign n37502 = n37501 ^ n37500 ^ n4331 ;
  assign n37503 = n33498 ^ n6111 ^ 1'b0 ;
  assign n37504 = n4060 ^ n441 ^ 1'b0 ;
  assign n37505 = n33632 ^ n4093 ^ 1'b0 ;
  assign n37506 = ~n37504 & n37505 ;
  assign n37507 = n2802 & n37506 ;
  assign n37508 = n28988 ^ n24885 ^ 1'b0 ;
  assign n37509 = n32469 & ~n37508 ;
  assign n37510 = n3844 | n9807 ;
  assign n37511 = n30118 | n37510 ;
  assign n37512 = n37511 ^ n32618 ^ n13342 ;
  assign n37513 = ( n11620 & n23430 ) | ( n11620 & ~n32700 ) | ( n23430 & ~n32700 ) ;
  assign n37514 = n5367 ^ n2349 ^ 1'b0 ;
  assign n37515 = n37514 ^ n15256 ^ n1352 ;
  assign n37516 = n21166 ^ n16804 ^ 1'b0 ;
  assign n37517 = ~n28635 & n32932 ;
  assign n37518 = n37517 ^ n6486 ^ 1'b0 ;
  assign n37519 = n6188 & n6831 ;
  assign n37520 = n37519 ^ n32133 ^ 1'b0 ;
  assign n37521 = n32953 ^ n23755 ^ 1'b0 ;
  assign n37522 = n16459 | n37521 ;
  assign n37523 = n21968 ^ x213 ^ 1'b0 ;
  assign n37524 = ( n875 & ~n3157 ) | ( n875 & n31980 ) | ( ~n3157 & n31980 ) ;
  assign n37525 = n11414 ^ n607 ^ 1'b0 ;
  assign n37526 = n37524 & ~n37525 ;
  assign n37527 = n37526 ^ n13556 ^ 1'b0 ;
  assign n37529 = n7909 & ~n14522 ;
  assign n37530 = n5966 & n37529 ;
  assign n37528 = n14601 ^ n7590 ^ 1'b0 ;
  assign n37531 = n37530 ^ n37528 ^ n10387 ;
  assign n37532 = ~x68 & n23015 ;
  assign n37533 = n21823 ^ n16680 ^ n16351 ;
  assign n37534 = n37533 ^ n15649 ^ 1'b0 ;
  assign n37535 = n35844 & n37534 ;
  assign n37536 = ~n26968 & n37535 ;
  assign n37537 = n14996 | n33929 ;
  assign n37538 = n37537 ^ n11467 ^ 1'b0 ;
  assign n37539 = n37227 ^ n28325 ^ n27494 ;
  assign n37542 = n6575 ^ n3707 ^ 1'b0 ;
  assign n37543 = n3946 | n37542 ;
  assign n37544 = ~n19193 & n37543 ;
  assign n37540 = ( n737 & ~n3992 ) | ( n737 & n6303 ) | ( ~n3992 & n6303 ) ;
  assign n37541 = n37540 ^ n2592 ^ 1'b0 ;
  assign n37545 = n37544 ^ n37541 ^ n24513 ;
  assign n37546 = ~n1311 & n14050 ;
  assign n37547 = n37546 ^ n35346 ^ n35096 ;
  assign n37548 = n13242 ^ n598 ^ 1'b0 ;
  assign n37549 = n37172 ^ n7369 ^ 1'b0 ;
  assign n37550 = n37060 ^ n20510 ^ n18531 ;
  assign n37551 = n6433 & ~n8105 ;
  assign n37552 = ( n4593 & n24740 ) | ( n4593 & n37551 ) | ( n24740 & n37551 ) ;
  assign n37553 = n37552 ^ n26708 ^ n4585 ;
  assign n37554 = x46 & n15398 ;
  assign n37555 = n37554 ^ n24961 ^ n1430 ;
  assign n37556 = ( n9500 & n13755 ) | ( n9500 & n18481 ) | ( n13755 & n18481 ) ;
  assign n37560 = n22983 ^ n19500 ^ n6644 ;
  assign n37557 = n4137 & ~n24109 ;
  assign n37558 = ~n16957 & n37557 ;
  assign n37559 = n37558 ^ n27325 ^ 1'b0 ;
  assign n37561 = n37560 ^ n37559 ^ n4816 ;
  assign n37562 = ( n27376 & ~n37556 ) | ( n27376 & n37561 ) | ( ~n37556 & n37561 ) ;
  assign n37563 = n16495 ^ n7831 ^ 1'b0 ;
  assign n37564 = n20353 | n37563 ;
  assign n37565 = ( n4450 & n5707 ) | ( n4450 & ~n22488 ) | ( n5707 & ~n22488 ) ;
  assign n37566 = n37565 ^ n23141 ^ 1'b0 ;
  assign n37567 = n37564 | n37566 ;
  assign n37568 = ( n1385 & ~n6143 ) | ( n1385 & n19483 ) | ( ~n6143 & n19483 ) ;
  assign n37569 = n37568 ^ n2201 ^ n2187 ;
  assign n37570 = n37569 ^ n24147 ^ n13859 ;
  assign n37571 = n8414 & n37570 ;
  assign n37572 = n1873 & n37571 ;
  assign n37573 = ( x248 & n19953 ) | ( x248 & n37572 ) | ( n19953 & n37572 ) ;
  assign n37574 = ~n7371 & n32922 ;
  assign n37575 = n23922 | n37574 ;
  assign n37576 = ( ~n1838 & n16412 ) | ( ~n1838 & n37384 ) | ( n16412 & n37384 ) ;
  assign n37577 = n3583 | n21533 ;
  assign n37578 = n37577 ^ n13655 ^ 1'b0 ;
  assign n37579 = n37578 ^ n18612 ^ 1'b0 ;
  assign n37580 = n9825 | n20336 ;
  assign n37581 = n10050 | n18187 ;
  assign n37582 = ( ~n31790 & n37580 ) | ( ~n31790 & n37581 ) | ( n37580 & n37581 ) ;
  assign n37583 = n2386 & ~n28022 ;
  assign n37584 = n5217 & n37583 ;
  assign n37585 = n37584 ^ n16049 ^ 1'b0 ;
  assign n37586 = n12417 | n37585 ;
  assign n37587 = n37586 ^ n8549 ^ 1'b0 ;
  assign n37588 = ~n4398 & n37587 ;
  assign n37589 = ( ~n1588 & n5352 ) | ( ~n1588 & n12895 ) | ( n5352 & n12895 ) ;
  assign n37590 = n5653 & ~n9554 ;
  assign n37591 = ~n831 & n37590 ;
  assign n37592 = ( n3694 & n5839 ) | ( n3694 & n11082 ) | ( n5839 & n11082 ) ;
  assign n37593 = n7127 | n26327 ;
  assign n37594 = n37592 & ~n37593 ;
  assign n37595 = n37594 ^ n27281 ^ 1'b0 ;
  assign n37596 = n6776 & ~n31286 ;
  assign n37597 = n37596 ^ n698 ^ 1'b0 ;
  assign n37599 = n1180 | n17489 ;
  assign n37600 = n3535 & ~n37599 ;
  assign n37598 = n24368 ^ n6128 ^ n5030 ;
  assign n37601 = n37600 ^ n37598 ^ 1'b0 ;
  assign n37602 = n6529 ^ n4338 ^ 1'b0 ;
  assign n37603 = ~n3563 & n37602 ;
  assign n37604 = ( n23022 & n30910 ) | ( n23022 & ~n37603 ) | ( n30910 & ~n37603 ) ;
  assign n37605 = ( n9363 & ~n37601 ) | ( n9363 & n37604 ) | ( ~n37601 & n37604 ) ;
  assign n37606 = n33202 ^ n16530 ^ n2867 ;
  assign n37607 = ~n8084 & n37606 ;
  assign n37608 = n37607 ^ n5951 ^ 1'b0 ;
  assign n37609 = n25887 & ~n37608 ;
  assign n37610 = n37609 ^ n13200 ^ n810 ;
  assign n37611 = n33967 ^ n1475 ^ 1'b0 ;
  assign n37612 = n6212 | n37611 ;
  assign n37613 = n26519 ^ n9534 ^ n6438 ;
  assign n37614 = n37613 ^ n12739 ^ 1'b0 ;
  assign n37615 = n11539 | n12912 ;
  assign n37616 = n37615 ^ n7291 ^ 1'b0 ;
  assign n37617 = n37616 ^ n24894 ^ 1'b0 ;
  assign n37618 = n37617 ^ n21682 ^ n6231 ;
  assign n37619 = n6117 & n37618 ;
  assign n37620 = n37619 ^ n32320 ^ 1'b0 ;
  assign n37625 = n12116 ^ n5579 ^ 1'b0 ;
  assign n37626 = n14052 & n37625 ;
  assign n37622 = ~n698 & n5427 ;
  assign n37623 = ~n11769 & n37622 ;
  assign n37621 = n6428 & n14988 ;
  assign n37624 = n37623 ^ n37621 ^ 1'b0 ;
  assign n37627 = n37626 ^ n37624 ^ n15238 ;
  assign n37628 = n15883 ^ n2374 ^ n2244 ;
  assign n37629 = ( n13915 & n18918 ) | ( n13915 & ~n36890 ) | ( n18918 & ~n36890 ) ;
  assign n37630 = n17342 ^ n6809 ^ 1'b0 ;
  assign n37631 = ~n17103 & n37630 ;
  assign n37632 = n30110 ^ n6373 ^ 1'b0 ;
  assign n37633 = n37631 & ~n37632 ;
  assign n37634 = n558 & n10270 ;
  assign n37635 = n37634 ^ n4947 ^ 1'b0 ;
  assign n37636 = ~n5199 & n37635 ;
  assign n37637 = n37636 ^ n3462 ^ 1'b0 ;
  assign n37638 = n4357 | n37637 ;
  assign n37639 = n34292 & ~n37638 ;
  assign n37640 = ~n22878 & n31254 ;
  assign n37641 = n37640 ^ n19837 ^ 1'b0 ;
  assign n37642 = n27118 ^ n17312 ^ n3332 ;
  assign n37643 = n15153 | n26999 ;
  assign n37644 = n13981 & n37643 ;
  assign n37647 = ( ~n7259 & n10633 ) | ( ~n7259 & n24377 ) | ( n10633 & n24377 ) ;
  assign n37648 = n20942 & ~n37647 ;
  assign n37645 = n12875 ^ n6219 ^ 1'b0 ;
  assign n37646 = n37645 ^ n22826 ^ n10540 ;
  assign n37649 = n37648 ^ n37646 ^ 1'b0 ;
  assign n37650 = ~n37644 & n37649 ;
  assign n37651 = n25079 ^ n15155 ^ 1'b0 ;
  assign n37652 = n30666 ^ n2662 ^ 1'b0 ;
  assign n37653 = ( n11434 & ~n37651 ) | ( n11434 & n37652 ) | ( ~n37651 & n37652 ) ;
  assign n37654 = n37156 ^ n22643 ^ 1'b0 ;
  assign n37655 = n25299 ^ n4350 ^ 1'b0 ;
  assign n37656 = n3041 | n37655 ;
  assign n37657 = ( n4566 & ~n37654 ) | ( n4566 & n37656 ) | ( ~n37654 & n37656 ) ;
  assign n37658 = n7067 & ~n35617 ;
  assign n37659 = n12910 & n37658 ;
  assign n37660 = n27851 ^ n17970 ^ 1'b0 ;
  assign n37661 = n18291 ^ n2502 ^ n1978 ;
  assign n37662 = n16348 & ~n23854 ;
  assign n37663 = n37662 ^ n37123 ^ 1'b0 ;
  assign n37664 = n10956 | n25927 ;
  assign n37665 = n23695 & ~n37664 ;
  assign n37666 = n22430 | n37665 ;
  assign n37667 = x117 | n37666 ;
  assign n37668 = ( n15496 & n19571 ) | ( n15496 & ~n37667 ) | ( n19571 & ~n37667 ) ;
  assign n37669 = ~n17203 & n33633 ;
  assign n37670 = n8976 & n37669 ;
  assign n37672 = n431 & ~n17585 ;
  assign n37673 = n37672 ^ n26679 ^ 1'b0 ;
  assign n37671 = n4243 | n13526 ;
  assign n37674 = n37673 ^ n37671 ^ 1'b0 ;
  assign n37675 = ( n16732 & ~n37670 ) | ( n16732 & n37674 ) | ( ~n37670 & n37674 ) ;
  assign n37676 = n27185 ^ n21159 ^ n13327 ;
  assign n37677 = n25033 ^ n15491 ^ 1'b0 ;
  assign n37678 = n37677 ^ n19476 ^ 1'b0 ;
  assign n37679 = n23777 | n37678 ;
  assign n37680 = n793 & ~n37679 ;
  assign n37681 = n37680 ^ n19059 ^ 1'b0 ;
  assign n37682 = n31705 ^ n26671 ^ 1'b0 ;
  assign n37683 = n37682 ^ n29426 ^ n7011 ;
  assign n37684 = n11876 ^ n10283 ^ 1'b0 ;
  assign n37685 = n37684 ^ n26329 ^ n17310 ;
  assign n37686 = n37685 ^ n17538 ^ n682 ;
  assign n37687 = n11621 ^ x171 ^ 1'b0 ;
  assign n37688 = n37687 ^ n32471 ^ n1158 ;
  assign n37689 = ~n22764 & n37688 ;
  assign n37690 = n1997 & ~n8889 ;
  assign n37691 = n3903 | n37690 ;
  assign n37692 = n37691 ^ n6857 ^ 1'b0 ;
  assign n37693 = n15163 | n35076 ;
  assign n37694 = n37693 ^ n34556 ^ 1'b0 ;
  assign n37695 = n1251 & n37694 ;
  assign n37696 = ~n1740 & n35974 ;
  assign n37697 = ~n12588 & n37696 ;
  assign n37698 = n26394 ^ n1187 ^ 1'b0 ;
  assign n37699 = n37697 | n37698 ;
  assign n37700 = n3117 & n6869 ;
  assign n37701 = ( ~n4083 & n28528 ) | ( ~n4083 & n37700 ) | ( n28528 & n37700 ) ;
  assign n37702 = n20945 | n37701 ;
  assign n37703 = n37702 ^ n36889 ^ 1'b0 ;
  assign n37704 = ~n22260 & n27496 ;
  assign n37705 = n37704 ^ n13841 ^ 1'b0 ;
  assign n37706 = ( n4695 & n12527 ) | ( n4695 & ~n34616 ) | ( n12527 & ~n34616 ) ;
  assign n37707 = n25225 ^ n2506 ^ 1'b0 ;
  assign n37708 = n37707 ^ n19456 ^ 1'b0 ;
  assign n37709 = n14998 & n37708 ;
  assign n37710 = ( n17122 & n23740 ) | ( n17122 & ~n24292 ) | ( n23740 & ~n24292 ) ;
  assign n37711 = n37710 ^ n35739 ^ 1'b0 ;
  assign n37712 = n37709 & ~n37711 ;
  assign n37713 = n16397 ^ n2135 ^ 1'b0 ;
  assign n37714 = n37713 ^ n30534 ^ 1'b0 ;
  assign n37715 = ~n11634 & n37714 ;
  assign n37716 = n8405 ^ n3427 ^ 1'b0 ;
  assign n37717 = ~n12254 & n37716 ;
  assign n37718 = n11193 & n24752 ;
  assign n37719 = ~n15788 & n22326 ;
  assign n37720 = n18285 ^ n16163 ^ 1'b0 ;
  assign n37721 = n11821 & n37720 ;
  assign n37722 = n37721 ^ n3168 ^ 1'b0 ;
  assign n37723 = n37722 ^ n20923 ^ n13642 ;
  assign n37724 = n2036 & ~n26042 ;
  assign n37725 = ~n33160 & n37724 ;
  assign n37726 = n14263 ^ n2860 ^ 1'b0 ;
  assign n37727 = ( n37723 & ~n37725 ) | ( n37723 & n37726 ) | ( ~n37725 & n37726 ) ;
  assign n37728 = ( n10372 & ~n19855 ) | ( n10372 & n37727 ) | ( ~n19855 & n37727 ) ;
  assign n37732 = n3767 & n32424 ;
  assign n37730 = n5219 ^ n2788 ^ n1046 ;
  assign n37731 = n17419 & ~n37730 ;
  assign n37733 = n37732 ^ n37731 ^ 1'b0 ;
  assign n37729 = n282 & ~n32460 ;
  assign n37734 = n37733 ^ n37729 ^ 1'b0 ;
  assign n37735 = n3748 | n12998 ;
  assign n37736 = ( n22063 & ~n37734 ) | ( n22063 & n37735 ) | ( ~n37734 & n37735 ) ;
  assign n37737 = n28441 ^ n12399 ^ 1'b0 ;
  assign n37738 = ( ~n2437 & n4455 ) | ( ~n2437 & n25359 ) | ( n4455 & n25359 ) ;
  assign n37739 = n24763 ^ n20821 ^ 1'b0 ;
  assign n37740 = ( n28511 & ~n37738 ) | ( n28511 & n37739 ) | ( ~n37738 & n37739 ) ;
  assign n37741 = n26986 ^ n634 ^ 1'b0 ;
  assign n37742 = ~n14436 & n37741 ;
  assign n37743 = n34291 | n37010 ;
  assign n37744 = n37743 ^ n4119 ^ 1'b0 ;
  assign n37745 = n37742 & ~n37744 ;
  assign n37746 = n31686 ^ n8405 ^ 1'b0 ;
  assign n37747 = n5012 | n37746 ;
  assign n37748 = n16504 ^ n2364 ^ 1'b0 ;
  assign n37749 = n30897 ^ n30468 ^ n25045 ;
  assign n37750 = n37749 ^ n5520 ^ 1'b0 ;
  assign n37751 = n30176 ^ n13279 ^ n4826 ;
  assign n37752 = n15767 ^ n4244 ^ 1'b0 ;
  assign n37753 = ~n19186 & n37752 ;
  assign n37754 = ~n6023 & n37753 ;
  assign n37755 = n5589 & n37754 ;
  assign n37756 = n18110 ^ n4259 ^ 1'b0 ;
  assign n37757 = ~n27875 & n37756 ;
  assign n37758 = n30834 ^ n15452 ^ n10943 ;
  assign n37759 = ~n11723 & n37758 ;
  assign n37760 = n37759 ^ n33492 ^ 1'b0 ;
  assign n37761 = ( n3942 & n16115 ) | ( n3942 & ~n37760 ) | ( n16115 & ~n37760 ) ;
  assign n37764 = ~n5246 & n6061 ;
  assign n37762 = n2267 ^ n1643 ^ 1'b0 ;
  assign n37763 = ~n8850 & n37762 ;
  assign n37765 = n37764 ^ n37763 ^ 1'b0 ;
  assign n37766 = n37765 ^ n18079 ^ n10979 ;
  assign n37767 = n13042 ^ n10653 ^ 1'b0 ;
  assign n37768 = n19835 & n37767 ;
  assign n37769 = n9724 & n37768 ;
  assign n37770 = n37769 ^ n9521 ^ 1'b0 ;
  assign n37771 = n26335 ^ n434 ^ 1'b0 ;
  assign n37772 = n9938 ^ n8502 ^ n7453 ;
  assign n37773 = n37772 ^ n11078 ^ 1'b0 ;
  assign n37774 = n13441 | n37773 ;
  assign n37775 = n7935 & n34620 ;
  assign n37777 = ~n5657 & n5929 ;
  assign n37778 = n37777 ^ n5052 ^ 1'b0 ;
  assign n37776 = n8786 | n30222 ;
  assign n37779 = n37778 ^ n37776 ^ 1'b0 ;
  assign n37780 = n37779 ^ n33130 ^ 1'b0 ;
  assign n37781 = ~n8802 & n37780 ;
  assign n37782 = ~n25224 & n37781 ;
  assign n37783 = ~n9933 & n37782 ;
  assign n37784 = n31929 ^ n2045 ^ 1'b0 ;
  assign n37785 = n2528 & n19993 ;
  assign n37786 = n23313 & ~n37785 ;
  assign n37787 = n33670 ^ n10461 ^ n10230 ;
  assign n37788 = ~n33093 & n33586 ;
  assign n37789 = ~n29884 & n37788 ;
  assign n37790 = n30549 & n37789 ;
  assign n37791 = ( n37786 & n37787 ) | ( n37786 & n37790 ) | ( n37787 & n37790 ) ;
  assign n37792 = n27631 ^ n13242 ^ 1'b0 ;
  assign n37793 = n37792 ^ n21900 ^ n21145 ;
  assign n37794 = n13999 ^ n3771 ^ 1'b0 ;
  assign n37795 = n11945 ^ n8056 ^ n7177 ;
  assign n37796 = n37795 ^ n11171 ^ 1'b0 ;
  assign n37797 = ~n18608 & n37796 ;
  assign n37798 = ~n1385 & n37797 ;
  assign n37799 = ( n2411 & n35740 ) | ( n2411 & ~n37649 ) | ( n35740 & ~n37649 ) ;
  assign n37800 = n27068 ^ n11348 ^ 1'b0 ;
  assign n37801 = n26648 ^ n9610 ^ 1'b0 ;
  assign n37802 = n7833 & ~n37801 ;
  assign n37803 = ~n34465 & n37802 ;
  assign n37804 = n10753 & n17556 ;
  assign n37805 = n37804 ^ n7696 ^ 1'b0 ;
  assign n37806 = n21288 ^ n8369 ^ 1'b0 ;
  assign n37807 = n7334 & n37806 ;
  assign n37812 = ~n7496 & n29472 ;
  assign n37813 = n3846 & n37812 ;
  assign n37814 = n37813 ^ n9076 ^ 1'b0 ;
  assign n37815 = n7748 | n8452 ;
  assign n37816 = n8041 & ~n37815 ;
  assign n37817 = ( n9910 & n37814 ) | ( n9910 & ~n37816 ) | ( n37814 & ~n37816 ) ;
  assign n37808 = n11689 & ~n13341 ;
  assign n37809 = n37808 ^ n12326 ^ 1'b0 ;
  assign n37810 = n37809 ^ n3701 ^ n1743 ;
  assign n37811 = ~n26592 & n37810 ;
  assign n37818 = n37817 ^ n37811 ^ 1'b0 ;
  assign n37819 = n23598 ^ n471 ^ 1'b0 ;
  assign n37820 = n13788 & n37819 ;
  assign n37821 = n37820 ^ n3889 ^ 1'b0 ;
  assign n37822 = n10898 & ~n11666 ;
  assign n37823 = ( n17875 & ~n20286 ) | ( n17875 & n23969 ) | ( ~n20286 & n23969 ) ;
  assign n37824 = ( ~n9941 & n11300 ) | ( ~n9941 & n24192 ) | ( n11300 & n24192 ) ;
  assign n37825 = n37824 ^ n20431 ^ n9727 ;
  assign n37826 = n345 & ~n12996 ;
  assign n37827 = n37826 ^ n35222 ^ 1'b0 ;
  assign n37828 = ~n22455 & n37827 ;
  assign n37829 = ( n15238 & ~n23265 ) | ( n15238 & n37828 ) | ( ~n23265 & n37828 ) ;
  assign n37832 = n19233 ^ n910 ^ 1'b0 ;
  assign n37833 = n11136 & n37832 ;
  assign n37834 = n5171 & n37833 ;
  assign n37830 = n16188 ^ n3177 ^ 1'b0 ;
  assign n37831 = n5126 & ~n37830 ;
  assign n37835 = n37834 ^ n37831 ^ n16392 ;
  assign n37836 = n8469 | n37464 ;
  assign n37837 = n25767 & ~n37836 ;
  assign n37838 = n36260 & n37837 ;
  assign n37839 = n33120 ^ n6814 ^ 1'b0 ;
  assign n37840 = n31823 ^ n5523 ^ n1870 ;
  assign n37841 = n37840 ^ n7869 ^ 1'b0 ;
  assign n37842 = ~n8978 & n37841 ;
  assign n37843 = n4695 ^ n4423 ^ n2611 ;
  assign n37844 = n29577 & ~n37843 ;
  assign n37845 = n2944 & ~n14109 ;
  assign n37846 = n19257 & n37845 ;
  assign n37847 = n37846 ^ n26938 ^ 1'b0 ;
  assign n37848 = n6328 | n35862 ;
  assign n37849 = n37848 ^ n13262 ^ 1'b0 ;
  assign n37850 = n7678 | n12755 ;
  assign n37851 = ( n2836 & n37849 ) | ( n2836 & n37850 ) | ( n37849 & n37850 ) ;
  assign n37852 = ~n11930 & n14359 ;
  assign n37853 = n37852 ^ n5972 ^ 1'b0 ;
  assign n37854 = n19174 ^ n1444 ^ 1'b0 ;
  assign n37855 = n37853 & n37854 ;
  assign n37856 = n8733 & n37855 ;
  assign n37857 = n15982 & n37856 ;
  assign n37858 = ( x42 & x207 ) | ( x42 & ~n20912 ) | ( x207 & ~n20912 ) ;
  assign n37859 = ( n24399 & n37857 ) | ( n24399 & ~n37858 ) | ( n37857 & ~n37858 ) ;
  assign n37860 = n19120 ^ n14396 ^ n4568 ;
  assign n37861 = ( n4107 & n8206 ) | ( n4107 & ~n37860 ) | ( n8206 & ~n37860 ) ;
  assign n37862 = n7016 | n37861 ;
  assign n37863 = n37862 ^ n8577 ^ 1'b0 ;
  assign n37864 = n7108 & n24674 ;
  assign n37865 = n3264 & ~n14053 ;
  assign n37866 = n10731 | n37865 ;
  assign n37867 = n11287 & ~n37866 ;
  assign n37868 = ~n26688 & n29349 ;
  assign n37869 = ( n2850 & n10577 ) | ( n2850 & n35475 ) | ( n10577 & n35475 ) ;
  assign n37870 = ( n6414 & n9485 ) | ( n6414 & ~n14587 ) | ( n9485 & ~n14587 ) ;
  assign n37871 = n9526 & ~n37870 ;
  assign n37872 = n37871 ^ n9093 ^ n4982 ;
  assign n37873 = n18101 | n18858 ;
  assign n37874 = n25278 & ~n37873 ;
  assign n37875 = n3453 | n37874 ;
  assign n37876 = n18148 & ~n37875 ;
  assign n37877 = n30321 | n37876 ;
  assign n37878 = n37877 ^ n16383 ^ 1'b0 ;
  assign n37879 = n21646 & n26875 ;
  assign n37880 = n13107 ^ n10482 ^ n6184 ;
  assign n37881 = ( n29312 & n35298 ) | ( n29312 & ~n37880 ) | ( n35298 & ~n37880 ) ;
  assign n37882 = n37881 ^ n32714 ^ n17485 ;
  assign n37883 = ~n36289 & n37882 ;
  assign n37884 = ( n2160 & n11030 ) | ( n2160 & ~n17154 ) | ( n11030 & ~n17154 ) ;
  assign n37885 = n37884 ^ n17083 ^ n934 ;
  assign n37886 = ( n7937 & ~n13969 ) | ( n7937 & n28244 ) | ( ~n13969 & n28244 ) ;
  assign n37887 = ( n3766 & n10267 ) | ( n3766 & ~n13679 ) | ( n10267 & ~n13679 ) ;
  assign n37889 = n35948 ^ n4790 ^ 1'b0 ;
  assign n37888 = n9697 | n13009 ;
  assign n37890 = n37889 ^ n37888 ^ 1'b0 ;
  assign n37891 = ~n3535 & n4001 ;
  assign n37892 = ~n17237 & n37891 ;
  assign n37893 = n9603 ^ n8390 ^ 1'b0 ;
  assign n37894 = ~n4345 & n37893 ;
  assign n37895 = ~n3001 & n37894 ;
  assign n37896 = n37895 ^ n30722 ^ 1'b0 ;
  assign n37897 = ~n268 & n36740 ;
  assign n37898 = n13216 ^ n10743 ^ 1'b0 ;
  assign n37899 = ( ~x220 & n499 ) | ( ~x220 & n37898 ) | ( n499 & n37898 ) ;
  assign n37900 = n37899 ^ n536 ^ 1'b0 ;
  assign n37901 = n37732 ^ n15223 ^ n8276 ;
  assign n37902 = ( n24120 & n36591 ) | ( n24120 & n37901 ) | ( n36591 & n37901 ) ;
  assign n37903 = x48 & n33866 ;
  assign n37904 = n37903 ^ n29304 ^ 1'b0 ;
  assign n37905 = ( n16025 & n37263 ) | ( n16025 & n37904 ) | ( n37263 & n37904 ) ;
  assign n37906 = ( n2406 & ~n10865 ) | ( n2406 & n25355 ) | ( ~n10865 & n25355 ) ;
  assign n37907 = n32867 ^ x61 ^ 1'b0 ;
  assign n37908 = ~n29867 & n30416 ;
  assign n37909 = ~n28663 & n37908 ;
  assign n37910 = n14973 | n26742 ;
  assign n37911 = n36964 | n37910 ;
  assign n37912 = n294 & n16537 ;
  assign n37913 = n30620 & n37912 ;
  assign n37914 = n37913 ^ n15477 ^ 1'b0 ;
  assign n37915 = n4589 ^ n3003 ^ 1'b0 ;
  assign n37916 = ( n36204 & n36949 ) | ( n36204 & n37915 ) | ( n36949 & n37915 ) ;
  assign n37917 = ~n6245 & n22071 ;
  assign n37918 = n30657 & ~n37917 ;
  assign n37919 = n37918 ^ n25095 ^ n2584 ;
  assign n37921 = n20353 ^ n15994 ^ n3906 ;
  assign n37920 = n6787 | n23305 ;
  assign n37922 = n37921 ^ n37920 ^ 1'b0 ;
  assign n37923 = n14164 ^ n9961 ^ 1'b0 ;
  assign n37924 = n12782 ^ n5991 ^ n5794 ;
  assign n37925 = n37923 | n37924 ;
  assign n37926 = n37925 ^ n28712 ^ 1'b0 ;
  assign n37927 = n22674 ^ n9701 ^ 1'b0 ;
  assign n37928 = n25003 & ~n37927 ;
  assign n37929 = n22914 & ~n27015 ;
  assign n37930 = n37477 ^ n12640 ^ 1'b0 ;
  assign n37931 = n37929 & ~n37930 ;
  assign n37932 = n10617 ^ n9814 ^ 1'b0 ;
  assign n37933 = n37932 ^ x182 ^ x133 ;
  assign n37934 = ~n17929 & n27163 ;
  assign n37935 = ~n1218 & n26483 ;
  assign n37936 = ( n748 & n5373 ) | ( n748 & n37935 ) | ( n5373 & n37935 ) ;
  assign n37937 = ( n5295 & ~n8495 ) | ( n5295 & n23251 ) | ( ~n8495 & n23251 ) ;
  assign n37938 = n37937 ^ n20096 ^ n4294 ;
  assign n37939 = n37938 ^ n12390 ^ 1'b0 ;
  assign n37940 = ~n13251 & n20592 ;
  assign n37941 = n37940 ^ n13689 ^ 1'b0 ;
  assign n37942 = n23406 ^ n10654 ^ 1'b0 ;
  assign n37943 = ~n6808 & n37942 ;
  assign n37944 = ( n4129 & n25340 ) | ( n4129 & n37943 ) | ( n25340 & n37943 ) ;
  assign n37945 = n37944 ^ n34816 ^ n7533 ;
  assign n37946 = n21129 ^ n10121 ^ 1'b0 ;
  assign n37947 = n37945 & n37946 ;
  assign n37948 = n4438 ^ n2994 ^ n2841 ;
  assign n37949 = ( ~n11261 & n17310 ) | ( ~n11261 & n21445 ) | ( n17310 & n21445 ) ;
  assign n37950 = n34642 ^ n14338 ^ x152 ;
  assign n37951 = n5877 ^ n1156 ^ 1'b0 ;
  assign n37952 = n18523 & ~n37951 ;
  assign n37953 = ~n27425 & n37952 ;
  assign n37959 = n33327 ^ n26653 ^ 1'b0 ;
  assign n37955 = n6796 ^ n4826 ^ 1'b0 ;
  assign n37954 = n18500 ^ n2565 ^ 1'b0 ;
  assign n37956 = n37955 ^ n37954 ^ n14520 ;
  assign n37957 = n26921 ^ n15137 ^ 1'b0 ;
  assign n37958 = n37956 | n37957 ;
  assign n37960 = n37959 ^ n37958 ^ 1'b0 ;
  assign n37966 = n25724 ^ n23238 ^ n455 ;
  assign n37964 = n1395 & ~n10665 ;
  assign n37965 = n19573 & n37964 ;
  assign n37962 = n28756 ^ n13964 ^ n2818 ;
  assign n37961 = n33015 ^ n22958 ^ n18623 ;
  assign n37963 = n37962 ^ n37961 ^ n37944 ;
  assign n37967 = n37966 ^ n37965 ^ n37963 ;
  assign n37968 = n7168 | n16064 ;
  assign n37969 = n37968 ^ n13001 ^ 1'b0 ;
  assign n37970 = ( n4597 & n24900 ) | ( n4597 & ~n30856 ) | ( n24900 & ~n30856 ) ;
  assign n37971 = ( n5390 & n37969 ) | ( n5390 & ~n37970 ) | ( n37969 & ~n37970 ) ;
  assign n37972 = n6629 & ~n36169 ;
  assign n37973 = ~n23185 & n37972 ;
  assign n37974 = ~n340 & n7191 ;
  assign n37975 = n37974 ^ n6641 ^ 1'b0 ;
  assign n37976 = n10730 & n32235 ;
  assign n37977 = ~n33695 & n37515 ;
  assign n37978 = ( n15820 & n18774 ) | ( n15820 & n32853 ) | ( n18774 & n32853 ) ;
  assign n37979 = n7688 | n10356 ;
  assign n37980 = n37979 ^ n5458 ^ 1'b0 ;
  assign n37981 = n37980 ^ n34350 ^ n16399 ;
  assign n37982 = n37981 ^ n21973 ^ 1'b0 ;
  assign n37983 = n12739 & n37982 ;
  assign n37984 = n871 | n7600 ;
  assign n37985 = n14859 ^ n11796 ^ 1'b0 ;
  assign n37986 = n15608 ^ n12978 ^ 1'b0 ;
  assign n37987 = n2816 & ~n37986 ;
  assign n37988 = ~n9014 & n37987 ;
  assign n37989 = ~n4850 & n37988 ;
  assign n37990 = n33743 ^ n14861 ^ 1'b0 ;
  assign n37991 = ( ~n4912 & n10733 ) | ( ~n4912 & n20452 ) | ( n10733 & n20452 ) ;
  assign n37992 = n37990 | n37991 ;
  assign n37993 = n17595 & n24985 ;
  assign n37994 = n12861 & n37993 ;
  assign n37995 = n23045 & n27971 ;
  assign n37996 = n10371 & n37995 ;
  assign n37997 = n4725 | n16914 ;
  assign n37998 = n37997 ^ n33331 ^ 1'b0 ;
  assign n37999 = n33040 ^ n6205 ^ 1'b0 ;
  assign n38000 = n37998 & n37999 ;
  assign n38001 = n9156 | n23463 ;
  assign n38002 = n38001 ^ n35777 ^ n20912 ;
  assign n38003 = n29871 ^ n3687 ^ 1'b0 ;
  assign n38004 = n14635 & n38003 ;
  assign n38005 = n4916 | n9094 ;
  assign n38006 = n16710 ^ n5050 ^ n3372 ;
  assign n38007 = n6928 | n10249 ;
  assign n38008 = n16548 & ~n38007 ;
  assign n38009 = n6752 | n38008 ;
  assign n38010 = n38009 ^ n8838 ^ 1'b0 ;
  assign n38011 = n38010 ^ n26772 ^ n15389 ;
  assign n38012 = ( n38005 & n38006 ) | ( n38005 & n38011 ) | ( n38006 & n38011 ) ;
  assign n38013 = n24085 ^ n21083 ^ n15271 ;
  assign n38014 = ~n36135 & n38013 ;
  assign n38015 = n16063 ^ n8856 ^ 1'b0 ;
  assign n38016 = n37603 & n38015 ;
  assign n38017 = n19218 & ~n38016 ;
  assign n38020 = n23141 ^ n15091 ^ 1'b0 ;
  assign n38021 = n26762 ^ n12755 ^ n9089 ;
  assign n38022 = ~n38020 & n38021 ;
  assign n38018 = n34041 ^ n14892 ^ 1'b0 ;
  assign n38019 = n38018 ^ n20118 ^ 1'b0 ;
  assign n38023 = n38022 ^ n38019 ^ 1'b0 ;
  assign n38024 = n13590 & n38023 ;
  assign n38025 = n31804 ^ n4912 ^ n4037 ;
  assign n38026 = n12032 | n13068 ;
  assign n38027 = ~n19642 & n23052 ;
  assign n38028 = n6394 & n38027 ;
  assign n38029 = n34817 | n38028 ;
  assign n38030 = n10595 & ~n38029 ;
  assign n38031 = n4473 & ~n20440 ;
  assign n38032 = n6030 ^ n990 ^ 1'b0 ;
  assign n38033 = ( n9262 & n16499 ) | ( n9262 & ~n38032 ) | ( n16499 & ~n38032 ) ;
  assign n38034 = ( n5326 & ~n23932 ) | ( n5326 & n29443 ) | ( ~n23932 & n29443 ) ;
  assign n38035 = n19473 ^ n11837 ^ 1'b0 ;
  assign n38036 = ~n10218 & n38035 ;
  assign n38037 = n38036 ^ n11319 ^ x51 ;
  assign n38038 = ( n2449 & n9705 ) | ( n2449 & ~n12591 ) | ( n9705 & ~n12591 ) ;
  assign n38039 = n38038 ^ n3409 ^ 1'b0 ;
  assign n38040 = n38039 ^ n9499 ^ 1'b0 ;
  assign n38041 = n893 & ~n38040 ;
  assign n38042 = ( n3717 & n7621 ) | ( n3717 & ~n38041 ) | ( n7621 & ~n38041 ) ;
  assign n38043 = ~n24471 & n29237 ;
  assign n38044 = n38043 ^ n18647 ^ n17827 ;
  assign n38045 = n18419 | n38044 ;
  assign n38046 = ( ~n3331 & n8390 ) | ( ~n3331 & n13167 ) | ( n8390 & n13167 ) ;
  assign n38047 = ( ~n9675 & n27895 ) | ( ~n9675 & n38046 ) | ( n27895 & n38046 ) ;
  assign n38048 = n38047 ^ n22353 ^ 1'b0 ;
  assign n38049 = n21071 ^ n1264 ^ 1'b0 ;
  assign n38050 = n23711 & ~n38049 ;
  assign n38051 = ( n1567 & ~n13692 ) | ( n1567 & n16917 ) | ( ~n13692 & n16917 ) ;
  assign n38053 = n12591 ^ n10100 ^ 1'b0 ;
  assign n38054 = ( n15598 & n37082 ) | ( n15598 & n38053 ) | ( n37082 & n38053 ) ;
  assign n38052 = n26266 ^ n24684 ^ n16375 ;
  assign n38055 = n38054 ^ n38052 ^ n10596 ;
  assign n38056 = n8630 | n38055 ;
  assign n38057 = n38056 ^ n18797 ^ 1'b0 ;
  assign n38058 = ( n15422 & n15605 ) | ( n15422 & ~n16316 ) | ( n15605 & ~n16316 ) ;
  assign n38059 = ( ~n9775 & n23474 ) | ( ~n9775 & n38058 ) | ( n23474 & n38058 ) ;
  assign n38060 = n25543 ^ n18156 ^ n16499 ;
  assign n38061 = n1776 | n38060 ;
  assign n38062 = n38061 ^ n21766 ^ 1'b0 ;
  assign n38063 = n16222 & ~n18535 ;
  assign n38064 = n4461 ^ n855 ^ 1'b0 ;
  assign n38065 = n8935 | n38064 ;
  assign n38066 = n20626 & ~n38065 ;
  assign n38067 = n38063 & n38066 ;
  assign n38068 = n16716 ^ n8448 ^ 1'b0 ;
  assign n38069 = n38067 | n38068 ;
  assign n38070 = n28658 ^ n8818 ^ 1'b0 ;
  assign n38071 = n5983 & n38070 ;
  assign n38072 = n22148 | n22918 ;
  assign n38073 = n21787 ^ n17628 ^ n12980 ;
  assign n38074 = n30133 ^ n3231 ^ 1'b0 ;
  assign n38075 = n6040 & n38074 ;
  assign n38076 = n38075 ^ n29273 ^ n2602 ;
  assign n38077 = ( n5064 & ~n35180 ) | ( n5064 & n38076 ) | ( ~n35180 & n38076 ) ;
  assign n38078 = n27523 ^ n26376 ^ 1'b0 ;
  assign n38079 = n11947 ^ n11482 ^ n9286 ;
  assign n38080 = n38079 ^ n23937 ^ 1'b0 ;
  assign n38081 = n31026 ^ n21371 ^ n10786 ;
  assign n38082 = n38081 ^ n32261 ^ 1'b0 ;
  assign n38083 = ~n10405 & n18191 ;
  assign n38084 = n32453 ^ n30564 ^ 1'b0 ;
  assign n38085 = ( n14826 & ~n38083 ) | ( n14826 & n38084 ) | ( ~n38083 & n38084 ) ;
  assign n38086 = ( ~n8793 & n14672 ) | ( ~n8793 & n20798 ) | ( n14672 & n20798 ) ;
  assign n38087 = n38086 ^ n34544 ^ n9136 ;
  assign n38089 = ~n8263 & n22220 ;
  assign n38088 = n27724 & n30406 ;
  assign n38090 = n38089 ^ n38088 ^ 1'b0 ;
  assign n38091 = n20887 ^ n2908 ^ n1790 ;
  assign n38092 = n5526 ^ n3457 ^ 1'b0 ;
  assign n38093 = n38091 & ~n38092 ;
  assign n38094 = ( ~n2549 & n11074 ) | ( ~n2549 & n19790 ) | ( n11074 & n19790 ) ;
  assign n38095 = ~n11287 & n38094 ;
  assign n38096 = n35342 ^ n27800 ^ n2299 ;
  assign n38097 = n16993 ^ n4284 ^ 1'b0 ;
  assign n38098 = ~n16044 & n38097 ;
  assign n38099 = n38098 ^ n11019 ^ 1'b0 ;
  assign n38100 = ~n33067 & n38099 ;
  assign n38101 = ( n16557 & n19511 ) | ( n16557 & n29605 ) | ( n19511 & n29605 ) ;
  assign n38102 = n11139 & ~n12425 ;
  assign n38103 = n38102 ^ n8513 ^ 1'b0 ;
  assign n38104 = n38103 ^ n4806 ^ 1'b0 ;
  assign n38105 = n21923 | n38104 ;
  assign n38106 = n11242 | n38105 ;
  assign n38107 = n38101 & ~n38106 ;
  assign n38108 = n7386 | n38107 ;
  assign n38109 = n8220 | n27379 ;
  assign n38110 = ( n6048 & n15256 ) | ( n6048 & ~n23219 ) | ( n15256 & ~n23219 ) ;
  assign n38111 = n14666 ^ n1934 ^ 1'b0 ;
  assign n38112 = n38110 & n38111 ;
  assign n38113 = n38112 ^ n13966 ^ 1'b0 ;
  assign n38114 = n19849 ^ n8290 ^ n4695 ;
  assign n38115 = n33726 ^ n16196 ^ n6326 ;
  assign n38116 = n17226 | n20459 ;
  assign n38117 = n38116 ^ n33572 ^ 1'b0 ;
  assign n38118 = ( n23644 & ~n25767 ) | ( n23644 & n33701 ) | ( ~n25767 & n33701 ) ;
  assign n38119 = n38118 ^ n14920 ^ 1'b0 ;
  assign n38120 = n29077 & ~n38119 ;
  assign n38121 = n28968 ^ n24846 ^ n14021 ;
  assign n38122 = ( n6753 & n10983 ) | ( n6753 & ~n11008 ) | ( n10983 & ~n11008 ) ;
  assign n38123 = ~n15837 & n31042 ;
  assign n38124 = n38123 ^ n10601 ^ 1'b0 ;
  assign n38125 = n38124 ^ n22306 ^ n10767 ;
  assign n38127 = ( n6138 & n20032 ) | ( n6138 & n33474 ) | ( n20032 & n33474 ) ;
  assign n38126 = n916 | n28308 ;
  assign n38128 = n38127 ^ n38126 ^ 1'b0 ;
  assign n38129 = n37441 ^ n24706 ^ n16953 ;
  assign n38130 = n38128 & ~n38129 ;
  assign n38131 = n38130 ^ n26056 ^ 1'b0 ;
  assign n38132 = n19724 ^ n8286 ^ 1'b0 ;
  assign n38133 = n38132 ^ n36972 ^ n4619 ;
  assign n38134 = ( n8675 & n13554 ) | ( n8675 & ~n28863 ) | ( n13554 & ~n28863 ) ;
  assign n38135 = n38134 ^ n18517 ^ n14880 ;
  assign n38136 = n29076 ^ n5917 ^ 1'b0 ;
  assign n38137 = ( n27654 & ~n38135 ) | ( n27654 & n38136 ) | ( ~n38135 & n38136 ) ;
  assign n38138 = n1634 | n31054 ;
  assign n38139 = n38138 ^ n37272 ^ 1'b0 ;
  assign n38140 = n15795 ^ n9583 ^ n4338 ;
  assign n38141 = n38140 ^ n957 ^ 1'b0 ;
  assign n38145 = n3841 | n29561 ;
  assign n38142 = n34018 ^ n3004 ^ 1'b0 ;
  assign n38143 = n5840 & ~n38142 ;
  assign n38144 = n38143 ^ n38013 ^ 1'b0 ;
  assign n38146 = n38145 ^ n38144 ^ n11767 ;
  assign n38148 = n15985 ^ n14467 ^ n11489 ;
  assign n38147 = n14710 & n16600 ;
  assign n38149 = n38148 ^ n38147 ^ 1'b0 ;
  assign n38150 = n12077 | n38149 ;
  assign n38151 = n22980 & ~n29468 ;
  assign n38152 = n38151 ^ n11750 ^ 1'b0 ;
  assign n38153 = n29026 ^ n9841 ^ n2536 ;
  assign n38154 = n18929 ^ n10418 ^ 1'b0 ;
  assign n38155 = n367 & ~n38154 ;
  assign n38156 = n15641 & ~n38155 ;
  assign n38161 = n3979 & n5866 ;
  assign n38162 = ~n3979 & n38161 ;
  assign n38163 = n6909 | n38162 ;
  assign n38159 = n23880 ^ n14265 ^ 1'b0 ;
  assign n38160 = n4517 & ~n38159 ;
  assign n38157 = n9488 & n18918 ;
  assign n38158 = ~n18918 & n38157 ;
  assign n38164 = n38163 ^ n38160 ^ n38158 ;
  assign n38165 = ( n11629 & n19933 ) | ( n11629 & ~n34747 ) | ( n19933 & ~n34747 ) ;
  assign n38166 = n19571 | n38165 ;
  assign n38167 = n6558 & ~n38166 ;
  assign n38168 = n38167 ^ n18924 ^ 1'b0 ;
  assign n38169 = n9403 ^ n759 ^ 1'b0 ;
  assign n38170 = n10225 | n38169 ;
  assign n38171 = n32160 ^ n32104 ^ 1'b0 ;
  assign n38172 = n8999 | n38171 ;
  assign n38173 = n12088 ^ n8945 ^ 1'b0 ;
  assign n38174 = ~n1915 & n12272 ;
  assign n38175 = ( n5712 & ~n18623 ) | ( n5712 & n24361 ) | ( ~n18623 & n24361 ) ;
  assign n38176 = n34892 ^ n34392 ^ 1'b0 ;
  assign n38177 = n26855 & ~n36268 ;
  assign n38178 = n26816 ^ n15943 ^ 1'b0 ;
  assign n38179 = n12157 & ~n25293 ;
  assign n38180 = n692 & n38179 ;
  assign n38181 = n8234 | n38180 ;
  assign n38182 = n26850 & ~n38181 ;
  assign n38183 = n38182 ^ n2805 ^ 1'b0 ;
  assign n38184 = ~n30497 & n38183 ;
  assign n38185 = n23962 ^ n23402 ^ 1'b0 ;
  assign n38186 = n38184 & ~n38185 ;
  assign n38187 = n3997 & ~n17718 ;
  assign n38188 = n38187 ^ n18800 ^ n7211 ;
  assign n38189 = ( n1124 & ~n20042 ) | ( n1124 & n38188 ) | ( ~n20042 & n38188 ) ;
  assign n38190 = n33423 ^ n21435 ^ 1'b0 ;
  assign n38194 = n18956 ^ n2786 ^ 1'b0 ;
  assign n38191 = ( n3682 & ~n11503 ) | ( n3682 & n12724 ) | ( ~n11503 & n12724 ) ;
  assign n38192 = n38191 ^ n12285 ^ 1'b0 ;
  assign n38193 = x205 & ~n38192 ;
  assign n38195 = n38194 ^ n38193 ^ n30053 ;
  assign n38196 = n24725 ^ n16214 ^ 1'b0 ;
  assign n38197 = n38196 ^ n35938 ^ n8256 ;
  assign n38198 = n26160 ^ n23242 ^ n12902 ;
  assign n38199 = n18049 & n38198 ;
  assign n38200 = ( n7310 & ~n7751 ) | ( n7310 & n8808 ) | ( ~n7751 & n8808 ) ;
  assign n38201 = ( n14509 & n18976 ) | ( n14509 & ~n38200 ) | ( n18976 & ~n38200 ) ;
  assign n38202 = ~n3599 & n18901 ;
  assign n38203 = n38202 ^ n36835 ^ 1'b0 ;
  assign n38204 = n7116 & n8531 ;
  assign n38205 = x63 & n3214 ;
  assign n38206 = n38205 ^ n23643 ^ 1'b0 ;
  assign n38207 = n38206 ^ n13758 ^ 1'b0 ;
  assign n38208 = n23536 & n38207 ;
  assign n38209 = ~n11337 & n11669 ;
  assign n38210 = ~n5128 & n38209 ;
  assign n38211 = n381 | n38210 ;
  assign n38212 = n9984 & n16502 ;
  assign n38213 = n38212 ^ n7238 ^ 1'b0 ;
  assign n38214 = n17419 & n38213 ;
  assign n38215 = ~n7986 & n38214 ;
  assign n38216 = n27210 | n38215 ;
  assign n38217 = n6096 & n20666 ;
  assign n38218 = ( n20640 & ~n38216 ) | ( n20640 & n38217 ) | ( ~n38216 & n38217 ) ;
  assign n38222 = n35501 ^ n3502 ^ 1'b0 ;
  assign n38223 = ~n18291 & n38222 ;
  assign n38224 = n38223 ^ n8726 ^ 1'b0 ;
  assign n38219 = ( n1941 & n10133 ) | ( n1941 & n29025 ) | ( n10133 & n29025 ) ;
  assign n38220 = n22111 ^ n16157 ^ n10129 ;
  assign n38221 = ( n17920 & ~n38219 ) | ( n17920 & n38220 ) | ( ~n38219 & n38220 ) ;
  assign n38225 = n38224 ^ n38221 ^ n10314 ;
  assign n38226 = n28318 ^ n25112 ^ n22257 ;
  assign n38227 = n2935 | n18000 ;
  assign n38228 = n2781 & ~n38227 ;
  assign n38229 = n12815 ^ n8573 ^ 1'b0 ;
  assign n38230 = n30819 ^ n25908 ^ 1'b0 ;
  assign n38231 = n38230 ^ n10248 ^ n9234 ;
  assign n38232 = ~n36990 & n38231 ;
  assign n38233 = ( ~n3154 & n10297 ) | ( ~n3154 & n11775 ) | ( n10297 & n11775 ) ;
  assign n38234 = n38233 ^ n26003 ^ n23648 ;
  assign n38235 = n3229 & n7733 ;
  assign n38236 = n38235 ^ n4707 ^ 1'b0 ;
  assign n38237 = n38236 ^ n21236 ^ n19526 ;
  assign n38238 = n5574 | n35922 ;
  assign n38239 = n8929 ^ n6132 ^ n2148 ;
  assign n38240 = n38239 ^ n15800 ^ 1'b0 ;
  assign n38241 = n17172 ^ n8613 ^ 1'b0 ;
  assign n38242 = n38241 ^ n31400 ^ n1068 ;
  assign n38243 = n6782 & n19605 ;
  assign n38244 = n2145 & n32234 ;
  assign n38245 = n16332 ^ n3032 ^ 1'b0 ;
  assign n38246 = n12516 & ~n38245 ;
  assign n38247 = ~n20060 & n35645 ;
  assign n38248 = ~n38246 & n38247 ;
  assign n38254 = n24910 ^ n20893 ^ n2854 ;
  assign n38249 = n12649 | n26581 ;
  assign n38250 = n38249 ^ n9853 ^ 1'b0 ;
  assign n38251 = ~n9700 & n38250 ;
  assign n38252 = ~n15682 & n38251 ;
  assign n38253 = n13383 & n38252 ;
  assign n38255 = n38254 ^ n38253 ^ n29969 ;
  assign n38256 = n38255 ^ n24500 ^ n9725 ;
  assign n38257 = n10223 ^ n6175 ^ 1'b0 ;
  assign n38258 = n5086 ^ n3341 ^ 1'b0 ;
  assign n38259 = n14377 & ~n38258 ;
  assign n38260 = n38257 & n38259 ;
  assign n38261 = ( n4965 & n17489 ) | ( n4965 & ~n38260 ) | ( n17489 & ~n38260 ) ;
  assign n38262 = n6565 & n38261 ;
  assign n38263 = n4945 & n38262 ;
  assign n38264 = n7050 & ~n38263 ;
  assign n38267 = ~n12847 & n35705 ;
  assign n38268 = n15666 & ~n38267 ;
  assign n38269 = n38268 ^ n8698 ^ 1'b0 ;
  assign n38270 = n38269 ^ n1681 ^ 1'b0 ;
  assign n38265 = ~n21421 & n24026 ;
  assign n38266 = ~n22301 & n38265 ;
  assign n38271 = n38270 ^ n38266 ^ n8254 ;
  assign n38272 = ~n15533 & n20508 ;
  assign n38273 = n13332 & ~n14755 ;
  assign n38274 = n38273 ^ n2557 ^ 1'b0 ;
  assign n38275 = ( n3264 & ~n30224 ) | ( n3264 & n38274 ) | ( ~n30224 & n38274 ) ;
  assign n38276 = n24387 ^ n12910 ^ 1'b0 ;
  assign n38277 = n38275 & n38276 ;
  assign n38278 = ( n2911 & ~n11584 ) | ( n2911 & n38277 ) | ( ~n11584 & n38277 ) ;
  assign n38279 = n19857 ^ n3136 ^ n1995 ;
  assign n38280 = n27705 ^ n17546 ^ 1'b0 ;
  assign n38281 = n15657 | n38280 ;
  assign n38282 = n798 & ~n2529 ;
  assign n38283 = n38282 ^ n3979 ^ 1'b0 ;
  assign n38284 = n22421 & ~n38283 ;
  assign n38285 = n19441 & n28304 ;
  assign n38286 = ~n2075 & n38285 ;
  assign n38287 = n38286 ^ n17433 ^ 1'b0 ;
  assign n38288 = n17682 ^ n4708 ^ 1'b0 ;
  assign n38289 = ( n3862 & ~n20361 ) | ( n3862 & n38288 ) | ( ~n20361 & n38288 ) ;
  assign n38290 = ( n16459 & ~n18008 ) | ( n16459 & n30179 ) | ( ~n18008 & n30179 ) ;
  assign n38291 = n38290 ^ n28214 ^ 1'b0 ;
  assign n38292 = n38291 ^ n36869 ^ 1'b0 ;
  assign n38293 = n29540 & n38292 ;
  assign n38294 = n38293 ^ n8663 ^ n4883 ;
  assign n38295 = n36670 ^ n7609 ^ 1'b0 ;
  assign n38296 = ( ~n10644 & n12684 ) | ( ~n10644 & n15630 ) | ( n12684 & n15630 ) ;
  assign n38297 = n18205 & n22847 ;
  assign n38298 = ( n2970 & ~n34242 ) | ( n2970 & n38297 ) | ( ~n34242 & n38297 ) ;
  assign n38299 = n32616 ^ n16559 ^ n6419 ;
  assign n38300 = n5702 ^ n1106 ^ 1'b0 ;
  assign n38301 = n2447 | n38300 ;
  assign n38302 = n7221 & ~n25856 ;
  assign n38303 = ~n38301 & n38302 ;
  assign n38304 = ~n38299 & n38303 ;
  assign n38305 = n4944 ^ n2422 ^ 1'b0 ;
  assign n38306 = n9290 & ~n38305 ;
  assign n38307 = n33156 ^ n12675 ^ n1397 ;
  assign n38308 = n16433 ^ n15943 ^ n1597 ;
  assign n38309 = ( ~n8907 & n37354 ) | ( ~n8907 & n38308 ) | ( n37354 & n38308 ) ;
  assign n38310 = ( n38306 & n38307 ) | ( n38306 & n38309 ) | ( n38307 & n38309 ) ;
  assign n38317 = n18283 & ~n31014 ;
  assign n38318 = ~n11986 & n38317 ;
  assign n38314 = n1342 & ~n19937 ;
  assign n38315 = n38314 ^ n19359 ^ 1'b0 ;
  assign n38316 = n38315 ^ n14151 ^ 1'b0 ;
  assign n38311 = ( n3323 & n15784 ) | ( n3323 & ~n17378 ) | ( n15784 & ~n17378 ) ;
  assign n38312 = n28855 | n38311 ;
  assign n38313 = n38312 ^ n17728 ^ n15308 ;
  assign n38319 = n38318 ^ n38316 ^ n38313 ;
  assign n38320 = n33730 ^ n14937 ^ 1'b0 ;
  assign n38321 = n19003 & n38320 ;
  assign n38322 = n38321 ^ n28793 ^ 1'b0 ;
  assign n38323 = n8495 & n38322 ;
  assign n38324 = n8199 & ~n21412 ;
  assign n38325 = n32143 ^ n13614 ^ 1'b0 ;
  assign n38326 = n38324 | n38325 ;
  assign n38327 = n4478 | n22981 ;
  assign n38328 = n38327 ^ n29630 ^ n29527 ;
  assign n38329 = n27485 ^ n7592 ^ 1'b0 ;
  assign n38330 = n1395 & n38329 ;
  assign n38331 = n17022 | n38330 ;
  assign n38332 = n11245 & n32651 ;
  assign n38333 = n38332 ^ n5687 ^ 1'b0 ;
  assign n38334 = n20645 | n22531 ;
  assign n38335 = n6274 ^ n6173 ^ n4464 ;
  assign n38336 = n38335 ^ n8328 ^ 1'b0 ;
  assign n38337 = n33799 ^ n25821 ^ 1'b0 ;
  assign n38338 = n38337 ^ n23930 ^ 1'b0 ;
  assign n38339 = n38336 & ~n38338 ;
  assign n38340 = n8671 | n30864 ;
  assign n38341 = n27732 & ~n38340 ;
  assign n38342 = ( n1734 & ~n13272 ) | ( n1734 & n26654 ) | ( ~n13272 & n26654 ) ;
  assign n38343 = n38342 ^ n21894 ^ n15258 ;
  assign n38344 = n28983 & n31919 ;
  assign n38345 = n18045 & ~n21329 ;
  assign n38346 = ~n18045 & n38345 ;
  assign n38347 = ( ~n34723 & n37233 ) | ( ~n34723 & n38346 ) | ( n37233 & n38346 ) ;
  assign n38348 = n31151 ^ n14486 ^ 1'b0 ;
  assign n38349 = n9205 & n38348 ;
  assign n38350 = n35685 ^ n19837 ^ 1'b0 ;
  assign n38351 = n25700 ^ n15085 ^ 1'b0 ;
  assign n38352 = n36923 & ~n38351 ;
  assign n38353 = n30310 ^ n15482 ^ 1'b0 ;
  assign n38354 = ~n18256 & n38353 ;
  assign n38355 = n34566 ^ n33502 ^ n21419 ;
  assign n38356 = n10781 ^ n6287 ^ n4732 ;
  assign n38357 = n38356 ^ n11212 ^ n10179 ;
  assign n38358 = n34946 ^ n12698 ^ 1'b0 ;
  assign n38359 = ~n38357 & n38358 ;
  assign n38360 = ~n611 & n10613 ;
  assign n38361 = n38360 ^ n4727 ^ 1'b0 ;
  assign n38362 = n23312 & ~n34912 ;
  assign n38363 = n38362 ^ n18811 ^ 1'b0 ;
  assign n38364 = n7510 & n23320 ;
  assign n38366 = ( n3887 & ~n8988 ) | ( n3887 & n16662 ) | ( ~n8988 & n16662 ) ;
  assign n38367 = n31791 & n38366 ;
  assign n38368 = n38367 ^ n14747 ^ 1'b0 ;
  assign n38365 = n4484 & n14793 ;
  assign n38369 = n38368 ^ n38365 ^ 1'b0 ;
  assign n38370 = n9169 & ~n38252 ;
  assign n38371 = ( n9695 & ~n17617 ) | ( n9695 & n21029 ) | ( ~n17617 & n21029 ) ;
  assign n38372 = ( n600 & ~n35292 ) | ( n600 & n38371 ) | ( ~n35292 & n38371 ) ;
  assign n38373 = ( n5323 & n9658 ) | ( n5323 & ~n38372 ) | ( n9658 & ~n38372 ) ;
  assign n38374 = n18765 & ~n19677 ;
  assign n38375 = n3837 | n37678 ;
  assign n38376 = x52 & ~n7547 ;
  assign n38377 = n20053 & n38376 ;
  assign n38378 = ( n5289 & n9803 ) | ( n5289 & ~n23040 ) | ( n9803 & ~n23040 ) ;
  assign n38379 = n3770 ^ n1611 ^ 1'b0 ;
  assign n38380 = n6441 & ~n7347 ;
  assign n38381 = n799 | n10184 ;
  assign n38382 = n38380 & ~n38381 ;
  assign n38383 = ( n895 & n9343 ) | ( n895 & n34040 ) | ( n9343 & n34040 ) ;
  assign n38384 = ( n625 & ~n38382 ) | ( n625 & n38383 ) | ( ~n38382 & n38383 ) ;
  assign n38385 = n25433 & n38384 ;
  assign n38386 = n38385 ^ n16748 ^ n3485 ;
  assign n38387 = n7161 | n18054 ;
  assign n38388 = n36949 ^ n10487 ^ 1'b0 ;
  assign n38389 = n3534 & n38388 ;
  assign n38390 = n31134 | n38389 ;
  assign n38391 = n6401 & n17614 ;
  assign n38392 = n38391 ^ n16325 ^ n550 ;
  assign n38393 = n9371 ^ n4139 ^ 1'b0 ;
  assign n38394 = n12048 | n38393 ;
  assign n38395 = n38394 ^ n15586 ^ 1'b0 ;
  assign n38396 = ( ~x156 & n3858 ) | ( ~x156 & n21036 ) | ( n3858 & n21036 ) ;
  assign n38397 = ( n3548 & n19967 ) | ( n3548 & ~n22678 ) | ( n19967 & ~n22678 ) ;
  assign n38398 = n38397 ^ n21724 ^ 1'b0 ;
  assign n38399 = n7146 ^ n7092 ^ 1'b0 ;
  assign n38400 = n31352 | n38399 ;
  assign n38401 = n20430 ^ n1075 ^ 1'b0 ;
  assign n38402 = n6480 | n38401 ;
  assign n38403 = n38402 ^ n6891 ^ 1'b0 ;
  assign n38404 = n38403 ^ n34364 ^ 1'b0 ;
  assign n38405 = n12618 & ~n38404 ;
  assign n38409 = ( ~n12426 & n31631 ) | ( ~n12426 & n34912 ) | ( n31631 & n34912 ) ;
  assign n38406 = n8996 ^ n2667 ^ 1'b0 ;
  assign n38407 = n38406 ^ n8304 ^ 1'b0 ;
  assign n38408 = n38407 ^ n3736 ^ n782 ;
  assign n38410 = n38409 ^ n38408 ^ 1'b0 ;
  assign n38411 = n2983 | n12048 ;
  assign n38412 = n340 & ~n38411 ;
  assign n38413 = n38412 ^ n37466 ^ n15001 ;
  assign n38414 = ~n20479 & n38086 ;
  assign n38415 = ( n22459 & ~n26968 ) | ( n22459 & n27259 ) | ( ~n26968 & n27259 ) ;
  assign n38416 = n38415 ^ n17060 ^ 1'b0 ;
  assign n38417 = ( ~n22269 & n33680 ) | ( ~n22269 & n38416 ) | ( n33680 & n38416 ) ;
  assign n38418 = n20791 ^ n7476 ^ n4419 ;
  assign n38419 = n495 ^ n284 ^ 1'b0 ;
  assign n38420 = n3975 & n38419 ;
  assign n38423 = n17958 ^ n5990 ^ 1'b0 ;
  assign n38424 = n4382 | n38423 ;
  assign n38421 = n15525 & ~n18780 ;
  assign n38422 = ~n7581 & n38421 ;
  assign n38425 = n38424 ^ n38422 ^ n16326 ;
  assign n38426 = n4432 | n9687 ;
  assign n38427 = ~n18781 & n38426 ;
  assign n38428 = n38425 | n38427 ;
  assign n38429 = n38420 | n38428 ;
  assign n38430 = ( ~n1748 & n27510 ) | ( ~n1748 & n38429 ) | ( n27510 & n38429 ) ;
  assign n38431 = n3110 & ~n8858 ;
  assign n38432 = n24197 & n38431 ;
  assign n38433 = n6421 & ~n32277 ;
  assign n38434 = ~n8475 & n38433 ;
  assign n38435 = n934 & n38434 ;
  assign n38436 = n7143 | n9161 ;
  assign n38437 = n38436 ^ n10819 ^ 1'b0 ;
  assign n38438 = n38437 ^ n24395 ^ n5251 ;
  assign n38439 = n34491 ^ n3175 ^ 1'b0 ;
  assign n38440 = n10314 & ~n38439 ;
  assign n38441 = ~n38438 & n38440 ;
  assign n38442 = n481 & ~n20483 ;
  assign n38443 = n38442 ^ n22523 ^ 1'b0 ;
  assign n38444 = n10631 & n20336 ;
  assign n38445 = n38444 ^ n17410 ^ 1'b0 ;
  assign n38446 = n38445 ^ n11278 ^ n3411 ;
  assign n38447 = ( n15169 & ~n26482 ) | ( n15169 & n30517 ) | ( ~n26482 & n30517 ) ;
  assign n38448 = ( n7211 & n8083 ) | ( n7211 & n14141 ) | ( n8083 & n14141 ) ;
  assign n38449 = ~n1933 & n38448 ;
  assign n38450 = ~n8896 & n38449 ;
  assign n38451 = n3120 & ~n38450 ;
  assign n38452 = n15282 & ~n17952 ;
  assign n38453 = n38452 ^ n20836 ^ 1'b0 ;
  assign n38454 = n4810 & ~n18361 ;
  assign n38455 = n15862 & n24005 ;
  assign n38456 = ~n8657 & n38455 ;
  assign n38457 = n4509 | n31139 ;
  assign n38458 = n38456 & ~n38457 ;
  assign n38459 = n20517 ^ n1883 ^ 1'b0 ;
  assign n38461 = n29378 ^ n4727 ^ x248 ;
  assign n38460 = n20991 | n28203 ;
  assign n38462 = n38461 ^ n38460 ^ n23274 ;
  assign n38463 = n34544 ^ n29824 ^ 1'b0 ;
  assign n38465 = n37584 ^ n3644 ^ n2529 ;
  assign n38466 = n27647 & n38465 ;
  assign n38464 = n27540 ^ n22306 ^ n12413 ;
  assign n38467 = n38466 ^ n38464 ^ n10647 ;
  assign n38468 = ( n1331 & ~n8098 ) | ( n1331 & n26636 ) | ( ~n8098 & n26636 ) ;
  assign n38469 = n38468 ^ n16252 ^ 1'b0 ;
  assign n38470 = n38469 ^ n9405 ^ 1'b0 ;
  assign n38471 = n36268 ^ n28733 ^ 1'b0 ;
  assign n38472 = n4459 | n19677 ;
  assign n38473 = n38472 ^ n5916 ^ 1'b0 ;
  assign n38474 = ( ~n790 & n27126 ) | ( ~n790 & n38473 ) | ( n27126 & n38473 ) ;
  assign n38475 = n6907 ^ n2249 ^ 1'b0 ;
  assign n38476 = n2040 & n38475 ;
  assign n38477 = n38476 ^ n1285 ^ 1'b0 ;
  assign n38478 = n28006 & n38477 ;
  assign n38479 = n38478 ^ n37112 ^ n23528 ;
  assign n38480 = ~n16960 & n21102 ;
  assign n38481 = ~n17652 & n38480 ;
  assign n38482 = n38481 ^ n22546 ^ 1'b0 ;
  assign n38483 = n597 & ~n21157 ;
  assign n38484 = ~n22232 & n38483 ;
  assign n38485 = n38484 ^ n27303 ^ 1'b0 ;
  assign n38486 = n38019 & ~n38485 ;
  assign n38487 = ( n13748 & ~n25204 ) | ( n13748 & n26768 ) | ( ~n25204 & n26768 ) ;
  assign n38488 = n38487 ^ n35781 ^ 1'b0 ;
  assign n38489 = n10873 & ~n38488 ;
  assign n38490 = n3301 & ~n20683 ;
  assign n38491 = n15943 | n17044 ;
  assign n38492 = n36996 | n38491 ;
  assign n38493 = n8858 | n38492 ;
  assign n38494 = n3756 | n30215 ;
  assign n38495 = ( n8278 & n10520 ) | ( n8278 & ~n34305 ) | ( n10520 & ~n34305 ) ;
  assign n38496 = n16310 ^ n5676 ^ 1'b0 ;
  assign n38497 = n19233 & ~n38496 ;
  assign n38498 = ~n18994 & n38497 ;
  assign n38499 = n6548 & ~n19180 ;
  assign n38500 = n38499 ^ n15175 ^ n13806 ;
  assign n38501 = n38500 ^ n28313 ^ n16720 ;
  assign n38502 = ( ~n4759 & n25179 ) | ( ~n4759 & n37624 ) | ( n25179 & n37624 ) ;
  assign n38503 = ( ~n4309 & n8717 ) | ( ~n4309 & n38315 ) | ( n8717 & n38315 ) ;
  assign n38504 = n32720 ^ n625 ^ 1'b0 ;
  assign n38505 = n21834 | n34936 ;
  assign n38506 = n38505 ^ n15271 ^ 1'b0 ;
  assign n38507 = n7415 ^ n3041 ^ 1'b0 ;
  assign n38508 = n20179 & n38507 ;
  assign n38509 = ( n18797 & n29395 ) | ( n18797 & n38508 ) | ( n29395 & n38508 ) ;
  assign n38510 = n18805 | n38509 ;
  assign n38511 = n38510 ^ n2117 ^ 1'b0 ;
  assign n38512 = n38506 & n38511 ;
  assign n38513 = ( n5874 & n20924 ) | ( n5874 & ~n29547 ) | ( n20924 & ~n29547 ) ;
  assign n38514 = ~n28414 & n38513 ;
  assign n38515 = ( n1912 & n26151 ) | ( n1912 & n35204 ) | ( n26151 & n35204 ) ;
  assign n38516 = n3616 & ~n12190 ;
  assign n38517 = n38516 ^ n8030 ^ 1'b0 ;
  assign n38518 = n38517 ^ n23633 ^ n21837 ;
  assign n38519 = ~n5541 & n13715 ;
  assign n38520 = ~n30770 & n38519 ;
  assign n38521 = n11656 ^ n7212 ^ n1743 ;
  assign n38522 = ( ~n5436 & n11840 ) | ( ~n5436 & n38521 ) | ( n11840 & n38521 ) ;
  assign n38523 = n38522 ^ n16860 ^ 1'b0 ;
  assign n38524 = ~n38520 & n38523 ;
  assign n38525 = n18840 & ~n22851 ;
  assign n38526 = n28256 & n38525 ;
  assign n38527 = n11156 ^ n6969 ^ x44 ;
  assign n38528 = n38527 ^ n27743 ^ 1'b0 ;
  assign n38529 = ( n5740 & n11400 ) | ( n5740 & n12353 ) | ( n11400 & n12353 ) ;
  assign n38530 = ( n29221 & n32761 ) | ( n29221 & ~n38529 ) | ( n32761 & ~n38529 ) ;
  assign n38531 = n7693 ^ n2846 ^ 1'b0 ;
  assign n38532 = n10371 ^ n4963 ^ 1'b0 ;
  assign n38533 = n22814 & ~n38532 ;
  assign n38534 = n38533 ^ n35214 ^ n10146 ;
  assign n38535 = n9724 & ~n13308 ;
  assign n38536 = n11227 & n38535 ;
  assign n38537 = n38536 ^ n8018 ^ 1'b0 ;
  assign n38538 = n16077 & ~n38537 ;
  assign n38539 = ~n8632 & n14936 ;
  assign n38540 = n38539 ^ n29560 ^ 1'b0 ;
  assign n38541 = n9288 ^ n6068 ^ 1'b0 ;
  assign n38542 = n25173 ^ n15438 ^ 1'b0 ;
  assign n38543 = n15792 & n38542 ;
  assign n38544 = n4557 ^ n551 ^ 1'b0 ;
  assign n38545 = n6683 | n38544 ;
  assign n38546 = n38543 | n38545 ;
  assign n38547 = ( n9868 & n38541 ) | ( n9868 & ~n38546 ) | ( n38541 & ~n38546 ) ;
  assign n38548 = n38547 ^ n14753 ^ n3858 ;
  assign n38549 = n20703 ^ n16555 ^ 1'b0 ;
  assign n38550 = n17952 | n38549 ;
  assign n38551 = n617 | n27799 ;
  assign n38552 = n14403 & ~n38551 ;
  assign n38553 = ( n21306 & ~n38550 ) | ( n21306 & n38552 ) | ( ~n38550 & n38552 ) ;
  assign n38554 = n8741 | n16187 ;
  assign n38555 = n38554 ^ n31347 ^ 1'b0 ;
  assign n38556 = n22688 ^ n20286 ^ n19324 ;
  assign n38557 = ( n13354 & ~n18642 ) | ( n13354 & n30107 ) | ( ~n18642 & n30107 ) ;
  assign n38558 = n38556 & ~n38557 ;
  assign n38559 = n15451 & n37595 ;
  assign n38560 = n28239 ^ n22385 ^ n21922 ;
  assign n38561 = n2402 & n11530 ;
  assign n38562 = n7485 & n38561 ;
  assign n38563 = n38562 ^ n25319 ^ n21344 ;
  assign n38564 = ( n24343 & n28223 ) | ( n24343 & n36295 ) | ( n28223 & n36295 ) ;
  assign n38565 = n8816 & n18992 ;
  assign n38566 = ~n18606 & n38565 ;
  assign n38567 = n38566 ^ n18226 ^ n9489 ;
  assign n38568 = n38567 ^ n18642 ^ 1'b0 ;
  assign n38569 = ~n3219 & n11527 ;
  assign n38570 = n38569 ^ n32226 ^ 1'b0 ;
  assign n38571 = n13604 ^ n3082 ^ 1'b0 ;
  assign n38572 = n38570 & ~n38571 ;
  assign n38573 = n9361 & n11116 ;
  assign n38574 = ~n3040 & n7291 ;
  assign n38575 = n8468 & n38574 ;
  assign n38576 = ~n2767 & n17477 ;
  assign n38577 = n20862 ^ n9747 ^ 1'b0 ;
  assign n38578 = ~n7801 & n38577 ;
  assign n38579 = n21675 ^ n20123 ^ n8933 ;
  assign n38580 = n25530 ^ n9658 ^ n3543 ;
  assign n38581 = n3568 ^ n938 ^ 1'b0 ;
  assign n38582 = n2384 & n38581 ;
  assign n38583 = n38582 ^ n580 ^ 1'b0 ;
  assign n38584 = n26348 | n38583 ;
  assign n38585 = n38580 | n38584 ;
  assign n38586 = ( n30381 & n32568 ) | ( n30381 & n38585 ) | ( n32568 & n38585 ) ;
  assign n38587 = n6227 ^ x42 ^ 1'b0 ;
  assign n38588 = n8981 & ~n38587 ;
  assign n38589 = n5493 & ~n22554 ;
  assign n38590 = ~n38588 & n38589 ;
  assign n38591 = n5097 ^ n4255 ^ 1'b0 ;
  assign n38592 = n30939 | n38591 ;
  assign n38596 = ( n8607 & n11897 ) | ( n8607 & ~n15327 ) | ( n11897 & ~n15327 ) ;
  assign n38597 = n38596 ^ n16838 ^ n8840 ;
  assign n38593 = n8463 ^ n3504 ^ 1'b0 ;
  assign n38594 = n38593 ^ n25536 ^ 1'b0 ;
  assign n38595 = n22116 & ~n38594 ;
  assign n38598 = n38597 ^ n38595 ^ n3794 ;
  assign n38599 = n38598 ^ n33609 ^ n29396 ;
  assign n38600 = ( n2078 & n23217 ) | ( n2078 & n37193 ) | ( n23217 & n37193 ) ;
  assign n38601 = n38600 ^ n30419 ^ n1900 ;
  assign n38602 = n6277 ^ n5640 ^ 1'b0 ;
  assign n38603 = n38602 ^ n16673 ^ n4247 ;
  assign n38604 = n38603 ^ n38427 ^ 1'b0 ;
  assign n38605 = ( ~n11990 & n23142 ) | ( ~n11990 & n27575 ) | ( n23142 & n27575 ) ;
  assign n38606 = n5982 ^ n1505 ^ 1'b0 ;
  assign n38607 = n2299 & n38606 ;
  assign n38608 = ( n25827 & n26372 ) | ( n25827 & ~n38607 ) | ( n26372 & ~n38607 ) ;
  assign n38609 = n22126 ^ n20231 ^ n2143 ;
  assign n38610 = ( n820 & ~n4036 ) | ( n820 & n14940 ) | ( ~n4036 & n14940 ) ;
  assign n38611 = n38610 ^ n24622 ^ 1'b0 ;
  assign n38612 = n38611 ^ n8085 ^ 1'b0 ;
  assign n38613 = ~n6245 & n19537 ;
  assign n38614 = n12967 & n38613 ;
  assign n38615 = n38614 ^ n22495 ^ n12620 ;
  assign n38616 = n22413 ^ n21883 ^ n2839 ;
  assign n38617 = ~n38615 & n38616 ;
  assign n38618 = ~n485 & n22888 ;
  assign n38619 = n5481 & n38618 ;
  assign n38620 = n1551 | n1834 ;
  assign n38621 = n38620 ^ n15570 ^ 1'b0 ;
  assign n38622 = n38621 ^ n4782 ^ 1'b0 ;
  assign n38623 = ~n38619 & n38622 ;
  assign n38624 = n18386 & n38623 ;
  assign n38625 = ~n14723 & n35924 ;
  assign n38626 = n23677 & n38625 ;
  assign n38627 = n7927 & n8725 ;
  assign n38628 = n5491 & n38627 ;
  assign n38629 = ( ~n4470 & n18892 ) | ( ~n4470 & n38628 ) | ( n18892 & n38628 ) ;
  assign n38630 = n5424 ^ n2775 ^ 1'b0 ;
  assign n38631 = n13785 & n38630 ;
  assign n38632 = n3697 & n38631 ;
  assign n38633 = n26466 & n38632 ;
  assign n38635 = n999 & n21500 ;
  assign n38634 = ~n2109 & n21404 ;
  assign n38636 = n38635 ^ n38634 ^ 1'b0 ;
  assign n38637 = ~n38316 & n38636 ;
  assign n38638 = ( n2758 & n23890 ) | ( n2758 & ~n35662 ) | ( n23890 & ~n35662 ) ;
  assign n38639 = n38638 ^ n20896 ^ n19666 ;
  assign n38640 = ( n4267 & n15047 ) | ( n4267 & n38639 ) | ( n15047 & n38639 ) ;
  assign n38641 = ( n7769 & n8486 ) | ( n7769 & ~n28010 ) | ( n8486 & ~n28010 ) ;
  assign n38642 = ( n3248 & n6815 ) | ( n3248 & ~n17614 ) | ( n6815 & ~n17614 ) ;
  assign n38643 = n38642 ^ n22702 ^ n4405 ;
  assign n38644 = n37725 ^ n25831 ^ n5111 ;
  assign n38645 = ( n15552 & n23731 ) | ( n15552 & ~n38644 ) | ( n23731 & ~n38644 ) ;
  assign n38646 = n38645 ^ n33062 ^ n23946 ;
  assign n38647 = n18028 ^ n10617 ^ n742 ;
  assign n38648 = ~n11929 & n38647 ;
  assign n38649 = n21060 ^ n10355 ^ n5793 ;
  assign n38650 = ( n15340 & ~n18373 ) | ( n15340 & n38649 ) | ( ~n18373 & n38649 ) ;
  assign n38651 = n17757 & ~n38650 ;
  assign n38652 = ~n5549 & n38651 ;
  assign n38653 = n35724 ^ n5177 ^ 1'b0 ;
  assign n38654 = ~n24708 & n25465 ;
  assign n38655 = n38654 ^ n21715 ^ n3138 ;
  assign n38659 = n5474 | n8975 ;
  assign n38660 = ( ~n24795 & n32354 ) | ( ~n24795 & n38659 ) | ( n32354 & n38659 ) ;
  assign n38656 = n12606 ^ n9534 ^ 1'b0 ;
  assign n38657 = n38656 ^ n36630 ^ 1'b0 ;
  assign n38658 = ~n10156 & n38657 ;
  assign n38661 = n38660 ^ n38658 ^ 1'b0 ;
  assign n38662 = n38655 & ~n38661 ;
  assign n38669 = ( n2602 & n9282 ) | ( n2602 & ~n13450 ) | ( n9282 & ~n13450 ) ;
  assign n38668 = n2761 | n25624 ;
  assign n38670 = n38669 ^ n38668 ^ 1'b0 ;
  assign n38663 = ( ~n426 & n2547 ) | ( ~n426 & n6209 ) | ( n2547 & n6209 ) ;
  assign n38664 = ( ~n4833 & n10370 ) | ( ~n4833 & n38663 ) | ( n10370 & n38663 ) ;
  assign n38665 = n15529 & ~n16021 ;
  assign n38666 = ~n38664 & n38665 ;
  assign n38667 = n38666 ^ n35745 ^ 1'b0 ;
  assign n38671 = n38670 ^ n38667 ^ n9798 ;
  assign n38672 = n8528 ^ n5357 ^ n3186 ;
  assign n38673 = ( ~n12334 & n14134 ) | ( ~n12334 & n28615 ) | ( n14134 & n28615 ) ;
  assign n38674 = n12447 & ~n38673 ;
  assign n38676 = n20620 ^ n2894 ^ 1'b0 ;
  assign n38675 = n6405 | n21841 ;
  assign n38677 = n38676 ^ n38675 ^ 1'b0 ;
  assign n38678 = n25318 & ~n38677 ;
  assign n38679 = n31840 ^ n3176 ^ 1'b0 ;
  assign n38680 = ~n25474 & n38679 ;
  assign n38681 = n12893 & n38680 ;
  assign n38682 = ~n7399 & n38681 ;
  assign n38685 = n13958 & n25545 ;
  assign n38683 = n9700 ^ n6778 ^ n1196 ;
  assign n38684 = x176 & n38683 ;
  assign n38686 = n38685 ^ n38684 ^ 1'b0 ;
  assign n38687 = n19831 | n27534 ;
  assign n38688 = n37097 ^ n19959 ^ n4504 ;
  assign n38689 = n12728 ^ n5804 ^ n3844 ;
  assign n38690 = n38689 ^ n1039 ^ x3 ;
  assign n38691 = n38188 ^ n36193 ^ 1'b0 ;
  assign n38692 = ( n8093 & ~n9887 ) | ( n8093 & n22160 ) | ( ~n9887 & n22160 ) ;
  assign n38693 = n578 ^ x10 ^ 1'b0 ;
  assign n38694 = n1749 & ~n38693 ;
  assign n38695 = n20646 | n23926 ;
  assign n38696 = n1786 & n34382 ;
  assign n38697 = n38696 ^ n38258 ^ 1'b0 ;
  assign n38702 = n1108 & ~n19855 ;
  assign n38703 = ~n16555 & n38702 ;
  assign n38698 = n7774 ^ n1061 ^ 1'b0 ;
  assign n38699 = n38698 ^ n7300 ^ n1662 ;
  assign n38700 = ~n26416 & n38699 ;
  assign n38701 = ~n37183 & n38700 ;
  assign n38704 = n38703 ^ n38701 ^ n28965 ;
  assign n38705 = n15214 ^ n12000 ^ 1'b0 ;
  assign n38706 = ~n36551 & n38705 ;
  assign n38707 = n12455 ^ n3440 ^ 1'b0 ;
  assign n38708 = n2782 & n38707 ;
  assign n38709 = n38708 ^ n11353 ^ 1'b0 ;
  assign n38710 = ( ~n27104 & n38706 ) | ( ~n27104 & n38709 ) | ( n38706 & n38709 ) ;
  assign n38711 = n2733 & n7396 ;
  assign n38712 = n15105 & n38711 ;
  assign n38713 = ( ~n20035 & n27256 ) | ( ~n20035 & n38712 ) | ( n27256 & n38712 ) ;
  assign n38714 = ( ~n747 & n2296 ) | ( ~n747 & n38713 ) | ( n2296 & n38713 ) ;
  assign n38715 = n14833 ^ n1604 ^ 1'b0 ;
  assign n38716 = n38715 ^ n25844 ^ n1497 ;
  assign n38717 = ( n7551 & n20625 ) | ( n7551 & ~n22835 ) | ( n20625 & ~n22835 ) ;
  assign n38718 = n38717 ^ n386 ^ 1'b0 ;
  assign n38719 = ~n15651 & n38718 ;
  assign n38720 = ( ~n9151 & n29943 ) | ( ~n9151 & n38719 ) | ( n29943 & n38719 ) ;
  assign n38721 = ~n25591 & n35541 ;
  assign n38722 = n780 & n38721 ;
  assign n38723 = ~n1039 & n2460 ;
  assign n38724 = n38723 ^ n35931 ^ 1'b0 ;
  assign n38726 = n13833 ^ n6382 ^ 1'b0 ;
  assign n38727 = ~n4669 & n38726 ;
  assign n38725 = n21465 & n25636 ;
  assign n38728 = n38727 ^ n38725 ^ 1'b0 ;
  assign n38730 = n3154 | n17574 ;
  assign n38729 = n26352 ^ n372 ^ 1'b0 ;
  assign n38731 = n38730 ^ n38729 ^ 1'b0 ;
  assign n38732 = n38731 ^ n7742 ^ 1'b0 ;
  assign n38733 = n16744 & ~n17379 ;
  assign n38736 = n5463 | n11483 ;
  assign n38734 = n4747 & ~n7318 ;
  assign n38735 = n38734 ^ n32848 ^ n7016 ;
  assign n38737 = n38736 ^ n38735 ^ n17729 ;
  assign n38738 = n24299 ^ n8134 ^ n7788 ;
  assign n38739 = n13535 ^ n1752 ^ 1'b0 ;
  assign n38740 = n1563 | n38739 ;
  assign n38741 = n18530 | n32736 ;
  assign n38746 = n8488 & n17928 ;
  assign n38747 = n38746 ^ n10228 ^ 1'b0 ;
  assign n38748 = n38747 ^ n11281 ^ 1'b0 ;
  assign n38749 = ~n32258 & n38748 ;
  assign n38742 = ( n4075 & n6800 ) | ( n4075 & n16195 ) | ( n6800 & n16195 ) ;
  assign n38743 = n38742 ^ n11770 ^ x100 ;
  assign n38744 = n38743 ^ n12203 ^ n5160 ;
  assign n38745 = n16262 & ~n38744 ;
  assign n38750 = n38749 ^ n38745 ^ 1'b0 ;
  assign n38751 = n12216 & n22761 ;
  assign n38752 = n38751 ^ n2241 ^ 1'b0 ;
  assign n38753 = ( ~n20055 & n34815 ) | ( ~n20055 & n38752 ) | ( n34815 & n38752 ) ;
  assign n38754 = n9814 | n15169 ;
  assign n38755 = n38754 ^ n30708 ^ 1'b0 ;
  assign n38756 = n38755 ^ n34339 ^ n7853 ;
  assign n38757 = n35503 ^ n26669 ^ 1'b0 ;
  assign n38758 = ~n2840 & n38757 ;
  assign n38759 = n5468 & ~n18323 ;
  assign n38760 = n38759 ^ n13499 ^ 1'b0 ;
  assign n38761 = n38760 ^ n25470 ^ 1'b0 ;
  assign n38762 = n38758 & ~n38761 ;
  assign n38763 = n29264 & n38762 ;
  assign n38764 = ( ~n5075 & n6142 ) | ( ~n5075 & n38763 ) | ( n6142 & n38763 ) ;
  assign n38765 = ( ~n35898 & n37175 ) | ( ~n35898 & n37417 ) | ( n37175 & n37417 ) ;
  assign n38771 = n9174 ^ n8088 ^ n3002 ;
  assign n38767 = n6237 & n9427 ;
  assign n38768 = n38767 ^ n19767 ^ 1'b0 ;
  assign n38769 = ( n16997 & ~n22915 ) | ( n16997 & n38768 ) | ( ~n22915 & n38768 ) ;
  assign n38766 = n5574 | n16836 ;
  assign n38770 = n38769 ^ n38766 ^ 1'b0 ;
  assign n38772 = n38771 ^ n38770 ^ n5532 ;
  assign n38773 = n38772 ^ n17807 ^ n9599 ;
  assign n38774 = n10201 & n21309 ;
  assign n38775 = n38774 ^ n18761 ^ 1'b0 ;
  assign n38776 = n31287 ^ n20679 ^ n19149 ;
  assign n38777 = n2077 & ~n35955 ;
  assign n38778 = n8120 | n9536 ;
  assign n38779 = n38778 ^ n32789 ^ 1'b0 ;
  assign n38780 = n17729 & ~n38779 ;
  assign n38781 = ~n20673 & n38780 ;
  assign n38782 = ~n25520 & n38781 ;
  assign n38788 = ~n777 & n1852 ;
  assign n38783 = n3840 | n4762 ;
  assign n38784 = n15572 & ~n38783 ;
  assign n38785 = n12205 & n12866 ;
  assign n38786 = n38785 ^ n1759 ^ 1'b0 ;
  assign n38787 = ~n38784 & n38786 ;
  assign n38789 = n38788 ^ n38787 ^ 1'b0 ;
  assign n38790 = n4158 & ~n13055 ;
  assign n38791 = ~n28408 & n38790 ;
  assign n38792 = ~n1121 & n15806 ;
  assign n38793 = n38792 ^ n26603 ^ 1'b0 ;
  assign n38794 = ( n261 & n16814 ) | ( n261 & ~n18531 ) | ( n16814 & ~n18531 ) ;
  assign n38795 = ~n3613 & n20869 ;
  assign n38796 = n38794 & n38795 ;
  assign n38797 = n38796 ^ n12843 ^ 1'b0 ;
  assign n38798 = ( n22675 & n22881 ) | ( n22675 & n38797 ) | ( n22881 & n38797 ) ;
  assign n38799 = n8304 | n29219 ;
  assign n38800 = n38799 ^ n4833 ^ 1'b0 ;
  assign n38801 = ( n12045 & n38180 ) | ( n12045 & n38800 ) | ( n38180 & n38800 ) ;
  assign n38802 = n38801 ^ n14273 ^ 1'b0 ;
  assign n38803 = n8578 ^ n1225 ^ n545 ;
  assign n38804 = n4126 ^ n3930 ^ x102 ;
  assign n38805 = n38804 ^ n31545 ^ n861 ;
  assign n38806 = n27882 ^ n15766 ^ 1'b0 ;
  assign n38807 = ~n9240 & n38806 ;
  assign n38808 = ~n9505 & n11544 ;
  assign n38809 = n5683 & ~n5842 ;
  assign n38810 = n38808 & n38809 ;
  assign n38811 = n11419 & n13556 ;
  assign n38812 = n406 | n36648 ;
  assign n38813 = n24881 | n29930 ;
  assign n38814 = n38813 ^ n4624 ^ 1'b0 ;
  assign n38815 = n5953 ^ n4261 ^ 1'b0 ;
  assign n38816 = n5451 & n38815 ;
  assign n38817 = ~n8813 & n38816 ;
  assign n38818 = n4423 & n38817 ;
  assign n38820 = ( n7750 & ~n25243 ) | ( n7750 & n33408 ) | ( ~n25243 & n33408 ) ;
  assign n38821 = n35919 & ~n38820 ;
  assign n38819 = n1269 & n13496 ;
  assign n38822 = n38821 ^ n38819 ^ 1'b0 ;
  assign n38824 = n11770 & ~n31996 ;
  assign n38825 = n38824 ^ n28726 ^ 1'b0 ;
  assign n38823 = n3769 & ~n25746 ;
  assign n38826 = n38825 ^ n38823 ^ 1'b0 ;
  assign n38827 = n9888 & n38826 ;
  assign n38828 = n28263 ^ n26781 ^ n18209 ;
  assign n38829 = ~n1412 & n19424 ;
  assign n38830 = n18505 & n38829 ;
  assign n38831 = ( n17776 & n26323 ) | ( n17776 & ~n38830 ) | ( n26323 & ~n38830 ) ;
  assign n38832 = n6474 | n23740 ;
  assign n38833 = ( n14688 & n25162 ) | ( n14688 & n38832 ) | ( n25162 & n38832 ) ;
  assign n38834 = n37723 ^ n26107 ^ n3504 ;
  assign n38835 = n8174 & ~n19985 ;
  assign n38836 = ~n38834 & n38835 ;
  assign n38837 = n499 & ~n19312 ;
  assign n38838 = n38837 ^ n10674 ^ 1'b0 ;
  assign n38839 = n3556 | n31468 ;
  assign n38840 = n32699 & ~n38839 ;
  assign n38841 = n26199 ^ n25663 ^ n8180 ;
  assign n38842 = n10678 & n21079 ;
  assign n38843 = ~n24154 & n38842 ;
  assign n38844 = n38843 ^ n17489 ^ n3575 ;
  assign n38845 = n15539 ^ n15081 ^ 1'b0 ;
  assign n38846 = n11851 ^ n4048 ^ 1'b0 ;
  assign n38847 = n5016 & ~n38846 ;
  assign n38848 = ( n7697 & n38845 ) | ( n7697 & n38847 ) | ( n38845 & n38847 ) ;
  assign n38849 = ~n14827 & n38848 ;
  assign n38851 = ( n3440 & n6785 ) | ( n3440 & n11087 ) | ( n6785 & n11087 ) ;
  assign n38850 = n23973 | n28366 ;
  assign n38852 = n38851 ^ n38850 ^ 1'b0 ;
  assign n38853 = n38852 ^ n34532 ^ n6829 ;
  assign n38854 = n10207 | n12974 ;
  assign n38855 = n524 & ~n12563 ;
  assign n38856 = n38855 ^ n23845 ^ n2961 ;
  assign n38857 = n23589 ^ n16485 ^ 1'b0 ;
  assign n38858 = n21554 & ~n26565 ;
  assign n38859 = ~n19196 & n38858 ;
  assign n38860 = n38859 ^ n3557 ^ 1'b0 ;
  assign n38862 = n25617 ^ n23848 ^ 1'b0 ;
  assign n38861 = n14677 | n19553 ;
  assign n38863 = n38862 ^ n38861 ^ 1'b0 ;
  assign n38864 = n4125 | n19726 ;
  assign n38865 = n15898 ^ n11741 ^ 1'b0 ;
  assign n38866 = n18568 & n38865 ;
  assign n38867 = ~n7790 & n38866 ;
  assign n38868 = n25349 ^ n1582 ^ 1'b0 ;
  assign n38869 = n38868 ^ n27883 ^ n3803 ;
  assign n38870 = n2506 & ~n9056 ;
  assign n38871 = n17385 & n38870 ;
  assign n38877 = n7724 & ~n12462 ;
  assign n38872 = n10411 ^ n3550 ^ 1'b0 ;
  assign n38873 = n16426 & n38872 ;
  assign n38874 = n38873 ^ n7006 ^ 1'b0 ;
  assign n38875 = n14249 | n38874 ;
  assign n38876 = n15980 & ~n38875 ;
  assign n38878 = n38877 ^ n38876 ^ 1'b0 ;
  assign n38879 = n17114 & ~n38878 ;
  assign n38880 = ( n5535 & ~n38871 ) | ( n5535 & n38879 ) | ( ~n38871 & n38879 ) ;
  assign n38881 = n4777 & ~n33588 ;
  assign n38882 = n38881 ^ n4713 ^ 1'b0 ;
  assign n38883 = ( ~n18729 & n30318 ) | ( ~n18729 & n38882 ) | ( n30318 & n38882 ) ;
  assign n38884 = ( n7941 & n29183 ) | ( n7941 & n38883 ) | ( n29183 & n38883 ) ;
  assign n38885 = n24320 ^ n23402 ^ n18330 ;
  assign n38886 = n12912 ^ n12800 ^ n9541 ;
  assign n38887 = n38886 ^ n16652 ^ 1'b0 ;
  assign n38888 = n29024 & n38887 ;
  assign n38894 = x3 & ~n13375 ;
  assign n38895 = n38894 ^ n17077 ^ n14052 ;
  assign n38896 = n19537 & n38895 ;
  assign n38890 = n5458 ^ n485 ^ 1'b0 ;
  assign n38891 = n11044 | n38890 ;
  assign n38889 = n37471 ^ n7617 ^ n3566 ;
  assign n38892 = n38891 ^ n38889 ^ 1'b0 ;
  assign n38893 = n7473 | n38892 ;
  assign n38897 = n38896 ^ n38893 ^ 1'b0 ;
  assign n38899 = n20836 & ~n29211 ;
  assign n38898 = n2666 | n3019 ;
  assign n38900 = n38899 ^ n38898 ^ 1'b0 ;
  assign n38901 = ( ~n266 & n12866 ) | ( ~n266 & n21420 ) | ( n12866 & n21420 ) ;
  assign n38902 = ~n26962 & n38901 ;
  assign n38903 = n38902 ^ n30673 ^ 1'b0 ;
  assign n38904 = x206 & ~n10155 ;
  assign n38905 = n38904 ^ n11722 ^ 1'b0 ;
  assign n38906 = n38905 ^ n9921 ^ 1'b0 ;
  assign n38907 = n2865 ^ n2236 ^ 1'b0 ;
  assign n38908 = ( ~n2004 & n25431 ) | ( ~n2004 & n38907 ) | ( n25431 & n38907 ) ;
  assign n38909 = n38908 ^ n22291 ^ n16121 ;
  assign n38910 = n19026 ^ n11350 ^ 1'b0 ;
  assign n38911 = n5059 & n38910 ;
  assign n38912 = n34662 ^ n16078 ^ 1'b0 ;
  assign n38913 = n13701 ^ n8140 ^ 1'b0 ;
  assign n38914 = n1801 & n38913 ;
  assign n38915 = ( n284 & n5639 ) | ( n284 & ~n10405 ) | ( n5639 & ~n10405 ) ;
  assign n38916 = n7801 & ~n38915 ;
  assign n38917 = n5946 | n38916 ;
  assign n38918 = n2306 & ~n38917 ;
  assign n38919 = n37284 ^ n36563 ^ 1'b0 ;
  assign n38921 = ( n2865 & ~n7080 ) | ( n2865 & n14474 ) | ( ~n7080 & n14474 ) ;
  assign n38920 = n36785 ^ n10774 ^ n1308 ;
  assign n38922 = n38921 ^ n38920 ^ n4553 ;
  assign n38923 = n30487 & n33756 ;
  assign n38924 = ( n4264 & ~n4473 ) | ( n4264 & n8884 ) | ( ~n4473 & n8884 ) ;
  assign n38925 = n38924 ^ n29458 ^ 1'b0 ;
  assign n38926 = ~n30876 & n38925 ;
  assign n38927 = n13186 & n34816 ;
  assign n38928 = n1552 & n38927 ;
  assign n38929 = n38928 ^ n394 ^ 1'b0 ;
  assign n38930 = n18414 | n37322 ;
  assign n38931 = x171 & n32760 ;
  assign n38932 = n27358 ^ n22479 ^ 1'b0 ;
  assign n38933 = n9978 | n38932 ;
  assign n38934 = n1958 & ~n38933 ;
  assign n38935 = n11215 & n38934 ;
  assign n38936 = n38935 ^ n18817 ^ 1'b0 ;
  assign n38937 = ~n6206 & n38936 ;
  assign n38938 = ~n2518 & n5951 ;
  assign n38939 = n38938 ^ n31241 ^ 1'b0 ;
  assign n38940 = n24169 & ~n33036 ;
  assign n38941 = n38940 ^ n36023 ^ 1'b0 ;
  assign n38942 = n15953 ^ n1037 ^ 1'b0 ;
  assign n38943 = n38942 ^ n27495 ^ 1'b0 ;
  assign n38944 = n8503 & n38943 ;
  assign n38947 = n3196 ^ n1385 ^ 1'b0 ;
  assign n38948 = n2043 | n38947 ;
  assign n38949 = n38948 ^ n28446 ^ 1'b0 ;
  assign n38945 = n13396 & ~n34288 ;
  assign n38946 = n10267 & n38945 ;
  assign n38950 = n38949 ^ n38946 ^ n20042 ;
  assign n38951 = ( n6534 & n11294 ) | ( n6534 & ~n11816 ) | ( n11294 & ~n11816 ) ;
  assign n38952 = n38951 ^ n27554 ^ n11117 ;
  assign n38953 = n30173 ^ n27667 ^ n13744 ;
  assign n38954 = n25660 ^ n6926 ^ n3484 ;
  assign n38955 = n330 & n1666 ;
  assign n38956 = ~n38954 & n38955 ;
  assign n38957 = n1732 & ~n4514 ;
  assign n38958 = n38957 ^ n30499 ^ 1'b0 ;
  assign n38959 = n28170 ^ n21222 ^ n20355 ;
  assign n38960 = n38959 ^ n30107 ^ 1'b0 ;
  assign n38961 = n5823 & ~n19786 ;
  assign n38962 = n38961 ^ n30521 ^ 1'b0 ;
  assign n38963 = n38962 ^ n13459 ^ 1'b0 ;
  assign n38964 = n38960 | n38963 ;
  assign n38965 = n11234 & ~n38964 ;
  assign n38966 = n8436 | n24162 ;
  assign n38967 = n38966 ^ n13635 ^ 1'b0 ;
  assign n38968 = ~n38424 & n38967 ;
  assign n38969 = n38968 ^ n18253 ^ n8465 ;
  assign n38970 = ( n21401 & n25139 ) | ( n21401 & n26655 ) | ( n25139 & n26655 ) ;
  assign n38971 = n6621 & ~n8818 ;
  assign n38972 = n734 & n38971 ;
  assign n38973 = n38972 ^ n32132 ^ 1'b0 ;
  assign n38974 = ( ~n27240 & n38970 ) | ( ~n27240 & n38973 ) | ( n38970 & n38973 ) ;
  assign n38975 = n22203 ^ n16693 ^ n11971 ;
  assign n38976 = n6390 & n9956 ;
  assign n38977 = ( ~n11339 & n23661 ) | ( ~n11339 & n38976 ) | ( n23661 & n38976 ) ;
  assign n38978 = n38977 ^ n36083 ^ 1'b0 ;
  assign n38979 = n21437 & ~n27087 ;
  assign n38980 = ~n1477 & n20851 ;
  assign n38981 = n38980 ^ n3939 ^ 1'b0 ;
  assign n38982 = n10468 & ~n26152 ;
  assign n38983 = n19134 | n34978 ;
  assign n38984 = n31365 | n38983 ;
  assign n38985 = n24095 ^ n23462 ^ n3504 ;
  assign n38986 = n38985 ^ n28037 ^ 1'b0 ;
  assign n38987 = n5699 | n26648 ;
  assign n38988 = n38987 ^ n802 ^ 1'b0 ;
  assign n38989 = n38988 ^ n38401 ^ n1430 ;
  assign n38990 = ( n6515 & n6998 ) | ( n6515 & ~n23689 ) | ( n6998 & ~n23689 ) ;
  assign n38991 = n28294 ^ n20155 ^ 1'b0 ;
  assign n38992 = n38990 & n38991 ;
  assign n38993 = ~n7154 & n26563 ;
  assign n38999 = ( n3315 & n5846 ) | ( n3315 & ~n12959 ) | ( n5846 & ~n12959 ) ;
  assign n39000 = n38999 ^ n15187 ^ n12801 ;
  assign n38997 = n773 | n21319 ;
  assign n38998 = n3953 & ~n38997 ;
  assign n38994 = ~n12670 & n18650 ;
  assign n38995 = ~n18650 & n38994 ;
  assign n38996 = ( n7433 & n19293 ) | ( n7433 & n38995 ) | ( n19293 & n38995 ) ;
  assign n39001 = n39000 ^ n38998 ^ n38996 ;
  assign n39002 = ( n462 & n22366 ) | ( n462 & n34835 ) | ( n22366 & n34835 ) ;
  assign n39003 = n7911 ^ n3323 ^ 1'b0 ;
  assign n39004 = n39003 ^ n32254 ^ 1'b0 ;
  assign n39005 = ~n9413 & n39004 ;
  assign n39006 = n31708 ^ n29985 ^ 1'b0 ;
  assign n39007 = n1099 & ~n39006 ;
  assign n39008 = n17922 & n39007 ;
  assign n39009 = n39008 ^ n6109 ^ 1'b0 ;
  assign n39010 = n10652 ^ n9730 ^ 1'b0 ;
  assign n39011 = n9559 ^ n3266 ^ 1'b0 ;
  assign n39012 = ~n15240 & n39011 ;
  assign n39013 = ( n13882 & n15030 ) | ( n13882 & ~n16462 ) | ( n15030 & ~n16462 ) ;
  assign n39014 = ~n15392 & n39013 ;
  assign n39015 = ( n1560 & ~n3843 ) | ( n1560 & n17728 ) | ( ~n3843 & n17728 ) ;
  assign n39016 = ( ~n7675 & n12900 ) | ( ~n7675 & n26201 ) | ( n12900 & n26201 ) ;
  assign n39017 = n7326 ^ n4731 ^ 1'b0 ;
  assign n39018 = n25968 & n32418 ;
  assign n39019 = n30153 ^ n28175 ^ n24833 ;
  assign n39020 = n32182 ^ n14561 ^ 1'b0 ;
  assign n39021 = n32476 & ~n39020 ;
  assign n39022 = n39021 ^ n25431 ^ n13477 ;
  assign n39023 = ( n6115 & n20856 ) | ( n6115 & ~n29130 ) | ( n20856 & ~n29130 ) ;
  assign n39024 = n11233 ^ n2197 ^ n1557 ;
  assign n39025 = ~n1590 & n39024 ;
  assign n39026 = ( n39022 & ~n39023 ) | ( n39022 & n39025 ) | ( ~n39023 & n39025 ) ;
  assign n39027 = n37137 ^ n4789 ^ 1'b0 ;
  assign n39028 = ~n18128 & n39027 ;
  assign n39029 = n12216 & ~n21052 ;
  assign n39030 = ~x52 & n39029 ;
  assign n39031 = n4503 | n20411 ;
  assign n39032 = n39031 ^ n10201 ^ 1'b0 ;
  assign n39033 = ( ~n4546 & n8239 ) | ( ~n4546 & n9964 ) | ( n8239 & n9964 ) ;
  assign n39034 = ( n5745 & n9989 ) | ( n5745 & ~n39033 ) | ( n9989 & ~n39033 ) ;
  assign n39035 = n33518 ^ n23949 ^ n23318 ;
  assign n39036 = n3945 & ~n8438 ;
  assign n39037 = n39036 ^ n26990 ^ n15994 ;
  assign n39038 = ( n11765 & ~n14199 ) | ( n11765 & n21596 ) | ( ~n14199 & n21596 ) ;
  assign n39039 = n36466 ^ n29472 ^ 1'b0 ;
  assign n39040 = ~n6434 & n9759 ;
  assign n39041 = n39040 ^ n16866 ^ 1'b0 ;
  assign n39042 = n39039 | n39041 ;
  assign n39043 = ( n8818 & ~n21177 ) | ( n8818 & n37802 ) | ( ~n21177 & n37802 ) ;
  assign n39044 = n2616 & n29353 ;
  assign n39045 = ~n29353 & n39044 ;
  assign n39046 = n12041 & ~n39045 ;
  assign n39047 = n39046 ^ n5242 ^ 1'b0 ;
  assign n39048 = ~n39043 & n39047 ;
  assign n39049 = n12879 ^ n10477 ^ 1'b0 ;
  assign n39050 = ( ~n22963 & n26324 ) | ( ~n22963 & n39049 ) | ( n26324 & n39049 ) ;
  assign n39051 = n39050 ^ n32842 ^ 1'b0 ;
  assign n39052 = n39048 & n39051 ;
  assign n39053 = n39052 ^ n21362 ^ 1'b0 ;
  assign n39054 = n7665 & ~n39053 ;
  assign n39055 = n17718 ^ n13112 ^ n662 ;
  assign n39056 = ( n17718 & n31169 ) | ( n17718 & ~n33868 ) | ( n31169 & ~n33868 ) ;
  assign n39057 = n13764 | n18106 ;
  assign n39058 = n39057 ^ n22677 ^ 1'b0 ;
  assign n39059 = n39058 ^ n14673 ^ 1'b0 ;
  assign n39060 = n11239 ^ n10270 ^ 1'b0 ;
  assign n39061 = n11646 & n39060 ;
  assign n39062 = n14117 | n14584 ;
  assign n39063 = n39062 ^ n2059 ^ 1'b0 ;
  assign n39064 = n2881 & ~n4383 ;
  assign n39065 = n39064 ^ n764 ^ 1'b0 ;
  assign n39066 = n39065 ^ n16378 ^ 1'b0 ;
  assign n39067 = ( n3865 & n17743 ) | ( n3865 & ~n39066 ) | ( n17743 & ~n39066 ) ;
  assign n39068 = ( n9168 & ~n12174 ) | ( n9168 & n32041 ) | ( ~n12174 & n32041 ) ;
  assign n39069 = n8403 ^ n2701 ^ 1'b0 ;
  assign n39070 = ( n9704 & n22081 ) | ( n9704 & n26002 ) | ( n22081 & n26002 ) ;
  assign n39071 = n18069 & n39070 ;
  assign n39072 = n31202 & ~n33690 ;
  assign n39073 = n39072 ^ n6413 ^ 1'b0 ;
  assign n39075 = ( n6380 & ~n6622 ) | ( n6380 & n7859 ) | ( ~n6622 & n7859 ) ;
  assign n39076 = ( ~n7638 & n28884 ) | ( ~n7638 & n39075 ) | ( n28884 & n39075 ) ;
  assign n39077 = n22006 ^ n2032 ^ 1'b0 ;
  assign n39078 = n39076 | n39077 ;
  assign n39074 = n21320 | n33388 ;
  assign n39079 = n39078 ^ n39074 ^ n10671 ;
  assign n39080 = ( n3761 & ~n6224 ) | ( n3761 & n16839 ) | ( ~n6224 & n16839 ) ;
  assign n39081 = n39080 ^ n6108 ^ n2549 ;
  assign n39082 = n39081 ^ n10571 ^ n468 ;
  assign n39083 = n39082 ^ n26192 ^ 1'b0 ;
  assign n39087 = n18370 ^ n9541 ^ n4327 ;
  assign n39084 = n9184 | n14531 ;
  assign n39085 = ( n29305 & n34309 ) | ( n29305 & ~n39084 ) | ( n34309 & ~n39084 ) ;
  assign n39086 = n32532 | n39085 ;
  assign n39088 = n39087 ^ n39086 ^ n32418 ;
  assign n39089 = ( n7797 & n25354 ) | ( n7797 & ~n34525 ) | ( n25354 & ~n34525 ) ;
  assign n39090 = ~n9997 & n31197 ;
  assign n39091 = n39090 ^ n2033 ^ 1'b0 ;
  assign n39092 = n1727 & n20816 ;
  assign n39093 = ( x189 & ~n16867 ) | ( x189 & n39092 ) | ( ~n16867 & n39092 ) ;
  assign n39094 = ( n18203 & n25605 ) | ( n18203 & n39093 ) | ( n25605 & n39093 ) ;
  assign n39095 = n2571 & ~n38063 ;
  assign n39096 = n39094 & n39095 ;
  assign n39099 = ~n17270 & n18114 ;
  assign n39100 = n39099 ^ x83 ^ 1'b0 ;
  assign n39098 = ( n1049 & n6575 ) | ( n1049 & ~n14856 ) | ( n6575 & ~n14856 ) ;
  assign n39101 = n39100 ^ n39098 ^ 1'b0 ;
  assign n39097 = ( ~n3250 & n14766 ) | ( ~n3250 & n30195 ) | ( n14766 & n30195 ) ;
  assign n39102 = n39101 ^ n39097 ^ n8494 ;
  assign n39103 = ( ~n1861 & n9725 ) | ( ~n1861 & n16143 ) | ( n9725 & n16143 ) ;
  assign n39104 = n24963 ^ n12116 ^ n2400 ;
  assign n39105 = ( n874 & n39103 ) | ( n874 & n39104 ) | ( n39103 & n39104 ) ;
  assign n39106 = n3664 | n10012 ;
  assign n39107 = ~n3101 & n4442 ;
  assign n39108 = n12401 & n39107 ;
  assign n39109 = n17250 & n21927 ;
  assign n39110 = n38865 ^ n4970 ^ x155 ;
  assign n39111 = ( n1826 & n2485 ) | ( n1826 & ~n21251 ) | ( n2485 & ~n21251 ) ;
  assign n39112 = n39111 ^ n32735 ^ 1'b0 ;
  assign n39113 = ~n33049 & n39112 ;
  assign n39114 = n39113 ^ n3385 ^ 1'b0 ;
  assign n39115 = n39110 | n39114 ;
  assign n39120 = n9552 & ~n9775 ;
  assign n39121 = n39120 ^ n11078 ^ 1'b0 ;
  assign n39119 = n25460 ^ n12998 ^ n324 ;
  assign n39116 = n36740 ^ n28270 ^ 1'b0 ;
  assign n39117 = ~n5509 & n7542 ;
  assign n39118 = ( ~n12899 & n39116 ) | ( ~n12899 & n39117 ) | ( n39116 & n39117 ) ;
  assign n39122 = n39121 ^ n39119 ^ n39118 ;
  assign n39123 = ~n5403 & n17597 ;
  assign n39124 = n39123 ^ n21225 ^ 1'b0 ;
  assign n39125 = n23470 ^ n8584 ^ n3441 ;
  assign n39126 = n31818 & ~n39125 ;
  assign n39127 = n1135 & ~n23954 ;
  assign n39128 = n39127 ^ n10207 ^ 1'b0 ;
  assign n39129 = n4959 | n13764 ;
  assign n39131 = ( n3157 & n5891 ) | ( n3157 & n8558 ) | ( n5891 & n8558 ) ;
  assign n39132 = n36397 ^ n11669 ^ 1'b0 ;
  assign n39133 = n39131 | n39132 ;
  assign n39130 = n2657 | n37861 ;
  assign n39134 = n39133 ^ n39130 ^ 1'b0 ;
  assign n39135 = n4970 & ~n26606 ;
  assign n39136 = ( ~n11027 & n27444 ) | ( ~n11027 & n39135 ) | ( n27444 & n39135 ) ;
  assign n39137 = n39136 ^ n16023 ^ 1'b0 ;
  assign n39138 = n10502 | n39137 ;
  assign n39139 = ~n31952 & n39138 ;
  assign n39140 = n34483 ^ n29410 ^ n11139 ;
  assign n39141 = ~n16464 & n17837 ;
  assign n39142 = n32015 & n39141 ;
  assign n39143 = ( n3266 & ~n38638 ) | ( n3266 & n39142 ) | ( ~n38638 & n39142 ) ;
  assign n39144 = n6379 | n23059 ;
  assign n39145 = n39144 ^ n14444 ^ 1'b0 ;
  assign n39146 = n31782 & ~n39145 ;
  assign n39147 = n15480 ^ n13133 ^ 1'b0 ;
  assign n39148 = ( ~n7973 & n20824 ) | ( ~n7973 & n21623 ) | ( n20824 & n21623 ) ;
  assign n39149 = ( n4068 & n20447 ) | ( n4068 & ~n39148 ) | ( n20447 & ~n39148 ) ;
  assign n39150 = n6311 | n39149 ;
  assign n39151 = n7670 & n15584 ;
  assign n39152 = ( ~n7323 & n11144 ) | ( ~n7323 & n25405 ) | ( n11144 & n25405 ) ;
  assign n39153 = n7118 & ~n39152 ;
  assign n39154 = n39153 ^ n20047 ^ 1'b0 ;
  assign n39155 = n23730 | n38521 ;
  assign n39156 = n36978 & ~n39155 ;
  assign n39157 = n11107 ^ n7226 ^ 1'b0 ;
  assign n39158 = n11237 & ~n39157 ;
  assign n39159 = ~n35457 & n39158 ;
  assign n39160 = n39159 ^ n28643 ^ 1'b0 ;
  assign n39161 = n18783 ^ n9607 ^ 1'b0 ;
  assign n39162 = n16548 | n39161 ;
  assign n39163 = n39162 ^ n19134 ^ 1'b0 ;
  assign n39164 = n22074 & n22546 ;
  assign n39165 = n39164 ^ n31974 ^ 1'b0 ;
  assign n39166 = n39165 ^ n11894 ^ 1'b0 ;
  assign n39169 = ( ~n6989 & n14917 ) | ( ~n6989 & n25504 ) | ( n14917 & n25504 ) ;
  assign n39167 = ~n14120 & n35994 ;
  assign n39168 = n22932 | n39167 ;
  assign n39170 = n39169 ^ n39168 ^ n19636 ;
  assign n39171 = ~n12952 & n13327 ;
  assign n39172 = ~n39170 & n39171 ;
  assign n39173 = n3420 & ~n6994 ;
  assign n39177 = n20120 ^ n9063 ^ 1'b0 ;
  assign n39174 = ~n1036 & n14818 ;
  assign n39175 = ~n8974 & n39174 ;
  assign n39176 = n15672 | n39175 ;
  assign n39178 = n39177 ^ n39176 ^ 1'b0 ;
  assign n39179 = ( ~n13508 & n13729 ) | ( ~n13508 & n17494 ) | ( n13729 & n17494 ) ;
  assign n39180 = n39178 & ~n39179 ;
  assign n39181 = ( n575 & ~n22105 ) | ( n575 & n24928 ) | ( ~n22105 & n24928 ) ;
  assign n39182 = n17614 ^ n1180 ^ 1'b0 ;
  assign n39184 = n32975 ^ n18615 ^ n9607 ;
  assign n39183 = ~n4737 & n24388 ;
  assign n39185 = n39184 ^ n39183 ^ 1'b0 ;
  assign n39186 = n13388 ^ n3977 ^ 1'b0 ;
  assign n39187 = n7057 & n39186 ;
  assign n39188 = n39187 ^ n15439 ^ 1'b0 ;
  assign n39189 = ~n4760 & n25915 ;
  assign n39190 = n28338 & n39189 ;
  assign n39191 = ( n5574 & n13461 ) | ( n5574 & n14844 ) | ( n13461 & n14844 ) ;
  assign n39192 = n38710 & ~n39191 ;
  assign n39193 = ~n28845 & n39192 ;
  assign n39194 = n30902 ^ n10745 ^ n8390 ;
  assign n39195 = n21152 & n22111 ;
  assign n39196 = n39195 ^ n9517 ^ 1'b0 ;
  assign n39197 = ~n16831 & n39196 ;
  assign n39198 = n6017 ^ n5270 ^ n742 ;
  assign n39199 = ( n39194 & ~n39197 ) | ( n39194 & n39198 ) | ( ~n39197 & n39198 ) ;
  assign n39200 = ( n19316 & n38581 ) | ( n19316 & ~n39199 ) | ( n38581 & ~n39199 ) ;
  assign n39201 = n11740 ^ n6606 ^ 1'b0 ;
  assign n39202 = n17430 & ~n37216 ;
  assign n39203 = n22674 ^ n2698 ^ 1'b0 ;
  assign n39204 = n17070 ^ n12871 ^ 1'b0 ;
  assign n39205 = n19352 & n39204 ;
  assign n39206 = ~n1834 & n5685 ;
  assign n39207 = n39206 ^ n4449 ^ 1'b0 ;
  assign n39208 = n39207 ^ n7869 ^ 1'b0 ;
  assign n39209 = n39208 ^ n20137 ^ n2256 ;
  assign n39210 = n27968 & n33746 ;
  assign n39211 = ( n1244 & n25167 ) | ( n1244 & n39210 ) | ( n25167 & n39210 ) ;
  assign n39212 = n7118 | n15288 ;
  assign n39213 = n11461 | n39212 ;
  assign n39214 = n29669 ^ n5324 ^ n2457 ;
  assign n39215 = n15087 | n39214 ;
  assign n39216 = n39213 | n39215 ;
  assign n39217 = n39216 ^ n10284 ^ n9674 ;
  assign n39218 = n4986 & ~n7301 ;
  assign n39219 = n39218 ^ n5660 ^ 1'b0 ;
  assign n39220 = n15328 ^ n14571 ^ 1'b0 ;
  assign n39221 = n29726 & n39220 ;
  assign n39222 = n26152 ^ n15386 ^ 1'b0 ;
  assign n39223 = n11220 | n39222 ;
  assign n39224 = n18245 | n24754 ;
  assign n39225 = n39223 & ~n39224 ;
  assign n39226 = n18770 & ~n32798 ;
  assign n39227 = ~n12750 & n28976 ;
  assign n39228 = n39227 ^ n31748 ^ 1'b0 ;
  assign n39229 = n39228 ^ n13569 ^ n6567 ;
  assign n39230 = n39229 ^ n10438 ^ n5660 ;
  assign n39231 = n32985 ^ n19707 ^ n12086 ;
  assign n39232 = n39231 ^ n19951 ^ n10562 ;
  assign n39233 = n28378 ^ n19974 ^ 1'b0 ;
  assign n39234 = n39233 ^ n9002 ^ 1'b0 ;
  assign n39235 = n20763 & ~n39234 ;
  assign n39236 = n31549 & n39235 ;
  assign n39237 = n39094 & n39236 ;
  assign n39239 = n7428 & n7634 ;
  assign n39240 = n39239 ^ n5081 ^ 1'b0 ;
  assign n39238 = n301 | n34187 ;
  assign n39241 = n39240 ^ n39238 ^ n36185 ;
  assign n39242 = ~n10505 & n39241 ;
  assign n39243 = n39242 ^ n21730 ^ 1'b0 ;
  assign n39244 = n16444 & n36915 ;
  assign n39249 = n26432 ^ n14958 ^ n14916 ;
  assign n39246 = n4201 ^ n1344 ^ 1'b0 ;
  assign n39247 = n17368 & n39246 ;
  assign n39245 = n979 | n15699 ;
  assign n39248 = n39247 ^ n39245 ^ n7895 ;
  assign n39250 = n39249 ^ n39248 ^ n31749 ;
  assign n39251 = n34931 | n36815 ;
  assign n39252 = n10914 & n28407 ;
  assign n39253 = n39252 ^ n13766 ^ 1'b0 ;
  assign n39254 = n30084 ^ n25275 ^ 1'b0 ;
  assign n39255 = ( ~n11117 & n13206 ) | ( ~n11117 & n14518 ) | ( n13206 & n14518 ) ;
  assign n39256 = ~n3745 & n39255 ;
  assign n39257 = n39254 & n39256 ;
  assign n39258 = ~n4307 & n28171 ;
  assign n39259 = ~n1436 & n39258 ;
  assign n39260 = n11857 | n25476 ;
  assign n39261 = n39260 ^ n20169 ^ 1'b0 ;
  assign n39262 = n19299 & n24571 ;
  assign n39263 = n39262 ^ n5299 ^ 1'b0 ;
  assign n39264 = n1112 & ~n39263 ;
  assign n39265 = n39264 ^ n34065 ^ 1'b0 ;
  assign n39266 = ( ~n9827 & n22443 ) | ( ~n9827 & n39265 ) | ( n22443 & n39265 ) ;
  assign n39267 = n12780 & ~n27939 ;
  assign n39268 = ~n7650 & n39267 ;
  assign n39269 = n3692 & ~n26438 ;
  assign n39270 = ~n22812 & n39269 ;
  assign n39271 = n29094 ^ n19994 ^ n4144 ;
  assign n39272 = ( ~n39268 & n39270 ) | ( ~n39268 & n39271 ) | ( n39270 & n39271 ) ;
  assign n39287 = n826 & ~n7950 ;
  assign n39288 = ~n3584 & n39287 ;
  assign n39289 = n12406 & ~n39288 ;
  assign n39282 = n865 & ~n1688 ;
  assign n39283 = n39282 ^ n6712 ^ 1'b0 ;
  assign n39284 = n39283 ^ n14188 ^ 1'b0 ;
  assign n39285 = n10448 | n39284 ;
  assign n39279 = ~n9965 & n15203 ;
  assign n39280 = n39279 ^ n11836 ^ 1'b0 ;
  assign n39273 = n2716 & n16392 ;
  assign n39274 = n15739 | n39273 ;
  assign n39275 = n10376 & n16831 ;
  assign n39276 = ( n9817 & n18089 ) | ( n9817 & ~n39275 ) | ( n18089 & ~n39275 ) ;
  assign n39277 = ( n2380 & ~n39274 ) | ( n2380 & n39276 ) | ( ~n39274 & n39276 ) ;
  assign n39278 = n34931 | n39277 ;
  assign n39281 = n39280 ^ n39278 ^ 1'b0 ;
  assign n39286 = n39285 ^ n39281 ^ n21852 ;
  assign n39290 = n39289 ^ n39286 ^ n5553 ;
  assign n39291 = ~n6254 & n6267 ;
  assign n39292 = ~n20444 & n39291 ;
  assign n39293 = n15392 & ~n39292 ;
  assign n39294 = n39293 ^ n16836 ^ 1'b0 ;
  assign n39295 = ( ~n6497 & n29494 ) | ( ~n6497 & n39294 ) | ( n29494 & n39294 ) ;
  assign n39296 = n15827 ^ n13288 ^ n8535 ;
  assign n39297 = n23704 & ~n39296 ;
  assign n39298 = n7774 | n14254 ;
  assign n39299 = n39298 ^ n8177 ^ 1'b0 ;
  assign n39300 = ~n18484 & n39299 ;
  assign n39301 = ( ~n2338 & n18338 ) | ( ~n2338 & n23837 ) | ( n18338 & n23837 ) ;
  assign n39302 = n13303 & ~n14398 ;
  assign n39303 = n2142 | n30257 ;
  assign n39304 = n21036 & ~n39303 ;
  assign n39305 = n39304 ^ n3366 ^ 1'b0 ;
  assign n39306 = n14313 ^ n6694 ^ 1'b0 ;
  assign n39307 = n29454 & ~n39306 ;
  assign n39308 = n13285 ^ n8201 ^ 1'b0 ;
  assign n39309 = n9882 | n39308 ;
  assign n39310 = n26934 ^ n23659 ^ 1'b0 ;
  assign n39311 = ~n17187 & n20885 ;
  assign n39312 = ~n28990 & n39311 ;
  assign n39316 = n25165 ^ n12640 ^ n10227 ;
  assign n39313 = x221 & n3216 ;
  assign n39314 = ~n1874 & n39313 ;
  assign n39315 = ( n7766 & ~n24993 ) | ( n7766 & n39314 ) | ( ~n24993 & n39314 ) ;
  assign n39317 = n39316 ^ n39315 ^ n6582 ;
  assign n39318 = n21849 | n39317 ;
  assign n39323 = n7321 ^ n3786 ^ n510 ;
  assign n39324 = n12657 & ~n39323 ;
  assign n39319 = n19940 ^ n1122 ^ 1'b0 ;
  assign n39320 = n39319 ^ n13822 ^ 1'b0 ;
  assign n39321 = n29124 | n39320 ;
  assign n39322 = n39321 ^ n14137 ^ n1582 ;
  assign n39325 = n39324 ^ n39322 ^ 1'b0 ;
  assign n39326 = n32763 & n32789 ;
  assign n39327 = ( ~n964 & n9588 ) | ( ~n964 & n10583 ) | ( n9588 & n10583 ) ;
  assign n39328 = n39327 ^ n11992 ^ n1524 ;
  assign n39329 = n28973 & n39328 ;
  assign n39330 = n30000 ^ n27146 ^ 1'b0 ;
  assign n39331 = n321 & ~n39330 ;
  assign n39332 = ~n4053 & n6878 ;
  assign n39333 = n39332 ^ n23496 ^ 1'b0 ;
  assign n39334 = ~n26998 & n38863 ;
  assign n39335 = n916 & n39334 ;
  assign n39336 = n2740 & n2814 ;
  assign n39337 = n31610 & n39336 ;
  assign n39338 = n9362 | n39337 ;
  assign n39339 = n14910 ^ n10085 ^ 1'b0 ;
  assign n39340 = n39339 ^ n3923 ^ 1'b0 ;
  assign n39341 = n24933 & n25186 ;
  assign n39342 = n39340 & n39341 ;
  assign n39343 = n39342 ^ n29907 ^ 1'b0 ;
  assign n39344 = n39338 | n39343 ;
  assign n39345 = ( n4710 & ~n24033 ) | ( n4710 & n37217 ) | ( ~n24033 & n37217 ) ;
  assign n39346 = ( n8474 & ~n12168 ) | ( n8474 & n22894 ) | ( ~n12168 & n22894 ) ;
  assign n39347 = ( n1791 & ~n2502 ) | ( n1791 & n3783 ) | ( ~n2502 & n3783 ) ;
  assign n39349 = n7700 & n19930 ;
  assign n39350 = n19152 & n39349 ;
  assign n39348 = ( ~n3371 & n7390 ) | ( ~n3371 & n22871 ) | ( n7390 & n22871 ) ;
  assign n39351 = n39350 ^ n39348 ^ n23081 ;
  assign n39352 = n11414 & ~n31941 ;
  assign n39353 = n29452 & n39352 ;
  assign n39354 = n16522 | n39353 ;
  assign n39355 = n39354 ^ n6869 ^ 1'b0 ;
  assign n39356 = n31533 ^ n25409 ^ n782 ;
  assign n39358 = n1075 | n14891 ;
  assign n39359 = n39358 ^ n6829 ^ 1'b0 ;
  assign n39357 = n7390 | n14750 ;
  assign n39360 = n39359 ^ n39357 ^ 1'b0 ;
  assign n39361 = n39360 ^ n13929 ^ 1'b0 ;
  assign n39362 = n16377 ^ n7028 ^ 1'b0 ;
  assign n39363 = ~n7944 & n39362 ;
  assign n39364 = n39363 ^ n32727 ^ n25686 ;
  assign n39365 = n20169 ^ n4930 ^ 1'b0 ;
  assign n39366 = n21732 & ~n39365 ;
  assign n39367 = n38760 ^ n21883 ^ 1'b0 ;
  assign n39368 = n14644 & ~n39367 ;
  assign n39369 = n32242 & n39368 ;
  assign n39370 = n1401 | n9980 ;
  assign n39371 = n18620 & n39370 ;
  assign n39372 = n22817 ^ n17837 ^ n9363 ;
  assign n39373 = ( n12244 & ~n19209 ) | ( n12244 & n20611 ) | ( ~n19209 & n20611 ) ;
  assign n39374 = ( n11804 & n20691 ) | ( n11804 & n36549 ) | ( n20691 & n36549 ) ;
  assign n39375 = n21683 & n39374 ;
  assign n39376 = n39375 ^ n35277 ^ 1'b0 ;
  assign n39377 = n22303 | n23872 ;
  assign n39378 = n6984 | n14776 ;
  assign n39379 = n25833 | n39378 ;
  assign n39380 = n16695 & n39379 ;
  assign n39381 = n20629 & n26016 ;
  assign n39382 = ~n19478 & n39381 ;
  assign n39383 = n11851 | n15460 ;
  assign n39384 = n39383 ^ n10691 ^ 1'b0 ;
  assign n39385 = n36540 ^ n26866 ^ n8343 ;
  assign n39386 = n39385 ^ n18873 ^ 1'b0 ;
  assign n39387 = n4141 ^ n2770 ^ 1'b0 ;
  assign n39388 = n32680 ^ n13864 ^ n8210 ;
  assign n39389 = ~n12364 & n21833 ;
  assign n39390 = n39389 ^ n19905 ^ n13916 ;
  assign n39391 = n39390 ^ n32380 ^ n12516 ;
  assign n39392 = ( ~n10957 & n37464 ) | ( ~n10957 & n38149 ) | ( n37464 & n38149 ) ;
  assign n39393 = n17325 & n39392 ;
  assign n39394 = n39393 ^ n10012 ^ 1'b0 ;
  assign n39395 = ( n15066 & ~n29109 ) | ( n15066 & n39394 ) | ( ~n29109 & n39394 ) ;
  assign n39396 = n34779 ^ n23163 ^ 1'b0 ;
  assign n39397 = n9475 ^ n326 ^ 1'b0 ;
  assign n39398 = n3730 & n24989 ;
  assign n39399 = n322 & n39398 ;
  assign n39400 = n10229 ^ n6515 ^ 1'b0 ;
  assign n39401 = ~n16839 & n39400 ;
  assign n39402 = ( n3294 & n8902 ) | ( n3294 & n21573 ) | ( n8902 & n21573 ) ;
  assign n39403 = ~n3462 & n10120 ;
  assign n39404 = ~n7917 & n39403 ;
  assign n39405 = n1533 & ~n11591 ;
  assign n39406 = n39405 ^ n18410 ^ 1'b0 ;
  assign n39407 = ( n39402 & n39404 ) | ( n39402 & ~n39406 ) | ( n39404 & ~n39406 ) ;
  assign n39408 = ~n13526 & n39407 ;
  assign n39409 = ~x11 & n39408 ;
  assign n39410 = n39409 ^ n14858 ^ 1'b0 ;
  assign n39411 = n32392 ^ n32384 ^ 1'b0 ;
  assign n39412 = n39411 ^ n23017 ^ n2270 ;
  assign n39413 = n4659 & ~n39412 ;
  assign n39414 = ( ~n30818 & n31864 ) | ( ~n30818 & n39413 ) | ( n31864 & n39413 ) ;
  assign n39415 = n12425 | n18488 ;
  assign n39416 = n34768 ^ n26352 ^ 1'b0 ;
  assign n39417 = n39415 & n39416 ;
  assign n39418 = ( n10489 & ~n20780 ) | ( n10489 & n39417 ) | ( ~n20780 & n39417 ) ;
  assign n39419 = n1024 | n11965 ;
  assign n39420 = n12053 ^ n2870 ^ 1'b0 ;
  assign n39421 = n8880 | n39420 ;
  assign n39422 = n39421 ^ n9247 ^ 1'b0 ;
  assign n39423 = n22010 & n39422 ;
  assign n39424 = n39419 & n39423 ;
  assign n39425 = n809 & ~n17263 ;
  assign n39426 = n21590 & n39425 ;
  assign n39427 = ~n21129 & n26471 ;
  assign n39428 = n39427 ^ n13022 ^ 1'b0 ;
  assign n39430 = n11590 | n15321 ;
  assign n39429 = n22101 | n34583 ;
  assign n39431 = n39430 ^ n39429 ^ 1'b0 ;
  assign n39432 = n39431 ^ n27708 ^ 1'b0 ;
  assign n39433 = n21653 & n38472 ;
  assign n39434 = ~n1574 & n21527 ;
  assign n39435 = n36668 ^ n4793 ^ 1'b0 ;
  assign n39436 = ~n24946 & n39435 ;
  assign n39437 = n39436 ^ n26811 ^ 1'b0 ;
  assign n39443 = ~n17224 & n31594 ;
  assign n39444 = n30001 & n39443 ;
  assign n39441 = n32805 ^ n13748 ^ 1'b0 ;
  assign n39438 = n4684 & ~n29686 ;
  assign n39439 = n39438 ^ n31515 ^ 1'b0 ;
  assign n39440 = n39439 ^ n2573 ^ n2428 ;
  assign n39442 = n39441 ^ n39440 ^ n16244 ;
  assign n39445 = n39444 ^ n39442 ^ n6464 ;
  assign n39446 = ( n311 & ~n39437 ) | ( n311 & n39445 ) | ( ~n39437 & n39445 ) ;
  assign n39447 = ~n6235 & n9726 ;
  assign n39448 = n6346 & n39447 ;
  assign n39449 = n1975 & ~n4005 ;
  assign n39450 = n3109 ^ n2040 ^ 1'b0 ;
  assign n39451 = ~n19805 & n39450 ;
  assign n39452 = ~n13227 & n39451 ;
  assign n39453 = n39452 ^ n12585 ^ 1'b0 ;
  assign n39454 = n1521 & ~n39453 ;
  assign n39455 = n28256 ^ n19326 ^ n1932 ;
  assign n39456 = ~n30009 & n39455 ;
  assign n39457 = n3441 & n14273 ;
  assign n39458 = ( n10031 & n15154 ) | ( n10031 & ~n22240 ) | ( n15154 & ~n22240 ) ;
  assign n39459 = n17490 | n39458 ;
  assign n39460 = n15976 ^ n12234 ^ 1'b0 ;
  assign n39461 = n23180 ^ n20247 ^ 1'b0 ;
  assign n39462 = n12859 & n39461 ;
  assign n39467 = n17484 ^ n3983 ^ 1'b0 ;
  assign n39463 = n1331 | n7117 ;
  assign n39464 = n6625 | n39463 ;
  assign n39465 = n39464 ^ n18868 ^ 1'b0 ;
  assign n39466 = ~n27780 & n39465 ;
  assign n39468 = n39467 ^ n39466 ^ 1'b0 ;
  assign n39469 = n39118 ^ n8791 ^ 1'b0 ;
  assign n39470 = n17084 & ~n39469 ;
  assign n39471 = n10242 | n22448 ;
  assign n39472 = n16444 ^ n9431 ^ n6860 ;
  assign n39473 = n16062 ^ n10841 ^ 1'b0 ;
  assign n39474 = ~n29270 & n39473 ;
  assign n39475 = ( x21 & n1066 ) | ( x21 & ~n5551 ) | ( n1066 & ~n5551 ) ;
  assign n39476 = ~n18937 & n39475 ;
  assign n39477 = n39476 ^ n19274 ^ 1'b0 ;
  assign n39478 = n8446 ^ n8091 ^ 1'b0 ;
  assign n39479 = n28074 ^ n26203 ^ n7163 ;
  assign n39480 = n11833 ^ n722 ^ 1'b0 ;
  assign n39481 = ~n34850 & n39480 ;
  assign n39482 = n24558 ^ n10816 ^ 1'b0 ;
  assign n39483 = ( n26674 & n39481 ) | ( n26674 & ~n39482 ) | ( n39481 & ~n39482 ) ;
  assign n39484 = n31622 & n39483 ;
  assign n39485 = n20831 ^ n11838 ^ n5222 ;
  assign n39486 = ~n2468 & n39485 ;
  assign n39487 = ~n24508 & n39486 ;
  assign n39488 = x209 | n6634 ;
  assign n39489 = n6562 | n39488 ;
  assign n39490 = n26954 & ~n39489 ;
  assign n39491 = n8500 ^ x154 ^ 1'b0 ;
  assign n39492 = n39491 ^ n28134 ^ n24321 ;
  assign n39493 = ( n4342 & n5744 ) | ( n4342 & n23118 ) | ( n5744 & n23118 ) ;
  assign n39494 = n26943 ^ n1491 ^ 1'b0 ;
  assign n39495 = ~n10009 & n39494 ;
  assign n39496 = ( n1539 & n29949 ) | ( n1539 & ~n39495 ) | ( n29949 & ~n39495 ) ;
  assign n39497 = n39496 ^ n21778 ^ n2617 ;
  assign n39498 = ~n11019 & n24158 ;
  assign n39500 = n37430 ^ n6860 ^ 1'b0 ;
  assign n39501 = ( n3878 & ~n17593 ) | ( n3878 & n39500 ) | ( ~n17593 & n39500 ) ;
  assign n39499 = n17747 & n35972 ;
  assign n39502 = n39501 ^ n39499 ^ 1'b0 ;
  assign n39504 = ~n1118 & n11702 ;
  assign n39503 = n16302 & n28305 ;
  assign n39505 = n39504 ^ n39503 ^ 1'b0 ;
  assign n39506 = n38820 ^ x10 ^ 1'b0 ;
  assign n39507 = n22578 ^ n13120 ^ 1'b0 ;
  assign n39508 = n4242 | n39507 ;
  assign n39509 = n17565 & ~n39508 ;
  assign n39510 = n39509 ^ n21360 ^ 1'b0 ;
  assign n39511 = ( n33019 & n39506 ) | ( n33019 & n39510 ) | ( n39506 & n39510 ) ;
  assign n39512 = n9297 ^ n7061 ^ n5342 ;
  assign n39513 = ~n2328 & n26261 ;
  assign n39514 = ~n9655 & n39513 ;
  assign n39515 = ( ~n16237 & n31430 ) | ( ~n16237 & n39514 ) | ( n31430 & n39514 ) ;
  assign n39516 = ~n3360 & n39515 ;
  assign n39517 = n6033 & n39516 ;
  assign n39518 = ( n25175 & ~n33312 ) | ( n25175 & n39517 ) | ( ~n33312 & n39517 ) ;
  assign n39519 = n8240 & ~n26323 ;
  assign n39520 = ~n15166 & n39519 ;
  assign n39521 = n15037 | n29664 ;
  assign n39522 = n39521 ^ n6771 ^ 1'b0 ;
  assign n39523 = n39522 ^ n37538 ^ n11613 ;
  assign n39524 = ~n3232 & n39523 ;
  assign n39525 = n39524 ^ n15109 ^ 1'b0 ;
  assign n39526 = n26732 | n31644 ;
  assign n39527 = n39526 ^ n39360 ^ 1'b0 ;
  assign n39528 = ~n4364 & n17088 ;
  assign n39529 = ~n7822 & n39528 ;
  assign n39530 = n18189 ^ n7757 ^ 1'b0 ;
  assign n39531 = ( n18367 & n25314 ) | ( n18367 & ~n39530 ) | ( n25314 & ~n39530 ) ;
  assign n39532 = n14026 & ~n39531 ;
  assign n39533 = n39529 & n39532 ;
  assign n39534 = n3462 & ~n9237 ;
  assign n39535 = n39534 ^ n14938 ^ 1'b0 ;
  assign n39536 = n6766 | n39535 ;
  assign n39537 = n39536 ^ n17883 ^ 1'b0 ;
  assign n39538 = n21683 & ~n39537 ;
  assign n39539 = n39538 ^ n11272 ^ 1'b0 ;
  assign n39540 = n38623 ^ n21242 ^ n5222 ;
  assign n39541 = ( ~n761 & n5274 ) | ( ~n761 & n18919 ) | ( n5274 & n18919 ) ;
  assign n39542 = n25243 & ~n39541 ;
  assign n39543 = n15684 ^ n13923 ^ n7021 ;
  assign n39544 = ( ~n6580 & n21393 ) | ( ~n6580 & n39543 ) | ( n21393 & n39543 ) ;
  assign n39545 = ( n1327 & n26991 ) | ( n1327 & n39544 ) | ( n26991 & n39544 ) ;
  assign n39546 = n24986 ^ n17974 ^ 1'b0 ;
  assign n39547 = n281 & n39546 ;
  assign n39548 = ( ~x113 & n18318 ) | ( ~x113 & n34319 ) | ( n18318 & n34319 ) ;
  assign n39549 = ( n30399 & n39547 ) | ( n30399 & ~n39548 ) | ( n39547 & ~n39548 ) ;
  assign n39550 = n25906 & n32490 ;
  assign n39551 = n39550 ^ n29064 ^ 1'b0 ;
  assign n39552 = n39551 ^ n18279 ^ 1'b0 ;
  assign n39553 = n32305 ^ n6083 ^ 1'b0 ;
  assign n39554 = n14093 & ~n25105 ;
  assign n39555 = ~n35237 & n39554 ;
  assign n39556 = n7873 | n31749 ;
  assign n39557 = n39556 ^ n9481 ^ 1'b0 ;
  assign n39558 = ( n5408 & ~n5674 ) | ( n5408 & n24052 ) | ( ~n5674 & n24052 ) ;
  assign n39559 = n27048 ^ n648 ^ 1'b0 ;
  assign n39560 = ( n15433 & n36102 ) | ( n15433 & n36431 ) | ( n36102 & n36431 ) ;
  assign n39561 = n7842 & n25783 ;
  assign n39562 = n35099 & n39561 ;
  assign n39563 = n21049 & n22331 ;
  assign n39564 = n39563 ^ n14749 ^ 1'b0 ;
  assign n39565 = n9961 & ~n11684 ;
  assign n39566 = n11859 & n39565 ;
  assign n39567 = ( ~n15659 & n27703 ) | ( ~n15659 & n34443 ) | ( n27703 & n34443 ) ;
  assign n39568 = n8783 | n9354 ;
  assign n39570 = n8272 & n9762 ;
  assign n39571 = n39570 ^ n18563 ^ 1'b0 ;
  assign n39569 = ~n26535 & n32397 ;
  assign n39572 = n39571 ^ n39569 ^ 1'b0 ;
  assign n39573 = n19028 & n39572 ;
  assign n39574 = ~n39568 & n39573 ;
  assign n39575 = n39574 ^ n21052 ^ n15649 ;
  assign n39576 = n1814 | n37365 ;
  assign n39577 = n4974 & ~n39576 ;
  assign n39578 = n13774 & ~n26764 ;
  assign n39579 = ~n3109 & n39578 ;
  assign n39580 = n39577 & n39579 ;
  assign n39581 = n1917 | n11954 ;
  assign n39582 = n39581 ^ n11958 ^ 1'b0 ;
  assign n39583 = ( n7568 & ~n12356 ) | ( n7568 & n16842 ) | ( ~n12356 & n16842 ) ;
  assign n39584 = n39583 ^ n19085 ^ n11959 ;
  assign n39585 = n19419 ^ n7117 ^ n2694 ;
  assign n39586 = ( ~n12937 & n21226 ) | ( ~n12937 & n39585 ) | ( n21226 & n39585 ) ;
  assign n39587 = n20294 ^ n12163 ^ n2372 ;
  assign n39588 = n1178 | n39587 ;
  assign n39589 = n5238 & ~n39588 ;
  assign n39590 = ( n21410 & n37733 ) | ( n21410 & ~n39589 ) | ( n37733 & ~n39589 ) ;
  assign n39591 = n17155 ^ n15496 ^ n6860 ;
  assign n39592 = n5208 & ~n25320 ;
  assign n39593 = n11022 & n39592 ;
  assign n39594 = n39593 ^ n8735 ^ 1'b0 ;
  assign n39595 = ( ~n31425 & n39591 ) | ( ~n31425 & n39594 ) | ( n39591 & n39594 ) ;
  assign n39596 = n23358 ^ n18899 ^ 1'b0 ;
  assign n39597 = ~n26474 & n39596 ;
  assign n39598 = n9015 ^ n5212 ^ 1'b0 ;
  assign n39599 = n39597 & ~n39598 ;
  assign n39600 = ~n30342 & n38089 ;
  assign n39601 = n10885 & n39600 ;
  assign n39602 = n27825 & n39601 ;
  assign n39603 = n22700 ^ n7209 ^ n2723 ;
  assign n39604 = n39603 ^ n32374 ^ 1'b0 ;
  assign n39605 = n7015 & n39604 ;
  assign n39606 = ~n3759 & n16116 ;
  assign n39607 = n17385 & n39606 ;
  assign n39608 = ( n12761 & n39605 ) | ( n12761 & ~n39607 ) | ( n39605 & ~n39607 ) ;
  assign n39609 = ( n1878 & n34786 ) | ( n1878 & n35801 ) | ( n34786 & n35801 ) ;
  assign n39614 = n9079 & ~n23946 ;
  assign n39611 = ~n1555 & n16363 ;
  assign n39612 = n5039 & n39611 ;
  assign n39610 = ~n9839 & n18462 ;
  assign n39613 = n39612 ^ n39610 ^ 1'b0 ;
  assign n39615 = n39614 ^ n39613 ^ n12043 ;
  assign n39616 = n24731 ^ n8614 ^ 1'b0 ;
  assign n39617 = ~n25928 & n31406 ;
  assign n39618 = n21680 | n35227 ;
  assign n39619 = n39618 ^ n13964 ^ 1'b0 ;
  assign n39620 = n39619 ^ n11272 ^ 1'b0 ;
  assign n39621 = ~n39617 & n39620 ;
  assign n39622 = n9254 ^ n8566 ^ 1'b0 ;
  assign n39623 = n20311 | n32456 ;
  assign n39624 = n13347 ^ n2755 ^ 1'b0 ;
  assign n39625 = n39623 | n39624 ;
  assign n39626 = n39622 & ~n39625 ;
  assign n39627 = n774 & ~n23973 ;
  assign n39628 = n3204 ^ n2050 ^ 1'b0 ;
  assign n39629 = ( n12564 & n32627 ) | ( n12564 & ~n38660 ) | ( n32627 & ~n38660 ) ;
  assign n39630 = n4404 & n39629 ;
  assign n39631 = n35900 ^ n7462 ^ 1'b0 ;
  assign n39632 = n23868 ^ n9804 ^ 1'b0 ;
  assign n39633 = n3619 ^ n3298 ^ n1543 ;
  assign n39634 = ( n2336 & n2682 ) | ( n2336 & ~n14915 ) | ( n2682 & ~n14915 ) ;
  assign n39635 = ( n14644 & n14936 ) | ( n14644 & n35251 ) | ( n14936 & n35251 ) ;
  assign n39636 = n29380 ^ n12930 ^ n6480 ;
  assign n39637 = n39636 ^ n26097 ^ 1'b0 ;
  assign n39638 = ~n1475 & n7972 ;
  assign n39640 = n20468 ^ n5313 ^ 1'b0 ;
  assign n39641 = ~n6335 & n39640 ;
  assign n39639 = n31133 ^ n21845 ^ n18975 ;
  assign n39642 = n39641 ^ n39639 ^ 1'b0 ;
  assign n39643 = ( ~n32286 & n39638 ) | ( ~n32286 & n39642 ) | ( n39638 & n39642 ) ;
  assign n39645 = n16703 ^ n15756 ^ n3167 ;
  assign n39644 = ~n3440 & n37231 ;
  assign n39646 = n39645 ^ n39644 ^ 1'b0 ;
  assign n39647 = n26909 ^ n15835 ^ 1'b0 ;
  assign n39648 = n642 | n1056 ;
  assign n39649 = n642 & ~n39648 ;
  assign n39650 = n444 & n633 ;
  assign n39651 = n39649 & n39650 ;
  assign n39652 = n1601 & ~n39651 ;
  assign n39653 = ~n1601 & n39652 ;
  assign n39654 = ( n977 & n1378 ) | ( n977 & ~n6737 ) | ( n1378 & ~n6737 ) ;
  assign n39655 = n11340 & n39654 ;
  assign n39656 = n39653 & n39655 ;
  assign n39657 = ( n25174 & n35254 ) | ( n25174 & ~n39656 ) | ( n35254 & ~n39656 ) ;
  assign n39658 = n18796 ^ n476 ^ 1'b0 ;
  assign n39659 = n6866 | n39658 ;
  assign n39660 = n8069 | n39659 ;
  assign n39661 = ( n23960 & n34551 ) | ( n23960 & ~n39660 ) | ( n34551 & ~n39660 ) ;
  assign n39662 = n10835 & ~n19207 ;
  assign n39663 = ~n1075 & n39662 ;
  assign n39664 = n39663 ^ n23985 ^ n13594 ;
  assign n39665 = n39664 ^ n15675 ^ 1'b0 ;
  assign n39667 = n10017 ^ x50 ^ 1'b0 ;
  assign n39666 = ~n5298 & n6878 ;
  assign n39668 = n39667 ^ n39666 ^ 1'b0 ;
  assign n39669 = n14021 & n14309 ;
  assign n39670 = ~n26060 & n26960 ;
  assign n39671 = ~n23401 & n39670 ;
  assign n39672 = n3063 & n15169 ;
  assign n39673 = n39672 ^ n27386 ^ n11411 ;
  assign n39674 = ~n2960 & n25872 ;
  assign n39675 = n32253 ^ n25295 ^ 1'b0 ;
  assign n39676 = n25624 ^ n5021 ^ n3964 ;
  assign n39677 = n8155 & n39676 ;
  assign n39678 = ~n9997 & n16084 ;
  assign n39679 = n28452 & n39678 ;
  assign n39680 = n2143 & n6474 ;
  assign n39681 = n39680 ^ n764 ^ 1'b0 ;
  assign n39682 = n39681 ^ n22398 ^ 1'b0 ;
  assign n39683 = ~n5325 & n39682 ;
  assign n39684 = n39683 ^ n7473 ^ 1'b0 ;
  assign n39685 = n10353 | n39684 ;
  assign n39687 = ( n7735 & n9583 ) | ( n7735 & n11459 ) | ( n9583 & n11459 ) ;
  assign n39686 = n9978 | n24664 ;
  assign n39688 = n39687 ^ n39686 ^ 1'b0 ;
  assign n39689 = n39688 ^ n29669 ^ n5080 ;
  assign n39692 = n13920 ^ n2354 ^ 1'b0 ;
  assign n39690 = ( n1433 & n19533 ) | ( n1433 & ~n34199 ) | ( n19533 & ~n34199 ) ;
  assign n39691 = ~n37474 & n39690 ;
  assign n39693 = n39692 ^ n39691 ^ 1'b0 ;
  assign n39694 = n34362 ^ n19485 ^ 1'b0 ;
  assign n39695 = n9851 & ~n11961 ;
  assign n39696 = n13681 | n20051 ;
  assign n39697 = n39696 ^ n28103 ^ 1'b0 ;
  assign n39698 = ~n4476 & n15309 ;
  assign n39699 = n39698 ^ n12970 ^ 1'b0 ;
  assign n39700 = n27350 ^ n23115 ^ 1'b0 ;
  assign n39701 = n39699 & ~n39700 ;
  assign n39702 = n10945 | n21571 ;
  assign n39703 = n4708 & ~n30138 ;
  assign n39704 = n39703 ^ n30602 ^ n8688 ;
  assign n39708 = n10786 ^ n2887 ^ 1'b0 ;
  assign n39706 = ( ~n3712 & n7647 ) | ( ~n3712 & n8739 ) | ( n7647 & n8739 ) ;
  assign n39705 = ( n2907 & n26984 ) | ( n2907 & ~n36569 ) | ( n26984 & ~n36569 ) ;
  assign n39707 = n39706 ^ n39705 ^ n18161 ;
  assign n39709 = n39708 ^ n39707 ^ n36097 ;
  assign n39710 = n39709 ^ n25204 ^ n17438 ;
  assign n39711 = n30653 ^ n9651 ^ 1'b0 ;
  assign n39712 = n866 & ~n39711 ;
  assign n39713 = n39712 ^ n19157 ^ n15585 ;
  assign n39714 = ( n617 & n3556 ) | ( n617 & ~n39713 ) | ( n3556 & ~n39713 ) ;
  assign n39715 = n12837 ^ n12812 ^ 1'b0 ;
  assign n39716 = n9309 & ~n39715 ;
  assign n39717 = n36451 & n39716 ;
  assign n39721 = n15251 ^ n14296 ^ n10403 ;
  assign n39722 = n39721 ^ n37943 ^ 1'b0 ;
  assign n39718 = ~n3043 & n21520 ;
  assign n39719 = n39718 ^ n12362 ^ 1'b0 ;
  assign n39720 = ~n24523 & n39719 ;
  assign n39723 = n39722 ^ n39720 ^ 1'b0 ;
  assign n39724 = n39723 ^ n12439 ^ 1'b0 ;
  assign n39725 = ~n39717 & n39724 ;
  assign n39731 = ( n5329 & n14812 ) | ( n5329 & n19105 ) | ( n14812 & n19105 ) ;
  assign n39726 = n2380 & n16412 ;
  assign n39727 = n39726 ^ n1672 ^ 1'b0 ;
  assign n39728 = n17708 ^ n14832 ^ n4725 ;
  assign n39729 = n39727 | n39728 ;
  assign n39730 = n31030 | n39729 ;
  assign n39732 = n39731 ^ n39730 ^ 1'b0 ;
  assign n39733 = n4648 ^ n414 ^ 1'b0 ;
  assign n39734 = ( ~n2749 & n4632 ) | ( ~n2749 & n39733 ) | ( n4632 & n39733 ) ;
  assign n39735 = ( n9161 & ~n10532 ) | ( n9161 & n23704 ) | ( ~n10532 & n23704 ) ;
  assign n39737 = n39406 ^ n32678 ^ n19665 ;
  assign n39736 = n32053 ^ n14790 ^ 1'b0 ;
  assign n39738 = n39737 ^ n39736 ^ n30571 ;
  assign n39739 = ~n6528 & n15404 ;
  assign n39740 = n25921 & n39739 ;
  assign n39741 = n29627 | n39740 ;
  assign n39742 = n27916 | n30975 ;
  assign n39743 = n25848 | n39742 ;
  assign n39744 = n39743 ^ n34974 ^ 1'b0 ;
  assign n39745 = ~n13092 & n35496 ;
  assign n39746 = n8735 ^ n4991 ^ 1'b0 ;
  assign n39747 = ~n11794 & n16674 ;
  assign n39748 = n39747 ^ n32637 ^ n22398 ;
  assign n39749 = n15410 & n38039 ;
  assign n39750 = ( n3301 & n11166 ) | ( n3301 & n16722 ) | ( n11166 & n16722 ) ;
  assign n39751 = ~n7321 & n39750 ;
  assign n39752 = n39751 ^ n16855 ^ 1'b0 ;
  assign n39755 = n32613 ^ n25032 ^ n21183 ;
  assign n39753 = n25401 ^ n14380 ^ 1'b0 ;
  assign n39754 = n28709 | n39753 ;
  assign n39756 = n39755 ^ n39754 ^ 1'b0 ;
  assign n39757 = n7156 & n39756 ;
  assign n39758 = n39757 ^ n20383 ^ 1'b0 ;
  assign n39759 = n36892 ^ n29758 ^ 1'b0 ;
  assign n39760 = n39322 ^ n9091 ^ n699 ;
  assign n39763 = x3 & ~n20627 ;
  assign n39764 = n39763 ^ n21729 ^ 1'b0 ;
  assign n39761 = ( n989 & ~n5882 ) | ( n989 & n23575 ) | ( ~n5882 & n23575 ) ;
  assign n39762 = ~n27089 & n39761 ;
  assign n39765 = n39764 ^ n39762 ^ n14701 ;
  assign n39766 = ( ~n31099 & n34382 ) | ( ~n31099 & n38439 ) | ( n34382 & n38439 ) ;
  assign n39767 = n25576 ^ n12373 ^ 1'b0 ;
  assign n39768 = n39767 ^ n9884 ^ 1'b0 ;
  assign n39769 = n39768 ^ n29734 ^ n23181 ;
  assign n39770 = n39769 ^ n14614 ^ 1'b0 ;
  assign n39771 = x93 & n21435 ;
  assign n39772 = n39771 ^ n2884 ^ 1'b0 ;
  assign n39773 = n7446 & ~n39772 ;
  assign n39774 = n12924 ^ n9492 ^ 1'b0 ;
  assign n39775 = n39773 | n39774 ;
  assign n39776 = ( n2460 & n9268 ) | ( n2460 & ~n22390 ) | ( n9268 & ~n22390 ) ;
  assign n39777 = ( ~n38960 & n39775 ) | ( ~n38960 & n39776 ) | ( n39775 & n39776 ) ;
  assign n39778 = n35407 ^ n4325 ^ 1'b0 ;
  assign n39779 = x83 & ~n39778 ;
  assign n39780 = n14425 ^ n9786 ^ n7761 ;
  assign n39781 = n1605 & ~n10225 ;
  assign n39782 = n39780 & n39781 ;
  assign n39783 = n2747 & n9100 ;
  assign n39784 = n7731 & n39783 ;
  assign n39785 = n39784 ^ n21231 ^ 1'b0 ;
  assign n39786 = n12993 & ~n26703 ;
  assign n39787 = n39786 ^ n684 ^ 1'b0 ;
  assign n39788 = ~n17301 & n39787 ;
  assign n39789 = n39788 ^ n1398 ^ 1'b0 ;
  assign n39790 = n39789 ^ n29533 ^ n17571 ;
  assign n39791 = n15832 & n27485 ;
  assign n39792 = n9554 & n39791 ;
  assign n39793 = n39792 ^ n30632 ^ n14769 ;
  assign n39794 = ( n6955 & n7167 ) | ( n6955 & n34364 ) | ( n7167 & n34364 ) ;
  assign n39795 = ( n17293 & n23230 ) | ( n17293 & ~n24284 ) | ( n23230 & ~n24284 ) ;
  assign n39796 = n38342 ^ n7881 ^ n838 ;
  assign n39797 = n10159 ^ n8217 ^ n1347 ;
  assign n39798 = n39797 ^ n10838 ^ 1'b0 ;
  assign n39799 = n35343 ^ n9495 ^ 1'b0 ;
  assign n39800 = n13388 & ~n39799 ;
  assign n39801 = n30086 ^ n28325 ^ 1'b0 ;
  assign n39802 = n22517 & n35931 ;
  assign n39803 = n39802 ^ n24377 ^ n7414 ;
  assign n39804 = n16901 & n19190 ;
  assign n39805 = n39804 ^ n6281 ^ 1'b0 ;
  assign n39806 = n39805 ^ n39551 ^ 1'b0 ;
  assign n39809 = n26251 & ~n37665 ;
  assign n39810 = n13430 & n39809 ;
  assign n39807 = n29881 ^ n5109 ^ 1'b0 ;
  assign n39808 = n19303 & n39807 ;
  assign n39811 = n39810 ^ n39808 ^ n14452 ;
  assign n39812 = n36209 ^ n3774 ^ 1'b0 ;
  assign n39813 = n1725 | n5141 ;
  assign n39814 = n39813 ^ n16136 ^ 1'b0 ;
  assign n39815 = n1644 & n39814 ;
  assign n39816 = n39815 ^ n22455 ^ n4774 ;
  assign n39817 = n39816 ^ n14639 ^ 1'b0 ;
  assign n39818 = n19198 & n39817 ;
  assign n39819 = n30427 ^ n821 ^ 1'b0 ;
  assign n39820 = n682 & ~n19785 ;
  assign n39821 = n23669 ^ n8992 ^ 1'b0 ;
  assign n39822 = ~n34854 & n39821 ;
  assign n39823 = n11780 | n22325 ;
  assign n39824 = n39823 ^ n7217 ^ 1'b0 ;
  assign n39825 = n473 & n39824 ;
  assign n39826 = ( n23660 & n31446 ) | ( n23660 & n38032 ) | ( n31446 & n38032 ) ;
  assign n39827 = n39825 | n39826 ;
  assign n39829 = n13447 ^ n6960 ^ n5681 ;
  assign n39830 = ( n8472 & n22257 ) | ( n8472 & n39829 ) | ( n22257 & n39829 ) ;
  assign n39828 = n26927 ^ n1159 ^ 1'b0 ;
  assign n39831 = n39830 ^ n39828 ^ 1'b0 ;
  assign n39832 = n12779 | n20721 ;
  assign n39833 = n10072 ^ n450 ^ 1'b0 ;
  assign n39834 = ~n39832 & n39833 ;
  assign n39835 = n3785 ^ n3764 ^ 1'b0 ;
  assign n39836 = ( n7928 & n18823 ) | ( n7928 & n38086 ) | ( n18823 & n38086 ) ;
  assign n39837 = n17559 & ~n18844 ;
  assign n39838 = n4148 & ~n39837 ;
  assign n39839 = n39838 ^ n12734 ^ n1558 ;
  assign n39840 = ~n12110 & n39839 ;
  assign n39841 = ( n3459 & n39836 ) | ( n3459 & n39840 ) | ( n39836 & n39840 ) ;
  assign n39842 = n23630 ^ n11244 ^ n8892 ;
  assign n39844 = n28781 ^ n1552 ^ 1'b0 ;
  assign n39845 = ~n25139 & n39844 ;
  assign n39843 = n9997 | n12313 ;
  assign n39846 = n39845 ^ n39843 ^ 1'b0 ;
  assign n39847 = n13549 ^ n5480 ^ n528 ;
  assign n39848 = n39847 ^ n8281 ^ n1876 ;
  assign n39849 = n39848 ^ n24507 ^ 1'b0 ;
  assign n39850 = n2169 & ~n9894 ;
  assign n39851 = n25864 | n38469 ;
  assign n39852 = ( n15972 & n17379 ) | ( n15972 & n39434 ) | ( n17379 & n39434 ) ;
  assign n39853 = ~n9816 & n33705 ;
  assign n39854 = n19926 ^ n7020 ^ 1'b0 ;
  assign n39855 = n3548 | n28490 ;
  assign n39856 = n39855 ^ n15101 ^ 1'b0 ;
  assign n39857 = ( n13963 & n29557 ) | ( n13963 & n39719 ) | ( n29557 & n39719 ) ;
  assign n39858 = n26336 ^ n5011 ^ 1'b0 ;
  assign n39859 = n2749 & n39858 ;
  assign n39860 = ~n22651 & n39859 ;
  assign n39861 = n16398 & n32907 ;
  assign n39862 = n19660 & n39861 ;
  assign n39863 = n10087 | n19653 ;
  assign n39864 = n39863 ^ n13924 ^ 1'b0 ;
  assign n39865 = ( n19027 & n28256 ) | ( n19027 & n39864 ) | ( n28256 & n39864 ) ;
  assign n39866 = n39865 ^ n32377 ^ 1'b0 ;
  assign n39867 = n34178 ^ n17534 ^ 1'b0 ;
  assign n39868 = n31524 ^ n28890 ^ n25032 ;
  assign n39869 = ( ~n5779 & n18360 ) | ( ~n5779 & n31533 ) | ( n18360 & n31533 ) ;
  assign n39870 = n20118 ^ n8411 ^ 1'b0 ;
  assign n39871 = x166 & n29334 ;
  assign n39872 = n4119 & n19034 ;
  assign n39873 = n39872 ^ n20046 ^ 1'b0 ;
  assign n39874 = n14585 | n39873 ;
  assign n39875 = x240 & n17137 ;
  assign n39876 = n32662 ^ n17607 ^ n5545 ;
  assign n39877 = ( n30941 & n39875 ) | ( n30941 & ~n39876 ) | ( n39875 & ~n39876 ) ;
  assign n39878 = n23281 | n35267 ;
  assign n39879 = n19244 ^ n11637 ^ 1'b0 ;
  assign n39880 = n7163 & ~n37025 ;
  assign n39881 = ~n10480 & n39880 ;
  assign n39893 = n14245 ^ n1558 ^ 1'b0 ;
  assign n39890 = n8785 & ~n32627 ;
  assign n39888 = x213 & n28618 ;
  assign n39889 = ~n10725 & n39888 ;
  assign n39891 = n39890 ^ n39889 ^ n6334 ;
  assign n39892 = n39891 ^ n14607 ^ n13757 ;
  assign n39894 = n39893 ^ n39892 ^ n2055 ;
  assign n39882 = n18354 ^ n15407 ^ n11641 ;
  assign n39883 = ( ~n600 & n11892 ) | ( ~n600 & n39882 ) | ( n11892 & n39882 ) ;
  assign n39884 = n39883 ^ n21577 ^ n16029 ;
  assign n39885 = n39884 ^ n37607 ^ 1'b0 ;
  assign n39886 = ~n10656 & n39885 ;
  assign n39887 = ~n4237 & n39886 ;
  assign n39895 = n39894 ^ n39887 ^ 1'b0 ;
  assign n39896 = n33855 ^ n4958 ^ 1'b0 ;
  assign n39897 = n39895 & n39896 ;
  assign n39898 = n10529 | n20372 ;
  assign n39899 = ( ~n1938 & n10195 ) | ( ~n1938 & n20911 ) | ( n10195 & n20911 ) ;
  assign n39900 = n4028 ^ n3126 ^ 1'b0 ;
  assign n39901 = n21890 | n39900 ;
  assign n39902 = ( n23184 & ~n30002 ) | ( n23184 & n39901 ) | ( ~n30002 & n39901 ) ;
  assign n39903 = ( n7050 & n8986 ) | ( n7050 & ~n14958 ) | ( n8986 & ~n14958 ) ;
  assign n39904 = n2466 & n4816 ;
  assign n39905 = n39904 ^ n24959 ^ n7968 ;
  assign n39906 = n39905 ^ n10442 ^ 1'b0 ;
  assign n39907 = ~n14594 & n39906 ;
  assign n39908 = ~n13527 & n39907 ;
  assign n39909 = n14226 & n29429 ;
  assign n39910 = ~n11795 & n39909 ;
  assign n39911 = ~n7061 & n15134 ;
  assign n39912 = n15722 ^ n1660 ^ 1'b0 ;
  assign n39913 = ( n796 & ~n28536 ) | ( n796 & n31571 ) | ( ~n28536 & n31571 ) ;
  assign n39914 = n25139 ^ n5863 ^ n4811 ;
  assign n39915 = n39914 ^ n19075 ^ n16161 ;
  assign n39917 = ( n5461 & ~n25127 ) | ( n5461 & n26302 ) | ( ~n25127 & n26302 ) ;
  assign n39916 = n18257 & ~n38368 ;
  assign n39918 = n39917 ^ n39916 ^ 1'b0 ;
  assign n39923 = ~n2655 & n7820 ;
  assign n39924 = ( ~n7539 & n13480 ) | ( ~n7539 & n39923 ) | ( n13480 & n39923 ) ;
  assign n39921 = n13828 ^ n5652 ^ n1323 ;
  assign n39919 = n2465 & ~n16566 ;
  assign n39920 = n39919 ^ n12484 ^ 1'b0 ;
  assign n39922 = n39921 ^ n39920 ^ n8628 ;
  assign n39925 = n39924 ^ n39922 ^ 1'b0 ;
  assign n39926 = n16401 & ~n34372 ;
  assign n39927 = n20818 ^ n12157 ^ n1251 ;
  assign n39928 = ( n3170 & n15484 ) | ( n3170 & ~n39927 ) | ( n15484 & ~n39927 ) ;
  assign n39929 = ( ~n1137 & n1290 ) | ( ~n1137 & n20276 ) | ( n1290 & n20276 ) ;
  assign n39930 = n39274 ^ n7342 ^ 1'b0 ;
  assign n39931 = n8229 & ~n39930 ;
  assign n39932 = ( n8813 & n39929 ) | ( n8813 & n39931 ) | ( n39929 & n39931 ) ;
  assign n39933 = n39932 ^ n17754 ^ n13296 ;
  assign n39934 = n33118 ^ n22855 ^ n9980 ;
  assign n39935 = ( n39928 & n39933 ) | ( n39928 & ~n39934 ) | ( n39933 & ~n39934 ) ;
  assign n39936 = ~n3528 & n18979 ;
  assign n39937 = n39936 ^ n16470 ^ 1'b0 ;
  assign n39938 = n20858 & n21754 ;
  assign n39939 = ( n6391 & n39937 ) | ( n6391 & n39938 ) | ( n39937 & n39938 ) ;
  assign n39941 = n5496 ^ n1328 ^ 1'b0 ;
  assign n39942 = n11157 & ~n39941 ;
  assign n39940 = n25948 & ~n30462 ;
  assign n39943 = n39942 ^ n39940 ^ 1'b0 ;
  assign n39944 = n19545 & ~n39943 ;
  assign n39945 = n26038 ^ n13552 ^ 1'b0 ;
  assign n39946 = n39944 & ~n39945 ;
  assign n39947 = ~n15734 & n26839 ;
  assign n39948 = ~n23448 & n39947 ;
  assign n39949 = n28937 ^ n14064 ^ n2395 ;
  assign n39950 = n39949 ^ n3138 ^ 1'b0 ;
  assign n39951 = ~n39948 & n39950 ;
  assign n39952 = n4257 & n8008 ;
  assign n39953 = n39952 ^ n21273 ^ 1'b0 ;
  assign n39954 = n39953 ^ n10170 ^ 1'b0 ;
  assign n39955 = n39954 ^ x119 ^ 1'b0 ;
  assign n39956 = n19540 | n39955 ;
  assign n39957 = n24564 | n39956 ;
  assign n39958 = n22227 ^ n12212 ^ 1'b0 ;
  assign n39959 = ~n15555 & n25648 ;
  assign n39960 = ~n11493 & n39959 ;
  assign n39961 = ~n6952 & n8533 ;
  assign n39962 = n39960 & n39961 ;
  assign n39965 = n26653 ^ n6949 ^ 1'b0 ;
  assign n39963 = ( n8325 & ~n29927 ) | ( n8325 & n36850 ) | ( ~n29927 & n36850 ) ;
  assign n39964 = ~n16026 & n39963 ;
  assign n39966 = n39965 ^ n39964 ^ 1'b0 ;
  assign n39967 = ( ~n30380 & n39962 ) | ( ~n30380 & n39966 ) | ( n39962 & n39966 ) ;
  assign n39974 = ( n15156 & n24690 ) | ( n15156 & n30350 ) | ( n24690 & n30350 ) ;
  assign n39968 = n6832 ^ n293 ^ 1'b0 ;
  assign n39969 = n11546 & n39968 ;
  assign n39970 = ~n6648 & n39969 ;
  assign n39971 = ~n7410 & n39970 ;
  assign n39972 = ( n971 & n31413 ) | ( n971 & ~n39971 ) | ( n31413 & ~n39971 ) ;
  assign n39973 = ~n13045 & n39972 ;
  assign n39975 = n39974 ^ n39973 ^ 1'b0 ;
  assign n39976 = n39975 ^ n32839 ^ n22921 ;
  assign n39978 = n13552 ^ n12907 ^ 1'b0 ;
  assign n39979 = n14389 | n39978 ;
  assign n39977 = ~n5583 & n6277 ;
  assign n39980 = n39979 ^ n39977 ^ n2861 ;
  assign n39981 = n37113 ^ n7735 ^ n5895 ;
  assign n39982 = n37579 ^ n34472 ^ 1'b0 ;
  assign n39983 = n5116 & n7428 ;
  assign n39984 = n39983 ^ n34988 ^ 1'b0 ;
  assign n39985 = n39984 ^ n19553 ^ 1'b0 ;
  assign n39986 = n8666 | n31770 ;
  assign n39987 = n21968 ^ n12323 ^ 1'b0 ;
  assign n39988 = ( n28152 & ~n32208 ) | ( n28152 & n36242 ) | ( ~n32208 & n36242 ) ;
  assign n39989 = n39987 | n39988 ;
  assign n39990 = n22744 ^ n16433 ^ 1'b0 ;
  assign n39991 = n3147 & n39990 ;
  assign n39992 = ( n2912 & ~n39989 ) | ( n2912 & n39991 ) | ( ~n39989 & n39991 ) ;
  assign n39993 = n37511 ^ n30219 ^ 1'b0 ;
  assign n39994 = n21698 & n39993 ;
  assign n39995 = n4139 & n7427 ;
  assign n39996 = n39995 ^ n3012 ^ 1'b0 ;
  assign n39997 = ~n24503 & n38473 ;
  assign n39998 = ~n39996 & n39997 ;
  assign n40002 = n23386 ^ n6220 ^ 1'b0 ;
  assign n40003 = ~n5585 & n40002 ;
  assign n40000 = n17700 & ~n24915 ;
  assign n40001 = n40000 ^ n34213 ^ n6615 ;
  assign n39999 = n8943 | n21893 ;
  assign n40004 = n40003 ^ n40001 ^ n39999 ;
  assign n40005 = n18710 ^ n10976 ^ n2960 ;
  assign n40006 = n40005 ^ n31837 ^ n6224 ;
  assign n40007 = ( n20053 & ~n25536 ) | ( n20053 & n30754 ) | ( ~n25536 & n30754 ) ;
  assign n40008 = n40007 ^ n16230 ^ 1'b0 ;
  assign n40009 = n5365 & n34975 ;
  assign n40010 = n40009 ^ n37054 ^ 1'b0 ;
  assign n40011 = n30133 ^ n6330 ^ 1'b0 ;
  assign n40012 = n32503 ^ n18259 ^ 1'b0 ;
  assign n40013 = n16049 ^ n11997 ^ 1'b0 ;
  assign n40014 = n27130 ^ n21457 ^ n11690 ;
  assign n40016 = x59 & ~n8286 ;
  assign n40017 = n40016 ^ n16277 ^ 1'b0 ;
  assign n40015 = n23544 & ~n38698 ;
  assign n40018 = n40017 ^ n40015 ^ 1'b0 ;
  assign n40019 = n40018 ^ n37339 ^ n35689 ;
  assign n40020 = n16699 & ~n37668 ;
  assign n40021 = n23749 ^ n13873 ^ 1'b0 ;
  assign n40022 = n21252 | n40021 ;
  assign n40023 = n2080 & ~n10027 ;
  assign n40024 = n40023 ^ n7217 ^ 1'b0 ;
  assign n40025 = n14585 | n15351 ;
  assign n40026 = n40024 & ~n40025 ;
  assign n40027 = n8263 | n32601 ;
  assign n40028 = n40026 & ~n40027 ;
  assign n40029 = ( ~n1406 & n16195 ) | ( ~n1406 & n23189 ) | ( n16195 & n23189 ) ;
  assign n40030 = n40029 ^ n32403 ^ n11925 ;
  assign n40031 = n40030 ^ n36781 ^ 1'b0 ;
  assign n40032 = n25906 ^ n9107 ^ 1'b0 ;
  assign n40033 = ~n15389 & n40032 ;
  assign n40034 = n21980 ^ n9137 ^ 1'b0 ;
  assign n40035 = n40034 ^ n25270 ^ n23561 ;
  assign n40036 = ( ~n9890 & n14464 ) | ( ~n9890 & n40035 ) | ( n14464 & n40035 ) ;
  assign n40037 = ( ~n4091 & n9556 ) | ( ~n4091 & n30112 ) | ( n9556 & n30112 ) ;
  assign n40038 = n40037 ^ n31083 ^ n30270 ;
  assign n40039 = n13828 ^ n4104 ^ 1'b0 ;
  assign n40042 = n2322 | n8564 ;
  assign n40040 = n19238 | n28879 ;
  assign n40041 = n40040 ^ n37831 ^ 1'b0 ;
  assign n40043 = n40042 ^ n40041 ^ 1'b0 ;
  assign n40044 = n40039 & n40043 ;
  assign n40045 = n19777 ^ n3513 ^ 1'b0 ;
  assign n40046 = n32415 ^ n22415 ^ n17129 ;
  assign n40047 = ~n9481 & n11272 ;
  assign n40048 = n40047 ^ n13457 ^ 1'b0 ;
  assign n40049 = n5579 | n40048 ;
  assign n40050 = n16738 & ~n40049 ;
  assign n40051 = n15821 ^ n1868 ^ 1'b0 ;
  assign n40052 = ~n10865 & n40051 ;
  assign n40053 = ~n11130 & n40052 ;
  assign n40054 = n40053 ^ n2218 ^ 1'b0 ;
  assign n40055 = n6468 ^ n1385 ^ 1'b0 ;
  assign n40056 = ( ~n9827 & n14492 ) | ( ~n9827 & n40055 ) | ( n14492 & n40055 ) ;
  assign n40057 = ~n13231 & n13535 ;
  assign n40058 = n2719 & n40057 ;
  assign n40059 = n3286 & ~n40058 ;
  assign n40060 = n40059 ^ n17541 ^ 1'b0 ;
  assign n40061 = n16526 ^ n5334 ^ 1'b0 ;
  assign n40062 = n40061 ^ n5493 ^ n1985 ;
  assign n40065 = n14646 ^ n13137 ^ n10461 ;
  assign n40063 = n18348 & ~n39617 ;
  assign n40064 = n40063 ^ n21505 ^ n15701 ;
  assign n40066 = n40065 ^ n40064 ^ 1'b0 ;
  assign n40067 = ( n11242 & n22095 ) | ( n11242 & n26761 ) | ( n22095 & n26761 ) ;
  assign n40068 = n8341 | n40067 ;
  assign n40069 = n9141 & ~n40068 ;
  assign n40070 = n25205 ^ n10630 ^ n7808 ;
  assign n40071 = n19049 ^ n2663 ^ 1'b0 ;
  assign n40072 = n40070 | n40071 ;
  assign n40073 = n29290 ^ n19923 ^ 1'b0 ;
  assign n40074 = n21154 | n38773 ;
  assign n40075 = n40073 | n40074 ;
  assign n40076 = n29029 ^ n20751 ^ n5687 ;
  assign n40077 = n32779 & ~n40076 ;
  assign n40078 = n22871 ^ n9399 ^ n774 ;
  assign n40079 = n40078 ^ n10793 ^ n5228 ;
  assign n40080 = n30626 ^ n14199 ^ 1'b0 ;
  assign n40081 = ~n10684 & n40080 ;
  assign n40082 = n483 & n8251 ;
  assign n40083 = n40082 ^ n34327 ^ n400 ;
  assign n40084 = n17033 | n29773 ;
  assign n40085 = n40084 ^ n14985 ^ n14513 ;
  assign n40086 = n4524 & ~n6626 ;
  assign n40087 = ~n3873 & n40086 ;
  assign n40088 = n40087 ^ n36804 ^ 1'b0 ;
  assign n40089 = n4401 & ~n5151 ;
  assign n40090 = ( ~n7888 & n12369 ) | ( ~n7888 & n16594 ) | ( n12369 & n16594 ) ;
  assign n40091 = n10282 & n40090 ;
  assign n40092 = n14134 ^ n8186 ^ 1'b0 ;
  assign n40093 = n38954 & n40092 ;
  assign n40094 = n26795 ^ n22216 ^ 1'b0 ;
  assign n40095 = n27780 & ~n38581 ;
  assign n40096 = n6928 | n40095 ;
  assign n40097 = n27565 ^ n409 ^ 1'b0 ;
  assign n40098 = ( ~n3844 & n7060 ) | ( ~n3844 & n40097 ) | ( n7060 & n40097 ) ;
  assign n40099 = n2274 & n32680 ;
  assign n40100 = ~n20897 & n40099 ;
  assign n40101 = ( n13579 & ~n40098 ) | ( n13579 & n40100 ) | ( ~n40098 & n40100 ) ;
  assign n40102 = n23574 ^ n13818 ^ 1'b0 ;
  assign n40103 = ( ~n733 & n2179 ) | ( ~n733 & n40102 ) | ( n2179 & n40102 ) ;
  assign n40104 = n15320 & n19318 ;
  assign n40105 = ~n8313 & n40104 ;
  assign n40106 = ( ~n3346 & n12442 ) | ( ~n3346 & n14199 ) | ( n12442 & n14199 ) ;
  assign n40107 = ( n16117 & n38915 ) | ( n16117 & ~n40106 ) | ( n38915 & ~n40106 ) ;
  assign n40108 = ~n7465 & n10773 ;
  assign n40109 = ~n40107 & n40108 ;
  assign n40110 = n16857 & ~n40109 ;
  assign n40111 = n40110 ^ n38316 ^ 1'b0 ;
  assign n40112 = n35213 ^ n6249 ^ 1'b0 ;
  assign n40113 = n2255 | n40112 ;
  assign n40114 = n22753 ^ n4300 ^ n2680 ;
  assign n40115 = n9217 ^ n3802 ^ 1'b0 ;
  assign n40116 = n40115 ^ n28738 ^ n6149 ;
  assign n40117 = n34589 ^ n30160 ^ n13694 ;
  assign n40118 = n17412 ^ n10088 ^ 1'b0 ;
  assign n40119 = ~n9288 & n40118 ;
  assign n40120 = n40119 ^ n13801 ^ 1'b0 ;
  assign n40121 = ~n35256 & n40120 ;
  assign n40122 = n4999 & ~n26944 ;
  assign n40123 = n32267 ^ n8856 ^ 1'b0 ;
  assign n40124 = n14564 & n40123 ;
  assign n40125 = n40124 ^ n1001 ^ 1'b0 ;
  assign n40126 = n18244 & ~n40125 ;
  assign n40127 = ~n12616 & n18032 ;
  assign n40128 = n977 & n40127 ;
  assign n40129 = n40128 ^ n20098 ^ n10767 ;
  assign n40131 = ( n1873 & n2987 ) | ( n1873 & n39883 ) | ( n2987 & n39883 ) ;
  assign n40130 = ~n483 & n12424 ;
  assign n40132 = n40131 ^ n40130 ^ 1'b0 ;
  assign n40134 = n23332 | n30107 ;
  assign n40133 = n13940 | n31642 ;
  assign n40135 = n40134 ^ n40133 ^ 1'b0 ;
  assign n40136 = n1173 & n39315 ;
  assign n40137 = ~n5607 & n40136 ;
  assign n40138 = ( n6624 & n14474 ) | ( n6624 & ~n30784 ) | ( n14474 & ~n30784 ) ;
  assign n40139 = n40138 ^ n11420 ^ n2370 ;
  assign n40140 = n14251 ^ n10920 ^ 1'b0 ;
  assign n40141 = n18318 & n40140 ;
  assign n40142 = n40141 ^ n16607 ^ 1'b0 ;
  assign n40143 = ~n40139 & n40142 ;
  assign n40144 = ( x116 & n15413 ) | ( x116 & n27119 ) | ( n15413 & n27119 ) ;
  assign n40145 = n20533 ^ n14785 ^ 1'b0 ;
  assign n40146 = x43 & ~n40145 ;
  assign n40147 = n40146 ^ n21943 ^ n5353 ;
  assign n40148 = ( n7342 & n27600 ) | ( n7342 & ~n40147 ) | ( n27600 & ~n40147 ) ;
  assign n40149 = n11084 & n28775 ;
  assign n40150 = n3670 & ~n40149 ;
  assign n40151 = n23254 & n40150 ;
  assign n40152 = n9341 & ~n17242 ;
  assign n40153 = n24712 & n40152 ;
  assign n40154 = n4257 & ~n6211 ;
  assign n40155 = n40154 ^ n12986 ^ 1'b0 ;
  assign n40156 = n33569 ^ n32272 ^ n9122 ;
  assign n40157 = n2287 & ~n12101 ;
  assign n40158 = ( n21835 & n40156 ) | ( n21835 & ~n40157 ) | ( n40156 & ~n40157 ) ;
  assign n40159 = n40158 ^ n14262 ^ 1'b0 ;
  assign n40160 = n13992 | n40159 ;
  assign n40161 = n10113 & n34712 ;
  assign n40162 = n40161 ^ n28594 ^ 1'b0 ;
  assign n40163 = ( ~n21743 & n30153 ) | ( ~n21743 & n36970 ) | ( n30153 & n36970 ) ;
  assign n40164 = n38200 ^ n13616 ^ n5002 ;
  assign n40165 = n11384 & n40164 ;
  assign n40166 = ~n27877 & n40165 ;
  assign n40167 = n7800 & n12493 ;
  assign n40168 = n4600 & n40167 ;
  assign n40169 = ( ~n1801 & n40166 ) | ( ~n1801 & n40168 ) | ( n40166 & n40168 ) ;
  assign n40170 = n28727 ^ n16164 ^ n8953 ;
  assign n40171 = n14506 ^ n11532 ^ n9387 ;
  assign n40172 = n40171 ^ n17070 ^ 1'b0 ;
  assign n40173 = ( n5989 & ~n40170 ) | ( n5989 & n40172 ) | ( ~n40170 & n40172 ) ;
  assign n40174 = n30643 ^ n20214 ^ 1'b0 ;
  assign n40175 = n40173 | n40174 ;
  assign n40176 = ( n3555 & n6589 ) | ( n3555 & ~n13310 ) | ( n6589 & ~n13310 ) ;
  assign n40177 = n40176 ^ n28165 ^ n19553 ;
  assign n40178 = n3208 | n25469 ;
  assign n40179 = ~n13553 & n31496 ;
  assign n40180 = n10477 | n33874 ;
  assign n40181 = n26802 | n40180 ;
  assign n40182 = ( n17220 & n32714 ) | ( n17220 & ~n40181 ) | ( n32714 & ~n40181 ) ;
  assign n40183 = n40179 & n40182 ;
  assign n40184 = n11335 ^ n6994 ^ 1'b0 ;
  assign n40185 = n40184 ^ n27703 ^ 1'b0 ;
  assign n40188 = n20706 & n21314 ;
  assign n40189 = n40188 ^ n11718 ^ 1'b0 ;
  assign n40186 = n20575 ^ n14728 ^ 1'b0 ;
  assign n40187 = n39240 & n40186 ;
  assign n40190 = n40189 ^ n40187 ^ n6973 ;
  assign n40191 = n18281 ^ n16683 ^ 1'b0 ;
  assign n40192 = n5130 | n40191 ;
  assign n40196 = n15217 ^ n3041 ^ n2463 ;
  assign n40194 = ( n2774 & n9084 ) | ( n2774 & n9380 ) | ( n9084 & n9380 ) ;
  assign n40193 = n14406 & n31365 ;
  assign n40195 = n40194 ^ n40193 ^ 1'b0 ;
  assign n40197 = n40196 ^ n40195 ^ n15283 ;
  assign n40198 = ( ~n19892 & n40192 ) | ( ~n19892 & n40197 ) | ( n40192 & n40197 ) ;
  assign n40199 = ( n11122 & ~n15658 ) | ( n11122 & n30135 ) | ( ~n15658 & n30135 ) ;
  assign n40200 = n25652 ^ n21971 ^ 1'b0 ;
  assign n40201 = ~n2151 & n40200 ;
  assign n40202 = ~n6364 & n40201 ;
  assign n40203 = n33734 ^ n3196 ^ 1'b0 ;
  assign n40204 = ~n33047 & n40203 ;
  assign n40205 = ( ~n6990 & n40202 ) | ( ~n6990 & n40204 ) | ( n40202 & n40204 ) ;
  assign n40206 = n40205 ^ n20831 ^ 1'b0 ;
  assign n40207 = n8702 & n24943 ;
  assign n40208 = n20352 & n40207 ;
  assign n40209 = n33468 ^ n30229 ^ n4304 ;
  assign n40210 = n4276 ^ n3129 ^ 1'b0 ;
  assign n40211 = n40209 | n40210 ;
  assign n40212 = n36763 | n40211 ;
  assign n40213 = n20055 ^ n18509 ^ 1'b0 ;
  assign n40214 = ~n9951 & n40213 ;
  assign n40215 = n4093 ^ n3337 ^ n2574 ;
  assign n40216 = n1652 | n12798 ;
  assign n40217 = n40216 ^ n5367 ^ n804 ;
  assign n40218 = n39703 ^ n22621 ^ 1'b0 ;
  assign n40219 = ~n4319 & n30941 ;
  assign n40220 = ~n17434 & n40219 ;
  assign n40221 = n40220 ^ n18247 ^ 1'b0 ;
  assign n40224 = n3362 ^ n261 ^ 1'b0 ;
  assign n40225 = n40224 ^ n4239 ^ 1'b0 ;
  assign n40222 = n12086 ^ n7308 ^ 1'b0 ;
  assign n40223 = n9859 & ~n40222 ;
  assign n40226 = n40225 ^ n40223 ^ 1'b0 ;
  assign n40227 = n19960 ^ n2519 ^ 1'b0 ;
  assign n40228 = n40227 ^ n29365 ^ n2966 ;
  assign n40229 = n13030 & ~n16180 ;
  assign n40230 = n40229 ^ n23427 ^ 1'b0 ;
  assign n40231 = n40230 ^ n8839 ^ n6194 ;
  assign n40232 = ( n5973 & ~n6782 ) | ( n5973 & n23111 ) | ( ~n6782 & n23111 ) ;
  assign n40233 = n8850 | n26535 ;
  assign n40234 = n40233 ^ n10563 ^ 1'b0 ;
  assign n40235 = n27137 | n38747 ;
  assign n40236 = n37414 & ~n40235 ;
  assign n40237 = n20372 ^ n18838 ^ 1'b0 ;
  assign n40238 = n40237 ^ n7522 ^ 1'b0 ;
  assign n40239 = ~n40236 & n40238 ;
  assign n40240 = ( n40232 & ~n40234 ) | ( n40232 & n40239 ) | ( ~n40234 & n40239 ) ;
  assign n40241 = n40240 ^ n28182 ^ n12125 ;
  assign n40242 = n40241 ^ n23243 ^ 1'b0 ;
  assign n40243 = n3824 ^ n3330 ^ 1'b0 ;
  assign n40244 = ( n10820 & n24979 ) | ( n10820 & ~n40243 ) | ( n24979 & ~n40243 ) ;
  assign n40245 = n27162 ^ n11212 ^ n8176 ;
  assign n40246 = ~n3496 & n17718 ;
  assign n40247 = ~n9726 & n40246 ;
  assign n40248 = n40247 ^ n3384 ^ 1'b0 ;
  assign n40249 = n18796 & ~n26139 ;
  assign n40250 = ~n13894 & n40249 ;
  assign n40251 = n10561 ^ n9096 ^ 1'b0 ;
  assign n40252 = n26488 ^ n15572 ^ 1'b0 ;
  assign n40253 = n35133 ^ n9851 ^ 1'b0 ;
  assign n40254 = n15276 & ~n40253 ;
  assign n40255 = ~n40252 & n40254 ;
  assign n40256 = n6019 ^ n1113 ^ 1'b0 ;
  assign n40257 = ~n4710 & n12883 ;
  assign n40258 = n40256 & n40257 ;
  assign n40259 = n40258 ^ n26990 ^ n10248 ;
  assign n40260 = n1314 & n13439 ;
  assign n40261 = ( n9945 & n34817 ) | ( n9945 & ~n40260 ) | ( n34817 & ~n40260 ) ;
  assign n40262 = n29573 ^ n5126 ^ 1'b0 ;
  assign n40263 = ~n28914 & n40262 ;
  assign n40264 = ( n6871 & n23010 ) | ( n6871 & n40263 ) | ( n23010 & n40263 ) ;
  assign n40265 = n19726 & n22168 ;
  assign n40266 = n40265 ^ n3931 ^ 1'b0 ;
  assign n40267 = n9189 ^ x171 ^ 1'b0 ;
  assign n40268 = n37779 | n40267 ;
  assign n40269 = n15434 & ~n40268 ;
  assign n40270 = ( n5444 & ~n7440 ) | ( n5444 & n37144 ) | ( ~n7440 & n37144 ) ;
  assign n40271 = ~n12242 & n19799 ;
  assign n40272 = n17225 & n40271 ;
  assign n40273 = ( n12897 & n40270 ) | ( n12897 & ~n40272 ) | ( n40270 & ~n40272 ) ;
  assign n40274 = ~n9065 & n21583 ;
  assign n40275 = ~n7122 & n40274 ;
  assign n40276 = n40275 ^ n15868 ^ 1'b0 ;
  assign n40277 = n40276 ^ n10860 ^ 1'b0 ;
  assign n40278 = ( ~n11140 & n13408 ) | ( ~n11140 & n29809 ) | ( n13408 & n29809 ) ;
  assign n40279 = n23782 | n40278 ;
  assign n40280 = ( n7158 & n14189 ) | ( n7158 & ~n20183 ) | ( n14189 & ~n20183 ) ;
  assign n40281 = ( n9542 & ~n31220 ) | ( n9542 & n40280 ) | ( ~n31220 & n40280 ) ;
  assign n40282 = n40281 ^ n26363 ^ n17489 ;
  assign n40283 = ( n27373 & ~n28643 ) | ( n27373 & n40282 ) | ( ~n28643 & n40282 ) ;
  assign n40284 = n23209 | n40138 ;
  assign n40285 = n14634 ^ n11837 ^ n1266 ;
  assign n40286 = ( n33125 & n37255 ) | ( n33125 & ~n40285 ) | ( n37255 & ~n40285 ) ;
  assign n40287 = n14201 ^ n13569 ^ 1'b0 ;
  assign n40288 = ( n40284 & n40286 ) | ( n40284 & n40287 ) | ( n40286 & n40287 ) ;
  assign n40289 = n3924 & n22033 ;
  assign n40290 = n40288 & n40289 ;
  assign n40291 = n29527 ^ n21346 ^ 1'b0 ;
  assign n40292 = ~n3946 & n8241 ;
  assign n40293 = n8779 & ~n18663 ;
  assign n40294 = n40293 ^ n15737 ^ 1'b0 ;
  assign n40295 = n15562 & n40294 ;
  assign n40296 = ~n40292 & n40295 ;
  assign n40297 = n13341 ^ n3330 ^ 1'b0 ;
  assign n40298 = n35290 & n40297 ;
  assign n40299 = n28704 ^ n7260 ^ 1'b0 ;
  assign n40300 = n40298 & n40299 ;
  assign n40307 = n6725 & n32453 ;
  assign n40308 = ~n12905 & n40307 ;
  assign n40301 = n23946 | n40267 ;
  assign n40302 = n13204 & ~n40301 ;
  assign n40303 = x142 & ~n10647 ;
  assign n40304 = n40303 ^ n23703 ^ 1'b0 ;
  assign n40305 = n40304 ^ n29211 ^ 1'b0 ;
  assign n40306 = ~n40302 & n40305 ;
  assign n40309 = n40308 ^ n40306 ^ 1'b0 ;
  assign n40310 = n40300 & ~n40309 ;
  assign n40311 = n13794 & ~n25120 ;
  assign n40312 = ( ~n7446 & n16640 ) | ( ~n7446 & n16964 ) | ( n16640 & n16964 ) ;
  assign n40313 = ~n21352 & n26266 ;
  assign n40314 = n40313 ^ n30265 ^ 1'b0 ;
  assign n40315 = ( n2899 & ~n40312 ) | ( n2899 & n40314 ) | ( ~n40312 & n40314 ) ;
  assign n40317 = n31180 ^ n9309 ^ n8802 ;
  assign n40318 = n5809 & ~n40317 ;
  assign n40319 = n4267 & n40318 ;
  assign n40320 = n40319 ^ n23973 ^ 1'b0 ;
  assign n40321 = ~n21105 & n40320 ;
  assign n40316 = n1222 | n22452 ;
  assign n40322 = n40321 ^ n40316 ^ 1'b0 ;
  assign n40323 = n21265 & ~n40322 ;
  assign n40324 = n25378 ^ n22468 ^ n1743 ;
  assign n40325 = n7707 | n32632 ;
  assign n40326 = n34303 ^ n10532 ^ 1'b0 ;
  assign n40327 = ~n32486 & n40326 ;
  assign n40328 = n26680 ^ n16213 ^ 1'b0 ;
  assign n40329 = n12489 & n40328 ;
  assign n40330 = n18657 ^ n6697 ^ 1'b0 ;
  assign n40331 = n28678 | n40330 ;
  assign n40332 = n7391 & ~n40331 ;
  assign n40333 = ~n3411 & n40332 ;
  assign n40334 = n32242 ^ n26565 ^ 1'b0 ;
  assign n40335 = ( ~n13410 & n38743 ) | ( ~n13410 & n39775 ) | ( n38743 & n39775 ) ;
  assign n40336 = ( ~n40333 & n40334 ) | ( ~n40333 & n40335 ) | ( n40334 & n40335 ) ;
  assign n40337 = n9442 ^ n6963 ^ 1'b0 ;
  assign n40338 = n21761 ^ n16601 ^ n5688 ;
  assign n40339 = n15588 ^ n3138 ^ n687 ;
  assign n40340 = ( n3498 & n28129 ) | ( n3498 & ~n40339 ) | ( n28129 & ~n40339 ) ;
  assign n40341 = ( n12090 & n14210 ) | ( n12090 & ~n25129 ) | ( n14210 & ~n25129 ) ;
  assign n40342 = n40341 ^ n21423 ^ 1'b0 ;
  assign n40343 = ( n1359 & n16101 ) | ( n1359 & ~n17936 ) | ( n16101 & ~n17936 ) ;
  assign n40344 = ~n2896 & n15002 ;
  assign n40345 = ~n40343 & n40344 ;
  assign n40346 = n5494 & n23458 ;
  assign n40347 = n4835 ^ n756 ^ x7 ;
  assign n40348 = n40347 ^ n30217 ^ n13763 ;
  assign n40349 = n24933 & n34145 ;
  assign n40350 = n18287 & n40349 ;
  assign n40351 = n40350 ^ n18230 ^ 1'b0 ;
  assign n40352 = n19928 ^ n12422 ^ n12283 ;
  assign n40353 = ( n16924 & ~n39367 ) | ( n16924 & n40352 ) | ( ~n39367 & n40352 ) ;
  assign n40354 = n32312 ^ n30657 ^ n15309 ;
  assign n40355 = n39607 ^ n12692 ^ 1'b0 ;
  assign n40356 = n8969 & ~n39893 ;
  assign n40357 = n40356 ^ n15180 ^ 1'b0 ;
  assign n40358 = n19227 ^ n7294 ^ 1'b0 ;
  assign n40359 = ~n24789 & n40358 ;
  assign n40360 = n34094 ^ n29669 ^ 1'b0 ;
  assign n40361 = ( x218 & n7306 ) | ( x218 & ~n17481 ) | ( n7306 & ~n17481 ) ;
  assign n40362 = ~n26542 & n37483 ;
  assign n40363 = n23059 & n40362 ;
  assign n40364 = ( n9825 & n14690 ) | ( n9825 & ~n34867 ) | ( n14690 & ~n34867 ) ;
  assign n40365 = ( n40361 & ~n40363 ) | ( n40361 & n40364 ) | ( ~n40363 & n40364 ) ;
  assign n40366 = ( n5864 & n14370 ) | ( n5864 & n16667 ) | ( n14370 & n16667 ) ;
  assign n40367 = n40366 ^ n35393 ^ 1'b0 ;
  assign n40368 = ~n1324 & n29535 ;
  assign n40369 = n40368 ^ n8503 ^ 1'b0 ;
  assign n40370 = n7540 & n40369 ;
  assign n40371 = n21639 ^ n2515 ^ 1'b0 ;
  assign n40372 = ~n26883 & n40371 ;
  assign n40373 = n34586 ^ n7296 ^ 1'b0 ;
  assign n40374 = n40372 & n40373 ;
  assign n40375 = n3499 & n40139 ;
  assign n40376 = ~n8369 & n22813 ;
  assign n40377 = n40376 ^ n10329 ^ 1'b0 ;
  assign n40378 = n31032 & n40377 ;
  assign n40379 = ( ~n7038 & n14304 ) | ( ~n7038 & n24569 ) | ( n14304 & n24569 ) ;
  assign n40380 = n40379 ^ n14270 ^ 1'b0 ;
  assign n40381 = ~n29136 & n32714 ;
  assign n40382 = ~n5164 & n40381 ;
  assign n40383 = n15240 | n35280 ;
  assign n40384 = n11227 & ~n40383 ;
  assign n40385 = n40384 ^ n14561 ^ n12912 ;
  assign n40386 = n22353 ^ n15969 ^ 1'b0 ;
  assign n40387 = ~n40385 & n40386 ;
  assign n40388 = ( ~n1779 & n10111 ) | ( ~n1779 & n12437 ) | ( n10111 & n12437 ) ;
  assign n40389 = n31158 ^ n10248 ^ x202 ;
  assign n40390 = n17445 & n40389 ;
  assign n40391 = ( ~n14275 & n18332 ) | ( ~n14275 & n34190 ) | ( n18332 & n34190 ) ;
  assign n40392 = n9551 | n27368 ;
  assign n40393 = n5226 & ~n13492 ;
  assign n40394 = n17401 ^ n17336 ^ 1'b0 ;
  assign n40395 = n40393 | n40394 ;
  assign n40396 = n4398 | n5334 ;
  assign n40397 = n40395 & ~n40396 ;
  assign n40398 = n40397 ^ n13226 ^ 1'b0 ;
  assign n40399 = ~n11100 & n30542 ;
  assign n40400 = ~n31868 & n40399 ;
  assign n40401 = ( n2687 & n17205 ) | ( n2687 & n20601 ) | ( n17205 & n20601 ) ;
  assign n40402 = n2305 & ~n40401 ;
  assign n40403 = n35472 ^ n23466 ^ n9262 ;
  assign n40404 = ~n12247 & n19438 ;
  assign n40405 = n40404 ^ n23772 ^ 1'b0 ;
  assign n40406 = n3402 & ~n15458 ;
  assign n40407 = n22094 ^ n15860 ^ 1'b0 ;
  assign n40408 = ~n24049 & n40407 ;
  assign n40409 = ( n2795 & n6030 ) | ( n2795 & ~n22987 ) | ( n6030 & ~n22987 ) ;
  assign n40410 = n7341 & n29971 ;
  assign n40411 = n40410 ^ n11724 ^ 1'b0 ;
  assign n40412 = ~n8959 & n40411 ;
  assign n40413 = ( n8882 & n13497 ) | ( n8882 & n40412 ) | ( n13497 & n40412 ) ;
  assign n40414 = ( ~n37450 & n40409 ) | ( ~n37450 & n40413 ) | ( n40409 & n40413 ) ;
  assign n40415 = n18850 & n21158 ;
  assign n40416 = n17643 & n40415 ;
  assign n40417 = ( n16797 & n19630 ) | ( n16797 & n40416 ) | ( n19630 & n40416 ) ;
  assign n40418 = n25155 ^ n8997 ^ n7810 ;
  assign n40420 = n12480 & n25117 ;
  assign n40419 = n19173 & ~n27607 ;
  assign n40421 = n40420 ^ n40419 ^ 1'b0 ;
  assign n40422 = ~n22205 & n36563 ;
  assign n40423 = n30770 & n35080 ;
  assign n40424 = n40423 ^ n18666 ^ n14546 ;
  assign n40425 = n27495 ^ n23266 ^ n1627 ;
  assign n40426 = n40425 ^ n30525 ^ 1'b0 ;
  assign n40427 = ( ~n9848 & n21282 ) | ( ~n9848 & n37450 ) | ( n21282 & n37450 ) ;
  assign n40428 = n29604 ^ n14641 ^ 1'b0 ;
  assign n40429 = n40428 ^ n18534 ^ n15128 ;
  assign n40430 = n11954 ^ n291 ^ 1'b0 ;
  assign n40431 = n26257 | n40430 ;
  assign n40432 = n10569 | n40431 ;
  assign n40433 = n24665 | n40432 ;
  assign n40434 = ~n29349 & n40122 ;
  assign n40435 = n40434 ^ n2752 ^ 1'b0 ;
  assign n40436 = n6829 | n24805 ;
  assign n40437 = ( n4648 & n8056 ) | ( n4648 & ~n21429 ) | ( n8056 & ~n21429 ) ;
  assign n40438 = n17427 ^ n14793 ^ n7398 ;
  assign n40440 = ~n8790 & n10613 ;
  assign n40439 = n7122 | n21476 ;
  assign n40441 = n40440 ^ n40439 ^ 1'b0 ;
  assign n40442 = ( n19086 & n27303 ) | ( n19086 & ~n37158 ) | ( n27303 & ~n37158 ) ;
  assign n40443 = n18992 & ~n20266 ;
  assign n40444 = ~n20514 & n40443 ;
  assign n40445 = ~n5409 & n40444 ;
  assign n40446 = ~n40442 & n40445 ;
  assign n40447 = n22172 ^ n5858 ^ n4830 ;
  assign n40448 = n18800 ^ n3752 ^ 1'b0 ;
  assign n40449 = n33582 & ~n40448 ;
  assign n40450 = n20626 & ~n40449 ;
  assign n40451 = n3854 & ~n20468 ;
  assign n40452 = n23240 ^ n19508 ^ 1'b0 ;
  assign n40454 = ( ~n7786 & n20076 ) | ( ~n7786 & n30278 ) | ( n20076 & n30278 ) ;
  assign n40453 = ~n6482 & n9146 ;
  assign n40455 = n40454 ^ n40453 ^ 1'b0 ;
  assign n40456 = n3748 & ~n39066 ;
  assign n40457 = n40456 ^ n4029 ^ 1'b0 ;
  assign n40458 = n17472 ^ n11770 ^ 1'b0 ;
  assign n40459 = n5804 & n40458 ;
  assign n40460 = ( n1475 & n1625 ) | ( n1475 & n40459 ) | ( n1625 & n40459 ) ;
  assign n40461 = n40460 ^ n18185 ^ 1'b0 ;
  assign n40462 = n38127 & ~n40461 ;
  assign n40463 = n35124 & n40462 ;
  assign n40464 = n9134 & ~n26109 ;
  assign n40465 = n24951 & ~n25151 ;
  assign n40466 = n14651 & n40465 ;
  assign n40467 = n16724 | n40466 ;
  assign n40468 = n40467 ^ n22965 ^ 1'b0 ;
  assign n40469 = n18848 & ~n33850 ;
  assign n40470 = n11603 | n13583 ;
  assign n40471 = n40470 ^ n11859 ^ 1'b0 ;
  assign n40472 = n29353 & n40471 ;
  assign n40473 = n21406 & ~n32890 ;
  assign n40474 = n24982 & ~n28538 ;
  assign n40478 = n17033 ^ n5889 ^ 1'b0 ;
  assign n40479 = n30240 & ~n40478 ;
  assign n40475 = n26088 ^ n16974 ^ 1'b0 ;
  assign n40476 = n22651 & n40475 ;
  assign n40477 = ~n17858 & n40476 ;
  assign n40480 = n40479 ^ n40477 ^ 1'b0 ;
  assign n40481 = n39699 ^ n10077 ^ 1'b0 ;
  assign n40482 = n9468 | n14974 ;
  assign n40483 = n40481 | n40482 ;
  assign n40484 = ~n4568 & n23087 ;
  assign n40485 = n12998 | n40484 ;
  assign n40486 = n40485 ^ n13848 ^ 1'b0 ;
  assign n40487 = n40486 ^ n35249 ^ n7666 ;
  assign n40488 = n15722 & n31459 ;
  assign n40489 = n40488 ^ n18620 ^ n3358 ;
  assign n40490 = n23073 ^ n14766 ^ 1'b0 ;
  assign n40491 = n40490 ^ n10675 ^ n6048 ;
  assign n40492 = n23677 ^ n10634 ^ 1'b0 ;
  assign n40493 = n690 & n9113 ;
  assign n40494 = n6353 & n40493 ;
  assign n40495 = n305 | n40494 ;
  assign n40496 = n5433 & ~n40495 ;
  assign n40497 = n40496 ^ n31094 ^ 1'b0 ;
  assign n40498 = n37567 | n40497 ;
  assign n40501 = ~n8598 & n31427 ;
  assign n40499 = n29738 ^ n17808 ^ n757 ;
  assign n40500 = n12047 & ~n40499 ;
  assign n40502 = n40501 ^ n40500 ^ 1'b0 ;
  assign n40503 = n30241 ^ n7852 ^ n7603 ;
  assign n40504 = n3901 & ~n11284 ;
  assign n40505 = n40504 ^ n11193 ^ 1'b0 ;
  assign n40506 = ( n4256 & ~n18298 ) | ( n4256 & n40505 ) | ( ~n18298 & n40505 ) ;
  assign n40507 = ~n1550 & n13750 ;
  assign n40508 = n40507 ^ n6683 ^ 1'b0 ;
  assign n40509 = ( n11612 & ~n39216 ) | ( n11612 & n40508 ) | ( ~n39216 & n40508 ) ;
  assign n40510 = n13540 | n30722 ;
  assign n40511 = n22079 ^ x122 ^ 1'b0 ;
  assign n40512 = n11389 & ~n40511 ;
  assign n40513 = n18683 ^ n8143 ^ 1'b0 ;
  assign n40514 = n40512 & n40513 ;
  assign n40515 = n19959 & n40514 ;
  assign n40516 = ~n1105 & n40515 ;
  assign n40517 = n40516 ^ n10202 ^ 1'b0 ;
  assign n40518 = n31049 & ~n40517 ;
  assign n40519 = n10842 ^ x83 ^ 1'b0 ;
  assign n40520 = n24529 & ~n40519 ;
  assign n40521 = n25571 & n40520 ;
  assign n40522 = ~n15610 & n40521 ;
  assign n40523 = ~n2468 & n2835 ;
  assign n40524 = ( n18323 & n18467 ) | ( n18323 & ~n24162 ) | ( n18467 & ~n24162 ) ;
  assign n40525 = n40524 ^ n18203 ^ n16300 ;
  assign n40526 = n40525 ^ n15988 ^ 1'b0 ;
  assign n40527 = n40523 | n40526 ;
  assign n40528 = n3162 | n5968 ;
  assign n40529 = ( n24641 & n36457 ) | ( n24641 & n40528 ) | ( n36457 & n40528 ) ;
  assign n40530 = n31923 ^ n24598 ^ 1'b0 ;
  assign n40531 = ( ~n32700 & n39629 ) | ( ~n32700 & n40530 ) | ( n39629 & n40530 ) ;
  assign n40532 = n30435 ^ n9146 ^ 1'b0 ;
  assign n40533 = n3087 & ~n40532 ;
  assign n40534 = n6178 | n40533 ;
  assign n40535 = n14525 ^ n13646 ^ 1'b0 ;
  assign n40537 = ( ~n449 & n2916 ) | ( ~n449 & n8214 ) | ( n2916 & n8214 ) ;
  assign n40536 = n7386 & ~n29674 ;
  assign n40538 = n40537 ^ n40536 ^ n5802 ;
  assign n40539 = n40535 & n40538 ;
  assign n40540 = n15067 & n24259 ;
  assign n40541 = ~n12777 & n40540 ;
  assign n40542 = n40541 ^ n22637 ^ 1'b0 ;
  assign n40543 = n14827 & ~n40542 ;
  assign n40544 = n40543 ^ n39974 ^ n33697 ;
  assign n40545 = n6819 & n40544 ;
  assign n40546 = ( n10166 & ~n17234 ) | ( n10166 & n28103 ) | ( ~n17234 & n28103 ) ;
  assign n40547 = n11673 & ~n40546 ;
  assign n40548 = n33735 & n40547 ;
  assign n40549 = n16131 ^ n12415 ^ 1'b0 ;
  assign n40550 = n25013 & n40549 ;
  assign n40551 = n8178 | n22389 ;
  assign n40552 = n6071 & n19665 ;
  assign n40553 = ~n27253 & n38743 ;
  assign n40554 = ( n14140 & n31431 ) | ( n14140 & n40553 ) | ( n31431 & n40553 ) ;
  assign n40555 = ( n2868 & n15835 ) | ( n2868 & ~n34544 ) | ( n15835 & ~n34544 ) ;
  assign n40556 = ~n14197 & n40555 ;
  assign n40557 = n40556 ^ n20473 ^ 1'b0 ;
  assign n40558 = n39440 ^ n31746 ^ n10605 ;
  assign n40559 = n40558 ^ n9091 ^ 1'b0 ;
  assign n40560 = n18492 ^ n7096 ^ 1'b0 ;
  assign n40561 = n27245 & n40560 ;
  assign n40562 = n3371 & n8165 ;
  assign n40563 = ~n15496 & n40562 ;
  assign n40564 = n21142 ^ n10657 ^ n1030 ;
  assign n40573 = ( n1162 & ~n8950 ) | ( n1162 & n17294 ) | ( ~n8950 & n17294 ) ;
  assign n40565 = n19535 & n37855 ;
  assign n40567 = ( n4589 & ~n15353 ) | ( n4589 & n17048 ) | ( ~n15353 & n17048 ) ;
  assign n40566 = n11313 ^ n5418 ^ n941 ;
  assign n40568 = n40567 ^ n40566 ^ 1'b0 ;
  assign n40569 = n40565 & n40568 ;
  assign n40570 = n40569 ^ n4976 ^ 1'b0 ;
  assign n40571 = n2554 & ~n40570 ;
  assign n40572 = n40571 ^ n30470 ^ n20164 ;
  assign n40574 = n40573 ^ n40572 ^ n4997 ;
  assign n40575 = n34469 ^ n16673 ^ n8357 ;
  assign n40576 = n29537 & n40575 ;
  assign n40577 = n26305 & n36819 ;
  assign n40578 = n40577 ^ n11959 ^ 1'b0 ;
  assign n40579 = n289 | n25941 ;
  assign n40580 = n40579 ^ n9517 ^ 1'b0 ;
  assign n40581 = n40578 | n40580 ;
  assign n40582 = n40581 ^ n4771 ^ 1'b0 ;
  assign n40583 = n37212 ^ n11018 ^ 1'b0 ;
  assign n40584 = n25313 ^ n4770 ^ 1'b0 ;
  assign n40585 = n40583 & ~n40584 ;
  assign n40586 = n23915 ^ n13237 ^ 1'b0 ;
  assign n40587 = n22264 ^ n865 ^ 1'b0 ;
  assign n40588 = ( n1754 & n13731 ) | ( n1754 & n36455 ) | ( n13731 & n36455 ) ;
  assign n40591 = n29024 ^ n2019 ^ 1'b0 ;
  assign n40589 = n7630 & n33313 ;
  assign n40590 = n20376 & n40589 ;
  assign n40592 = n40591 ^ n40590 ^ n8090 ;
  assign n40593 = ( n1351 & ~n6074 ) | ( n1351 & n39772 ) | ( ~n6074 & n39772 ) ;
  assign n40594 = n11803 | n40593 ;
  assign n40595 = n410 & ~n40594 ;
  assign n40596 = n2771 & n7700 ;
  assign n40597 = n5833 | n15680 ;
  assign n40598 = n8159 | n40597 ;
  assign n40599 = ( n783 & n7608 ) | ( n783 & n40598 ) | ( n7608 & n40598 ) ;
  assign n40600 = n40599 ^ n26173 ^ n6620 ;
  assign n40601 = n12363 & ~n40600 ;
  assign n40602 = ( ~x211 & n473 ) | ( ~x211 & n3109 ) | ( n473 & n3109 ) ;
  assign n40603 = n40602 ^ n26501 ^ 1'b0 ;
  assign n40604 = n12834 ^ n2503 ^ 1'b0 ;
  assign n40605 = ~n11118 & n40604 ;
  assign n40606 = ( n4952 & ~n12125 ) | ( n4952 & n16394 ) | ( ~n12125 & n16394 ) ;
  assign n40607 = n8111 | n23111 ;
  assign n40608 = n2484 & ~n40607 ;
  assign n40609 = ~n1247 & n5085 ;
  assign n40610 = n5763 & n40609 ;
  assign n40611 = ( n20573 & ~n40608 ) | ( n20573 & n40610 ) | ( ~n40608 & n40610 ) ;
  assign n40612 = ~n15428 & n35994 ;
  assign n40613 = n40612 ^ n26008 ^ 1'b0 ;
  assign n40614 = ( n4224 & n25908 ) | ( n4224 & n40613 ) | ( n25908 & n40613 ) ;
  assign n40615 = n40614 ^ n392 ^ 1'b0 ;
  assign n40620 = ( ~n9043 & n10929 ) | ( ~n9043 & n15749 ) | ( n10929 & n15749 ) ;
  assign n40618 = n21320 ^ n10386 ^ 1'b0 ;
  assign n40619 = n40618 ^ n32254 ^ n22075 ;
  assign n40621 = n40620 ^ n40619 ^ 1'b0 ;
  assign n40616 = n35530 & ~n35875 ;
  assign n40617 = n40616 ^ n20689 ^ 1'b0 ;
  assign n40622 = n40621 ^ n40617 ^ n20445 ;
  assign n40623 = n10282 & ~n11190 ;
  assign n40624 = n17947 & ~n34211 ;
  assign n40625 = n40624 ^ n15023 ^ 1'b0 ;
  assign n40626 = n36755 & ~n40625 ;
  assign n40627 = n16357 ^ n10761 ^ 1'b0 ;
  assign n40628 = n1301 & n40627 ;
  assign n40630 = ( n6860 & n25295 ) | ( n6860 & ~n26458 ) | ( n25295 & ~n26458 ) ;
  assign n40629 = n35684 ^ n24549 ^ n3116 ;
  assign n40631 = n40630 ^ n40629 ^ n25108 ;
  assign n40632 = ( n23526 & n25104 ) | ( n23526 & ~n39118 ) | ( n25104 & ~n39118 ) ;
  assign n40633 = n14546 ^ x185 ^ 1'b0 ;
  assign n40634 = n31748 | n40633 ;
  assign n40635 = n13201 ^ n2071 ^ n1482 ;
  assign n40636 = ( n4553 & ~n27474 ) | ( n4553 & n40635 ) | ( ~n27474 & n40635 ) ;
  assign n40637 = n40636 ^ n814 ^ 1'b0 ;
  assign n40638 = n21226 & ~n40637 ;
  assign n40641 = n12660 ^ n357 ^ 1'b0 ;
  assign n40642 = n32714 & ~n40641 ;
  assign n40639 = n4655 ^ n1508 ^ 1'b0 ;
  assign n40640 = n40639 ^ n28961 ^ n7522 ;
  assign n40643 = n40642 ^ n40640 ^ n32370 ;
  assign n40644 = n9856 ^ n8972 ^ 1'b0 ;
  assign n40645 = n40643 | n40644 ;
  assign n40646 = n11644 | n29548 ;
  assign n40647 = n40646 ^ n11727 ^ 1'b0 ;
  assign n40648 = n3541 & ~n40647 ;
  assign n40649 = n40648 ^ n31425 ^ 1'b0 ;
  assign n40650 = n11794 ^ n2982 ^ 1'b0 ;
  assign n40651 = n40650 ^ n27457 ^ n6755 ;
  assign n40652 = n1583 & ~n40651 ;
  assign n40653 = n8653 & n40652 ;
  assign n40654 = n11316 | n32275 ;
  assign n40655 = n9064 & n40654 ;
  assign n40656 = ( ~n2529 & n39908 ) | ( ~n2529 & n40655 ) | ( n39908 & n40655 ) ;
  assign n40657 = ~n4323 & n9447 ;
  assign n40658 = n11168 ^ n8986 ^ 1'b0 ;
  assign n40659 = n27965 & n40658 ;
  assign n40660 = ( n9271 & n40657 ) | ( n9271 & ~n40659 ) | ( n40657 & ~n40659 ) ;
  assign n40661 = ~n8199 & n19518 ;
  assign n40662 = n8069 & n21034 ;
  assign n40663 = n34833 ^ n33051 ^ 1'b0 ;
  assign n40664 = n18570 | n40663 ;
  assign n40665 = n3346 & n6979 ;
  assign n40666 = n6577 & n40665 ;
  assign n40667 = n40664 & n40666 ;
  assign n40668 = n11984 ^ n8707 ^ 1'b0 ;
  assign n40670 = n40508 ^ n939 ^ 1'b0 ;
  assign n40671 = n20477 & n40670 ;
  assign n40669 = n16707 & n19810 ;
  assign n40672 = n40671 ^ n40669 ^ 1'b0 ;
  assign n40673 = ( ~n20833 & n40668 ) | ( ~n20833 & n40672 ) | ( n40668 & n40672 ) ;
  assign n40674 = ( n4538 & ~n7079 ) | ( n4538 & n10391 ) | ( ~n7079 & n10391 ) ;
  assign n40675 = n13305 & ~n32848 ;
  assign n40676 = ~n769 & n40675 ;
  assign n40677 = n14120 & ~n24194 ;
  assign n40678 = n32491 ^ n28129 ^ 1'b0 ;
  assign n40679 = n40677 & ~n40678 ;
  assign n40687 = n35604 ^ n13617 ^ 1'b0 ;
  assign n40684 = n10686 | n13585 ;
  assign n40685 = n40684 ^ n8319 ^ 1'b0 ;
  assign n40686 = n4127 & ~n40685 ;
  assign n40688 = n40687 ^ n40686 ^ n17038 ;
  assign n40680 = n21572 ^ n4260 ^ 1'b0 ;
  assign n40681 = n29965 & n40680 ;
  assign n40682 = ~n1305 & n40681 ;
  assign n40683 = n25532 & n40682 ;
  assign n40689 = n40688 ^ n40683 ^ n13970 ;
  assign n40690 = n33605 ^ n15616 ^ n3806 ;
  assign n40691 = ( n21071 & ~n31773 ) | ( n21071 & n38239 ) | ( ~n31773 & n38239 ) ;
  assign n40693 = n13697 ^ n13571 ^ 1'b0 ;
  assign n40694 = n40693 ^ n21408 ^ n3928 ;
  assign n40695 = n17084 & n40694 ;
  assign n40696 = n18957 & ~n40695 ;
  assign n40697 = ~n8001 & n40696 ;
  assign n40692 = n34473 ^ n20196 ^ n2279 ;
  assign n40698 = n40697 ^ n40692 ^ 1'b0 ;
  assign n40699 = n35700 ^ n34365 ^ n28622 ;
  assign n40700 = n25587 ^ n19473 ^ 1'b0 ;
  assign n40701 = ~n36223 & n37991 ;
  assign n40702 = n40701 ^ n15375 ^ 1'b0 ;
  assign n40703 = n23125 ^ n7123 ^ n847 ;
  assign n40709 = n1315 & ~n21046 ;
  assign n40710 = n21046 & n40709 ;
  assign n40711 = n40710 ^ n6644 ^ 1'b0 ;
  assign n40712 = n40711 ^ n26734 ^ n13580 ;
  assign n40704 = n2986 | n12425 ;
  assign n40705 = n12425 & ~n40704 ;
  assign n40706 = n615 | n40705 ;
  assign n40707 = ~n16325 & n33859 ;
  assign n40708 = n40706 & n40707 ;
  assign n40713 = n40712 ^ n40708 ^ 1'b0 ;
  assign n40714 = n12452 ^ n7678 ^ 1'b0 ;
  assign n40715 = n40713 & n40714 ;
  assign n40717 = ( ~n1461 & n4346 ) | ( ~n1461 & n39987 ) | ( n4346 & n39987 ) ;
  assign n40716 = n9890 & ~n29134 ;
  assign n40718 = n40717 ^ n40716 ^ 1'b0 ;
  assign n40719 = n1901 & n2980 ;
  assign n40720 = ( n10841 & ~n11691 ) | ( n10841 & n30998 ) | ( ~n11691 & n30998 ) ;
  assign n40722 = n6121 ^ n5932 ^ 1'b0 ;
  assign n40721 = n8137 ^ n6299 ^ n1342 ;
  assign n40723 = n40722 ^ n40721 ^ n2906 ;
  assign n40724 = ( x86 & n15075 ) | ( x86 & ~n16193 ) | ( n15075 & ~n16193 ) ;
  assign n40725 = n40724 ^ n23098 ^ n18366 ;
  assign n40726 = n40725 ^ n20781 ^ n8913 ;
  assign n40727 = n2764 | n22325 ;
  assign n40728 = n40727 ^ n24662 ^ n5188 ;
  assign n40729 = ~n20371 & n40728 ;
  assign n40730 = n40729 ^ n7492 ^ 1'b0 ;
  assign n40731 = ( n7503 & n33711 ) | ( n7503 & ~n40730 ) | ( n33711 & ~n40730 ) ;
  assign n40732 = ( n3513 & n3738 ) | ( n3513 & n9917 ) | ( n3738 & n9917 ) ;
  assign n40733 = n1891 | n14771 ;
  assign n40734 = ( n14633 & n39223 ) | ( n14633 & n40733 ) | ( n39223 & n40733 ) ;
  assign n40735 = ( ~n9246 & n40732 ) | ( ~n9246 & n40734 ) | ( n40732 & n40734 ) ;
  assign n40736 = ( n21790 & n40731 ) | ( n21790 & n40735 ) | ( n40731 & n40735 ) ;
  assign n40737 = n9368 & n23015 ;
  assign n40738 = ~n34164 & n40737 ;
  assign n40739 = n32253 ^ n6068 ^ n1359 ;
  assign n40740 = ( n28757 & n33460 ) | ( n28757 & n40739 ) | ( n33460 & n40739 ) ;
  assign n40741 = n24151 & ~n40740 ;
  assign n40742 = n40741 ^ n34726 ^ 1'b0 ;
  assign n40743 = n2427 ^ n1697 ^ 1'b0 ;
  assign n40744 = ~n6434 & n40743 ;
  assign n40745 = n40744 ^ n11659 ^ 1'b0 ;
  assign n40746 = n2783 & n23647 ;
  assign n40747 = n40739 ^ n10520 ^ n5129 ;
  assign n40748 = n40747 ^ n24503 ^ n18157 ;
  assign n40749 = n7971 ^ n3325 ^ 1'b0 ;
  assign n40750 = n26495 & ~n40749 ;
  assign n40751 = n40750 ^ n40364 ^ n7953 ;
  assign n40752 = n40751 ^ n26846 ^ n7595 ;
  assign n40753 = n8740 & ~n40752 ;
  assign n40754 = ~n40748 & n40753 ;
  assign n40755 = ( ~n9363 & n20548 ) | ( ~n9363 & n24020 ) | ( n20548 & n24020 ) ;
  assign n40756 = n4996 & ~n18061 ;
  assign n40757 = n40756 ^ n37487 ^ 1'b0 ;
  assign n40758 = n6755 & n18963 ;
  assign n40759 = n40758 ^ n14916 ^ 1'b0 ;
  assign n40760 = n28341 ^ n19778 ^ 1'b0 ;
  assign n40761 = n1289 & ~n40760 ;
  assign n40762 = n40761 ^ n8622 ^ 1'b0 ;
  assign n40763 = n7489 | n40762 ;
  assign n40764 = n40759 | n40763 ;
  assign n40765 = n40764 ^ n16378 ^ 1'b0 ;
  assign n40766 = n14328 ^ n10179 ^ n4989 ;
  assign n40767 = n40766 ^ n35541 ^ n29777 ;
  assign n40768 = n21156 & ~n33837 ;
  assign n40770 = n14013 ^ n2667 ^ 1'b0 ;
  assign n40771 = ~n31987 & n40770 ;
  assign n40769 = n3964 & ~n17673 ;
  assign n40772 = n40771 ^ n40769 ^ 1'b0 ;
  assign n40773 = n36521 & ~n40772 ;
  assign n40774 = ~n18550 & n40773 ;
  assign n40775 = n21403 ^ n6874 ^ 1'b0 ;
  assign n40776 = n7300 & n40775 ;
  assign n40777 = n40776 ^ n27547 ^ n22504 ;
  assign n40778 = n25274 ^ n8898 ^ 1'b0 ;
  assign n40779 = n40778 ^ n12615 ^ 1'b0 ;
  assign n40780 = n40777 & ~n40779 ;
  assign n40782 = ( n4080 & ~n7704 ) | ( n4080 & n10885 ) | ( ~n7704 & n10885 ) ;
  assign n40781 = n2444 & n19884 ;
  assign n40783 = n40782 ^ n40781 ^ 1'b0 ;
  assign n40786 = ( n431 & n1180 ) | ( n431 & ~n23575 ) | ( n1180 & ~n23575 ) ;
  assign n40784 = n31543 ^ n8142 ^ 1'b0 ;
  assign n40785 = n6874 | n40784 ;
  assign n40787 = n40786 ^ n40785 ^ 1'b0 ;
  assign n40788 = n40783 & n40787 ;
  assign n40789 = n13359 ^ n4852 ^ 1'b0 ;
  assign n40790 = n16131 & ~n40789 ;
  assign n40791 = ( n21375 & n32712 ) | ( n21375 & ~n40790 ) | ( n32712 & ~n40790 ) ;
  assign n40792 = n31916 ^ n5204 ^ n2765 ;
  assign n40793 = n16802 ^ n14741 ^ n1385 ;
  assign n40794 = n40792 & n40793 ;
  assign n40795 = n18549 | n18673 ;
  assign n40796 = n14665 ^ n2803 ^ 1'b0 ;
  assign n40797 = n40795 & n40796 ;
  assign n40798 = ( n2596 & n29209 ) | ( n2596 & ~n40797 ) | ( n29209 & ~n40797 ) ;
  assign n40799 = n34002 ^ n7283 ^ 1'b0 ;
  assign n40800 = ~n38415 & n40799 ;
  assign n40801 = ( n19610 & n20343 ) | ( n19610 & n40800 ) | ( n20343 & n40800 ) ;
  assign n40802 = ( n17729 & n27110 ) | ( n17729 & n30929 ) | ( n27110 & n30929 ) ;
  assign n40803 = ~n4110 & n15786 ;
  assign n40804 = n2682 & ~n7248 ;
  assign n40805 = n40804 ^ n5485 ^ 1'b0 ;
  assign n40806 = n2509 | n40805 ;
  assign n40807 = n40803 | n40806 ;
  assign n40808 = n15771 | n35384 ;
  assign n40809 = n40808 ^ n19146 ^ 1'b0 ;
  assign n40810 = ( n6634 & ~n15548 ) | ( n6634 & n40809 ) | ( ~n15548 & n40809 ) ;
  assign n40811 = n32993 & ~n40810 ;
  assign n40812 = ~n34543 & n40811 ;
  assign n40813 = n16121 | n20936 ;
  assign n40814 = n40813 ^ n17289 ^ 1'b0 ;
  assign n40815 = n19098 & ~n33118 ;
  assign n40816 = n40815 ^ n6780 ^ 1'b0 ;
  assign n40817 = n16667 ^ n13915 ^ 1'b0 ;
  assign n40819 = n26119 | n30645 ;
  assign n40818 = ( n9926 & ~n14316 ) | ( n9926 & n23762 ) | ( ~n14316 & n23762 ) ;
  assign n40820 = n40819 ^ n40818 ^ n14491 ;
  assign n40821 = n34040 ^ n14507 ^ n3250 ;
  assign n40822 = n7678 & ~n23137 ;
  assign n40823 = ( n7596 & n11330 ) | ( n7596 & n13710 ) | ( n11330 & n13710 ) ;
  assign n40824 = ( ~n8465 & n31088 ) | ( ~n8465 & n40823 ) | ( n31088 & n40823 ) ;
  assign n40825 = n40824 ^ n11325 ^ 1'b0 ;
  assign n40826 = n40822 | n40825 ;
  assign n40827 = n2445 | n17009 ;
  assign n40828 = n40827 ^ n33572 ^ 1'b0 ;
  assign n40829 = n6000 & ~n19279 ;
  assign n40830 = n40829 ^ n24541 ^ 1'b0 ;
  assign n40831 = n15906 & n32738 ;
  assign n40832 = n29502 ^ n6092 ^ n3323 ;
  assign n40833 = n9542 & n29703 ;
  assign n40834 = ~n5021 & n40833 ;
  assign n40835 = n40834 ^ n14050 ^ 1'b0 ;
  assign n40836 = n40835 ^ n8109 ^ 1'b0 ;
  assign n40837 = ~n28647 & n40836 ;
  assign n40838 = n16952 ^ n15174 ^ 1'b0 ;
  assign n40839 = n40166 ^ n23263 ^ n1646 ;
  assign n40840 = n12222 | n40839 ;
  assign n40841 = n40840 ^ n19577 ^ 1'b0 ;
  assign n40842 = n33312 & n40841 ;
  assign n40843 = n14259 ^ n10650 ^ n3656 ;
  assign n40844 = n842 & ~n8632 ;
  assign n40845 = n40844 ^ n33929 ^ 1'b0 ;
  assign n40846 = n24033 & ~n40845 ;
  assign n40847 = n25218 & ~n40846 ;
  assign n40848 = n5909 & ~n10399 ;
  assign n40849 = n4557 & ~n14195 ;
  assign n40850 = n40849 ^ n12908 ^ 1'b0 ;
  assign n40851 = ( n3298 & n40848 ) | ( n3298 & n40850 ) | ( n40848 & n40850 ) ;
  assign n40852 = n40851 ^ n1908 ^ 1'b0 ;
  assign n40853 = n11261 ^ n3946 ^ 1'b0 ;
  assign n40854 = ~n8653 & n40853 ;
  assign n40855 = n40854 ^ n19476 ^ n10514 ;
  assign n40856 = ( n9956 & ~n9991 ) | ( n9956 & n40855 ) | ( ~n9991 & n40855 ) ;
  assign n40857 = ~n22564 & n40856 ;
  assign n40858 = ~n550 & n40857 ;
  assign n40863 = n12733 ^ n2369 ^ n1542 ;
  assign n40862 = n32023 ^ n27792 ^ 1'b0 ;
  assign n40859 = n11542 & ~n15440 ;
  assign n40860 = n40859 ^ n25744 ^ 1'b0 ;
  assign n40861 = ( ~n11996 & n30546 ) | ( ~n11996 & n40860 ) | ( n30546 & n40860 ) ;
  assign n40864 = n40863 ^ n40862 ^ n40861 ;
  assign n40865 = ~n19026 & n25071 ;
  assign n40866 = n10922 | n15315 ;
  assign n40867 = n39339 & ~n40866 ;
  assign n40870 = ( n8894 & n19143 ) | ( n8894 & ~n26895 ) | ( n19143 & ~n26895 ) ;
  assign n40868 = n2841 | n20848 ;
  assign n40869 = n24083 | n40868 ;
  assign n40871 = n40870 ^ n40869 ^ n6068 ;
  assign n40872 = n22042 ^ n5019 ^ n2887 ;
  assign n40873 = ( n5631 & ~n20736 ) | ( n5631 & n21986 ) | ( ~n20736 & n21986 ) ;
  assign n40874 = ( ~n27663 & n40872 ) | ( ~n27663 & n40873 ) | ( n40872 & n40873 ) ;
  assign n40878 = n5474 & ~n23460 ;
  assign n40875 = n16262 ^ n8768 ^ 1'b0 ;
  assign n40876 = n26209 ^ n2226 ^ 1'b0 ;
  assign n40877 = n40875 & n40876 ;
  assign n40879 = n40878 ^ n40877 ^ n8236 ;
  assign n40880 = n40879 ^ n24023 ^ 1'b0 ;
  assign n40881 = n30701 | n37104 ;
  assign n40882 = n6788 | n40881 ;
  assign n40884 = ~n2127 & n9249 ;
  assign n40885 = ~n35282 & n40884 ;
  assign n40886 = n40885 ^ n24907 ^ x44 ;
  assign n40887 = n2994 ^ n1104 ^ 1'b0 ;
  assign n40888 = n19533 & ~n40887 ;
  assign n40889 = n40886 & n40888 ;
  assign n40883 = n3368 & n9033 ;
  assign n40890 = n40889 ^ n40883 ^ 1'b0 ;
  assign n40891 = n39617 ^ n38460 ^ n14462 ;
  assign n40892 = ( n8297 & ~n15830 ) | ( n8297 & n16195 ) | ( ~n15830 & n16195 ) ;
  assign n40893 = n35355 | n37817 ;
  assign n40894 = ~n2595 & n13548 ;
  assign n40895 = n31440 ^ n21000 ^ n14520 ;
  assign n40896 = n3692 & n18474 ;
  assign n40897 = ~n33313 & n40896 ;
  assign n40898 = n11155 ^ n8956 ^ 1'b0 ;
  assign n40899 = n40898 ^ n22535 ^ 1'b0 ;
  assign n40900 = n34938 ^ n20404 ^ 1'b0 ;
  assign n40901 = n9242 ^ n3923 ^ n3030 ;
  assign n40902 = ~n11815 & n13951 ;
  assign n40903 = ( ~n2968 & n30738 ) | ( ~n2968 & n33074 ) | ( n30738 & n33074 ) ;
  assign n40904 = ( n40901 & n40902 ) | ( n40901 & n40903 ) | ( n40902 & n40903 ) ;
  assign n40905 = n4923 ^ n4741 ^ 1'b0 ;
  assign n40906 = n1939 & n40905 ;
  assign n40907 = ( n5401 & ~n9635 ) | ( n5401 & n40906 ) | ( ~n9635 & n40906 ) ;
  assign n40908 = ( n8529 & n13940 ) | ( n8529 & n40907 ) | ( n13940 & n40907 ) ;
  assign n40909 = n20636 ^ n7169 ^ 1'b0 ;
  assign n40910 = n11326 & n15465 ;
  assign n40911 = n40910 ^ n3669 ^ 1'b0 ;
  assign n40912 = n25475 ^ n22732 ^ n13668 ;
  assign n40913 = n6878 ^ n3960 ^ 1'b0 ;
  assign n40914 = n14448 & n25858 ;
  assign n40915 = n40914 ^ n6270 ^ 1'b0 ;
  assign n40916 = ( n20362 & ~n40913 ) | ( n20362 & n40915 ) | ( ~n40913 & n40915 ) ;
  assign n40917 = ( n25566 & n32432 ) | ( n25566 & ~n34910 ) | ( n32432 & ~n34910 ) ;
  assign n40918 = n30960 ^ n23291 ^ 1'b0 ;
  assign n40919 = ( ~n25235 & n40917 ) | ( ~n25235 & n40918 ) | ( n40917 & n40918 ) ;
  assign n40920 = n34164 ^ n1417 ^ 1'b0 ;
  assign n40921 = n40920 ^ n18993 ^ 1'b0 ;
  assign n40924 = ~n5381 & n5524 ;
  assign n40925 = n22402 & n28643 ;
  assign n40926 = n40924 & n40925 ;
  assign n40922 = n3641 & ~n12660 ;
  assign n40923 = n38460 & ~n40922 ;
  assign n40927 = n40926 ^ n40923 ^ 1'b0 ;
  assign n40928 = n22492 & ~n25642 ;
  assign n40929 = n9034 | n13048 ;
  assign n40930 = n40928 & ~n40929 ;
  assign n40934 = ~n5349 & n9996 ;
  assign n40935 = n10759 & n40934 ;
  assign n40931 = n1468 & n1885 ;
  assign n40932 = n40931 ^ n421 ^ 1'b0 ;
  assign n40933 = ( n2781 & n8247 ) | ( n2781 & n40932 ) | ( n8247 & n40932 ) ;
  assign n40936 = n40935 ^ n40933 ^ x24 ;
  assign n40937 = n30536 ^ n30445 ^ n15810 ;
  assign n40938 = n17819 ^ n17719 ^ 1'b0 ;
  assign n40939 = n31501 | n40938 ;
  assign n40940 = n511 & n38135 ;
  assign n40941 = n40940 ^ n20168 ^ 1'b0 ;
  assign n40942 = n9067 & ~n16462 ;
  assign n40943 = n40942 ^ n4256 ^ 1'b0 ;
  assign n40946 = n2173 & ~n34223 ;
  assign n40944 = n23505 ^ n9853 ^ n324 ;
  assign n40945 = n40944 ^ n28026 ^ n13898 ;
  assign n40947 = n40946 ^ n40945 ^ n15109 ;
  assign n40948 = n16663 ^ n4597 ^ 1'b0 ;
  assign n40949 = ~n325 & n40948 ;
  assign n40950 = ~n29295 & n40949 ;
  assign n40951 = n8810 & ~n34262 ;
  assign n40952 = n31458 | n40951 ;
  assign n40953 = ~n30425 & n35265 ;
  assign n40954 = ~n3095 & n40953 ;
  assign n40955 = n29839 & n40954 ;
  assign n40956 = n5257 & n7821 ;
  assign n40957 = ( n4041 & n16252 ) | ( n4041 & n23477 ) | ( n16252 & n23477 ) ;
  assign n40958 = n32665 ^ n10653 ^ n4342 ;
  assign n40962 = n35883 ^ n19190 ^ n1963 ;
  assign n40959 = n6254 | n13428 ;
  assign n40960 = n40959 ^ n7331 ^ 1'b0 ;
  assign n40961 = n40960 ^ n19867 ^ 1'b0 ;
  assign n40963 = n40962 ^ n40961 ^ n19819 ;
  assign n40964 = ~n2476 & n23417 ;
  assign n40965 = ~n1901 & n40964 ;
  assign n40966 = n39372 ^ n24659 ^ 1'b0 ;
  assign n40967 = n40965 | n40966 ;
  assign n40969 = n11823 ^ n8573 ^ n1672 ;
  assign n40968 = n13476 & n24916 ;
  assign n40970 = n40969 ^ n40968 ^ 1'b0 ;
  assign n40971 = ~n33196 & n40970 ;
  assign n40972 = n40971 ^ n5006 ^ 1'b0 ;
  assign n40973 = n27704 ^ n16322 ^ 1'b0 ;
  assign n40974 = ~n1176 & n40973 ;
  assign n40976 = ~n8824 & n36835 ;
  assign n40977 = n40976 ^ n2276 ^ 1'b0 ;
  assign n40975 = n1223 & ~n18795 ;
  assign n40978 = n40977 ^ n40975 ^ 1'b0 ;
  assign n40979 = n777 | n16506 ;
  assign n40980 = n18641 & ~n40979 ;
  assign n40981 = ( ~n6333 & n18048 ) | ( ~n6333 & n19324 ) | ( n18048 & n19324 ) ;
  assign n40982 = n40981 ^ n1305 ^ 1'b0 ;
  assign n40983 = n14834 | n31937 ;
  assign n40984 = n40982 | n40983 ;
  assign n40985 = n37616 ^ n16629 ^ 1'b0 ;
  assign n40986 = ( ~n14463 & n19844 ) | ( ~n14463 & n40985 ) | ( n19844 & n40985 ) ;
  assign n40987 = ( ~x49 & n30826 ) | ( ~x49 & n38257 ) | ( n30826 & n38257 ) ;
  assign n40988 = n602 & ~n40987 ;
  assign n40989 = n7151 & ~n30702 ;
  assign n40990 = ~n22561 & n40989 ;
  assign n40991 = n4300 & n34475 ;
  assign n40992 = n40990 & n40991 ;
  assign n40993 = n32990 ^ n10571 ^ 1'b0 ;
  assign n40994 = n27598 | n32240 ;
  assign n40995 = n18614 & ~n40994 ;
  assign n40996 = n421 & ~n21515 ;
  assign n40998 = ( ~n18750 & n23054 ) | ( ~n18750 & n40851 ) | ( n23054 & n40851 ) ;
  assign n40997 = n33298 & ~n35462 ;
  assign n40999 = n40998 ^ n40997 ^ 1'b0 ;
  assign n41000 = n12420 & n28164 ;
  assign n41001 = n10139 & ~n41000 ;
  assign n41002 = n41001 ^ n35181 ^ 1'b0 ;
  assign n41003 = n22528 & ~n35870 ;
  assign n41004 = n18662 & ~n41003 ;
  assign n41005 = ~n7238 & n41004 ;
  assign n41006 = x148 & ~n41005 ;
  assign n41007 = n26939 ^ n14533 ^ 1'b0 ;
  assign n41008 = n41007 ^ n8861 ^ 1'b0 ;
  assign n41009 = n13888 ^ n13000 ^ n796 ;
  assign n41010 = n31850 ^ n10846 ^ 1'b0 ;
  assign n41011 = ( n6551 & n14397 ) | ( n6551 & ~n23016 ) | ( n14397 & ~n23016 ) ;
  assign n41012 = n31508 ^ n20559 ^ 1'b0 ;
  assign n41013 = n15359 & n41012 ;
  assign n41014 = ( n15020 & ~n16958 ) | ( n15020 & n17808 ) | ( ~n16958 & n17808 ) ;
  assign n41015 = n41014 ^ n32828 ^ n27515 ;
  assign n41016 = n2030 & ~n8614 ;
  assign n41017 = n13383 & n41016 ;
  assign n41018 = ( ~n23923 & n27342 ) | ( ~n23923 & n41017 ) | ( n27342 & n41017 ) ;
  assign n41019 = n19006 ^ n18801 ^ n15344 ;
  assign n41020 = n3055 & n41019 ;
  assign n41021 = ~n11462 & n40743 ;
  assign n41022 = n2470 & n41021 ;
  assign n41023 = n35444 ^ n11303 ^ 1'b0 ;
  assign n41024 = ( n8854 & n41022 ) | ( n8854 & ~n41023 ) | ( n41022 & ~n41023 ) ;
  assign n41025 = n2149 & ~n22688 ;
  assign n41026 = n41025 ^ n8904 ^ 1'b0 ;
  assign n41027 = ( n15104 & ~n20206 ) | ( n15104 & n41026 ) | ( ~n20206 & n41026 ) ;
  assign n41028 = n15797 & ~n32142 ;
  assign n41029 = n12331 & n41028 ;
  assign n41030 = n41029 ^ n18070 ^ n16961 ;
  assign n41031 = n41030 ^ n18977 ^ n11883 ;
  assign n41032 = n41031 ^ n14284 ^ 1'b0 ;
  assign n41033 = n19244 ^ n9743 ^ n7182 ;
  assign n41034 = n41033 ^ n5866 ^ 1'b0 ;
  assign n41035 = n41032 & n41034 ;
  assign n41036 = n13894 & ~n29002 ;
  assign n41037 = ~n29343 & n41036 ;
  assign n41039 = n16663 & n17176 ;
  assign n41040 = n7110 & n41039 ;
  assign n41038 = n1067 & ~n1331 ;
  assign n41041 = n41040 ^ n41038 ^ 1'b0 ;
  assign n41042 = ~n24813 & n29551 ;
  assign n41043 = n41042 ^ n14052 ^ 1'b0 ;
  assign n41046 = x34 & n39275 ;
  assign n41044 = n23217 ^ n8809 ^ 1'b0 ;
  assign n41045 = n7030 | n41044 ;
  assign n41047 = n41046 ^ n41045 ^ n14292 ;
  assign n41048 = n7464 & ~n12820 ;
  assign n41049 = ( n19229 & ~n23318 ) | ( n19229 & n38556 ) | ( ~n23318 & n38556 ) ;
  assign n41050 = n10314 & ~n12607 ;
  assign n41051 = n41050 ^ n13344 ^ 1'b0 ;
  assign n41052 = n22405 | n26823 ;
  assign n41053 = n533 & n20306 ;
  assign n41054 = ( n28834 & ~n41052 ) | ( n28834 & n41053 ) | ( ~n41052 & n41053 ) ;
  assign n41055 = n609 | n19640 ;
  assign n41056 = n41055 ^ n13161 ^ 1'b0 ;
  assign n41057 = n34762 & ~n41056 ;
  assign n41058 = ~n41054 & n41057 ;
  assign n41060 = n1571 & ~n29877 ;
  assign n41059 = n10826 | n13335 ;
  assign n41061 = n41060 ^ n41059 ^ 1'b0 ;
  assign n41062 = n21686 ^ n18474 ^ 1'b0 ;
  assign n41063 = n41062 ^ n33615 ^ n3683 ;
  assign n41064 = ( n20974 & n27417 ) | ( n20974 & n30026 ) | ( n27417 & n30026 ) ;
  assign n41065 = n1666 & n38131 ;
  assign n41066 = n41065 ^ n22595 ^ 1'b0 ;
  assign n41067 = n31662 ^ n4081 ^ 1'b0 ;
  assign n41068 = n3750 & n41067 ;
  assign n41069 = ( n8902 & n11460 ) | ( n8902 & ~n41068 ) | ( n11460 & ~n41068 ) ;
  assign n41070 = n41069 ^ n1996 ^ 1'b0 ;
  assign n41071 = ~n1258 & n26227 ;
  assign n41072 = ~n41070 & n41071 ;
  assign n41073 = n1879 & n36295 ;
  assign n41074 = n35410 ^ n21687 ^ n15998 ;
  assign n41075 = ( n8711 & ~n23281 ) | ( n8711 & n27993 ) | ( ~n23281 & n27993 ) ;
  assign n41076 = ( ~n23980 & n41074 ) | ( ~n23980 & n41075 ) | ( n41074 & n41075 ) ;
  assign n41077 = n17379 ^ n7119 ^ n4554 ;
  assign n41078 = n17141 & n41077 ;
  assign n41079 = ( ~n7174 & n10921 ) | ( ~n7174 & n15917 ) | ( n10921 & n15917 ) ;
  assign n41080 = n4231 & n41079 ;
  assign n41081 = n37935 & ~n41080 ;
  assign n41082 = n41081 ^ n20751 ^ 1'b0 ;
  assign n41083 = n20112 | n27259 ;
  assign n41084 = n2965 | n41083 ;
  assign n41085 = n41084 ^ n10820 ^ 1'b0 ;
  assign n41086 = n4737 | n31483 ;
  assign n41087 = n41086 ^ n16439 ^ 1'b0 ;
  assign n41088 = n3479 ^ n1374 ^ 1'b0 ;
  assign n41089 = n35982 | n41088 ;
  assign n41090 = n13464 & ~n41089 ;
  assign n41093 = n15548 ^ n5299 ^ n4740 ;
  assign n41091 = n26159 ^ n14332 ^ n9745 ;
  assign n41092 = n2820 & ~n41091 ;
  assign n41094 = n41093 ^ n41092 ^ 1'b0 ;
  assign n41095 = ~n4100 & n41094 ;
  assign n41096 = ( n16774 & ~n17302 ) | ( n16774 & n39761 ) | ( ~n17302 & n39761 ) ;
  assign n41097 = n37048 ^ n29509 ^ 1'b0 ;
  assign n41099 = ( n5797 & n22195 ) | ( n5797 & n36582 ) | ( n22195 & n36582 ) ;
  assign n41100 = ( n4232 & n8433 ) | ( n4232 & n41099 ) | ( n8433 & n41099 ) ;
  assign n41101 = n41100 ^ n29699 ^ n5789 ;
  assign n41098 = n19938 | n26562 ;
  assign n41102 = n41101 ^ n41098 ^ 1'b0 ;
  assign n41103 = n1101 ^ n919 ^ 1'b0 ;
  assign n41104 = ~n24599 & n41103 ;
  assign n41105 = n41104 ^ n20574 ^ 1'b0 ;
  assign n41106 = n17618 ^ n8735 ^ 1'b0 ;
  assign n41107 = ~n19049 & n41106 ;
  assign n41108 = n41107 ^ n9177 ^ 1'b0 ;
  assign n41110 = n3742 & ~n9552 ;
  assign n41111 = n41110 ^ n10775 ^ 1'b0 ;
  assign n41112 = n40331 | n41111 ;
  assign n41109 = ( n1039 & ~n11609 ) | ( n1039 & n20196 ) | ( ~n11609 & n20196 ) ;
  assign n41113 = n41112 ^ n41109 ^ 1'b0 ;
  assign n41114 = ( n11409 & n13264 ) | ( n11409 & ~n13800 ) | ( n13264 & ~n13800 ) ;
  assign n41115 = n41114 ^ n30393 ^ 1'b0 ;
  assign n41116 = ~n284 & n41115 ;
  assign n41117 = n36781 ^ n27054 ^ x144 ;
  assign n41118 = n7377 ^ n2700 ^ 1'b0 ;
  assign n41119 = n11724 & ~n13191 ;
  assign n41120 = n17827 & n24293 ;
  assign n41121 = n37504 & n41120 ;
  assign n41122 = n24729 ^ n8230 ^ 1'b0 ;
  assign n41123 = n33137 ^ n32879 ^ n30110 ;
  assign n41124 = ( n5371 & ~n10926 ) | ( n5371 & n14485 ) | ( ~n10926 & n14485 ) ;
  assign n41125 = ( n6428 & n25700 ) | ( n6428 & n41124 ) | ( n25700 & n41124 ) ;
  assign n41126 = n38600 ^ n6543 ^ 1'b0 ;
  assign n41127 = n41125 & n41126 ;
  assign n41128 = n28082 & n41127 ;
  assign n41129 = ( n4767 & ~n8992 ) | ( n4767 & n41128 ) | ( ~n8992 & n41128 ) ;
  assign n41130 = ( n322 & n8169 ) | ( n322 & ~n26083 ) | ( n8169 & ~n26083 ) ;
  assign n41131 = n4283 & ~n39965 ;
  assign n41132 = ~n11622 & n41131 ;
  assign n41133 = ( n2768 & n34676 ) | ( n2768 & ~n41132 ) | ( n34676 & ~n41132 ) ;
  assign n41134 = n41130 | n41133 ;
  assign n41135 = n33637 ^ n5627 ^ 1'b0 ;
  assign n41136 = n18767 & ~n41135 ;
  assign n41137 = ~n34415 & n36870 ;
  assign n41138 = n332 & ~n13260 ;
  assign n41139 = ( ~n2326 & n38408 ) | ( ~n2326 & n41138 ) | ( n38408 & n41138 ) ;
  assign n41140 = n41139 ^ n2980 ^ 1'b0 ;
  assign n41141 = n14163 | n41140 ;
  assign n41142 = n27696 ^ n5568 ^ 1'b0 ;
  assign n41143 = n26273 ^ n4232 ^ 1'b0 ;
  assign n41144 = ~n41066 & n41143 ;
  assign n41145 = ~n41142 & n41144 ;
  assign n41146 = n7421 & n35850 ;
  assign n41147 = ~n14717 & n41146 ;
  assign n41152 = n18571 ^ n9352 ^ 1'b0 ;
  assign n41153 = ~n2924 & n41152 ;
  assign n41148 = n36065 ^ n7637 ^ 1'b0 ;
  assign n41149 = n2712 & n41148 ;
  assign n41150 = n41149 ^ n22147 ^ 1'b0 ;
  assign n41151 = ~n27616 & n41150 ;
  assign n41154 = n41153 ^ n41151 ^ 1'b0 ;
  assign n41158 = n22151 ^ n9921 ^ n7280 ;
  assign n41156 = n17175 | n22297 ;
  assign n41157 = n41156 ^ n25783 ^ 1'b0 ;
  assign n41159 = n41158 ^ n41157 ^ n21062 ;
  assign n41160 = n33729 ^ n20005 ^ 1'b0 ;
  assign n41161 = n41159 & ~n41160 ;
  assign n41155 = ~n19205 & n26367 ;
  assign n41162 = n41161 ^ n41155 ^ 1'b0 ;
  assign n41163 = ( n16691 & n29368 ) | ( n16691 & ~n41162 ) | ( n29368 & ~n41162 ) ;
  assign n41164 = ( n1127 & ~n1632 ) | ( n1127 & n12101 ) | ( ~n1632 & n12101 ) ;
  assign n41165 = ~n2362 & n16412 ;
  assign n41166 = ( n11302 & n41164 ) | ( n11302 & ~n41165 ) | ( n41164 & ~n41165 ) ;
  assign n41167 = n33265 & n38793 ;
  assign n41168 = n9238 & n22303 ;
  assign n41169 = n41168 ^ n1758 ^ 1'b0 ;
  assign n41170 = n14458 & n41169 ;
  assign n41171 = n7551 | n31281 ;
  assign n41172 = n41171 ^ n14776 ^ n12348 ;
  assign n41173 = n41172 ^ n5982 ^ 1'b0 ;
  assign n41174 = n26613 ^ n10442 ^ 1'b0 ;
  assign n41175 = n41173 & ~n41174 ;
  assign n41176 = n29455 ^ n23323 ^ 1'b0 ;
  assign n41177 = ~n5476 & n41176 ;
  assign n41178 = ~n13539 & n37279 ;
  assign n41179 = n41178 ^ n20817 ^ 1'b0 ;
  assign n41180 = n41179 ^ n22332 ^ n3586 ;
  assign n41183 = n8327 | n8604 ;
  assign n41184 = n8327 & ~n41183 ;
  assign n41181 = n16658 & n16675 ;
  assign n41182 = ~n16675 & n41181 ;
  assign n41185 = n41184 ^ n41182 ^ n23213 ;
  assign n41186 = n34642 ^ n14638 ^ 1'b0 ;
  assign n41187 = n1986 & n41186 ;
  assign n41188 = n18556 & n24304 ;
  assign n41189 = ( n899 & n16665 ) | ( n899 & ~n28727 ) | ( n16665 & ~n28727 ) ;
  assign n41190 = n41189 ^ n13464 ^ 1'b0 ;
  assign n41191 = n41190 ^ n33478 ^ n16711 ;
  assign n41192 = ~n10928 & n16901 ;
  assign n41193 = n41192 ^ n12897 ^ 1'b0 ;
  assign n41195 = n5951 & ~n6915 ;
  assign n41194 = x153 & n7754 ;
  assign n41196 = n41195 ^ n41194 ^ n6362 ;
  assign n41199 = ~n284 & n23052 ;
  assign n41200 = n41199 ^ n22167 ^ 1'b0 ;
  assign n41197 = n28592 ^ n1524 ^ 1'b0 ;
  assign n41198 = n25753 & n41197 ;
  assign n41201 = n41200 ^ n41198 ^ n11339 ;
  assign n41202 = n3067 & n4142 ;
  assign n41203 = n41202 ^ n3032 ^ 1'b0 ;
  assign n41204 = n41203 ^ n30081 ^ 1'b0 ;
  assign n41205 = n35958 & n41204 ;
  assign n41206 = n41205 ^ n40499 ^ n12457 ;
  assign n41207 = n6757 & n9278 ;
  assign n41208 = n33201 ^ n25519 ^ n8503 ;
  assign n41209 = ( x195 & n39080 ) | ( x195 & n41208 ) | ( n39080 & n41208 ) ;
  assign n41210 = ( n12147 & n13327 ) | ( n12147 & ~n40664 ) | ( n13327 & ~n40664 ) ;
  assign n41212 = n4501 & ~n10028 ;
  assign n41213 = ~n17565 & n41212 ;
  assign n41211 = ( n1669 & ~n4260 ) | ( n1669 & n5570 ) | ( ~n4260 & n5570 ) ;
  assign n41214 = n41213 ^ n41211 ^ n6819 ;
  assign n41215 = n41214 ^ n7815 ^ 1'b0 ;
  assign n41216 = n41210 & n41215 ;
  assign n41217 = n6584 | n27626 ;
  assign n41218 = n21443 ^ n18815 ^ n14044 ;
  assign n41219 = n34712 ^ n24457 ^ n23684 ;
  assign n41220 = n36937 ^ n5415 ^ 1'b0 ;
  assign n41221 = n33872 ^ n21698 ^ 1'b0 ;
  assign n41222 = n41221 ^ n6854 ^ n1315 ;
  assign n41223 = n31004 ^ n15701 ^ n11248 ;
  assign n41224 = n14606 & n24893 ;
  assign n41225 = ~n9762 & n41224 ;
  assign n41226 = ( n11901 & n22092 ) | ( n11901 & n41225 ) | ( n22092 & n41225 ) ;
  assign n41227 = n17165 ^ n4617 ^ 1'b0 ;
  assign n41228 = n24135 & ~n41227 ;
  assign n41229 = n41228 ^ n35185 ^ 1'b0 ;
  assign n41230 = n6288 & n12902 ;
  assign n41231 = n41230 ^ n7771 ^ 1'b0 ;
  assign n41233 = ~n17932 & n18008 ;
  assign n41232 = n9143 & n10116 ;
  assign n41234 = n41233 ^ n41232 ^ 1'b0 ;
  assign n41235 = n15167 & ~n41234 ;
  assign n41236 = x66 & ~n13322 ;
  assign n41237 = ~n40017 & n41236 ;
  assign n41238 = n5923 ^ n1926 ^ 1'b0 ;
  assign n41239 = ~n26732 & n41238 ;
  assign n41240 = n3905 | n41239 ;
  assign n41241 = ( n17378 & ~n25417 ) | ( n17378 & n30488 ) | ( ~n25417 & n30488 ) ;
  assign n41242 = ~n1278 & n2233 ;
  assign n41243 = n41242 ^ n40352 ^ n2828 ;
  assign n41244 = n9563 & n10546 ;
  assign n41245 = n2914 | n4235 ;
  assign n41246 = n3266 & ~n41245 ;
  assign n41247 = n2134 | n27428 ;
  assign n41248 = n41247 ^ n39946 ^ 1'b0 ;
  assign n41249 = ~n13548 & n41248 ;
  assign n41250 = ~n9972 & n11532 ;
  assign n41251 = ~n4471 & n41250 ;
  assign n41252 = n14051 ^ n8319 ^ n3536 ;
  assign n41253 = ( n6128 & ~n24982 ) | ( n6128 & n41252 ) | ( ~n24982 & n41252 ) ;
  assign n41254 = ~n41251 & n41253 ;
  assign n41256 = n25314 ^ n13289 ^ n9904 ;
  assign n41255 = n6878 ^ x117 ^ 1'b0 ;
  assign n41257 = n41256 ^ n41255 ^ 1'b0 ;
  assign n41258 = n41257 ^ n13553 ^ 1'b0 ;
  assign n41259 = ( n6342 & n25104 ) | ( n6342 & ~n36919 ) | ( n25104 & ~n36919 ) ;
  assign n41260 = ( n13027 & n24163 ) | ( n13027 & ~n41259 ) | ( n24163 & ~n41259 ) ;
  assign n41261 = n10873 & n11810 ;
  assign n41262 = n15413 & n41261 ;
  assign n41263 = n16312 | n41262 ;
  assign n41264 = n41263 ^ n16878 ^ n7879 ;
  assign n41265 = n40018 ^ n5476 ^ n681 ;
  assign n41266 = n41265 ^ n16081 ^ n4243 ;
  assign n41267 = n6853 & ~n25576 ;
  assign n41269 = n5263 & n29921 ;
  assign n41268 = ~n3932 & n5365 ;
  assign n41270 = n41269 ^ n41268 ^ n14710 ;
  assign n41271 = n41270 ^ n32792 ^ n13369 ;
  assign n41272 = ~n16609 & n35503 ;
  assign n41273 = ~n8984 & n41272 ;
  assign n41274 = n41273 ^ n18606 ^ 1'b0 ;
  assign n41275 = n22129 | n41274 ;
  assign n41276 = n12455 & ~n13810 ;
  assign n41277 = n35892 & ~n41276 ;
  assign n41278 = ~n33225 & n41277 ;
  assign n41279 = n40640 ^ n6871 ^ 1'b0 ;
  assign n41280 = n40960 & n41279 ;
  assign n41281 = n19579 ^ n19458 ^ 1'b0 ;
  assign n41282 = n618 & ~n41281 ;
  assign n41283 = n23840 ^ n7404 ^ 1'b0 ;
  assign n41284 = n6672 & n29103 ;
  assign n41285 = n32247 ^ n31972 ^ 1'b0 ;
  assign n41286 = n25713 & ~n41285 ;
  assign n41287 = ( n12753 & ~n21379 ) | ( n12753 & n29443 ) | ( ~n21379 & n29443 ) ;
  assign n41288 = ~n10065 & n19281 ;
  assign n41289 = n18214 & n41288 ;
  assign n41290 = n41287 & n41289 ;
  assign n41291 = n13495 | n28250 ;
  assign n41295 = ( n3545 & n5799 ) | ( n3545 & n20686 ) | ( n5799 & n20686 ) ;
  assign n41292 = n32343 ^ n28894 ^ n17371 ;
  assign n41293 = n41292 ^ n28006 ^ 1'b0 ;
  assign n41294 = n17580 & n41293 ;
  assign n41296 = n41295 ^ n41294 ^ 1'b0 ;
  assign n41297 = n2236 & ~n12925 ;
  assign n41298 = n31213 ^ n477 ^ 1'b0 ;
  assign n41299 = n7121 | n41298 ;
  assign n41300 = n12507 | n18642 ;
  assign n41301 = ( n36047 & ~n41299 ) | ( n36047 & n41300 ) | ( ~n41299 & n41300 ) ;
  assign n41302 = ~n3992 & n25850 ;
  assign n41303 = ~n37786 & n41302 ;
  assign n41304 = n41303 ^ n30144 ^ 1'b0 ;
  assign n41305 = n20904 & ~n41109 ;
  assign n41306 = n39915 ^ n32848 ^ 1'b0 ;
  assign n41307 = n21519 & ~n41306 ;
  assign n41308 = ~n6347 & n7726 ;
  assign n41309 = ~n14578 & n41308 ;
  assign n41310 = n41309 ^ n4052 ^ 1'b0 ;
  assign n41311 = n12893 & ~n41310 ;
  assign n41312 = n41311 ^ n6399 ^ 1'b0 ;
  assign n41313 = n17647 ^ n8551 ^ n826 ;
  assign n41314 = n5615 | n17662 ;
  assign n41315 = ( n8569 & n41313 ) | ( n8569 & ~n41314 ) | ( n41313 & ~n41314 ) ;
  assign n41316 = n13289 ^ n7410 ^ 1'b0 ;
  assign n41317 = n25302 ^ n17643 ^ n1347 ;
  assign n41318 = n10114 & ~n13321 ;
  assign n41319 = n41318 ^ n15279 ^ 1'b0 ;
  assign n41320 = n21584 | n37020 ;
  assign n41321 = n41320 ^ n6924 ^ 1'b0 ;
  assign n41322 = n28179 ^ n11304 ^ 1'b0 ;
  assign n41323 = n41322 ^ n38220 ^ 1'b0 ;
  assign n41324 = ~n38103 & n41323 ;
  assign n41326 = ( ~n1489 & n7957 ) | ( ~n1489 & n15281 ) | ( n7957 & n15281 ) ;
  assign n41325 = n12447 & ~n12507 ;
  assign n41327 = n41326 ^ n41325 ^ 1'b0 ;
  assign n41328 = n11872 | n41327 ;
  assign n41329 = n28879 & ~n41328 ;
  assign n41330 = ( n1508 & ~n8303 ) | ( n1508 & n28440 ) | ( ~n8303 & n28440 ) ;
  assign n41331 = n12121 & n41330 ;
  assign n41332 = ( n1538 & n3818 ) | ( n1538 & n17200 ) | ( n3818 & n17200 ) ;
  assign n41333 = ( n25617 & ~n35940 ) | ( n25617 & n41332 ) | ( ~n35940 & n41332 ) ;
  assign n41334 = n1181 & ~n1787 ;
  assign n41337 = n13316 | n34265 ;
  assign n41338 = n4350 & ~n41337 ;
  assign n41335 = n17201 & n23825 ;
  assign n41336 = n41335 ^ n7222 ^ 1'b0 ;
  assign n41339 = n41338 ^ n41336 ^ n4886 ;
  assign n41340 = ( n8984 & n18666 ) | ( n8984 & n41339 ) | ( n18666 & n41339 ) ;
  assign n41341 = n9814 | n36049 ;
  assign n41342 = n41341 ^ n34480 ^ 1'b0 ;
  assign n41344 = n14148 ^ n1118 ^ 1'b0 ;
  assign n41343 = n7805 & n31520 ;
  assign n41345 = n41344 ^ n41343 ^ 1'b0 ;
  assign n41350 = n32245 ^ n3713 ^ 1'b0 ;
  assign n41346 = n32953 ^ n7154 ^ n3087 ;
  assign n41347 = n41346 ^ n2476 ^ 1'b0 ;
  assign n41348 = n5299 & n41347 ;
  assign n41349 = n31076 & n41348 ;
  assign n41351 = n41350 ^ n41349 ^ n17198 ;
  assign n41352 = ( ~n23901 & n31726 ) | ( ~n23901 & n37286 ) | ( n31726 & n37286 ) ;
  assign n41354 = n1643 | n22688 ;
  assign n41355 = n41354 ^ n537 ^ 1'b0 ;
  assign n41353 = n34645 ^ n4688 ^ 1'b0 ;
  assign n41356 = n41355 ^ n41353 ^ n9489 ;
  assign n41357 = n40224 ^ n32814 ^ 1'b0 ;
  assign n41358 = n28380 ^ n21049 ^ 1'b0 ;
  assign n41359 = n40647 | n41358 ;
  assign n41360 = n1430 ^ n790 ^ 1'b0 ;
  assign n41361 = ( n8671 & n8708 ) | ( n8671 & n9943 ) | ( n8708 & n9943 ) ;
  assign n41362 = n41361 ^ n27039 ^ 1'b0 ;
  assign n41363 = n41360 & ~n41362 ;
  assign n41364 = n3062 ^ n584 ^ 1'b0 ;
  assign n41365 = ( n3745 & n8904 ) | ( n3745 & ~n19640 ) | ( n8904 & ~n19640 ) ;
  assign n41366 = n41365 ^ n14565 ^ 1'b0 ;
  assign n41367 = n15855 ^ n5785 ^ 1'b0 ;
  assign n41368 = n4851 & ~n6340 ;
  assign n41369 = n41368 ^ n4281 ^ 1'b0 ;
  assign n41370 = n24597 & n41369 ;
  assign n41371 = n41370 ^ n7913 ^ n2714 ;
  assign n41372 = ( n5639 & n35649 ) | ( n5639 & ~n41371 ) | ( n35649 & ~n41371 ) ;
  assign n41373 = ( n7542 & n41367 ) | ( n7542 & n41372 ) | ( n41367 & n41372 ) ;
  assign n41374 = ( n2880 & ~n31234 ) | ( n2880 & n36130 ) | ( ~n31234 & n36130 ) ;
  assign n41375 = ( ~n626 & n4124 ) | ( ~n626 & n6468 ) | ( n4124 & n6468 ) ;
  assign n41376 = n41375 ^ n16042 ^ n6626 ;
  assign n41377 = ~n17349 & n21281 ;
  assign n41378 = n41377 ^ n40731 ^ 1'b0 ;
  assign n41379 = ( ~n11200 & n18120 ) | ( ~n11200 & n41378 ) | ( n18120 & n41378 ) ;
  assign n41380 = n4155 | n25848 ;
  assign n41381 = ( n6753 & n16412 ) | ( n6753 & n22453 ) | ( n16412 & n22453 ) ;
  assign n41382 = ( ~n16784 & n22272 ) | ( ~n16784 & n31777 ) | ( n22272 & n31777 ) ;
  assign n41383 = n15466 ^ n10482 ^ 1'b0 ;
  assign n41384 = n16070 & n41383 ;
  assign n41385 = n4946 & ~n7166 ;
  assign n41386 = ~n3324 & n41385 ;
  assign n41387 = n41386 ^ n13000 ^ 1'b0 ;
  assign n41388 = n41384 | n41387 ;
  assign n41389 = ~n26850 & n38460 ;
  assign n41390 = ~n15190 & n41389 ;
  assign n41391 = ( n6326 & n20486 ) | ( n6326 & ~n41390 ) | ( n20486 & ~n41390 ) ;
  assign n41392 = ~n12801 & n25541 ;
  assign n41393 = ~n9771 & n41392 ;
  assign n41394 = n41391 & ~n41393 ;
  assign n41395 = ( n29925 & ~n30235 ) | ( n29925 & n35113 ) | ( ~n30235 & n35113 ) ;
  assign n41396 = n24316 & ~n36760 ;
  assign n41397 = ~n40869 & n41396 ;
  assign n41398 = n9902 ^ n6615 ^ 1'b0 ;
  assign n41399 = n17485 & n41398 ;
  assign n41400 = n15835 ^ n4805 ^ x122 ;
  assign n41401 = n19363 ^ n16570 ^ n7475 ;
  assign n41402 = n15727 ^ n14091 ^ n13648 ;
  assign n41403 = n8325 & n31529 ;
  assign n41404 = ~n41402 & n41403 ;
  assign n41405 = ( n22592 & n33132 ) | ( n22592 & n41404 ) | ( n33132 & n41404 ) ;
  assign n41406 = n33973 ^ n13214 ^ 1'b0 ;
  assign n41409 = ~n774 & n14852 ;
  assign n41410 = n41409 ^ n37716 ^ 1'b0 ;
  assign n41407 = n37551 ^ n23910 ^ n9655 ;
  assign n41408 = n41407 ^ n34703 ^ 1'b0 ;
  assign n41411 = n41410 ^ n41408 ^ 1'b0 ;
  assign n41412 = n21489 ^ n13157 ^ 1'b0 ;
  assign n41413 = n29204 & n37524 ;
  assign n41414 = n481 & n9032 ;
  assign n41415 = n41414 ^ n22321 ^ 1'b0 ;
  assign n41416 = n20663 & n41415 ;
  assign n41417 = ( n5512 & n10834 ) | ( n5512 & n14652 ) | ( n10834 & n14652 ) ;
  assign n41420 = n40722 ^ n17047 ^ 1'b0 ;
  assign n41418 = n39441 ^ n11849 ^ n11075 ;
  assign n41419 = ~n9378 & n41418 ;
  assign n41421 = n41420 ^ n41419 ^ n25966 ;
  assign n41422 = n29064 ^ n19363 ^ 1'b0 ;
  assign n41423 = n3425 ^ x244 ^ 1'b0 ;
  assign n41424 = n1356 & n7192 ;
  assign n41425 = n29859 ^ n13689 ^ 1'b0 ;
  assign n41426 = ~n39593 & n41425 ;
  assign n41427 = n41426 ^ n22835 ^ 1'b0 ;
  assign n41428 = n33572 ^ n26885 ^ n5706 ;
  assign n41429 = n41428 ^ n37760 ^ 1'b0 ;
  assign n41430 = n3617 ^ n2705 ^ 1'b0 ;
  assign n41431 = n12830 | n41430 ;
  assign n41432 = ( ~n12433 & n34319 ) | ( ~n12433 & n37790 ) | ( n34319 & n37790 ) ;
  assign n41433 = n21082 & ~n25489 ;
  assign n41434 = ~n41432 & n41433 ;
  assign n41435 = ~n38652 & n40602 ;
  assign n41436 = n12472 & n24570 ;
  assign n41437 = n41436 ^ n6722 ^ 1'b0 ;
  assign n41438 = n41437 ^ n38149 ^ 1'b0 ;
  assign n41439 = n41173 ^ n36775 ^ n4473 ;
  assign n41440 = ( n2229 & n6770 ) | ( n2229 & n13963 ) | ( n6770 & n13963 ) ;
  assign n41441 = n41440 ^ n10461 ^ n10107 ;
  assign n41442 = n3666 & ~n13313 ;
  assign n41443 = n41442 ^ n34690 ^ 1'b0 ;
  assign n41444 = n41443 ^ n21225 ^ n962 ;
  assign n41445 = n35723 ^ n5415 ^ 1'b0 ;
  assign n41446 = ~n21666 & n41445 ;
  assign n41447 = n7795 ^ n5526 ^ n3285 ;
  assign n41448 = n41447 ^ n4826 ^ 1'b0 ;
  assign n41449 = n41448 ^ n24461 ^ 1'b0 ;
  assign n41450 = ( n4828 & ~n15670 ) | ( n4828 & n33752 ) | ( ~n15670 & n33752 ) ;
  assign n41451 = n41450 ^ n35562 ^ n28301 ;
  assign n41452 = ( n9299 & n20532 ) | ( n9299 & ~n30643 ) | ( n20532 & ~n30643 ) ;
  assign n41453 = n3569 & ~n15800 ;
  assign n41454 = ~n16841 & n41453 ;
  assign n41455 = n41454 ^ n10655 ^ 1'b0 ;
  assign n41456 = ( n20556 & n22083 ) | ( n20556 & n32761 ) | ( n22083 & n32761 ) ;
  assign n41457 = n9798 & ~n23039 ;
  assign n41458 = n41457 ^ n27239 ^ 1'b0 ;
  assign n41459 = ~n35396 & n41458 ;
  assign n41460 = n27127 ^ n20588 ^ n8364 ;
  assign n41461 = n41460 ^ n7296 ^ 1'b0 ;
  assign n41462 = ~n4749 & n41461 ;
  assign n41463 = n7020 | n23125 ;
  assign n41464 = n41463 ^ n24158 ^ 1'b0 ;
  assign n41465 = ( n7935 & ~n35613 ) | ( n7935 & n41464 ) | ( ~n35613 & n41464 ) ;
  assign n41466 = ( ~n5685 & n13398 ) | ( ~n5685 & n39748 ) | ( n13398 & n39748 ) ;
  assign n41467 = ( ~n23900 & n32159 ) | ( ~n23900 & n40187 ) | ( n32159 & n40187 ) ;
  assign n41468 = ~n4310 & n10002 ;
  assign n41471 = ~n14853 & n15682 ;
  assign n41469 = n27048 ^ n23419 ^ 1'b0 ;
  assign n41470 = n1589 & ~n41469 ;
  assign n41472 = n41471 ^ n41470 ^ n38380 ;
  assign n41473 = ~n5638 & n6940 ;
  assign n41474 = ( n15418 & n40431 ) | ( n15418 & ~n41473 ) | ( n40431 & ~n41473 ) ;
  assign n41475 = ~n17574 & n41474 ;
  assign n41476 = n25819 & n41475 ;
  assign n41477 = ( n1464 & ~n3765 ) | ( n1464 & n7682 ) | ( ~n3765 & n7682 ) ;
  assign n41478 = n1214 & n17848 ;
  assign n41479 = n41477 & n41478 ;
  assign n41480 = ~n30491 & n39681 ;
  assign n41481 = n41480 ^ n7395 ^ 1'b0 ;
  assign n41482 = n10563 ^ n8375 ^ 1'b0 ;
  assign n41483 = ~n31204 & n41482 ;
  assign n41487 = ( ~n12798 & n18505 ) | ( ~n12798 & n34251 ) | ( n18505 & n34251 ) ;
  assign n41484 = n7336 & ~n8971 ;
  assign n41485 = ( n9298 & n22188 ) | ( n9298 & ~n41484 ) | ( n22188 & ~n41484 ) ;
  assign n41486 = n6301 & ~n41485 ;
  assign n41488 = n41487 ^ n41486 ^ 1'b0 ;
  assign n41490 = ( n13024 & ~n13241 ) | ( n13024 & n24002 ) | ( ~n13241 & n24002 ) ;
  assign n41489 = ~n6394 & n17671 ;
  assign n41491 = n41490 ^ n41489 ^ 1'b0 ;
  assign n41492 = ( n5508 & n23910 ) | ( n5508 & n30231 ) | ( n23910 & n30231 ) ;
  assign n41494 = n14804 & n17614 ;
  assign n41493 = n10848 & ~n32456 ;
  assign n41495 = n41494 ^ n41493 ^ n9911 ;
  assign n41497 = n15405 ^ n14940 ^ 1'b0 ;
  assign n41496 = n4989 & ~n18667 ;
  assign n41498 = n41497 ^ n41496 ^ n27195 ;
  assign n41499 = n41498 ^ n2790 ^ 1'b0 ;
  assign n41500 = n31216 ^ n23371 ^ 1'b0 ;
  assign n41501 = n22817 & ~n41500 ;
  assign n41502 = ~n4045 & n34135 ;
  assign n41503 = ~n5265 & n41502 ;
  assign n41504 = n8797 & ~n21012 ;
  assign n41505 = n6038 & n41504 ;
  assign n41506 = n22339 | n41505 ;
  assign n41507 = n41503 & ~n41506 ;
  assign n41508 = n29280 | n41282 ;
  assign n41509 = n639 & ~n12570 ;
  assign n41510 = n13832 & n26956 ;
  assign n41511 = ~n26853 & n41510 ;
  assign n41512 = n21281 & ~n41511 ;
  assign n41513 = n41512 ^ n1375 ^ 1'b0 ;
  assign n41514 = n14116 ^ n6382 ^ n4351 ;
  assign n41515 = n19262 ^ n7693 ^ n1196 ;
  assign n41516 = n32632 ^ n30643 ^ n1527 ;
  assign n41517 = n18334 & ~n27110 ;
  assign n41518 = n2709 & n41517 ;
  assign n41519 = n30934 ^ n27276 ^ 1'b0 ;
  assign n41520 = n6228 | n41519 ;
  assign n41521 = n15968 ^ n10211 ^ n2087 ;
  assign n41522 = n41521 ^ n15607 ^ n7717 ;
  assign n41523 = n19289 | n41522 ;
  assign n41524 = ( n20285 & n23674 ) | ( n20285 & ~n25563 ) | ( n23674 & ~n25563 ) ;
  assign n41525 = n30845 ^ n8621 ^ n5146 ;
  assign n41526 = ( n18676 & n22799 ) | ( n18676 & n41525 ) | ( n22799 & n41525 ) ;
  assign n41527 = ~n9561 & n23332 ;
  assign n41528 = n18306 & ~n29460 ;
  assign n41529 = n41528 ^ n16117 ^ 1'b0 ;
  assign n41530 = ~n4253 & n10309 ;
  assign n41531 = n41530 ^ n14905 ^ 1'b0 ;
  assign n41532 = n1662 & n41531 ;
  assign n41533 = ~n24228 & n41532 ;
  assign n41534 = n2011 & n39372 ;
  assign n41535 = n34295 ^ n333 ^ 1'b0 ;
  assign n41536 = n1738 & n14764 ;
  assign n41537 = n15285 ^ x66 ^ 1'b0 ;
  assign n41538 = ( n39216 & n41536 ) | ( n39216 & ~n41537 ) | ( n41536 & ~n41537 ) ;
  assign n41539 = n12528 ^ n11503 ^ n7579 ;
  assign n41540 = n3271 & ~n11230 ;
  assign n41541 = ~n331 & n41540 ;
  assign n41542 = n22022 ^ n16200 ^ 1'b0 ;
  assign n41543 = ~n41541 & n41542 ;
  assign n41544 = ( n18355 & n41539 ) | ( n18355 & n41543 ) | ( n41539 & n41543 ) ;
  assign n41545 = n19571 ^ n12289 ^ 1'b0 ;
  assign n41546 = n41545 ^ n19124 ^ n11674 ;
  assign n41547 = n16193 & ~n21583 ;
  assign n41548 = ~n4384 & n29348 ;
  assign n41549 = n28772 & ~n41548 ;
  assign n41550 = n41549 ^ n30297 ^ 1'b0 ;
  assign n41551 = n26629 ^ n15653 ^ 1'b0 ;
  assign n41552 = n409 | n35710 ;
  assign n41553 = n20592 | n20606 ;
  assign n41554 = ( n18789 & n22717 ) | ( n18789 & n41553 ) | ( n22717 & n41553 ) ;
  assign n41555 = n41554 ^ n13548 ^ 1'b0 ;
  assign n41556 = ~n11440 & n41555 ;
  assign n41557 = n41556 ^ n14129 ^ 1'b0 ;
  assign n41558 = n7083 ^ n6490 ^ 1'b0 ;
  assign n41559 = n32258 | n40499 ;
  assign n41560 = ( n21807 & n41558 ) | ( n21807 & ~n41559 ) | ( n41558 & ~n41559 ) ;
  assign n41561 = n41557 | n41560 ;
  assign n41562 = n13039 ^ n12871 ^ 1'b0 ;
  assign n41563 = n11427 & n41562 ;
  assign n41564 = ~n24666 & n36896 ;
  assign n41565 = ( n20229 & n41563 ) | ( n20229 & ~n41564 ) | ( n41563 & ~n41564 ) ;
  assign n41566 = n31860 ^ n16330 ^ n15762 ;
  assign n41567 = n15172 | n34961 ;
  assign n41568 = n41567 ^ n7867 ^ n1354 ;
  assign n41569 = n3056 | n23703 ;
  assign n41570 = n8983 | n22982 ;
  assign n41571 = n41569 | n41570 ;
  assign n41572 = n13039 ^ n2153 ^ n1482 ;
  assign n41573 = ( n1989 & ~n18563 ) | ( n1989 & n34687 ) | ( ~n18563 & n34687 ) ;
  assign n41574 = n11747 & n20326 ;
  assign n41575 = n3483 | n30933 ;
  assign n41576 = n41574 | n41575 ;
  assign n41577 = n21171 ^ n1591 ^ 1'b0 ;
  assign n41578 = n4942 & ~n41577 ;
  assign n41579 = n15660 ^ n4008 ^ 1'b0 ;
  assign n41580 = n37031 & ~n41579 ;
  assign n41581 = ~n9787 & n33894 ;
  assign n41582 = ~n23814 & n41581 ;
  assign n41583 = ( ~n10623 & n30015 ) | ( ~n10623 & n41582 ) | ( n30015 & n41582 ) ;
  assign n41584 = n37318 ^ n13335 ^ 1'b0 ;
  assign n41585 = ~n11062 & n24027 ;
  assign n41586 = n41585 ^ n29064 ^ 1'b0 ;
  assign n41587 = n41586 ^ n23101 ^ 1'b0 ;
  assign n41588 = n7367 | n41587 ;
  assign n41589 = n12496 | n31861 ;
  assign n41590 = n26706 | n41589 ;
  assign n41591 = n41590 ^ n17813 ^ 1'b0 ;
  assign n41592 = ( ~n41584 & n41588 ) | ( ~n41584 & n41591 ) | ( n41588 & n41591 ) ;
  assign n41593 = n18375 & ~n32275 ;
  assign n41594 = n17252 ^ n12722 ^ n9540 ;
  assign n41595 = n26839 ^ n6374 ^ 1'b0 ;
  assign n41596 = ( n20940 & n38852 ) | ( n20940 & ~n40665 ) | ( n38852 & ~n40665 ) ;
  assign n41597 = n16481 & ~n41596 ;
  assign n41598 = ~n4868 & n9103 ;
  assign n41599 = n41598 ^ n19419 ^ 1'b0 ;
  assign n41600 = n20305 & ~n41599 ;
  assign n41601 = n41600 ^ n2347 ^ 1'b0 ;
  assign n41602 = n36993 ^ n33055 ^ 1'b0 ;
  assign n41603 = n1018 & ~n41056 ;
  assign n41604 = n41603 ^ n32721 ^ 1'b0 ;
  assign n41605 = n4828 | n12446 ;
  assign n41606 = n29007 & ~n41605 ;
  assign n41607 = n26198 ^ n20303 ^ 1'b0 ;
  assign n41608 = n41607 ^ n25559 ^ n6296 ;
  assign n41612 = ( n2917 & ~n8156 ) | ( n2917 & n8423 ) | ( ~n8156 & n8423 ) ;
  assign n41609 = n6115 & ~n15864 ;
  assign n41610 = ~n593 & n41609 ;
  assign n41611 = n41610 ^ n13742 ^ 1'b0 ;
  assign n41613 = n41612 ^ n41611 ^ n15410 ;
  assign n41614 = n41613 ^ n35309 ^ n17672 ;
  assign n41615 = n10290 | n36534 ;
  assign n41616 = n23474 ^ n14683 ^ 1'b0 ;
  assign n41617 = n35476 | n41616 ;
  assign n41618 = ~n24280 & n24951 ;
  assign n41619 = ~n4182 & n41618 ;
  assign n41621 = ( n4968 & n11185 ) | ( n4968 & ~n27679 ) | ( n11185 & ~n27679 ) ;
  assign n41620 = n799 | n24335 ;
  assign n41622 = n41621 ^ n41620 ^ 1'b0 ;
  assign n41623 = n32991 | n33427 ;
  assign n41624 = n9398 & n41623 ;
  assign n41625 = n30930 ^ n9385 ^ 1'b0 ;
  assign n41626 = n24430 | n41625 ;
  assign n41627 = n14929 | n41626 ;
  assign n41628 = n41627 ^ n9218 ^ 1'b0 ;
  assign n41629 = n26187 ^ n15283 ^ 1'b0 ;
  assign n41630 = ~n3330 & n41629 ;
  assign n41631 = ( n9633 & ~n16208 ) | ( n9633 & n29087 ) | ( ~n16208 & n29087 ) ;
  assign n41632 = n41631 ^ n34589 ^ n13886 ;
  assign n41633 = n41632 ^ n20504 ^ n506 ;
  assign n41634 = n6312 & n16823 ;
  assign n41635 = ~n31938 & n41634 ;
  assign n41636 = ( n7935 & n9651 ) | ( n7935 & ~n18896 ) | ( n9651 & ~n18896 ) ;
  assign n41637 = ~n13791 & n41636 ;
  assign n41638 = ( n6641 & n19643 ) | ( n6641 & ~n41637 ) | ( n19643 & ~n41637 ) ;
  assign n41639 = n8027 | n9448 ;
  assign n41640 = n41639 ^ n26882 ^ 1'b0 ;
  assign n41641 = n14109 ^ n9334 ^ 1'b0 ;
  assign n41642 = n38875 ^ n6411 ^ x99 ;
  assign n41643 = n12030 & ~n41642 ;
  assign n41644 = n16387 & n17237 ;
  assign n41645 = n41644 ^ n32238 ^ 1'b0 ;
  assign n41646 = n35474 ^ n12884 ^ 1'b0 ;
  assign n41647 = n41645 | n41646 ;
  assign n41648 = n24417 ^ n2076 ^ 1'b0 ;
  assign n41649 = ~n9700 & n15183 ;
  assign n41650 = n41649 ^ n21519 ^ n3846 ;
  assign n41651 = n32927 ^ n21871 ^ n11062 ;
  assign n41652 = ~n6541 & n9960 ;
  assign n41653 = ~n33419 & n41652 ;
  assign n41654 = ~n17796 & n17861 ;
  assign n41655 = n41654 ^ n33644 ^ 1'b0 ;
  assign n41656 = n1120 | n29372 ;
  assign n41657 = n20595 & ~n41656 ;
  assign n41658 = ( n11741 & ~n31834 ) | ( n11741 & n34839 ) | ( ~n31834 & n34839 ) ;
  assign n41659 = n4095 & ~n18101 ;
  assign n41661 = n14764 ^ n13175 ^ 1'b0 ;
  assign n41662 = n29535 & ~n41661 ;
  assign n41660 = n9570 | n21248 ;
  assign n41663 = n41662 ^ n41660 ^ 1'b0 ;
  assign n41666 = n2305 | n41017 ;
  assign n41667 = n41666 ^ n21617 ^ 1'b0 ;
  assign n41664 = ~n13579 & n18083 ;
  assign n41665 = n36551 & ~n41664 ;
  assign n41668 = n41667 ^ n41665 ^ 1'b0 ;
  assign n41670 = n3782 | n39195 ;
  assign n41669 = ~n9587 & n31404 ;
  assign n41671 = n41670 ^ n41669 ^ 1'b0 ;
  assign n41673 = n36721 ^ n10709 ^ 1'b0 ;
  assign n41674 = n34081 & n41673 ;
  assign n41672 = n11866 ^ n3933 ^ n1786 ;
  assign n41675 = n41674 ^ n41672 ^ 1'b0 ;
  assign n41676 = n32397 ^ n8860 ^ 1'b0 ;
  assign n41677 = n40505 ^ n10498 ^ 1'b0 ;
  assign n41678 = ~n41676 & n41677 ;
  assign n41679 = n41678 ^ n28304 ^ n27825 ;
  assign n41680 = ( n12434 & n21555 ) | ( n12434 & n31049 ) | ( n21555 & n31049 ) ;
  assign n41681 = n34533 ^ n9509 ^ n6553 ;
  assign n41682 = ( n5251 & ~n7160 ) | ( n5251 & n19097 ) | ( ~n7160 & n19097 ) ;
  assign n41683 = n41682 ^ n9522 ^ 1'b0 ;
  assign n41684 = n30240 & ~n41683 ;
  assign n41686 = n23494 ^ n15155 ^ 1'b0 ;
  assign n41687 = n24401 | n41686 ;
  assign n41688 = n41687 ^ n27275 ^ n7215 ;
  assign n41685 = ~n14656 & n40321 ;
  assign n41689 = n41688 ^ n41685 ^ 1'b0 ;
  assign n41690 = ~n543 & n33522 ;
  assign n41691 = n41690 ^ n32568 ^ 1'b0 ;
  assign n41692 = ~n11285 & n11766 ;
  assign n41693 = n41692 ^ n28907 ^ 1'b0 ;
  assign n41694 = n41693 ^ n37738 ^ n17648 ;
  assign n41695 = ( n4335 & ~n6413 ) | ( n4335 & n41694 ) | ( ~n6413 & n41694 ) ;
  assign n41696 = ( n22117 & n24558 ) | ( n22117 & ~n31779 ) | ( n24558 & ~n31779 ) ;
  assign n41697 = n40317 ^ n33656 ^ 1'b0 ;
  assign n41698 = n40848 ^ n14401 ^ n13561 ;
  assign n41699 = ( ~n18917 & n19676 ) | ( ~n18917 & n41698 ) | ( n19676 & n41698 ) ;
  assign n41700 = n41699 ^ n36169 ^ n30939 ;
  assign n41701 = ~n6617 & n19176 ;
  assign n41702 = ~n1787 & n24570 ;
  assign n41703 = n26152 | n31129 ;
  assign n41704 = n41702 | n41703 ;
  assign n41705 = n23682 ^ n21751 ^ 1'b0 ;
  assign n41706 = n4819 & n41705 ;
  assign n41707 = ( ~n14932 & n15269 ) | ( ~n14932 & n15673 ) | ( n15269 & n15673 ) ;
  assign n41708 = n22238 | n41707 ;
  assign n41709 = ( n1984 & n14762 ) | ( n1984 & ~n30413 ) | ( n14762 & ~n30413 ) ;
  assign n41710 = ~n32727 & n41709 ;
  assign n41711 = ( n1695 & ~n6869 ) | ( n1695 & n7152 ) | ( ~n6869 & n7152 ) ;
  assign n41712 = ( n6397 & n10173 ) | ( n6397 & n41711 ) | ( n10173 & n41711 ) ;
  assign n41713 = n38550 ^ n14473 ^ 1'b0 ;
  assign n41714 = ~n7963 & n41713 ;
  assign n41715 = ( n6282 & ~n41712 ) | ( n6282 & n41714 ) | ( ~n41712 & n41714 ) ;
  assign n41716 = n40241 ^ n16650 ^ 1'b0 ;
  assign n41717 = ( ~n14401 & n28286 ) | ( ~n14401 & n30521 ) | ( n28286 & n30521 ) ;
  assign n41718 = n41717 ^ n15986 ^ 1'b0 ;
  assign n41719 = n16413 ^ n8056 ^ n1986 ;
  assign n41720 = n13431 ^ n4763 ^ 1'b0 ;
  assign n41721 = n8408 ^ n7163 ^ n813 ;
  assign n41722 = n1566 & n41721 ;
  assign n41723 = n41720 & n41722 ;
  assign n41724 = ~n27429 & n41723 ;
  assign n41725 = n31640 | n34118 ;
  assign n41726 = n41725 ^ n31704 ^ 1'b0 ;
  assign n41727 = n12140 ^ n6038 ^ 1'b0 ;
  assign n41728 = n1192 & n41727 ;
  assign n41729 = n36047 ^ n2019 ^ 1'b0 ;
  assign n41730 = ( n18810 & ~n20747 ) | ( n18810 & n36799 ) | ( ~n20747 & n36799 ) ;
  assign n41731 = ( n7790 & n21544 ) | ( n7790 & ~n23470 ) | ( n21544 & ~n23470 ) ;
  assign n41732 = n3752 & ~n6178 ;
  assign n41733 = n18029 & n28018 ;
  assign n41734 = ~n10071 & n41733 ;
  assign n41735 = ~n1346 & n18888 ;
  assign n41736 = n19910 ^ n9030 ^ 1'b0 ;
  assign n41737 = n15128 | n20526 ;
  assign n41738 = n41737 ^ n6213 ^ 1'b0 ;
  assign n41739 = n41738 ^ n39932 ^ n38473 ;
  assign n41740 = ( n27936 & n31722 ) | ( n27936 & ~n34890 ) | ( n31722 & ~n34890 ) ;
  assign n41741 = n12963 & n20907 ;
  assign n41742 = n41741 ^ n1348 ^ 1'b0 ;
  assign n41743 = n18305 & ~n41742 ;
  assign n41744 = n13643 & ~n19831 ;
  assign n41745 = n41744 ^ n18403 ^ 1'b0 ;
  assign n41746 = ~n11440 & n20765 ;
  assign n41747 = ~n41745 & n41746 ;
  assign n41748 = n7216 & ~n9615 ;
  assign n41749 = n23676 & n41748 ;
  assign n41750 = n4349 & ~n41749 ;
  assign n41751 = n41750 ^ n18029 ^ 1'b0 ;
  assign n41752 = n38038 ^ n25016 ^ n21327 ;
  assign n41753 = n41751 | n41752 ;
  assign n41754 = n13039 | n41753 ;
  assign n41755 = n39768 ^ n9856 ^ 1'b0 ;
  assign n41756 = n41006 | n41755 ;
  assign n41757 = n8622 | n21488 ;
  assign n41758 = ~n3704 & n5367 ;
  assign n41759 = ( n25917 & n40304 ) | ( n25917 & n41758 ) | ( n40304 & n41758 ) ;
  assign n41760 = n38942 ^ n7733 ^ 1'b0 ;
  assign n41761 = n37343 ^ n10588 ^ n9087 ;
  assign n41762 = n41761 ^ n33722 ^ n7707 ;
  assign n41764 = ( n326 & n3980 ) | ( n326 & ~n20888 ) | ( n3980 & ~n20888 ) ;
  assign n41763 = n12540 & ~n17788 ;
  assign n41765 = n41764 ^ n41763 ^ 1'b0 ;
  assign n41766 = n34341 ^ n28599 ^ n14932 ;
  assign n41767 = n568 & n10623 ;
  assign n41768 = n41767 ^ n259 ^ 1'b0 ;
  assign n41769 = n41768 ^ n4219 ^ 1'b0 ;
  assign n41770 = n41766 & n41769 ;
  assign n41771 = ( ~n6423 & n10542 ) | ( ~n6423 & n38008 ) | ( n10542 & n38008 ) ;
  assign n41772 = ( n19665 & ~n20206 ) | ( n19665 & n41771 ) | ( ~n20206 & n41771 ) ;
  assign n41773 = ( ~n12092 & n19322 ) | ( ~n12092 & n25882 ) | ( n19322 & n25882 ) ;
  assign n41774 = ( n4102 & n8705 ) | ( n4102 & ~n27249 ) | ( n8705 & ~n27249 ) ;
  assign n41775 = ( n32908 & ~n41773 ) | ( n32908 & n41774 ) | ( ~n41773 & n41774 ) ;
  assign n41777 = n8108 | n22799 ;
  assign n41778 = n41777 ^ n7870 ^ 1'b0 ;
  assign n41776 = n3898 | n5334 ;
  assign n41779 = n41778 ^ n41776 ^ 1'b0 ;
  assign n41780 = n29474 ^ n29071 ^ n7208 ;
  assign n41781 = n37950 ^ n27985 ^ 1'b0 ;
  assign n41782 = n7604 & ~n41781 ;
  assign n41783 = ~n5876 & n39402 ;
  assign n41785 = n2423 & n5066 ;
  assign n41786 = n41785 ^ n14607 ^ 1'b0 ;
  assign n41784 = n32946 & n34686 ;
  assign n41787 = n41786 ^ n41784 ^ 1'b0 ;
  assign n41788 = n1879 | n14639 ;
  assign n41789 = n21114 | n41788 ;
  assign n41790 = n41789 ^ n26408 ^ n21148 ;
  assign n41793 = ( n5803 & n10644 ) | ( n5803 & ~n24086 ) | ( n10644 & ~n24086 ) ;
  assign n41792 = ( ~n2985 & n4375 ) | ( ~n2985 & n12524 ) | ( n4375 & n12524 ) ;
  assign n41791 = n23953 & n24694 ;
  assign n41794 = n41793 ^ n41792 ^ n41791 ;
  assign n41795 = ( n20897 & n28320 ) | ( n20897 & n33647 ) | ( n28320 & n33647 ) ;
  assign n41796 = ( ~n4924 & n10389 ) | ( ~n4924 & n22550 ) | ( n10389 & n22550 ) ;
  assign n41797 = n13051 | n25867 ;
  assign n41798 = n22602 | n41797 ;
  assign n41799 = ( n5057 & ~n31587 ) | ( n5057 & n41798 ) | ( ~n31587 & n41798 ) ;
  assign n41800 = n3209 & ~n19233 ;
  assign n41801 = n41800 ^ n1074 ^ 1'b0 ;
  assign n41802 = n19861 & n41801 ;
  assign n41803 = ~n2365 & n41802 ;
  assign n41804 = n6204 & n8568 ;
  assign n41805 = n41803 & n41804 ;
  assign n41806 = n27037 ^ n1475 ^ n1380 ;
  assign n41807 = ~n33889 & n41806 ;
  assign n41808 = ( n1624 & n7792 ) | ( n1624 & n35532 ) | ( n7792 & n35532 ) ;
  assign n41809 = n4376 & ~n10048 ;
  assign n41810 = ~n7388 & n41809 ;
  assign n41811 = n41810 ^ n34303 ^ 1'b0 ;
  assign n41812 = n1682 & n30673 ;
  assign n41813 = ( n5510 & n23610 ) | ( n5510 & n35775 ) | ( n23610 & n35775 ) ;
  assign n41814 = n33956 ^ n28175 ^ 1'b0 ;
  assign n41815 = n24659 & n41814 ;
  assign n41816 = n1354 & n41815 ;
  assign n41817 = ~n41813 & n41816 ;
  assign n41818 = ~n3042 & n39892 ;
  assign n41819 = ~n39036 & n41818 ;
  assign n41820 = n21707 ^ n11760 ^ n10777 ;
  assign n41821 = n6722 | n41820 ;
  assign n41822 = n8964 & ~n41821 ;
  assign n41824 = n2960 ^ n992 ^ 1'b0 ;
  assign n41823 = n36374 ^ n31339 ^ 1'b0 ;
  assign n41825 = n41824 ^ n41823 ^ n25044 ;
  assign n41826 = n2704 | n12277 ;
  assign n41827 = ( n329 & ~n1018 ) | ( n329 & n3757 ) | ( ~n1018 & n3757 ) ;
  assign n41828 = n41827 ^ n27758 ^ 1'b0 ;
  assign n41829 = ~n14742 & n41828 ;
  assign n41830 = ( n1538 & n12775 ) | ( n1538 & ~n41829 ) | ( n12775 & ~n41829 ) ;
  assign n41831 = ( n8709 & n12598 ) | ( n8709 & n23105 ) | ( n12598 & n23105 ) ;
  assign n41832 = n3878 & n24996 ;
  assign n41833 = n19999 & ~n41832 ;
  assign n41834 = n12507 ^ n11787 ^ 1'b0 ;
  assign n41835 = n18778 & n41834 ;
  assign n41836 = ~n3055 & n41835 ;
  assign n41837 = n4401 & n29181 ;
  assign n41838 = n23478 | n28336 ;
  assign n41839 = n41838 ^ n11954 ^ 1'b0 ;
  assign n41840 = ( n4666 & ~n29795 ) | ( n4666 & n41758 ) | ( ~n29795 & n41758 ) ;
  assign n41841 = ~n5678 & n14640 ;
  assign n41842 = n41841 ^ n16697 ^ 1'b0 ;
  assign n41843 = ( n7145 & n24499 ) | ( n7145 & ~n41842 ) | ( n24499 & ~n41842 ) ;
  assign n41844 = n41843 ^ n31899 ^ n24126 ;
  assign n41845 = ( n28011 & n41840 ) | ( n28011 & n41844 ) | ( n41840 & n41844 ) ;
  assign n41846 = n10281 & ~n14614 ;
  assign n41847 = n5880 | n41846 ;
  assign n41848 = n12135 & ~n41847 ;
  assign n41849 = n14873 ^ n7993 ^ n2712 ;
  assign n41850 = ( n12107 & ~n39360 ) | ( n12107 & n41849 ) | ( ~n39360 & n41849 ) ;
  assign n41851 = n3829 & n41850 ;
  assign n41852 = n10844 & n41851 ;
  assign n41853 = n21554 & n30305 ;
  assign n41854 = n707 | n19275 ;
  assign n41855 = n22812 ^ n15867 ^ 1'b0 ;
  assign n41856 = n29910 ^ n23402 ^ n22518 ;
  assign n41857 = n3651 & n18862 ;
  assign n41858 = n41857 ^ n10570 ^ 1'b0 ;
  assign n41859 = n37091 ^ n9790 ^ 1'b0 ;
  assign n41860 = n1422 & n23957 ;
  assign n41861 = n37111 ^ n30392 ^ n6723 ;
  assign n41862 = n41761 ^ n5294 ^ x154 ;
  assign n41863 = n40982 ^ n31107 ^ x174 ;
  assign n41864 = n31896 & n38406 ;
  assign n41865 = n11013 | n12807 ;
  assign n41866 = n20209 ^ n17325 ^ 1'b0 ;
  assign n41867 = n41865 | n41866 ;
  assign n41868 = n41867 ^ n36687 ^ 1'b0 ;
  assign n41869 = n3320 & ~n7806 ;
  assign n41870 = n3290 & ~n41869 ;
  assign n41871 = n18090 & n41870 ;
  assign n41872 = n37981 ^ n1287 ^ 1'b0 ;
  assign n41873 = n36565 & n41872 ;
  assign n41874 = n480 | n16982 ;
  assign n41875 = n27557 & n41874 ;
  assign n41876 = n13430 & n35664 ;
  assign n41877 = n1099 & ~n5177 ;
  assign n41879 = ~n789 & n22595 ;
  assign n41880 = n41879 ^ n7449 ^ 1'b0 ;
  assign n41881 = n6315 ^ n2252 ^ 1'b0 ;
  assign n41882 = n41880 & ~n41881 ;
  assign n41878 = n18497 ^ n7889 ^ 1'b0 ;
  assign n41883 = n41882 ^ n41878 ^ n15579 ;
  assign n41884 = n6058 & n22888 ;
  assign n41885 = ~n7211 & n41884 ;
  assign n41886 = n3712 & ~n21238 ;
  assign n41887 = n9024 & n41886 ;
  assign n41888 = n7801 & ~n41887 ;
  assign n41889 = n41888 ^ n24702 ^ 1'b0 ;
  assign n41890 = n28998 ^ n18929 ^ n4256 ;
  assign n41891 = n25783 ^ n3070 ^ n1882 ;
  assign n41892 = n26880 & n41891 ;
  assign n41893 = ( ~n2856 & n4102 ) | ( ~n2856 & n17803 ) | ( n4102 & n17803 ) ;
  assign n41894 = ( n9469 & n41892 ) | ( n9469 & n41893 ) | ( n41892 & n41893 ) ;
  assign n41895 = n1483 & n20733 ;
  assign n41896 = n41895 ^ n8191 ^ 1'b0 ;
  assign n41897 = n1318 & ~n18698 ;
  assign n41898 = n41896 & n41897 ;
  assign n41900 = n41269 ^ n3923 ^ n1475 ;
  assign n41899 = n19657 ^ n3765 ^ 1'b0 ;
  assign n41901 = n41900 ^ n41899 ^ 1'b0 ;
  assign n41902 = n35796 ^ n33674 ^ n6906 ;
  assign n41903 = ( n15123 & ~n24959 ) | ( n15123 & n38293 ) | ( ~n24959 & n38293 ) ;
  assign n41904 = ( n14443 & n30986 ) | ( n14443 & n37898 ) | ( n30986 & n37898 ) ;
  assign n41905 = ( ~n24446 & n26912 ) | ( ~n24446 & n41904 ) | ( n26912 & n41904 ) ;
  assign n41906 = n41905 ^ n16100 ^ n13059 ;
  assign n41907 = n1961 ^ n1822 ^ 1'b0 ;
  assign n41908 = n41907 ^ n30189 ^ 1'b0 ;
  assign n41909 = n13246 | n29409 ;
  assign n41910 = n41909 ^ n11532 ^ 1'b0 ;
  assign n41912 = n14691 | n19556 ;
  assign n41911 = n24397 ^ n11575 ^ n10223 ;
  assign n41913 = n41912 ^ n41911 ^ n4435 ;
  assign n41914 = n41910 & ~n41913 ;
  assign n41915 = n32306 ^ n13552 ^ n13382 ;
  assign n41916 = n41915 ^ n11302 ^ n7873 ;
  assign n41917 = n15623 | n41916 ;
  assign n41918 = n11784 ^ n1964 ^ 1'b0 ;
  assign n41919 = n28143 ^ x245 ^ x128 ;
  assign n41920 = n17607 & n41919 ;
  assign n41921 = n7382 & n29176 ;
  assign n41922 = n33912 ^ n3783 ^ 1'b0 ;
  assign n41923 = n12880 & ~n41922 ;
  assign n41925 = n37165 ^ n33822 ^ 1'b0 ;
  assign n41926 = n4488 & n41925 ;
  assign n41924 = n38420 ^ n3975 ^ 1'b0 ;
  assign n41927 = n41926 ^ n41924 ^ n38990 ;
  assign n41928 = ( n15136 & ~n16327 ) | ( n15136 & n20141 ) | ( ~n16327 & n20141 ) ;
  assign n41929 = n15828 ^ n8735 ^ 1'b0 ;
  assign n41932 = n18746 ^ n14073 ^ 1'b0 ;
  assign n41930 = n14885 ^ n8214 ^ 1'b0 ;
  assign n41931 = ~n21335 & n41930 ;
  assign n41933 = n41932 ^ n41931 ^ 1'b0 ;
  assign n41934 = n12803 & ~n36437 ;
  assign n41935 = ~n4932 & n41934 ;
  assign n41936 = n25205 ^ n16317 ^ n326 ;
  assign n41937 = n32453 ^ n17822 ^ n6235 ;
  assign n41938 = ( ~n26549 & n41936 ) | ( ~n26549 & n41937 ) | ( n41936 & n41937 ) ;
  assign n41939 = n2127 & n8835 ;
  assign n41940 = ( ~n374 & n17354 ) | ( ~n374 & n39233 ) | ( n17354 & n39233 ) ;
  assign n41941 = n17489 ^ n14749 ^ n9275 ;
  assign n41942 = n643 & n5313 ;
  assign n41943 = n41942 ^ n20204 ^ n9872 ;
  assign n41944 = n13428 ^ n12528 ^ 1'b0 ;
  assign n41945 = n41944 ^ n15929 ^ 1'b0 ;
  assign n41946 = ~n8396 & n41945 ;
  assign n41947 = n24338 ^ n23290 ^ 1'b0 ;
  assign n41948 = n18017 & ~n41947 ;
  assign n41949 = n16931 ^ n3162 ^ 1'b0 ;
  assign n41950 = n23458 | n27775 ;
  assign n41951 = ( n10443 & n24833 ) | ( n10443 & n41950 ) | ( n24833 & n41950 ) ;
  assign n41954 = ( ~x118 & n12823 ) | ( ~x118 & n15016 ) | ( n12823 & n15016 ) ;
  assign n41955 = n41954 ^ n12142 ^ 1'b0 ;
  assign n41953 = ( n5355 & n21976 ) | ( n5355 & ~n23063 ) | ( n21976 & ~n23063 ) ;
  assign n41952 = n23181 & n34544 ;
  assign n41956 = n41955 ^ n41953 ^ n41952 ;
  assign n41957 = ~n4036 & n6076 ;
  assign n41958 = n25512 | n29580 ;
  assign n41959 = n41957 & ~n41958 ;
  assign n41960 = ( n5466 & ~n20508 ) | ( n5466 & n41959 ) | ( ~n20508 & n41959 ) ;
  assign n41961 = ( n7360 & n35299 ) | ( n7360 & n41960 ) | ( n35299 & n41960 ) ;
  assign n41962 = ~n1444 & n22914 ;
  assign n41963 = n41962 ^ n6934 ^ 1'b0 ;
  assign n41964 = n41963 ^ n33647 ^ n25361 ;
  assign n41965 = n11574 ^ n6000 ^ n4450 ;
  assign n41966 = n8707 ^ n8651 ^ 1'b0 ;
  assign n41967 = ( n11637 & n34266 ) | ( n11637 & n41966 ) | ( n34266 & n41966 ) ;
  assign n41968 = ( n8373 & ~n41965 ) | ( n8373 & n41967 ) | ( ~n41965 & n41967 ) ;
  assign n41969 = n9015 ^ n5712 ^ 1'b0 ;
  assign n41970 = n37343 & ~n41969 ;
  assign n41971 = ( n40109 & n41968 ) | ( n40109 & n41970 ) | ( n41968 & n41970 ) ;
  assign n41972 = n13165 & ~n34458 ;
  assign n41973 = n41972 ^ n29325 ^ 1'b0 ;
  assign n41974 = ( n22042 & ~n22662 ) | ( n22042 & n28695 ) | ( ~n22662 & n28695 ) ;
  assign n41975 = ( n10002 & ~n19518 ) | ( n10002 & n41974 ) | ( ~n19518 & n41974 ) ;
  assign n41976 = n10201 & ~n41975 ;
  assign n41977 = n3112 & n26300 ;
  assign n41978 = n14821 ^ n13149 ^ n8701 ;
  assign n41979 = ~n13670 & n41978 ;
  assign n41980 = ~n6087 & n41979 ;
  assign n41981 = n2936 | n3348 ;
  assign n41982 = n2389 | n16860 ;
  assign n41983 = n41982 ^ n3802 ^ 1'b0 ;
  assign n41984 = n41981 & ~n41983 ;
  assign n41985 = ~n2211 & n41984 ;
  assign n41987 = n5082 & n6630 ;
  assign n41988 = n41987 ^ n16234 ^ 1'b0 ;
  assign n41986 = n6780 | n25191 ;
  assign n41989 = n41988 ^ n41986 ^ 1'b0 ;
  assign n41990 = n34990 & n41989 ;
  assign n41991 = n1808 & n22208 ;
  assign n41992 = n41991 ^ n30286 ^ 1'b0 ;
  assign n41993 = n41992 ^ n33117 ^ n15899 ;
  assign n41994 = ( n21353 & n31148 ) | ( n21353 & ~n39104 ) | ( n31148 & ~n39104 ) ;
  assign n41995 = n22607 ^ n9250 ^ n4638 ;
  assign n41996 = n14279 ^ n2525 ^ 1'b0 ;
  assign n41997 = n20173 & ~n41996 ;
  assign n41998 = ( n11564 & n25645 ) | ( n11564 & ~n41997 ) | ( n25645 & ~n41997 ) ;
  assign n41999 = n11217 ^ n7135 ^ 1'b0 ;
  assign n42000 = n30856 | n41999 ;
  assign n42001 = n20103 & n22628 ;
  assign n42002 = n42000 & n42001 ;
  assign n42003 = ~n7207 & n25657 ;
  assign n42004 = ~n31263 & n42003 ;
  assign n42005 = n8386 & n12489 ;
  assign n42006 = n21967 & n42005 ;
  assign n42007 = n21497 | n42006 ;
  assign n42008 = n32043 ^ n10759 ^ 1'b0 ;
  assign n42009 = n14086 & n42008 ;
  assign n42010 = ( n11306 & n13051 ) | ( n11306 & n42009 ) | ( n13051 & n42009 ) ;
  assign n42011 = n19632 ^ n4548 ^ 1'b0 ;
  assign n42012 = n42011 ^ n33726 ^ n13591 ;
  assign n42013 = ( n2858 & n17105 ) | ( n2858 & n29195 ) | ( n17105 & n29195 ) ;
  assign n42014 = n25228 ^ n24085 ^ n4747 ;
  assign n42015 = n5931 & ~n7770 ;
  assign n42016 = n5524 | n32971 ;
  assign n42017 = n42015 | n42016 ;
  assign n42018 = n42017 ^ n41558 ^ n30167 ;
  assign n42019 = ~n42014 & n42018 ;
  assign n42020 = n15281 ^ n6930 ^ 1'b0 ;
  assign n42021 = n3208 | n33670 ;
  assign n42022 = n28208 & n42021 ;
  assign n42023 = ~n42020 & n42022 ;
  assign n42024 = n42023 ^ n22156 ^ 1'b0 ;
  assign n42025 = n1828 & n42024 ;
  assign n42026 = n5857 & n13791 ;
  assign n42027 = n7112 | n17669 ;
  assign n42028 = ( n32220 & n42026 ) | ( n32220 & ~n42027 ) | ( n42026 & ~n42027 ) ;
  assign n42029 = n20069 ^ n8519 ^ 1'b0 ;
  assign n42030 = n12937 | n42029 ;
  assign n42031 = ~n19994 & n42030 ;
  assign n42032 = n42031 ^ n34587 ^ n33367 ;
  assign n42033 = n867 | n6335 ;
  assign n42034 = ( n16547 & ~n31966 ) | ( n16547 & n38717 ) | ( ~n31966 & n38717 ) ;
  assign n42035 = ( n29969 & ~n35096 ) | ( n29969 & n42034 ) | ( ~n35096 & n42034 ) ;
  assign n42036 = n4715 ^ n757 ^ 1'b0 ;
  assign n42037 = n16330 | n42036 ;
  assign n42039 = ( ~n10307 & n32637 ) | ( ~n10307 & n34081 ) | ( n32637 & n34081 ) ;
  assign n42038 = ~n19676 & n38865 ;
  assign n42040 = n42039 ^ n42038 ^ 1'b0 ;
  assign n42041 = ~n34510 & n42040 ;
  assign n42042 = n42041 ^ n26890 ^ 1'b0 ;
  assign n42043 = n5183 & n41592 ;
  assign n42044 = n42043 ^ n9752 ^ 1'b0 ;
  assign n42045 = n800 & ~n9969 ;
  assign n42046 = n42045 ^ n4642 ^ 1'b0 ;
  assign n42047 = n42046 ^ n32807 ^ 1'b0 ;
  assign n42050 = n1279 | n9636 ;
  assign n42051 = n42050 ^ n26984 ^ n15254 ;
  assign n42048 = ~n3289 & n35979 ;
  assign n42049 = n39235 & ~n42048 ;
  assign n42052 = n42051 ^ n42049 ^ n6231 ;
  assign n42053 = n3109 & n22602 ;
  assign n42054 = n42053 ^ n21158 ^ 1'b0 ;
  assign n42055 = n42054 ^ n2073 ^ 1'b0 ;
  assign n42056 = n35302 ^ n11811 ^ n7981 ;
  assign n42058 = n14953 & ~n19570 ;
  assign n42059 = n42058 ^ n12737 ^ 1'b0 ;
  assign n42057 = n27533 ^ n10840 ^ 1'b0 ;
  assign n42060 = n42059 ^ n42057 ^ n2707 ;
  assign n42061 = n3688 & n6342 ;
  assign n42062 = ~n8606 & n42061 ;
  assign n42063 = ~n8919 & n42062 ;
  assign n42064 = n42063 ^ n27844 ^ 1'b0 ;
  assign n42065 = n28549 ^ n22259 ^ 1'b0 ;
  assign n42066 = n2251 & ~n42065 ;
  assign n42067 = n8088 ^ n3469 ^ 1'b0 ;
  assign n42068 = n17191 | n42067 ;
  assign n42069 = n42068 ^ n26792 ^ 1'b0 ;
  assign n42070 = n1475 | n29548 ;
  assign n42071 = n18559 & ~n42070 ;
  assign n42072 = n42071 ^ n33883 ^ n2074 ;
  assign n42073 = n16101 ^ n15361 ^ n2103 ;
  assign n42074 = x137 & n1867 ;
  assign n42075 = n1897 & ~n17433 ;
  assign n42076 = n42075 ^ n40822 ^ 1'b0 ;
  assign n42077 = n8122 & ~n42076 ;
  assign n42078 = n31485 ^ n17743 ^ 1'b0 ;
  assign n42079 = n23738 ^ n18773 ^ 1'b0 ;
  assign n42080 = n42078 & ~n42079 ;
  assign n42081 = ~n3617 & n12428 ;
  assign n42082 = n42081 ^ n13832 ^ 1'b0 ;
  assign n42083 = n9786 & ~n42082 ;
  assign n42084 = n5757 | n42083 ;
  assign n42085 = n3495 | n42084 ;
  assign n42086 = n40693 ^ n488 ^ 1'b0 ;
  assign n42087 = n5887 | n42086 ;
  assign n42088 = n33723 & ~n42087 ;
  assign n42089 = ( ~n30248 & n39389 ) | ( ~n30248 & n42088 ) | ( n39389 & n42088 ) ;
  assign n42090 = n28271 ^ n25256 ^ n14042 ;
  assign n42091 = ( ~n16847 & n35158 ) | ( ~n16847 & n42090 ) | ( n35158 & n42090 ) ;
  assign n42096 = n18071 ^ n6816 ^ n4086 ;
  assign n42097 = ( n22631 & ~n27086 ) | ( n22631 & n42096 ) | ( ~n27086 & n42096 ) ;
  assign n42098 = n42097 ^ n9137 ^ 1'b0 ;
  assign n42099 = ( n8840 & n35361 ) | ( n8840 & ~n42098 ) | ( n35361 & ~n42098 ) ;
  assign n42095 = ~n6384 & n30180 ;
  assign n42100 = n42099 ^ n42095 ^ 1'b0 ;
  assign n42092 = n32782 ^ n12631 ^ 1'b0 ;
  assign n42093 = n6048 & n42092 ;
  assign n42094 = n10042 & n42093 ;
  assign n42101 = n42100 ^ n42094 ^ 1'b0 ;
  assign n42102 = ~n11765 & n17703 ;
  assign n42103 = n42102 ^ n40790 ^ 1'b0 ;
  assign n42104 = n42103 ^ n5510 ^ 1'b0 ;
  assign n42105 = n23661 ^ n12230 ^ 1'b0 ;
  assign n42106 = n18252 | n42105 ;
  assign n42107 = n8754 ^ n5440 ^ 1'b0 ;
  assign n42108 = n42107 ^ n6265 ^ 1'b0 ;
  assign n42110 = ( n5062 & n17676 ) | ( n5062 & ~n22031 ) | ( n17676 & ~n22031 ) ;
  assign n42111 = ( n3168 & n14381 ) | ( n3168 & n42110 ) | ( n14381 & n42110 ) ;
  assign n42109 = n9256 & n21882 ;
  assign n42112 = n42111 ^ n42109 ^ 1'b0 ;
  assign n42113 = n20085 ^ n11937 ^ x221 ;
  assign n42114 = n20797 | n42113 ;
  assign n42115 = n14344 & ~n19415 ;
  assign n42116 = n42115 ^ n13154 ^ 1'b0 ;
  assign n42117 = ~n3498 & n42116 ;
  assign n42118 = n42117 ^ n20191 ^ 1'b0 ;
  assign n42119 = ( n1010 & n4793 ) | ( n1010 & n13394 ) | ( n4793 & n13394 ) ;
  assign n42120 = n42119 ^ n4552 ^ 1'b0 ;
  assign n42121 = ( n38129 & ~n42118 ) | ( n38129 & n42120 ) | ( ~n42118 & n42120 ) ;
  assign n42122 = n27800 ^ n12507 ^ n9972 ;
  assign n42123 = n42122 ^ n34266 ^ n17623 ;
  assign n42124 = ( ~n838 & n30886 ) | ( ~n838 & n42123 ) | ( n30886 & n42123 ) ;
  assign n42125 = n23611 ^ n1181 ^ 1'b0 ;
  assign n42126 = n42125 ^ n41768 ^ n23736 ;
  assign n42127 = ( x116 & n715 ) | ( x116 & n22888 ) | ( n715 & n22888 ) ;
  assign n42128 = n42127 ^ n39837 ^ n31587 ;
  assign n42129 = n42128 ^ n18640 ^ x67 ;
  assign n42131 = n7136 & n10963 ;
  assign n42130 = n22072 ^ n19306 ^ n12116 ;
  assign n42132 = n42131 ^ n42130 ^ n12622 ;
  assign n42133 = n10921 & n42132 ;
  assign n42134 = n42133 ^ n23898 ^ 1'b0 ;
  assign n42135 = n42134 ^ n20986 ^ 1'b0 ;
  assign n42136 = n23337 & n42135 ;
  assign n42137 = n19687 ^ n5850 ^ 1'b0 ;
  assign n42138 = n20986 & ~n42137 ;
  assign n42139 = n41052 ^ n7952 ^ n2220 ;
  assign n42140 = n35779 ^ n26474 ^ 1'b0 ;
  assign n42141 = n1579 | n42140 ;
  assign n42142 = n42141 ^ n19236 ^ n13534 ;
  assign n42143 = n2113 & n12602 ;
  assign n42144 = n20690 | n25564 ;
  assign n42145 = n42143 | n42144 ;
  assign n42146 = n42145 ^ n27993 ^ n11435 ;
  assign n42147 = ( n2711 & n34250 ) | ( n2711 & ~n42146 ) | ( n34250 & ~n42146 ) ;
  assign n42148 = ( n1016 & n4044 ) | ( n1016 & n22607 ) | ( n4044 & n22607 ) ;
  assign n42149 = n42148 ^ n39731 ^ n38663 ;
  assign n42150 = n32638 ^ n5581 ^ 1'b0 ;
  assign n42151 = n22649 | n42150 ;
  assign n42152 = n19174 ^ n1859 ^ 1'b0 ;
  assign n42153 = n11671 & ~n42152 ;
  assign n42154 = n4850 | n17354 ;
  assign n42155 = n42154 ^ n7538 ^ 1'b0 ;
  assign n42156 = n12446 ^ n12181 ^ 1'b0 ;
  assign n42157 = n8122 & ~n42156 ;
  assign n42158 = n24729 & n37474 ;
  assign n42159 = ( n34391 & ~n42157 ) | ( n34391 & n42158 ) | ( ~n42157 & n42158 ) ;
  assign n42160 = n1705 & ~n6081 ;
  assign n42161 = ( n1338 & n4757 ) | ( n1338 & n42160 ) | ( n4757 & n42160 ) ;
  assign n42162 = n17874 | n42161 ;
  assign n42163 = n1315 | n28620 ;
  assign n42164 = n18705 & n36191 ;
  assign n42165 = ~n37618 & n42164 ;
  assign n42166 = ~n13382 & n27029 ;
  assign n42167 = n42166 ^ n5671 ^ 1'b0 ;
  assign n42168 = n38805 ^ n17870 ^ 1'b0 ;
  assign n42169 = ( n1028 & n10829 ) | ( n1028 & n25759 ) | ( n10829 & n25759 ) ;
  assign n42170 = n42169 ^ n17846 ^ n2122 ;
  assign n42171 = ( n15906 & ~n19425 ) | ( n15906 & n42170 ) | ( ~n19425 & n42170 ) ;
  assign n42172 = n35836 | n36534 ;
  assign n42173 = n6438 & ~n17270 ;
  assign n42174 = n42173 ^ n35657 ^ n23738 ;
  assign n42175 = n14546 ^ n7788 ^ 1'b0 ;
  assign n42176 = ( ~n3030 & n10518 ) | ( ~n3030 & n10978 ) | ( n10518 & n10978 ) ;
  assign n42177 = ~n42175 & n42176 ;
  assign n42178 = n42177 ^ n21028 ^ 1'b0 ;
  assign n42179 = n3844 & ~n42178 ;
  assign n42180 = x135 & ~n17175 ;
  assign n42181 = n42180 ^ n15337 ^ 1'b0 ;
  assign n42182 = n23209 & n42181 ;
  assign n42183 = ~n20539 & n38699 ;
  assign n42184 = n42182 & n42183 ;
  assign n42185 = ~n37414 & n39039 ;
  assign n42186 = n34245 ^ n16691 ^ 1'b0 ;
  assign n42187 = n42185 & ~n42186 ;
  assign n42188 = n12096 | n34739 ;
  assign n42189 = n42188 ^ n27720 ^ 1'b0 ;
  assign n42190 = ( n3578 & n13826 ) | ( n3578 & n17986 ) | ( n13826 & n17986 ) ;
  assign n42191 = n42190 ^ n16291 ^ 1'b0 ;
  assign n42192 = n3859 & n42191 ;
  assign n42195 = ( n5757 & n14402 ) | ( n5757 & ~n22560 ) | ( n14402 & ~n22560 ) ;
  assign n42193 = ~n3361 & n9182 ;
  assign n42194 = n42193 ^ n13749 ^ n13133 ;
  assign n42196 = n42195 ^ n42194 ^ 1'b0 ;
  assign n42197 = n12801 ^ n9349 ^ 1'b0 ;
  assign n42198 = n42197 ^ n35940 ^ n5508 ;
  assign n42199 = n19984 & ~n20633 ;
  assign n42200 = n42199 ^ n1285 ^ 1'b0 ;
  assign n42201 = n33660 & ~n42200 ;
  assign n42202 = ~n42198 & n42201 ;
  assign n42203 = n42196 | n42202 ;
  assign n42204 = n6714 & n25418 ;
  assign n42205 = n42204 ^ n9702 ^ 1'b0 ;
  assign n42206 = n6804 & n42205 ;
  assign n42207 = ( ~n25382 & n27794 ) | ( ~n25382 & n28164 ) | ( n27794 & n28164 ) ;
  assign n42208 = ( n2540 & n42206 ) | ( n2540 & ~n42207 ) | ( n42206 & ~n42207 ) ;
  assign n42209 = n32368 ^ n5853 ^ 1'b0 ;
  assign n42210 = n11878 & ~n42209 ;
  assign n42211 = n40457 ^ n29891 ^ 1'b0 ;
  assign n42212 = n22675 ^ n18772 ^ 1'b0 ;
  assign n42213 = ~n15448 & n42212 ;
  assign n42214 = n21653 ^ n12356 ^ 1'b0 ;
  assign n42215 = n17371 & ~n42214 ;
  assign n42216 = n18913 & n42215 ;
  assign n42217 = n42216 ^ n22003 ^ 1'b0 ;
  assign n42218 = n5466 & ~n12003 ;
  assign n42219 = n9912 & n42218 ;
  assign n42220 = n10540 ^ n2841 ^ 1'b0 ;
  assign n42221 = ( ~n9246 & n23140 ) | ( ~n9246 & n37710 ) | ( n23140 & n37710 ) ;
  assign n42222 = ( n2795 & n42220 ) | ( n2795 & ~n42221 ) | ( n42220 & ~n42221 ) ;
  assign n42223 = n33947 & ~n36385 ;
  assign n42224 = ~n12101 & n17848 ;
  assign n42225 = n42224 ^ n23349 ^ n9559 ;
  assign n42227 = ~n4364 & n17476 ;
  assign n42228 = n8645 & n42227 ;
  assign n42229 = n42228 ^ n30897 ^ 1'b0 ;
  assign n42226 = n12060 ^ n7755 ^ 1'b0 ;
  assign n42230 = n42229 ^ n42226 ^ n22397 ;
  assign n42231 = n2270 | n37544 ;
  assign n42232 = n42231 ^ n29322 ^ 1'b0 ;
  assign n42234 = ~n5689 & n7701 ;
  assign n42233 = ~n12076 & n27674 ;
  assign n42235 = n42234 ^ n42233 ^ 1'b0 ;
  assign n42236 = n42232 | n42235 ;
  assign n42239 = n2571 & n19729 ;
  assign n42237 = n18903 ^ n17175 ^ 1'b0 ;
  assign n42238 = ~n13897 & n42237 ;
  assign n42240 = n42239 ^ n42238 ^ n30286 ;
  assign n42241 = n4304 & ~n5263 ;
  assign n42242 = ~n4787 & n42241 ;
  assign n42243 = n11325 | n42242 ;
  assign n42244 = n42243 ^ n12571 ^ 1'b0 ;
  assign n42245 = n8265 | n11793 ;
  assign n42246 = ( ~n3156 & n5840 ) | ( ~n3156 & n42245 ) | ( n5840 & n42245 ) ;
  assign n42247 = n42246 ^ n11067 ^ 1'b0 ;
  assign n42248 = n42244 & n42247 ;
  assign n42249 = ~n19620 & n42248 ;
  assign n42250 = ( n2646 & ~n30258 ) | ( n2646 & n42249 ) | ( ~n30258 & n42249 ) ;
  assign n42251 = n21868 ^ n18287 ^ n5482 ;
  assign n42252 = ( ~n16248 & n21911 ) | ( ~n16248 & n39092 ) | ( n21911 & n39092 ) ;
  assign n42253 = n12575 & n24934 ;
  assign n42254 = ~n9814 & n42253 ;
  assign n42255 = x173 & ~n21509 ;
  assign n42256 = ( n22992 & n32525 ) | ( n22992 & n35915 ) | ( n32525 & n35915 ) ;
  assign n42257 = n28577 ^ n15389 ^ n8382 ;
  assign n42258 = n4895 & n14072 ;
  assign n42259 = n42258 ^ n17556 ^ 1'b0 ;
  assign n42260 = n23448 ^ n12931 ^ n266 ;
  assign n42261 = n5579 | n42260 ;
  assign n42262 = n9094 & ~n42261 ;
  assign n42263 = n38094 ^ n22726 ^ 1'b0 ;
  assign n42264 = n20617 & ~n42263 ;
  assign n42265 = ( ~n2985 & n3510 ) | ( ~n2985 & n16823 ) | ( n3510 & n16823 ) ;
  assign n42266 = n5602 & n42265 ;
  assign n42267 = n29129 | n37665 ;
  assign n42268 = ~n2870 & n9519 ;
  assign n42269 = n42267 & n42268 ;
  assign n42270 = ( n33351 & n42266 ) | ( n33351 & ~n42269 ) | ( n42266 & ~n42269 ) ;
  assign n42271 = n3791 & ~n12380 ;
  assign n42272 = ( n1550 & n6776 ) | ( n1550 & ~n42271 ) | ( n6776 & ~n42271 ) ;
  assign n42273 = ( x40 & ~n6658 ) | ( x40 & n17074 ) | ( ~n6658 & n17074 ) ;
  assign n42274 = n42273 ^ n32483 ^ n22366 ;
  assign n42275 = n42274 ^ n12478 ^ 1'b0 ;
  assign n42276 = ~n1372 & n18932 ;
  assign n42277 = n42276 ^ n20486 ^ 1'b0 ;
  assign n42278 = n22177 & n32731 ;
  assign n42279 = ( ~n22903 & n42277 ) | ( ~n22903 & n42278 ) | ( n42277 & n42278 ) ;
  assign n42280 = n21850 | n41273 ;
  assign n42281 = n42280 ^ n33237 ^ 1'b0 ;
  assign n42282 = n21110 & ~n38999 ;
  assign n42283 = n30447 & n42282 ;
  assign n42284 = n42283 ^ n41786 ^ n12442 ;
  assign n42285 = n27154 & ~n42284 ;
  assign n42286 = n33246 ^ n17447 ^ 1'b0 ;
  assign n42287 = n14432 & ~n42286 ;
  assign n42288 = ~n25517 & n42287 ;
  assign n42289 = ~n10144 & n25550 ;
  assign n42290 = n42289 ^ n38252 ^ n21027 ;
  assign n42291 = n42290 ^ n16961 ^ 1'b0 ;
  assign n42292 = n24221 ^ n17120 ^ n17025 ;
  assign n42293 = n14973 | n16160 ;
  assign n42294 = n42293 ^ n21647 ^ 1'b0 ;
  assign n42295 = n42294 ^ n13179 ^ n3105 ;
  assign n42296 = n33830 ^ n20749 ^ 1'b0 ;
  assign n42297 = n20031 | n42296 ;
  assign n42298 = n42297 ^ n27469 ^ n15598 ;
  assign n42299 = n37623 ^ n33367 ^ 1'b0 ;
  assign n42301 = ( ~x132 & n980 ) | ( ~x132 & n10178 ) | ( n980 & n10178 ) ;
  assign n42302 = ( ~n17441 & n23135 ) | ( ~n17441 & n42301 ) | ( n23135 & n42301 ) ;
  assign n42300 = n9859 & ~n23141 ;
  assign n42303 = n42302 ^ n42300 ^ 1'b0 ;
  assign n42304 = n23324 ^ n17410 ^ n10142 ;
  assign n42305 = n27832 ^ n23285 ^ 1'b0 ;
  assign n42306 = ( n1353 & n7650 ) | ( n1353 & ~n40840 ) | ( n7650 & ~n40840 ) ;
  assign n42307 = n36763 ^ n27306 ^ 1'b0 ;
  assign n42308 = ~n25281 & n42307 ;
  assign n42309 = ( n19106 & n41505 ) | ( n19106 & ~n42308 ) | ( n41505 & ~n42308 ) ;
  assign n42310 = n42309 ^ n12972 ^ 1'b0 ;
  assign n42311 = n9839 ^ n8114 ^ n471 ;
  assign n42312 = ~n8175 & n34784 ;
  assign n42313 = n42312 ^ n30294 ^ 1'b0 ;
  assign n42314 = n10979 & ~n24415 ;
  assign n42315 = n9650 ^ n5281 ^ 1'b0 ;
  assign n42316 = n26036 & ~n42315 ;
  assign n42317 = n873 | n1396 ;
  assign n42318 = n42317 ^ n16593 ^ 1'b0 ;
  assign n42319 = n42318 ^ n7978 ^ 1'b0 ;
  assign n42320 = n41623 & n42319 ;
  assign n42321 = ( n3703 & n5490 ) | ( n3703 & ~n41776 ) | ( n5490 & ~n41776 ) ;
  assign n42322 = n20106 & ~n28658 ;
  assign n42323 = n6090 & n42322 ;
  assign n42324 = n42323 ^ n35395 ^ n18757 ;
  assign n42325 = n10706 ^ n1068 ^ 1'b0 ;
  assign n42326 = n10126 & n24240 ;
  assign n42327 = ~n42325 & n42326 ;
  assign n42328 = n7280 & n42327 ;
  assign n42329 = n42328 ^ n32729 ^ 1'b0 ;
  assign n42330 = n14214 ^ n2265 ^ 1'b0 ;
  assign n42331 = n25034 & n42330 ;
  assign n42332 = n5367 & ~n24014 ;
  assign n42333 = n42332 ^ n36730 ^ 1'b0 ;
  assign n42334 = n3104 & n17676 ;
  assign n42335 = ( n4701 & n35048 ) | ( n4701 & n37956 ) | ( n35048 & n37956 ) ;
  assign n42336 = ( n6483 & n16724 ) | ( n6483 & n42335 ) | ( n16724 & n42335 ) ;
  assign n42337 = n42336 ^ n38899 ^ 1'b0 ;
  assign n42338 = n42334 | n42337 ;
  assign n42344 = n18438 ^ n8757 ^ x59 ;
  assign n42345 = ( n21161 & n32513 ) | ( n21161 & n42344 ) | ( n32513 & n42344 ) ;
  assign n42346 = n42345 ^ n11150 ^ 1'b0 ;
  assign n42341 = n10238 ^ n9305 ^ n7957 ;
  assign n42339 = n23882 ^ n19945 ^ 1'b0 ;
  assign n42340 = n13648 & n42339 ;
  assign n42342 = n42341 ^ n42340 ^ n4808 ;
  assign n42343 = ( n27605 & n32322 ) | ( n27605 & n42342 ) | ( n32322 & n42342 ) ;
  assign n42347 = n42346 ^ n42343 ^ n27243 ;
  assign n42353 = n3541 | n34118 ;
  assign n42354 = n5508 & ~n42353 ;
  assign n42348 = ( n9975 & n17891 ) | ( n9975 & n28804 ) | ( n17891 & n28804 ) ;
  assign n42349 = n18351 ^ n10647 ^ 1'b0 ;
  assign n42350 = n29364 & ~n42349 ;
  assign n42351 = ~n42348 & n42350 ;
  assign n42352 = n10916 & n42351 ;
  assign n42355 = n42354 ^ n42352 ^ n12931 ;
  assign n42356 = n12301 ^ n9817 ^ n6408 ;
  assign n42357 = n42356 ^ n38469 ^ n1377 ;
  assign n42363 = n10667 ^ n8762 ^ 1'b0 ;
  assign n42364 = ( ~n5682 & n6765 ) | ( ~n5682 & n42363 ) | ( n6765 & n42363 ) ;
  assign n42365 = n42364 ^ n35612 ^ n27626 ;
  assign n42358 = n9910 ^ n1557 ^ 1'b0 ;
  assign n42359 = n42107 & n42358 ;
  assign n42360 = ~n6587 & n42359 ;
  assign n42361 = n867 & n42360 ;
  assign n42362 = n32415 | n42361 ;
  assign n42366 = n42365 ^ n42362 ^ 1'b0 ;
  assign n42367 = n29835 ^ n27655 ^ 1'b0 ;
  assign n42368 = n12631 & n42367 ;
  assign n42372 = n14866 | n18761 ;
  assign n42369 = ~n10929 & n25408 ;
  assign n42370 = n42369 ^ n877 ^ 1'b0 ;
  assign n42371 = n9108 | n42370 ;
  assign n42373 = n42372 ^ n42371 ^ n33565 ;
  assign n42374 = n10126 & n19566 ;
  assign n42375 = n42374 ^ n23836 ^ n8984 ;
  assign n42376 = ( n5357 & n20389 ) | ( n5357 & ~n21036 ) | ( n20389 & ~n21036 ) ;
  assign n42377 = n42376 ^ n33544 ^ n2314 ;
  assign n42378 = n20659 ^ n20432 ^ n7716 ;
  assign n42379 = n31523 ^ n11171 ^ 1'b0 ;
  assign n42380 = n20434 & n42379 ;
  assign n42381 = n18725 & n42380 ;
  assign n42382 = ~n12659 & n42381 ;
  assign n42383 = ( n3803 & ~n5435 ) | ( n3803 & n9693 ) | ( ~n5435 & n9693 ) ;
  assign n42384 = n37141 ^ n4947 ^ 1'b0 ;
  assign n42385 = n42383 | n42384 ;
  assign n42386 = n12130 ^ n3122 ^ n281 ;
  assign n42387 = n42386 ^ n38933 ^ 1'b0 ;
  assign n42388 = n32561 ^ n18911 ^ n2785 ;
  assign n42389 = n9234 & n12391 ;
  assign n42390 = n42389 ^ n40254 ^ n21165 ;
  assign n42391 = n42390 ^ n41139 ^ n27279 ;
  assign n42393 = n3858 | n6955 ;
  assign n42394 = n42393 ^ n455 ^ 1'b0 ;
  assign n42395 = n42394 ^ n22587 ^ 1'b0 ;
  assign n42396 = ~n2203 & n42395 ;
  assign n42397 = n640 & n14721 ;
  assign n42398 = ~n42396 & n42397 ;
  assign n42392 = ( ~n9920 & n13180 ) | ( ~n9920 & n25342 ) | ( n13180 & n25342 ) ;
  assign n42399 = n42398 ^ n42392 ^ 1'b0 ;
  assign n42400 = n17104 ^ n17089 ^ 1'b0 ;
  assign n42401 = n38384 & ~n42400 ;
  assign n42402 = n14569 ^ n12595 ^ 1'b0 ;
  assign n42403 = n15956 ^ n6110 ^ n5306 ;
  assign n42404 = n18833 | n25011 ;
  assign n42405 = n6451 & ~n42404 ;
  assign n42406 = n14847 & ~n17675 ;
  assign n42407 = n14395 & n42406 ;
  assign n42408 = n24368 ^ n14906 ^ 1'b0 ;
  assign n42409 = n2421 & n42408 ;
  assign n42410 = n508 & n5060 ;
  assign n42411 = ~n2989 & n42410 ;
  assign n42412 = n42409 | n42411 ;
  assign n42413 = n4007 ^ n2510 ^ 1'b0 ;
  assign n42414 = n9155 & ~n42413 ;
  assign n42415 = n16271 ^ n2659 ^ 1'b0 ;
  assign n42416 = n2710 & ~n42415 ;
  assign n42417 = ( n4090 & n42414 ) | ( n4090 & n42416 ) | ( n42414 & n42416 ) ;
  assign n42418 = n2168 & n31067 ;
  assign n42419 = n42418 ^ n8647 ^ 1'b0 ;
  assign n42420 = n3652 & n42419 ;
  assign n42422 = n27083 ^ n19050 ^ 1'b0 ;
  assign n42421 = n5535 ^ n4740 ^ 1'b0 ;
  assign n42423 = n42422 ^ n42421 ^ n31145 ;
  assign n42424 = ~n10913 & n42423 ;
  assign n42425 = n7678 & n42424 ;
  assign n42426 = n8341 | n25050 ;
  assign n42427 = n42426 ^ n4893 ^ 1'b0 ;
  assign n42428 = n16120 ^ n3898 ^ n3074 ;
  assign n42429 = n6153 & ~n42428 ;
  assign n42430 = n16500 ^ n6835 ^ n2563 ;
  assign n42431 = ( n11080 & ~n11747 ) | ( n11080 & n20942 ) | ( ~n11747 & n20942 ) ;
  assign n42432 = n40530 ^ n19228 ^ 1'b0 ;
  assign n42433 = n15084 | n25188 ;
  assign n42434 = n6320 & ~n13991 ;
  assign n42435 = n42434 ^ x181 ^ 1'b0 ;
  assign n42436 = n42435 ^ n15706 ^ n2823 ;
  assign n42441 = n21186 ^ n971 ^ 1'b0 ;
  assign n42440 = ( ~n7708 & n12532 ) | ( ~n7708 & n28350 ) | ( n12532 & n28350 ) ;
  assign n42442 = n42441 ^ n42440 ^ n4697 ;
  assign n42443 = n42442 ^ n13057 ^ 1'b0 ;
  assign n42437 = ( ~n7743 & n11400 ) | ( ~n7743 & n40659 ) | ( n11400 & n40659 ) ;
  assign n42438 = n42437 ^ n13406 ^ n12610 ;
  assign n42439 = x213 & n42438 ;
  assign n42444 = n42443 ^ n42439 ^ 1'b0 ;
  assign n42445 = ~n660 & n4076 ;
  assign n42446 = n42445 ^ n22944 ^ 1'b0 ;
  assign n42447 = n42446 ^ n34848 ^ 1'b0 ;
  assign n42448 = n7067 & ~n42447 ;
  assign n42454 = n33130 ^ n16448 ^ 1'b0 ;
  assign n42455 = ~n5381 & n42454 ;
  assign n42456 = n42455 ^ n10753 ^ 1'b0 ;
  assign n42450 = ~n5899 & n15133 ;
  assign n42451 = n12594 & n42450 ;
  assign n42452 = ( ~n8533 & n36167 ) | ( ~n8533 & n42451 ) | ( n36167 & n42451 ) ;
  assign n42453 = n35168 & ~n42452 ;
  assign n42457 = n42456 ^ n42453 ^ 1'b0 ;
  assign n42458 = n42457 ^ n41109 ^ n2336 ;
  assign n42449 = n5826 & ~n12444 ;
  assign n42459 = n42458 ^ n42449 ^ 1'b0 ;
  assign n42460 = n31097 ^ n28164 ^ n5259 ;
  assign n42461 = n4002 ^ n2113 ^ 1'b0 ;
  assign n42462 = ~n8382 & n42461 ;
  assign n42463 = n42462 ^ n1173 ^ 1'b0 ;
  assign n42464 = ~n19209 & n31611 ;
  assign n42465 = n7086 & ~n42464 ;
  assign n42466 = n18517 ^ n2470 ^ 1'b0 ;
  assign n42467 = ~n9701 & n13609 ;
  assign n42468 = n24343 & n42467 ;
  assign n42469 = n36233 | n42468 ;
  assign n42470 = n18606 | n42469 ;
  assign n42471 = ( n1524 & n5523 ) | ( n1524 & ~n31001 ) | ( n5523 & ~n31001 ) ;
  assign n42472 = n22658 ^ n21041 ^ n15213 ;
  assign n42473 = n42472 ^ n11507 ^ 1'b0 ;
  assign n42474 = n42473 ^ n38988 ^ n26931 ;
  assign n42475 = n1101 & ~n42474 ;
  assign n42476 = n30733 & n34187 ;
  assign n42477 = n37604 ^ n6683 ^ 1'b0 ;
  assign n42478 = n29622 | n36012 ;
  assign n42479 = n5183 | n42478 ;
  assign n42480 = n17602 | n22514 ;
  assign n42481 = n19280 | n42480 ;
  assign n42482 = n23053 ^ n1280 ^ 1'b0 ;
  assign n42483 = n8560 | n8719 ;
  assign n42484 = n42483 ^ n27598 ^ n21138 ;
  assign n42485 = n42484 ^ n10013 ^ n602 ;
  assign n42486 = ( n9635 & n25200 ) | ( n9635 & ~n39241 ) | ( n25200 & ~n39241 ) ;
  assign n42487 = n9472 ^ n6330 ^ 1'b0 ;
  assign n42488 = ~n15269 & n42487 ;
  assign n42489 = n42488 ^ n20393 ^ 1'b0 ;
  assign n42490 = n22607 & ~n42489 ;
  assign n42491 = n23901 | n30650 ;
  assign n42492 = n42491 ^ n41310 ^ 1'b0 ;
  assign n42493 = n11408 | n41496 ;
  assign n42494 = n17871 ^ n4471 ^ 1'b0 ;
  assign n42495 = ( n6841 & n9449 ) | ( n6841 & ~n20035 ) | ( n9449 & ~n20035 ) ;
  assign n42496 = ~n42494 & n42495 ;
  assign n42497 = n42496 ^ n13011 ^ 1'b0 ;
  assign n42499 = ~n20717 & n22896 ;
  assign n42500 = n38067 | n42499 ;
  assign n42498 = n15815 & n24948 ;
  assign n42501 = n42500 ^ n42498 ^ 1'b0 ;
  assign n42502 = ( ~n11478 & n42497 ) | ( ~n11478 & n42501 ) | ( n42497 & n42501 ) ;
  assign n42503 = n41033 ^ n31165 ^ 1'b0 ;
  assign n42504 = n20609 ^ n2903 ^ 1'b0 ;
  assign n42505 = n25967 | n42504 ;
  assign n42506 = n7810 & ~n42505 ;
  assign n42507 = n23372 | n42506 ;
  assign n42508 = n42507 ^ n35032 ^ 1'b0 ;
  assign n42509 = n42508 ^ n21189 ^ 1'b0 ;
  assign n42510 = n5827 & n41715 ;
  assign n42511 = n19806 ^ n3247 ^ 1'b0 ;
  assign n42512 = n42511 ^ n15181 ^ 1'b0 ;
  assign n42513 = n12659 & ~n42512 ;
  assign n42514 = ~n3050 & n19615 ;
  assign n42515 = n11849 & ~n33668 ;
  assign n42516 = n42515 ^ n16951 ^ 1'b0 ;
  assign n42517 = n42516 ^ n3369 ^ 1'b0 ;
  assign n42518 = n14782 & ~n22987 ;
  assign n42519 = n42518 ^ n25074 ^ 1'b0 ;
  assign n42520 = ~n26757 & n38139 ;
  assign n42521 = ~n4382 & n6804 ;
  assign n42522 = n8053 & n42521 ;
  assign n42523 = ~n11075 & n42522 ;
  assign n42524 = n8210 & ~n23144 ;
  assign n42525 = n10131 & n10188 ;
  assign n42526 = n42525 ^ n39097 ^ 1'b0 ;
  assign n42527 = n12538 & ~n29825 ;
  assign n42528 = ( n5510 & n13561 ) | ( n5510 & ~n14583 ) | ( n13561 & ~n14583 ) ;
  assign n42529 = ( n5070 & ~n36928 ) | ( n5070 & n42528 ) | ( ~n36928 & n42528 ) ;
  assign n42530 = ( ~n1112 & n8973 ) | ( ~n1112 & n18108 ) | ( n8973 & n18108 ) ;
  assign n42531 = n42530 ^ n33723 ^ n20064 ;
  assign n42533 = n16935 ^ n1114 ^ 1'b0 ;
  assign n42534 = n2575 & n42533 ;
  assign n42532 = n992 & ~n3599 ;
  assign n42535 = n42534 ^ n42532 ^ 1'b0 ;
  assign n42537 = n37199 ^ n1385 ^ 1'b0 ;
  assign n42538 = n25459 & ~n42537 ;
  assign n42536 = ~n6905 & n17887 ;
  assign n42539 = n42538 ^ n42536 ^ 1'b0 ;
  assign n42543 = n21555 ^ n14824 ^ n4596 ;
  assign n42541 = n602 | n4270 ;
  assign n42542 = n42541 ^ n2220 ^ 1'b0 ;
  assign n42540 = ( n3054 & n29414 ) | ( n3054 & ~n36211 ) | ( n29414 & ~n36211 ) ;
  assign n42544 = n42543 ^ n42542 ^ n42540 ;
  assign n42545 = n8475 ^ n562 ^ 1'b0 ;
  assign n42546 = ( n10391 & n36969 ) | ( n10391 & ~n42545 ) | ( n36969 & ~n42545 ) ;
  assign n42547 = ( n608 & n14173 ) | ( n608 & n25861 ) | ( n14173 & n25861 ) ;
  assign n42548 = n12437 ^ n4796 ^ 1'b0 ;
  assign n42549 = n20082 & n42548 ;
  assign n42550 = n42549 ^ n1538 ^ 1'b0 ;
  assign n42551 = n42550 ^ n20784 ^ n15645 ;
  assign n42552 = ~n2299 & n3757 ;
  assign n42553 = n14469 & n24434 ;
  assign n42554 = n42552 & n42553 ;
  assign n42555 = n33864 ^ n21582 ^ 1'b0 ;
  assign n42556 = n9553 & ~n25519 ;
  assign n42557 = n42556 ^ n3279 ^ 1'b0 ;
  assign n42558 = n637 & n41221 ;
  assign n42559 = ~n17721 & n42558 ;
  assign n42560 = n29583 ^ n19736 ^ 1'b0 ;
  assign n42561 = ~n13331 & n42560 ;
  assign n42562 = n12042 ^ n10538 ^ n329 ;
  assign n42563 = n13566 | n42562 ;
  assign n42564 = n42563 ^ n39753 ^ 1'b0 ;
  assign n42565 = n39504 ^ n20961 ^ n14632 ;
  assign n42566 = n35818 & ~n37584 ;
  assign n42567 = n31236 & n42566 ;
  assign n42568 = n26032 ^ n2593 ^ 1'b0 ;
  assign n42569 = n38241 ^ n18151 ^ 1'b0 ;
  assign n42570 = n26528 | n40198 ;
  assign n42571 = n42569 & ~n42570 ;
  assign n42572 = n1457 & n4124 ;
  assign n42573 = n42572 ^ n36683 ^ 1'b0 ;
  assign n42574 = n24547 ^ n6600 ^ 1'b0 ;
  assign n42575 = n29696 ^ n6461 ^ n3008 ;
  assign n42576 = n13854 ^ n3226 ^ 1'b0 ;
  assign n42577 = n3940 & ~n42576 ;
  assign n42578 = n42577 ^ n8727 ^ n6692 ;
  assign n42579 = n42578 ^ n11136 ^ n4337 ;
  assign n42580 = n14611 & ~n23588 ;
  assign n42581 = n42580 ^ n22518 ^ n8536 ;
  assign n42582 = n10329 ^ n1953 ^ n1871 ;
  assign n42583 = n42582 ^ n42340 ^ 1'b0 ;
  assign n42584 = n42583 ^ n12219 ^ 1'b0 ;
  assign n42585 = ( n3110 & n12308 ) | ( n3110 & n22592 ) | ( n12308 & n22592 ) ;
  assign n42586 = n13723 ^ n1349 ^ 1'b0 ;
  assign n42587 = n42585 & ~n42586 ;
  assign n42588 = ~n14331 & n21187 ;
  assign n42589 = n42588 ^ n30733 ^ 1'b0 ;
  assign n42590 = n11018 ^ n4700 ^ 1'b0 ;
  assign n42591 = ( n12019 & n25899 ) | ( n12019 & n38046 ) | ( n25899 & n38046 ) ;
  assign n42592 = n36800 ^ n13236 ^ n1617 ;
  assign n42593 = n5253 ^ n1385 ^ 1'b0 ;
  assign n42594 = n6301 & n42593 ;
  assign n42595 = n42594 ^ n28806 ^ n3840 ;
  assign n42596 = n42595 ^ n10093 ^ n1934 ;
  assign n42597 = ~n31414 & n42596 ;
  assign n42598 = ~n10317 & n42597 ;
  assign n42599 = n28583 ^ n9358 ^ 1'b0 ;
  assign n42600 = n24522 & ~n42599 ;
  assign n42601 = n18878 ^ n13419 ^ 1'b0 ;
  assign n42602 = ( n1932 & ~n28397 ) | ( n1932 & n36785 ) | ( ~n28397 & n36785 ) ;
  assign n42603 = n42602 ^ n18284 ^ n4556 ;
  assign n42604 = n18156 ^ n10456 ^ n1265 ;
  assign n42605 = n42604 ^ n23107 ^ 1'b0 ;
  assign n42606 = ~n31323 & n42605 ;
  assign n42607 = ( n1102 & n8176 ) | ( n1102 & ~n8605 ) | ( n8176 & ~n8605 ) ;
  assign n42608 = ~n16127 & n18144 ;
  assign n42609 = n42607 & n42608 ;
  assign n42610 = n5605 & n37839 ;
  assign n42611 = ~n16772 & n42610 ;
  assign n42612 = n11341 ^ n722 ^ 1'b0 ;
  assign n42613 = ~n445 & n42612 ;
  assign n42614 = ( n13163 & n28292 ) | ( n13163 & ~n42613 ) | ( n28292 & ~n42613 ) ;
  assign n42615 = n37474 ^ n37054 ^ n16648 ;
  assign n42616 = n631 | n15736 ;
  assign n42617 = ( n26504 & ~n42436 ) | ( n26504 & n42616 ) | ( ~n42436 & n42616 ) ;
  assign n42618 = n40822 ^ n12334 ^ 1'b0 ;
  assign n42619 = x232 & ~n36282 ;
  assign n42620 = n42619 ^ n25952 ^ 1'b0 ;
  assign n42621 = n24831 ^ n19146 ^ 1'b0 ;
  assign n42622 = n8828 | n42621 ;
  assign n42623 = n41139 ^ n32644 ^ 1'b0 ;
  assign n42624 = ( n7160 & n19091 ) | ( n7160 & ~n42623 ) | ( n19091 & ~n42623 ) ;
  assign n42625 = n31431 ^ n18992 ^ 1'b0 ;
  assign n42626 = ( n2818 & ~n12140 ) | ( n2818 & n18317 ) | ( ~n12140 & n18317 ) ;
  assign n42627 = n42626 ^ n5443 ^ n2139 ;
  assign n42628 = n9079 | n42494 ;
  assign n42629 = n12155 ^ n10150 ^ 1'b0 ;
  assign n42630 = ~n28443 & n42629 ;
  assign n42631 = n3165 | n25819 ;
  assign n42632 = n42631 ^ n40265 ^ 1'b0 ;
  assign n42634 = n11565 & ~n13645 ;
  assign n42633 = n14584 & n22629 ;
  assign n42635 = n42634 ^ n42633 ^ 1'b0 ;
  assign n42636 = ( ~n4562 & n5945 ) | ( ~n4562 & n16480 ) | ( n5945 & n16480 ) ;
  assign n42637 = n42636 ^ n5996 ^ 1'b0 ;
  assign n42638 = n13127 & ~n42637 ;
  assign n42639 = n36885 ^ n5014 ^ 1'b0 ;
  assign n42640 = ~n21890 & n42639 ;
  assign n42641 = n27157 ^ n1808 ^ 1'b0 ;
  assign n42642 = n14516 | n25531 ;
  assign n42643 = n42642 ^ n26114 ^ n7304 ;
  assign n42644 = n1164 | n30267 ;
  assign n42645 = n42644 ^ n16060 ^ 1'b0 ;
  assign n42646 = n29374 ^ n11166 ^ 1'b0 ;
  assign n42647 = n42646 ^ n14155 ^ 1'b0 ;
  assign n42648 = n4429 & ~n19157 ;
  assign n42649 = ~n695 & n42648 ;
  assign n42650 = n10585 & ~n42649 ;
  assign n42651 = n22166 ^ n17718 ^ 1'b0 ;
  assign n42652 = n38604 & n42651 ;
  assign n42653 = n23886 ^ n21435 ^ n20486 ;
  assign n42654 = n9468 | n42653 ;
  assign n42655 = n42654 ^ n34272 ^ 1'b0 ;
  assign n42656 = n6281 | n14117 ;
  assign n42657 = n7902 & ~n8771 ;
  assign n42658 = ~n26464 & n42657 ;
  assign n42659 = n1775 & n11018 ;
  assign n42660 = n42659 ^ n2944 ^ 1'b0 ;
  assign n42661 = ~n42658 & n42660 ;
  assign n42662 = ( n10283 & ~n42656 ) | ( n10283 & n42661 ) | ( ~n42656 & n42661 ) ;
  assign n42663 = n11503 & n29113 ;
  assign n42664 = n2680 & ~n4032 ;
  assign n42665 = n42663 & n42664 ;
  assign n42666 = n42665 ^ n20706 ^ n11723 ;
  assign n42667 = ( ~n31626 & n35115 ) | ( ~n31626 & n38263 ) | ( n35115 & n38263 ) ;
  assign n42668 = n1848 | n15368 ;
  assign n42669 = n42668 ^ n19492 ^ 1'b0 ;
  assign n42670 = n28118 ^ n5730 ^ 1'b0 ;
  assign n42671 = n11247 & n42670 ;
  assign n42672 = n16221 ^ n8383 ^ n5387 ;
  assign n42673 = n42672 ^ n14443 ^ 1'b0 ;
  assign n42674 = n35541 & ~n42673 ;
  assign n42675 = ( n13022 & n14931 ) | ( n13022 & ~n32263 ) | ( n14931 & ~n32263 ) ;
  assign n42676 = ~n21261 & n42675 ;
  assign n42677 = ~n30062 & n42676 ;
  assign n42678 = n31750 ^ n13082 ^ 1'b0 ;
  assign n42679 = ~n42677 & n42678 ;
  assign n42680 = ~n5744 & n42015 ;
  assign n42681 = n42680 ^ n19874 ^ 1'b0 ;
  assign n42682 = n42681 ^ n28295 ^ n26075 ;
  assign n42683 = n22937 & n42682 ;
  assign n42684 = n40276 ^ n29172 ^ 1'b0 ;
  assign n42685 = n26755 ^ n9824 ^ n8606 ;
  assign n42686 = n40599 ^ n5359 ^ 1'b0 ;
  assign n42687 = ( n2523 & n28103 ) | ( n2523 & ~n41410 ) | ( n28103 & ~n41410 ) ;
  assign n42688 = n39761 & n39893 ;
  assign n42689 = n11261 & n40655 ;
  assign n42690 = ~n39772 & n42689 ;
  assign n42691 = ( ~n12278 & n12607 ) | ( ~n12278 & n36923 ) | ( n12607 & n36923 ) ;
  assign n42692 = n5554 & ~n6499 ;
  assign n42695 = n11108 ^ n8707 ^ 1'b0 ;
  assign n42696 = n42695 ^ n18810 ^ n9941 ;
  assign n42693 = n21826 ^ n21666 ^ n8613 ;
  assign n42694 = ( n14170 & n14207 ) | ( n14170 & n42693 ) | ( n14207 & n42693 ) ;
  assign n42697 = n42696 ^ n42694 ^ n29439 ;
  assign n42698 = ~n9486 & n25538 ;
  assign n42699 = ( ~x131 & n16552 ) | ( ~x131 & n42698 ) | ( n16552 & n42698 ) ;
  assign n42700 = n690 & ~n24339 ;
  assign n42701 = n42700 ^ n13524 ^ 1'b0 ;
  assign n42702 = ( ~n791 & n42699 ) | ( ~n791 & n42701 ) | ( n42699 & n42701 ) ;
  assign n42703 = n39082 ^ n6097 ^ 1'b0 ;
  assign n42704 = n42703 ^ n28414 ^ n4048 ;
  assign n42705 = n17647 & ~n22436 ;
  assign n42706 = n1934 & ~n2215 ;
  assign n42707 = ( ~n10181 & n10919 ) | ( ~n10181 & n42706 ) | ( n10919 & n42706 ) ;
  assign n42708 = ( n8038 & ~n27289 ) | ( n8038 & n34678 ) | ( ~n27289 & n34678 ) ;
  assign n42709 = n3721 & ~n42708 ;
  assign n42710 = n42707 & n42709 ;
  assign n42711 = n13195 & n20546 ;
  assign n42712 = ~n23434 & n42711 ;
  assign n42713 = n7263 & ~n42712 ;
  assign n42714 = n5699 & n42713 ;
  assign n42715 = n11735 & ~n33567 ;
  assign n42716 = ~n29819 & n42715 ;
  assign n42717 = n30600 ^ n9413 ^ n1680 ;
  assign n42718 = n10922 ^ x33 ^ 1'b0 ;
  assign n42719 = n42717 & n42718 ;
  assign n42720 = n6375 | n9069 ;
  assign n42721 = n42720 ^ n6757 ^ 1'b0 ;
  assign n42722 = n1352 & ~n13780 ;
  assign n42723 = n13002 | n36309 ;
  assign n42724 = n21882 | n42723 ;
  assign n42725 = ( n421 & n7064 ) | ( n421 & ~n38972 ) | ( n7064 & ~n38972 ) ;
  assign n42726 = n42725 ^ n31645 ^ n5762 ;
  assign n42727 = ( n26896 & ~n42724 ) | ( n26896 & n42726 ) | ( ~n42724 & n42726 ) ;
  assign n42728 = ( n9452 & n10151 ) | ( n9452 & n20392 ) | ( n10151 & n20392 ) ;
  assign n42729 = n23258 ^ n19972 ^ 1'b0 ;
  assign n42730 = n18292 & ~n42729 ;
  assign n42731 = n42728 & n42730 ;
  assign n42732 = ( n27568 & ~n38267 ) | ( n27568 & n42731 ) | ( ~n38267 & n42731 ) ;
  assign n42733 = n40593 ^ n841 ^ 1'b0 ;
  assign n42734 = n3528 & ~n7007 ;
  assign n42735 = n29576 ^ n28066 ^ 1'b0 ;
  assign n42736 = n9091 & ~n42735 ;
  assign n42737 = x54 & n6615 ;
  assign n42738 = n9787 & n42737 ;
  assign n42739 = n42738 ^ n15862 ^ 1'b0 ;
  assign n42740 = n11330 | n42739 ;
  assign n42741 = n30925 | n42740 ;
  assign n42742 = n42736 | n42741 ;
  assign n42743 = n16159 | n27996 ;
  assign n42744 = n11816 ^ n9397 ^ n3605 ;
  assign n42745 = n42744 ^ n9578 ^ n445 ;
  assign n42746 = n42745 ^ n11872 ^ n3310 ;
  assign n42747 = n29643 ^ n19709 ^ n17609 ;
  assign n42748 = n6912 & ~n12583 ;
  assign n42749 = n42748 ^ n7220 ^ 1'b0 ;
  assign n42750 = n11968 | n42749 ;
  assign n42751 = n13777 & ~n42750 ;
  assign n42752 = ( n3796 & n42747 ) | ( n3796 & n42751 ) | ( n42747 & n42751 ) ;
  assign n42753 = ~n17929 & n39485 ;
  assign n42754 = ~n13388 & n42753 ;
  assign n42755 = n42754 ^ n15174 ^ n13187 ;
  assign n42756 = n42755 ^ n40578 ^ n39826 ;
  assign n42757 = n6145 & n12675 ;
  assign n42758 = n42757 ^ n3721 ^ 1'b0 ;
  assign n42759 = n42758 ^ n12300 ^ 1'b0 ;
  assign n42760 = n42759 ^ n27071 ^ n3930 ;
  assign n42761 = ( n11111 & ~n23979 ) | ( n11111 & n42760 ) | ( ~n23979 & n42760 ) ;
  assign n42762 = ( n5880 & ~n32853 ) | ( n5880 & n42761 ) | ( ~n32853 & n42761 ) ;
  assign n42763 = ~n10682 & n34631 ;
  assign n42764 = n42763 ^ n7973 ^ 1'b0 ;
  assign n42765 = n594 | n42764 ;
  assign n42766 = n29696 ^ n9572 ^ 1'b0 ;
  assign n42767 = ( n5254 & n17585 ) | ( n5254 & ~n18994 ) | ( n17585 & ~n18994 ) ;
  assign n42768 = n20102 | n42767 ;
  assign n42769 = n42766 & ~n42768 ;
  assign n42770 = n4256 & ~n13524 ;
  assign n42771 = n42770 ^ n28778 ^ 1'b0 ;
  assign n42772 = n42771 ^ n15753 ^ n2559 ;
  assign n42773 = n40403 & ~n42772 ;
  assign n42774 = ~n2878 & n23805 ;
  assign n42775 = ~n17757 & n42774 ;
  assign n42776 = n1181 & ~n9266 ;
  assign n42777 = n42776 ^ n25532 ^ n18624 ;
  assign n42778 = n41560 | n42777 ;
  assign n42779 = n18811 | n42778 ;
  assign n42780 = n42779 ^ n9180 ^ 1'b0 ;
  assign n42781 = n8614 ^ n7374 ^ 1'b0 ;
  assign n42782 = n42781 ^ n8854 ^ 1'b0 ;
  assign n42783 = n18172 & ~n42782 ;
  assign n42784 = n3121 & n42783 ;
  assign n42785 = ~n40598 & n42784 ;
  assign n42786 = n42785 ^ n6258 ^ n4378 ;
  assign n42787 = n20630 ^ n6825 ^ 1'b0 ;
  assign n42788 = ( n11909 & n35692 ) | ( n11909 & ~n42787 ) | ( n35692 & ~n42787 ) ;
  assign n42789 = n13219 & n14425 ;
  assign n42790 = n42789 ^ n15532 ^ 1'b0 ;
  assign n42791 = n42788 & ~n42790 ;
  assign n42792 = ( n2083 & ~n8063 ) | ( n2083 & n8175 ) | ( ~n8063 & n8175 ) ;
  assign n42793 = n42792 ^ n11492 ^ 1'b0 ;
  assign n42794 = ~n13252 & n24484 ;
  assign n42795 = n42794 ^ n39004 ^ 1'b0 ;
  assign n42797 = n21043 ^ n3031 ^ n898 ;
  assign n42796 = x109 & n28049 ;
  assign n42798 = n42797 ^ n42796 ^ 1'b0 ;
  assign n42799 = n32990 ^ n21572 ^ 1'b0 ;
  assign n42800 = n14602 & n26775 ;
  assign n42801 = ~n2432 & n42800 ;
  assign n42802 = n42801 ^ n41273 ^ 1'b0 ;
  assign n42803 = n30295 ^ n23848 ^ 1'b0 ;
  assign n42804 = ( n686 & ~n3168 ) | ( n686 & n42803 ) | ( ~n3168 & n42803 ) ;
  assign n42805 = ( ~n1588 & n11348 ) | ( ~n1588 & n41806 ) | ( n11348 & n41806 ) ;
  assign n42806 = ( n10903 & n11196 ) | ( n10903 & n42805 ) | ( n11196 & n42805 ) ;
  assign n42807 = n42806 ^ n39319 ^ 1'b0 ;
  assign n42808 = n37665 ^ n37499 ^ n24351 ;
  assign n42809 = n11809 ^ n8910 ^ 1'b0 ;
  assign n42810 = n9590 & n36887 ;
  assign n42811 = n19306 & n42810 ;
  assign n42812 = ( n11606 & n12593 ) | ( n11606 & ~n42811 ) | ( n12593 & ~n42811 ) ;
  assign n42813 = ~n42809 & n42812 ;
  assign n42814 = ~n5563 & n42813 ;
  assign n42816 = n30206 ^ n13169 ^ 1'b0 ;
  assign n42815 = n4759 & ~n11227 ;
  assign n42817 = n42816 ^ n42815 ^ 1'b0 ;
  assign n42818 = n19940 ^ n2506 ^ 1'b0 ;
  assign n42819 = n42817 & n42818 ;
  assign n42820 = n10177 & ~n15977 ;
  assign n42821 = n42820 ^ n4762 ^ 1'b0 ;
  assign n42822 = n42821 ^ n19205 ^ n11802 ;
  assign n42823 = ( n7375 & n37707 ) | ( n7375 & n42822 ) | ( n37707 & n42822 ) ;
  assign n42824 = n17310 & n34544 ;
  assign n42825 = ( n5912 & n18233 ) | ( n5912 & ~n42506 ) | ( n18233 & ~n42506 ) ;
  assign n42828 = n2201 & n7902 ;
  assign n42829 = ~n2201 & n42828 ;
  assign n42830 = n9364 & n9623 ;
  assign n42831 = n42829 & n42830 ;
  assign n42832 = n8913 & n8924 ;
  assign n42833 = n42831 & n42832 ;
  assign n42826 = n5751 & n19651 ;
  assign n42827 = n42826 ^ n32891 ^ n18853 ;
  assign n42834 = n42833 ^ n42827 ^ n31708 ;
  assign n42835 = n35771 ^ n26051 ^ 1'b0 ;
  assign n42836 = n17170 ^ n6304 ^ 1'b0 ;
  assign n42837 = n10478 | n20550 ;
  assign n42838 = n42836 | n42837 ;
  assign n42839 = n19244 & n28152 ;
  assign n42840 = n15614 & ~n42839 ;
  assign n42841 = n42840 ^ n4538 ^ 1'b0 ;
  assign n42842 = n42841 ^ n7107 ^ 1'b0 ;
  assign n42843 = n22079 | n42842 ;
  assign n42844 = n24069 ^ n20254 ^ 1'b0 ;
  assign n42845 = ( n7538 & n20802 ) | ( n7538 & ~n26270 ) | ( n20802 & ~n26270 ) ;
  assign n42846 = n26914 ^ n24086 ^ 1'b0 ;
  assign n42847 = n11565 & ~n42846 ;
  assign n42848 = n42847 ^ n32093 ^ x48 ;
  assign n42849 = n8884 ^ n8737 ^ n5017 ;
  assign n42850 = n4827 & ~n22012 ;
  assign n42851 = n42850 ^ n16575 ^ 1'b0 ;
  assign n42852 = n26674 ^ n4137 ^ n1049 ;
  assign n42853 = n36090 & n42852 ;
  assign n42854 = ~n12194 & n42853 ;
  assign n42856 = n7314 & n27009 ;
  assign n42855 = n9238 & n30360 ;
  assign n42857 = n42856 ^ n42855 ^ 1'b0 ;
  assign n42859 = n12551 ^ n11940 ^ n4025 ;
  assign n42858 = ~n11212 & n17296 ;
  assign n42860 = n42859 ^ n42858 ^ 1'b0 ;
  assign n42863 = n29939 ^ n11401 ^ 1'b0 ;
  assign n42864 = n2127 & ~n42863 ;
  assign n42861 = n28970 ^ n8421 ^ 1'b0 ;
  assign n42862 = n2086 & ~n42861 ;
  assign n42865 = n42864 ^ n42862 ^ 1'b0 ;
  assign n42866 = n16650 ^ n14600 ^ n930 ;
  assign n42867 = n19375 & ~n42866 ;
  assign n42868 = n6918 & n21367 ;
  assign n42869 = n34715 ^ n5233 ^ n5183 ;
  assign n42870 = n5316 | n12203 ;
  assign n42871 = n42870 ^ n7126 ^ 1'b0 ;
  assign n42872 = n42871 ^ n23477 ^ x10 ;
  assign n42873 = n15113 | n31490 ;
  assign n42874 = n36255 ^ n14499 ^ 1'b0 ;
  assign n42875 = n15347 ^ n1539 ^ 1'b0 ;
  assign n42876 = ( n39613 & n42874 ) | ( n39613 & ~n42875 ) | ( n42874 & ~n42875 ) ;
  assign n42877 = ~n31621 & n42876 ;
  assign n42878 = n33312 ^ n12988 ^ 1'b0 ;
  assign n42879 = n25482 | n42878 ;
  assign n42880 = n4404 | n8405 ;
  assign n42881 = n42880 ^ n8063 ^ 1'b0 ;
  assign n42882 = ( ~n8290 & n29146 ) | ( ~n8290 & n42881 ) | ( n29146 & n42881 ) ;
  assign n42883 = n28314 ^ n17407 ^ 1'b0 ;
  assign n42886 = n10332 | n29165 ;
  assign n42884 = n11242 ^ n477 ^ 1'b0 ;
  assign n42885 = n30297 | n42884 ;
  assign n42887 = n42886 ^ n42885 ^ 1'b0 ;
  assign n42888 = ( n7395 & n17000 ) | ( n7395 & n25639 ) | ( n17000 & n25639 ) ;
  assign n42889 = n15713 ^ n15528 ^ 1'b0 ;
  assign n42890 = n14258 | n42889 ;
  assign n42891 = ( ~n24411 & n42888 ) | ( ~n24411 & n42890 ) | ( n42888 & n42890 ) ;
  assign n42894 = n7203 & n34729 ;
  assign n42895 = n42894 ^ n6068 ^ 1'b0 ;
  assign n42896 = n42895 ^ n4733 ^ 1'b0 ;
  assign n42897 = ~n8716 & n42896 ;
  assign n42898 = n8913 ^ n4202 ^ 1'b0 ;
  assign n42899 = n42897 & ~n42898 ;
  assign n42892 = ( n14533 & n22814 ) | ( n14533 & ~n36449 ) | ( n22814 & ~n36449 ) ;
  assign n42893 = n10815 & n42892 ;
  assign n42900 = n42899 ^ n42893 ^ 1'b0 ;
  assign n42901 = n15080 & ~n17179 ;
  assign n42902 = n42901 ^ n25129 ^ 1'b0 ;
  assign n42903 = ( ~n5402 & n15892 ) | ( ~n5402 & n18796 ) | ( n15892 & n18796 ) ;
  assign n42904 = ~n3281 & n42903 ;
  assign n42905 = n27470 ^ n19201 ^ 1'b0 ;
  assign n42906 = n42904 | n42905 ;
  assign n42907 = ( n10623 & n35558 ) | ( n10623 & n37730 ) | ( n35558 & n37730 ) ;
  assign n42908 = ( n26512 & n31373 ) | ( n26512 & n35353 ) | ( n31373 & n35353 ) ;
  assign n42909 = n12400 & ~n22264 ;
  assign n42910 = n42909 ^ n17439 ^ n5123 ;
  assign n42911 = n21755 & n42910 ;
  assign n42912 = n28264 ^ n13021 ^ 1'b0 ;
  assign n42914 = n36201 ^ n1311 ^ 1'b0 ;
  assign n42913 = ~n9213 & n33400 ;
  assign n42915 = n42914 ^ n42913 ^ 1'b0 ;
  assign n42916 = ~n5502 & n8921 ;
  assign n42917 = ( n634 & ~n13619 ) | ( n634 & n19393 ) | ( ~n13619 & n19393 ) ;
  assign n42918 = ( ~x25 & n20962 ) | ( ~x25 & n24067 ) | ( n20962 & n24067 ) ;
  assign n42919 = n42918 ^ n14094 ^ 1'b0 ;
  assign n42920 = n6216 | n42919 ;
  assign n42921 = n42920 ^ n26934 ^ 1'b0 ;
  assign n42922 = ( n3175 & ~n12147 ) | ( n3175 & n26040 ) | ( ~n12147 & n26040 ) ;
  assign n42923 = n12869 ^ n10189 ^ 1'b0 ;
  assign n42924 = ( n8087 & ~n42922 ) | ( n8087 & n42923 ) | ( ~n42922 & n42923 ) ;
  assign n42925 = ~n13023 & n22303 ;
  assign n42926 = n42925 ^ n19940 ^ 1'b0 ;
  assign n42927 = n42926 ^ n9220 ^ n4416 ;
  assign n42928 = ~n757 & n42927 ;
  assign n42929 = n42928 ^ n28055 ^ 1'b0 ;
  assign n42930 = ~n15828 & n20611 ;
  assign n42931 = n42930 ^ n23498 ^ 1'b0 ;
  assign n42932 = ( n42924 & n42929 ) | ( n42924 & ~n42931 ) | ( n42929 & ~n42931 ) ;
  assign n42933 = n24450 ^ n23543 ^ n22828 ;
  assign n42934 = ~n780 & n36167 ;
  assign n42935 = n31400 & n42934 ;
  assign n42936 = n7731 & ~n16982 ;
  assign n42937 = n18838 ^ n11250 ^ 1'b0 ;
  assign n42938 = ~n5233 & n42937 ;
  assign n42939 = ( n1745 & n42936 ) | ( n1745 & n42938 ) | ( n42936 & n42938 ) ;
  assign n42940 = ( n10077 & ~n42935 ) | ( n10077 & n42939 ) | ( ~n42935 & n42939 ) ;
  assign n42941 = ~n12638 & n42940 ;
  assign n42942 = ~n40226 & n42941 ;
  assign n42943 = n16623 ^ n14712 ^ 1'b0 ;
  assign n42944 = n6889 ^ n3151 ^ 1'b0 ;
  assign n42945 = n21537 ^ n4591 ^ 1'b0 ;
  assign n42946 = n17685 & ~n42945 ;
  assign n42947 = ( n6252 & n9385 ) | ( n6252 & n12757 ) | ( n9385 & n12757 ) ;
  assign n42948 = n22282 | n42947 ;
  assign n42949 = n2614 & ~n42607 ;
  assign n42950 = n42949 ^ n30929 ^ 1'b0 ;
  assign n42951 = ~n42948 & n42950 ;
  assign n42952 = ~n42141 & n42951 ;
  assign n42953 = ( n14042 & n42946 ) | ( n14042 & n42952 ) | ( n42946 & n42952 ) ;
  assign n42954 = n27792 & n42953 ;
  assign n42955 = ~n42944 & n42954 ;
  assign n42956 = ( ~n6589 & n11766 ) | ( ~n6589 & n17872 ) | ( n11766 & n17872 ) ;
  assign n42957 = n16887 & ~n19520 ;
  assign n42958 = n42957 ^ n33752 ^ 1'b0 ;
  assign n42959 = n26323 | n42958 ;
  assign n42960 = ( n2747 & n10271 ) | ( n2747 & n37991 ) | ( n10271 & n37991 ) ;
  assign n42961 = n14472 ^ n9710 ^ n3730 ;
  assign n42962 = n42961 ^ n31060 ^ 1'b0 ;
  assign n42963 = n9961 ^ n5981 ^ 1'b0 ;
  assign n42964 = n40873 & ~n42963 ;
  assign n42965 = ( n812 & n4881 ) | ( n812 & n34003 ) | ( n4881 & n34003 ) ;
  assign n42966 = n38647 ^ n9067 ^ 1'b0 ;
  assign n42967 = n31270 & n42966 ;
  assign n42968 = n42967 ^ n32635 ^ n22118 ;
  assign n42969 = n42968 ^ n14067 ^ 1'b0 ;
  assign n42970 = n42965 & ~n42969 ;
  assign n42971 = n14636 | n26354 ;
  assign n42972 = n38307 & ~n42971 ;
  assign n42973 = n5557 ^ n1844 ^ 1'b0 ;
  assign n42974 = n17321 & n42973 ;
  assign n42975 = ( ~n23046 & n23759 ) | ( ~n23046 & n42974 ) | ( n23759 & n42974 ) ;
  assign n42976 = ( n448 & n12242 ) | ( n448 & n25679 ) | ( n12242 & n25679 ) ;
  assign n42977 = n20850 ^ n7200 ^ n1171 ;
  assign n42978 = ~n4677 & n42977 ;
  assign n42979 = ~n9130 & n42978 ;
  assign n42980 = n6197 & n25276 ;
  assign n42981 = n3790 & n11434 ;
  assign n42982 = ( n3571 & n42457 ) | ( n3571 & n42981 ) | ( n42457 & n42981 ) ;
  assign n42983 = n2203 ^ n2132 ^ 1'b0 ;
  assign n42984 = ~n2394 & n42983 ;
  assign n42985 = n13414 & n15682 ;
  assign n42986 = ~n42984 & n42985 ;
  assign n42987 = ~n340 & n22492 ;
  assign n42988 = ~n16030 & n42987 ;
  assign n42989 = n17984 | n25882 ;
  assign n42990 = n12081 | n42989 ;
  assign n42991 = n6646 ^ n4809 ^ 1'b0 ;
  assign n42992 = n42990 & n42991 ;
  assign n42993 = n14613 ^ n9075 ^ 1'b0 ;
  assign n42994 = n358 & n42993 ;
  assign n42995 = n2835 | n42994 ;
  assign n42996 = ( n5901 & n31400 ) | ( n5901 & n33538 ) | ( n31400 & n33538 ) ;
  assign n42997 = n42996 ^ n29502 ^ n2686 ;
  assign n42998 = n42997 ^ n10322 ^ n6229 ;
  assign n42999 = n12929 ^ n11576 ^ 1'b0 ;
  assign n43000 = ~n21849 & n41004 ;
  assign n43001 = n43000 ^ n21807 ^ 1'b0 ;
  assign n43002 = ( n25692 & n26228 ) | ( n25692 & ~n43001 ) | ( n26228 & ~n43001 ) ;
  assign n43003 = ~n6068 & n11222 ;
  assign n43004 = n43003 ^ x66 ^ 1'b0 ;
  assign n43005 = ( ~n8942 & n19744 ) | ( ~n8942 & n43004 ) | ( n19744 & n43004 ) ;
  assign n43006 = n12817 ^ n2411 ^ n1454 ;
  assign n43007 = n43006 ^ n19773 ^ 1'b0 ;
  assign n43008 = n9606 & n43007 ;
  assign n43009 = n43008 ^ x81 ^ 1'b0 ;
  assign n43011 = n38124 ^ n36146 ^ n18460 ;
  assign n43010 = n24346 ^ n14432 ^ n8176 ;
  assign n43012 = n43011 ^ n43010 ^ n37913 ;
  assign n43013 = n11838 | n17370 ;
  assign n43014 = n12564 & n43013 ;
  assign n43015 = n15333 ^ n14341 ^ 1'b0 ;
  assign n43016 = n33875 | n43015 ;
  assign n43020 = n14992 ^ n8110 ^ 1'b0 ;
  assign n43017 = n1323 & n26294 ;
  assign n43018 = ~n22035 & n43017 ;
  assign n43019 = n8695 & ~n43018 ;
  assign n43021 = n43020 ^ n43019 ^ 1'b0 ;
  assign n43022 = n21519 & n40459 ;
  assign n43023 = n43022 ^ n8612 ^ 1'b0 ;
  assign n43024 = n21131 ^ n11492 ^ 1'b0 ;
  assign n43025 = n42506 ^ n36667 ^ n23258 ;
  assign n43026 = n33563 ^ n15596 ^ 1'b0 ;
  assign n43027 = n40743 ^ n33097 ^ n5532 ;
  assign n43028 = n31394 ^ n23422 ^ 1'b0 ;
  assign n43029 = ~n43027 & n43028 ;
  assign n43030 = n10816 & ~n13252 ;
  assign n43031 = ( n21797 & n26400 ) | ( n21797 & ~n40556 ) | ( n26400 & ~n40556 ) ;
  assign n43032 = ( ~n19393 & n43030 ) | ( ~n19393 & n43031 ) | ( n43030 & n43031 ) ;
  assign n43033 = n2244 & ~n43032 ;
  assign n43034 = n40333 ^ n21059 ^ n18684 ;
  assign n43035 = n43034 ^ n26942 ^ 1'b0 ;
  assign n43036 = n13127 & ~n37004 ;
  assign n43037 = n25982 ^ n9452 ^ n2555 ;
  assign n43038 = n813 | n4904 ;
  assign n43039 = n9858 | n29033 ;
  assign n43040 = n6297 | n32822 ;
  assign n43041 = n43040 ^ n39353 ^ n16906 ;
  assign n43046 = n8050 & n12519 ;
  assign n43047 = n43046 ^ n20689 ^ n5809 ;
  assign n43042 = x79 & n40454 ;
  assign n43043 = n43042 ^ n11463 ^ 1'b0 ;
  assign n43044 = n43043 ^ n32560 ^ 1'b0 ;
  assign n43045 = n1480 | n43044 ;
  assign n43048 = n43047 ^ n43045 ^ n5660 ;
  assign n43049 = n10991 ^ n4688 ^ 1'b0 ;
  assign n43050 = n16689 & ~n43049 ;
  assign n43051 = n43050 ^ n6730 ^ 1'b0 ;
  assign n43052 = n43051 ^ n20144 ^ n2386 ;
  assign n43053 = n406 & n41553 ;
  assign n43054 = n43053 ^ n19675 ^ n18124 ;
  assign n43055 = n33246 | n43054 ;
  assign n43056 = n966 & n2341 ;
  assign n43057 = n43056 ^ n22966 ^ 1'b0 ;
  assign n43058 = n39733 & ~n43057 ;
  assign n43060 = n2017 & n19822 ;
  assign n43059 = n16548 | n34678 ;
  assign n43061 = n43060 ^ n43059 ^ 1'b0 ;
  assign n43062 = ~n11699 & n33857 ;
  assign n43063 = n11518 | n12223 ;
  assign n43064 = n43063 ^ n24169 ^ n8390 ;
  assign n43065 = n31504 ^ n12685 ^ 1'b0 ;
  assign n43066 = ~n38880 & n42675 ;
  assign n43067 = ~n10161 & n20305 ;
  assign n43068 = n14270 & n43067 ;
  assign n43069 = n31151 | n41189 ;
  assign n43070 = n20315 & n43069 ;
  assign n43071 = n43070 ^ n27895 ^ 1'b0 ;
  assign n43072 = n7721 | n11132 ;
  assign n43073 = ( ~n9963 & n24401 ) | ( ~n9963 & n43072 ) | ( n24401 & n43072 ) ;
  assign n43074 = n3286 & ~n15066 ;
  assign n43075 = ~n11461 & n43074 ;
  assign n43076 = n43075 ^ n28134 ^ n14446 ;
  assign n43077 = ( ~n1855 & n16873 ) | ( ~n1855 & n19795 ) | ( n16873 & n19795 ) ;
  assign n43078 = ~n10028 & n11560 ;
  assign n43079 = ~n18623 & n33655 ;
  assign n43080 = ( n43077 & ~n43078 ) | ( n43077 & n43079 ) | ( ~n43078 & n43079 ) ;
  assign n43081 = n43080 ^ n18800 ^ n12549 ;
  assign n43082 = n37662 ^ n28733 ^ 1'b0 ;
  assign n43083 = ( n22741 & n40489 ) | ( n22741 & n43082 ) | ( n40489 & n43082 ) ;
  assign n43084 = n11820 ^ n810 ^ 1'b0 ;
  assign n43085 = n40803 ^ n1660 ^ 1'b0 ;
  assign n43086 = n12147 & ~n43085 ;
  assign n43087 = ~n3133 & n29447 ;
  assign n43088 = n43087 ^ n8076 ^ 1'b0 ;
  assign n43089 = n40822 ^ n12341 ^ 1'b0 ;
  assign n43090 = n30020 ^ n25469 ^ n9994 ;
  assign n43091 = n36151 ^ n14722 ^ 1'b0 ;
  assign n43092 = ~n9965 & n43091 ;
  assign n43093 = n19091 ^ n9497 ^ 1'b0 ;
  assign n43094 = n37106 & n43093 ;
  assign n43095 = n43094 ^ n43001 ^ n27076 ;
  assign n43096 = n22559 ^ n2104 ^ 1'b0 ;
  assign n43097 = n9661 & n43096 ;
  assign n43098 = n17926 ^ n11115 ^ 1'b0 ;
  assign n43099 = n43097 & n43098 ;
  assign n43100 = ~n1438 & n43099 ;
  assign n43101 = n2843 | n43100 ;
  assign n43102 = n2908 ^ n1631 ^ 1'b0 ;
  assign n43103 = n2031 & ~n9827 ;
  assign n43104 = n43103 ^ n29839 ^ 1'b0 ;
  assign n43105 = n11083 & ~n32789 ;
  assign n43106 = ~n24646 & n43105 ;
  assign n43107 = n5387 & n30010 ;
  assign n43108 = ~n32714 & n43107 ;
  assign n43109 = ( n22302 & ~n43106 ) | ( n22302 & n43108 ) | ( ~n43106 & n43108 ) ;
  assign n43110 = ( n5872 & ~n24527 ) | ( n5872 & n27515 ) | ( ~n24527 & n27515 ) ;
  assign n43111 = n43110 ^ n31800 ^ 1'b0 ;
  assign n43112 = n20286 ^ n13020 ^ n5038 ;
  assign n43114 = n12130 & n19204 ;
  assign n43115 = ~n640 & n43114 ;
  assign n43113 = n24571 & n34190 ;
  assign n43116 = n43115 ^ n43113 ^ 1'b0 ;
  assign n43117 = n4353 | n32772 ;
  assign n43118 = n43117 ^ n35575 ^ 1'b0 ;
  assign n43119 = n34085 ^ n18098 ^ 1'b0 ;
  assign n43120 = n40797 & ~n43119 ;
  assign n43121 = n5725 ^ n2216 ^ 1'b0 ;
  assign n43122 = n13536 | n43121 ;
  assign n43123 = n40483 & ~n43122 ;
  assign n43124 = ~n43120 & n43123 ;
  assign n43126 = ( n11107 & n20282 ) | ( n11107 & n24194 ) | ( n20282 & n24194 ) ;
  assign n43125 = n15806 ^ x7 ^ 1'b0 ;
  assign n43127 = n43126 ^ n43125 ^ n7741 ;
  assign n43128 = n30044 ^ n19386 ^ 1'b0 ;
  assign n43129 = n28270 ^ n23909 ^ 1'b0 ;
  assign n43130 = n17808 | n43129 ;
  assign n43131 = ( n11997 & n18323 ) | ( n11997 & ~n26966 ) | ( n18323 & ~n26966 ) ;
  assign n43132 = ~n43130 & n43131 ;
  assign n43133 = n43132 ^ n30965 ^ 1'b0 ;
  assign n43134 = n41310 | n43133 ;
  assign n43135 = ( n3828 & ~n43128 ) | ( n3828 & n43134 ) | ( ~n43128 & n43134 ) ;
  assign n43136 = n24481 & ~n37175 ;
  assign n43139 = n17629 & n21209 ;
  assign n43140 = n43139 ^ n28005 ^ n1971 ;
  assign n43137 = n19322 | n23913 ;
  assign n43138 = ~n18252 & n43137 ;
  assign n43141 = n43140 ^ n43138 ^ 1'b0 ;
  assign n43146 = n7644 ^ n4098 ^ 1'b0 ;
  assign n43143 = n13039 | n38947 ;
  assign n43144 = n43143 ^ x192 ^ 1'b0 ;
  assign n43142 = n8237 | n11496 ;
  assign n43145 = n43144 ^ n43142 ^ 1'b0 ;
  assign n43147 = n43146 ^ n43145 ^ n3167 ;
  assign n43148 = ~n22244 & n43147 ;
  assign n43149 = n43148 ^ n18659 ^ 1'b0 ;
  assign n43150 = ~n305 & n21921 ;
  assign n43151 = n13488 ^ n11829 ^ 1'b0 ;
  assign n43152 = n7644 & n43151 ;
  assign n43153 = ~n6679 & n43152 ;
  assign n43154 = n41418 ^ n1093 ^ 1'b0 ;
  assign n43155 = n13588 ^ n7796 ^ n5295 ;
  assign n43156 = n25526 & ~n28752 ;
  assign n43157 = ~n21459 & n43156 ;
  assign n43158 = ( n1006 & ~n43155 ) | ( n1006 & n43157 ) | ( ~n43155 & n43157 ) ;
  assign n43159 = n9112 ^ n5895 ^ 1'b0 ;
  assign n43160 = n40523 ^ n11910 ^ 1'b0 ;
  assign n43161 = n12879 | n43160 ;
  assign n43162 = n27343 ^ n23104 ^ n12117 ;
  assign n43163 = n43161 | n43162 ;
  assign n43164 = n5112 & ~n36695 ;
  assign n43165 = n43164 ^ n11616 ^ n4589 ;
  assign n43166 = n26354 ^ n7466 ^ 1'b0 ;
  assign n43167 = n29400 & n43166 ;
  assign n43168 = ( n4004 & n14652 ) | ( n4004 & n43167 ) | ( n14652 & n43167 ) ;
  assign n43169 = ( ~n42736 & n43165 ) | ( ~n42736 & n43168 ) | ( n43165 & n43168 ) ;
  assign n43170 = n42859 ^ n24754 ^ 1'b0 ;
  assign n43171 = ~n43169 & n43170 ;
  assign n43173 = n30380 ^ n22126 ^ 1'b0 ;
  assign n43172 = n9399 & ~n15285 ;
  assign n43174 = n43173 ^ n43172 ^ n3905 ;
  assign n43175 = n8613 & n17875 ;
  assign n43176 = ( ~n21399 & n25190 ) | ( ~n21399 & n43175 ) | ( n25190 & n43175 ) ;
  assign n43177 = ( n18287 & n41981 ) | ( n18287 & n43176 ) | ( n41981 & n43176 ) ;
  assign n43178 = n16995 | n33519 ;
  assign n43179 = n19099 | n43178 ;
  assign n43180 = n8751 ^ n8301 ^ 1'b0 ;
  assign n43181 = ~n19928 & n43180 ;
  assign n43182 = n17982 | n43181 ;
  assign n43183 = n24189 | n43182 ;
  assign n43184 = n43179 & ~n43183 ;
  assign n43185 = ( ~n12933 & n14298 ) | ( ~n12933 & n22975 ) | ( n14298 & n22975 ) ;
  assign n43186 = n9079 ^ n736 ^ 1'b0 ;
  assign n43187 = ~n6549 & n43186 ;
  assign n43188 = n9765 | n10330 ;
  assign n43189 = n43188 ^ n15037 ^ 1'b0 ;
  assign n43190 = ~n25299 & n26248 ;
  assign n43191 = n6931 & n43190 ;
  assign n43192 = n7503 & ~n7678 ;
  assign n43193 = n7022 & n43192 ;
  assign n43195 = n12160 & ~n29312 ;
  assign n43196 = n23204 & n43195 ;
  assign n43194 = n20571 ^ n14493 ^ 1'b0 ;
  assign n43197 = n43196 ^ n43194 ^ n5561 ;
  assign n43198 = ( n20038 & n28545 ) | ( n20038 & n43197 ) | ( n28545 & n43197 ) ;
  assign n43199 = n14680 | n15949 ;
  assign n43200 = n43199 ^ n14618 ^ 1'b0 ;
  assign n43201 = n30895 | n43200 ;
  assign n43202 = n43201 ^ n23707 ^ 1'b0 ;
  assign n43203 = ( n2825 & n25995 ) | ( n2825 & ~n43202 ) | ( n25995 & ~n43202 ) ;
  assign n43204 = n21052 ^ n4514 ^ n3581 ;
  assign n43205 = ( n14833 & n19671 ) | ( n14833 & n24773 ) | ( n19671 & n24773 ) ;
  assign n43206 = n33773 ^ n22807 ^ 1'b0 ;
  assign n43207 = n22984 & ~n43206 ;
  assign n43208 = ( n15915 & n33839 ) | ( n15915 & ~n34749 ) | ( n33839 & ~n34749 ) ;
  assign n43209 = ( n28392 & n43207 ) | ( n28392 & n43208 ) | ( n43207 & n43208 ) ;
  assign n43210 = n18533 | n38820 ;
  assign n43211 = n43210 ^ n6672 ^ 1'b0 ;
  assign n43212 = n18519 ^ n716 ^ 1'b0 ;
  assign n43213 = ~n10487 & n19841 ;
  assign n43214 = ~n43212 & n43213 ;
  assign n43215 = n13398 & ~n21269 ;
  assign n43216 = n43215 ^ n10841 ^ 1'b0 ;
  assign n43217 = ~n9397 & n43216 ;
  assign n43218 = n43217 ^ n15661 ^ 1'b0 ;
  assign n43219 = n43218 ^ n10852 ^ 1'b0 ;
  assign n43220 = n10671 ^ n4876 ^ 1'b0 ;
  assign n43221 = n23929 ^ n23076 ^ 1'b0 ;
  assign n43222 = ( n1988 & ~n43220 ) | ( n1988 & n43221 ) | ( ~n43220 & n43221 ) ;
  assign n43223 = n43222 ^ n15506 ^ 1'b0 ;
  assign n43224 = n43223 ^ n16050 ^ 1'b0 ;
  assign n43225 = n10774 ^ n3692 ^ 1'b0 ;
  assign n43226 = n8965 ^ n1309 ^ 1'b0 ;
  assign n43227 = ~n1971 & n43226 ;
  assign n43228 = n11000 | n36197 ;
  assign n43229 = n43227 | n43228 ;
  assign n43230 = ~n37607 & n43229 ;
  assign n43231 = n18918 ^ n14653 ^ n10740 ;
  assign n43232 = ( n12391 & n15074 ) | ( n12391 & ~n43231 ) | ( n15074 & ~n43231 ) ;
  assign n43233 = n19815 ^ n15867 ^ 1'b0 ;
  assign n43234 = n27433 & ~n43233 ;
  assign n43235 = ( n33312 & ~n43232 ) | ( n33312 & n43234 ) | ( ~n43232 & n43234 ) ;
  assign n43236 = n22395 ^ n16824 ^ 1'b0 ;
  assign n43237 = n35393 ^ n4021 ^ n1184 ;
  assign n43238 = n43237 ^ n4059 ^ 1'b0 ;
  assign n43239 = n13412 & n43238 ;
  assign n43240 = n42892 ^ n3004 ^ 1'b0 ;
  assign n43241 = n43239 & n43240 ;
  assign n43242 = n3085 & n13103 ;
  assign n43243 = n43242 ^ n10655 ^ 1'b0 ;
  assign n43244 = n13925 | n43243 ;
  assign n43245 = n32574 | n43244 ;
  assign n43246 = n3202 | n7998 ;
  assign n43247 = n43246 ^ n14284 ^ 1'b0 ;
  assign n43248 = n43247 ^ n637 ^ 1'b0 ;
  assign n43249 = n7473 & n43248 ;
  assign n43250 = n41262 ^ n25217 ^ 1'b0 ;
  assign n43251 = n43250 ^ n40651 ^ n39256 ;
  assign n43252 = n34410 ^ n3404 ^ n1961 ;
  assign n43253 = ( n22944 & ~n26639 ) | ( n22944 & n37041 ) | ( ~n26639 & n37041 ) ;
  assign n43254 = ~n17739 & n29378 ;
  assign n43255 = ( n11437 & n21852 ) | ( n11437 & n22631 ) | ( n21852 & n22631 ) ;
  assign n43256 = n42196 ^ n9229 ^ 1'b0 ;
  assign n43257 = n5092 & n12217 ;
  assign n43259 = n13114 | n24526 ;
  assign n43260 = n43259 ^ n15608 ^ 1'b0 ;
  assign n43258 = ~n16390 & n16711 ;
  assign n43261 = n43260 ^ n43258 ^ n7463 ;
  assign n43262 = n41159 ^ n41150 ^ 1'b0 ;
  assign n43263 = ( ~n10258 & n13494 ) | ( ~n10258 & n19167 ) | ( n13494 & n19167 ) ;
  assign n43264 = n32400 ^ n10403 ^ 1'b0 ;
  assign n43265 = n15232 | n28188 ;
  assign n43266 = n43265 ^ n12862 ^ 1'b0 ;
  assign n43267 = n20231 ^ n6837 ^ 1'b0 ;
  assign n43268 = ~n11871 & n25058 ;
  assign n43269 = ( n7437 & n23626 ) | ( n7437 & ~n33542 ) | ( n23626 & ~n33542 ) ;
  assign n43270 = ( n14548 & n42781 ) | ( n14548 & n43269 ) | ( n42781 & n43269 ) ;
  assign n43271 = n33327 ^ n25635 ^ 1'b0 ;
  assign n43272 = ~n43270 & n43271 ;
  assign n43273 = n43272 ^ n29227 ^ n13655 ;
  assign n43274 = ( ~n11771 & n26823 ) | ( ~n11771 & n30202 ) | ( n26823 & n30202 ) ;
  assign n43275 = n35415 | n35829 ;
  assign n43276 = n43275 ^ n35838 ^ n9295 ;
  assign n43277 = n12726 ^ n5051 ^ 1'b0 ;
  assign n43278 = n29789 | n43277 ;
  assign n43279 = n12688 | n18250 ;
  assign n43280 = ( n15687 & n21965 ) | ( n15687 & n24396 ) | ( n21965 & n24396 ) ;
  assign n43281 = n515 & ~n43280 ;
  assign n43282 = ~n6427 & n43281 ;
  assign n43283 = n43279 | n43282 ;
  assign n43284 = n25744 ^ n24192 ^ n13789 ;
  assign n43285 = n43284 ^ n3113 ^ 1'b0 ;
  assign n43286 = ~n11246 & n43285 ;
  assign n43287 = ( n2986 & ~n25974 ) | ( n2986 & n43286 ) | ( ~n25974 & n43286 ) ;
  assign n43288 = n19762 ^ n7444 ^ 1'b0 ;
  assign n43289 = n43288 ^ n42277 ^ n36012 ;
  assign n43290 = ~n10910 & n43289 ;
  assign n43291 = n13393 ^ n9448 ^ n471 ;
  assign n43292 = ( n2368 & n8824 ) | ( n2368 & n9701 ) | ( n8824 & n9701 ) ;
  assign n43293 = ~n9463 & n24974 ;
  assign n43294 = n43293 ^ n16005 ^ 1'b0 ;
  assign n43295 = n43294 ^ n9506 ^ n4452 ;
  assign n43296 = n20507 | n32516 ;
  assign n43297 = n43296 ^ n492 ^ 1'b0 ;
  assign n43298 = n7184 ^ x67 ^ 1'b0 ;
  assign n43299 = n26430 ^ n26131 ^ 1'b0 ;
  assign n43300 = n43298 & n43299 ;
  assign n43301 = ( n1226 & n23414 ) | ( n1226 & ~n37238 ) | ( n23414 & ~n37238 ) ;
  assign n43302 = n43301 ^ n14766 ^ 1'b0 ;
  assign n43303 = ~n8692 & n43302 ;
  assign n43304 = ( n1405 & ~n23882 ) | ( n1405 & n30738 ) | ( ~n23882 & n30738 ) ;
  assign n43305 = n13882 & ~n21078 ;
  assign n43306 = n14672 & n43305 ;
  assign n43307 = n43304 | n43306 ;
  assign n43308 = ( n1910 & n15638 ) | ( n1910 & n43307 ) | ( n15638 & n43307 ) ;
  assign n43309 = n27474 | n43308 ;
  assign n43310 = n19028 ^ n14633 ^ n2260 ;
  assign n43311 = n30542 ^ n15816 ^ 1'b0 ;
  assign n43312 = n39707 ^ n36527 ^ n4827 ;
  assign n43313 = ~n2735 & n34033 ;
  assign n43314 = ( n9876 & n11809 ) | ( n9876 & n25541 ) | ( n11809 & n25541 ) ;
  assign n43315 = n43314 ^ n12919 ^ 1'b0 ;
  assign n43316 = n26538 ^ n7910 ^ 1'b0 ;
  assign n43317 = ~n43315 & n43316 ;
  assign n43318 = n24948 & ~n41471 ;
  assign n43322 = n11623 ^ n2771 ^ 1'b0 ;
  assign n43319 = n3466 & ~n17096 ;
  assign n43320 = ~n42205 & n43319 ;
  assign n43321 = n38336 & ~n43320 ;
  assign n43323 = n43322 ^ n43321 ^ 1'b0 ;
  assign n43324 = n22039 ^ n18811 ^ 1'b0 ;
  assign n43325 = ~n43323 & n43324 ;
  assign n43326 = n18482 ^ n7814 ^ 1'b0 ;
  assign n43327 = n36779 ^ n21317 ^ n1932 ;
  assign n43328 = n7758 ^ n2796 ^ 1'b0 ;
  assign n43329 = n33400 ^ n23363 ^ n18479 ;
  assign n43330 = ( n4217 & n9553 ) | ( n4217 & n29067 ) | ( n9553 & n29067 ) ;
  assign n43331 = n23376 ^ n4803 ^ 1'b0 ;
  assign n43332 = n43331 ^ n24287 ^ 1'b0 ;
  assign n43333 = ( ~n10613 & n43330 ) | ( ~n10613 & n43332 ) | ( n43330 & n43332 ) ;
  assign n43334 = n22761 & n43333 ;
  assign n43335 = n9780 & ~n33758 ;
  assign n43336 = n43335 ^ n27206 ^ 1'b0 ;
  assign n43337 = n21784 & ~n39849 ;
  assign n43338 = n30049 ^ n11209 ^ n947 ;
  assign n43339 = n26257 & ~n43338 ;
  assign n43340 = n26457 ^ n7318 ^ 1'b0 ;
  assign n43341 = ~n2886 & n43340 ;
  assign n43342 = n43341 ^ n41157 ^ n31823 ;
  assign n43343 = n43342 ^ n33919 ^ n15362 ;
  assign n43344 = ( ~n1811 & n19973 ) | ( ~n1811 & n31137 ) | ( n19973 & n31137 ) ;
  assign n43345 = n20136 ^ n4950 ^ 1'b0 ;
  assign n43346 = n12117 | n43345 ;
  assign n43347 = n35113 ^ n11495 ^ n11007 ;
  assign n43348 = n21429 & ~n43347 ;
  assign n43349 = n7043 & n43348 ;
  assign n43350 = n35866 ^ n18144 ^ n6294 ;
  assign n43351 = n43350 ^ n15973 ^ 1'b0 ;
  assign n43352 = ( n43346 & n43349 ) | ( n43346 & n43351 ) | ( n43349 & n43351 ) ;
  assign n43353 = n3225 & n37431 ;
  assign n43354 = n43353 ^ n17601 ^ 1'b0 ;
  assign n43357 = n14325 ^ n10936 ^ 1'b0 ;
  assign n43355 = n19612 ^ n7719 ^ 1'b0 ;
  assign n43356 = n488 & n43355 ;
  assign n43358 = n43357 ^ n43356 ^ n9643 ;
  assign n43359 = n10173 & n43358 ;
  assign n43360 = n43354 & ~n43359 ;
  assign n43361 = ~n1217 & n29497 ;
  assign n43362 = n28894 & n43361 ;
  assign n43363 = n15724 ^ n686 ^ 1'b0 ;
  assign n43364 = n34318 & n43363 ;
  assign n43365 = n41410 ^ n11025 ^ 1'b0 ;
  assign n43366 = n6800 & ~n31290 ;
  assign n43367 = n43366 ^ n38795 ^ 1'b0 ;
  assign n43368 = n42245 ^ n21825 ^ n5301 ;
  assign n43369 = n33370 ^ n20710 ^ n4289 ;
  assign n43370 = n12617 ^ n4852 ^ 1'b0 ;
  assign n43371 = n2925 & n23184 ;
  assign n43372 = n30012 & n43371 ;
  assign n43373 = n19033 ^ n2208 ^ 1'b0 ;
  assign n43374 = n41477 | n43373 ;
  assign n43375 = n23164 ^ n5625 ^ 1'b0 ;
  assign n43376 = n35189 | n43375 ;
  assign n43377 = n10569 | n17960 ;
  assign n43378 = n43377 ^ n27799 ^ n14625 ;
  assign n43379 = ( n1823 & n27844 ) | ( n1823 & n36097 ) | ( n27844 & n36097 ) ;
  assign n43380 = n39169 ^ n8247 ^ 1'b0 ;
  assign n43381 = ( ~n6445 & n8727 ) | ( ~n6445 & n32258 ) | ( n8727 & n32258 ) ;
  assign n43382 = n17320 | n43381 ;
  assign n43383 = n14648 | n36958 ;
  assign n43384 = n43383 ^ n16744 ^ 1'b0 ;
  assign n43385 = ~n6345 & n11327 ;
  assign n43386 = ~n20179 & n43385 ;
  assign n43387 = ~n997 & n3301 ;
  assign n43388 = ~n5003 & n43387 ;
  assign n43389 = n43388 ^ n2723 ^ 1'b0 ;
  assign n43390 = n8450 & ~n17568 ;
  assign n43391 = n43390 ^ n7803 ^ 1'b0 ;
  assign n43392 = n21225 ^ n11858 ^ n4455 ;
  assign n43393 = ( n2425 & n34566 ) | ( n2425 & ~n40131 ) | ( n34566 & ~n40131 ) ;
  assign n43394 = ( n13676 & ~n19995 ) | ( n13676 & n43393 ) | ( ~n19995 & n43393 ) ;
  assign n43395 = n7600 & n12803 ;
  assign n43396 = n43395 ^ n22675 ^ 1'b0 ;
  assign n43397 = ( n40728 & n41966 ) | ( n40728 & ~n43396 ) | ( n41966 & ~n43396 ) ;
  assign n43398 = n43397 ^ n914 ^ 1'b0 ;
  assign n43399 = n12847 ^ n8179 ^ 1'b0 ;
  assign n43400 = ~n23695 & n43399 ;
  assign n43401 = ~n43399 & n43400 ;
  assign n43402 = n7203 & n14021 ;
  assign n43403 = ~n7203 & n43402 ;
  assign n43404 = n3212 | n43403 ;
  assign n43405 = n3212 & ~n43404 ;
  assign n43406 = n43405 ^ n26045 ^ 1'b0 ;
  assign n43407 = ~n43401 & n43406 ;
  assign n43408 = n21869 ^ n19620 ^ 1'b0 ;
  assign n43409 = n9658 & ~n43408 ;
  assign n43410 = n29522 ^ n1674 ^ 1'b0 ;
  assign n43411 = ~n16507 & n43410 ;
  assign n43412 = n43108 ^ n8124 ^ 1'b0 ;
  assign n43413 = ~n22053 & n43412 ;
  assign n43414 = n43413 ^ n2571 ^ 1'b0 ;
  assign n43415 = n43414 ^ n37938 ^ n30190 ;
  assign n43420 = ( n8597 & n9139 ) | ( n8597 & ~n12069 ) | ( n9139 & ~n12069 ) ;
  assign n43416 = n279 | n5763 ;
  assign n43417 = n43416 ^ n7770 ^ 1'b0 ;
  assign n43418 = n16736 & n23447 ;
  assign n43419 = n43417 & n43418 ;
  assign n43421 = n43420 ^ n43419 ^ n9910 ;
  assign n43422 = n6428 & ~n15365 ;
  assign n43423 = n16222 & n43422 ;
  assign n43424 = ( ~n2931 & n12977 ) | ( ~n2931 & n24138 ) | ( n12977 & n24138 ) ;
  assign n43425 = n41882 ^ n1056 ^ 1'b0 ;
  assign n43426 = n30481 & n43425 ;
  assign n43427 = ( n1427 & n6425 ) | ( n1427 & n34226 ) | ( n6425 & n34226 ) ;
  assign n43428 = ~n10911 & n43427 ;
  assign n43429 = n2571 | n43428 ;
  assign n43430 = n24776 ^ n22557 ^ n4592 ;
  assign n43431 = n26000 ^ n19663 ^ n14706 ;
  assign n43432 = n35129 ^ n12733 ^ 1'b0 ;
  assign n43433 = n35439 ^ x152 ^ 1'b0 ;
  assign n43434 = ( n10659 & n37865 ) | ( n10659 & ~n43433 ) | ( n37865 & ~n43433 ) ;
  assign n43435 = n29534 ^ n7270 ^ 1'b0 ;
  assign n43436 = n2444 & ~n10432 ;
  assign n43438 = ( ~n7579 & n24388 ) | ( ~n7579 & n38145 ) | ( n24388 & n38145 ) ;
  assign n43437 = n1211 | n9328 ;
  assign n43439 = n43438 ^ n43437 ^ 1'b0 ;
  assign n43440 = n2080 & ~n4183 ;
  assign n43441 = n43440 ^ n33561 ^ 1'b0 ;
  assign n43442 = ( ~n25501 & n31737 ) | ( ~n25501 & n43441 ) | ( n31737 & n43441 ) ;
  assign n43443 = n28036 ^ n9703 ^ 1'b0 ;
  assign n43444 = n43442 | n43443 ;
  assign n43445 = n22037 ^ n3765 ^ 1'b0 ;
  assign n43446 = n7626 & ~n43445 ;
  assign n43447 = n14735 ^ n14686 ^ n9172 ;
  assign n43448 = n3813 & ~n13137 ;
  assign n43449 = n43448 ^ n29765 ^ 1'b0 ;
  assign n43450 = ( n677 & ~n4435 ) | ( n677 & n43449 ) | ( ~n4435 & n43449 ) ;
  assign n43451 = n23749 & n34167 ;
  assign n43452 = n17183 | n43451 ;
  assign n43453 = ~n13115 & n13987 ;
  assign n43454 = n9190 & ~n30543 ;
  assign n43455 = n33305 ^ n8924 ^ 1'b0 ;
  assign n43456 = n43455 ^ n11326 ^ 1'b0 ;
  assign n43457 = ~n5994 & n7317 ;
  assign n43458 = n15394 & ~n43457 ;
  assign n43460 = ~n10026 & n13075 ;
  assign n43461 = n43460 ^ n14872 ^ 1'b0 ;
  assign n43462 = n29976 ^ n7564 ^ n3127 ;
  assign n43463 = n8295 & ~n43462 ;
  assign n43464 = ( n4215 & ~n43461 ) | ( n4215 & n43463 ) | ( ~n43461 & n43463 ) ;
  assign n43459 = n7221 & n41288 ;
  assign n43465 = n43464 ^ n43459 ^ 1'b0 ;
  assign n43466 = n25791 | n43465 ;
  assign n43467 = n13819 & ~n35527 ;
  assign n43468 = ~n3561 & n43467 ;
  assign n43469 = n8458 | n9250 ;
  assign n43470 = n43468 & ~n43469 ;
  assign n43471 = ~n6150 & n7270 ;
  assign n43472 = n34397 ^ n19369 ^ 1'b0 ;
  assign n43473 = n13412 & ~n43472 ;
  assign n43474 = n43473 ^ n15777 ^ 1'b0 ;
  assign n43475 = n43474 ^ n26518 ^ n24597 ;
  assign n43476 = n24527 ^ n645 ^ 1'b0 ;
  assign n43477 = n43476 ^ n32830 ^ 1'b0 ;
  assign n43478 = ( n8769 & ~n11150 ) | ( n8769 & n13233 ) | ( ~n11150 & n13233 ) ;
  assign n43479 = ( ~n4741 & n42569 ) | ( ~n4741 & n43478 ) | ( n42569 & n43478 ) ;
  assign n43480 = n29478 ^ n26042 ^ n15995 ;
  assign n43481 = ( ~n7177 & n39603 ) | ( ~n7177 & n43480 ) | ( n39603 & n43480 ) ;
  assign n43482 = n15632 ^ n11095 ^ 1'b0 ;
  assign n43483 = n30182 ^ n23645 ^ n4748 ;
  assign n43484 = ~n33944 & n43483 ;
  assign n43485 = n378 & ~n42693 ;
  assign n43486 = n43484 | n43485 ;
  assign n43490 = n20338 ^ n10076 ^ n6793 ;
  assign n43487 = n21401 | n33634 ;
  assign n43488 = n11072 & ~n43487 ;
  assign n43489 = n19650 & ~n43488 ;
  assign n43491 = n43490 ^ n43489 ^ 1'b0 ;
  assign n43492 = n15203 ^ n10517 ^ 1'b0 ;
  assign n43493 = n23019 & n39996 ;
  assign n43494 = n43076 & n43493 ;
  assign n43495 = ( n28887 & n42267 ) | ( n28887 & ~n43494 ) | ( n42267 & ~n43494 ) ;
  assign n43496 = n5767 & n31947 ;
  assign n43497 = n12276 ^ n2397 ^ 1'b0 ;
  assign n43498 = n16927 ^ n7473 ^ 1'b0 ;
  assign n43499 = n9661 & n43498 ;
  assign n43500 = ( n8364 & n12728 ) | ( n8364 & n43499 ) | ( n12728 & n43499 ) ;
  assign n43501 = n14010 ^ x18 ^ 1'b0 ;
  assign n43502 = n20579 & ~n43501 ;
  assign n43503 = n43502 ^ n28743 ^ n16982 ;
  assign n43504 = n3171 | n12302 ;
  assign n43505 = ~n16074 & n43504 ;
  assign n43506 = n24198 ^ n18680 ^ n7300 ;
  assign n43507 = n4720 ^ n785 ^ 1'b0 ;
  assign n43508 = n43507 ^ n41173 ^ n25639 ;
  assign n43509 = n37145 ^ n31427 ^ 1'b0 ;
  assign n43514 = n26519 ^ n19565 ^ 1'b0 ;
  assign n43510 = n16273 | n18838 ;
  assign n43511 = n43510 ^ n21831 ^ 1'b0 ;
  assign n43512 = ( ~n11374 & n30313 ) | ( ~n11374 & n43511 ) | ( n30313 & n43511 ) ;
  assign n43513 = n43512 ^ n9722 ^ n3717 ;
  assign n43515 = n43514 ^ n43513 ^ 1'b0 ;
  assign n43516 = n9423 & n43515 ;
  assign n43517 = n15959 & ~n30925 ;
  assign n43518 = n43517 ^ n38478 ^ 1'b0 ;
  assign n43519 = ( ~n9449 & n27659 ) | ( ~n9449 & n36041 ) | ( n27659 & n36041 ) ;
  assign n43520 = n21158 & ~n43519 ;
  assign n43521 = n43520 ^ n34757 ^ 1'b0 ;
  assign n43522 = n13969 ^ n8940 ^ n1057 ;
  assign n43523 = n43522 ^ n41309 ^ n23283 ;
  assign n43524 = n22696 ^ n14050 ^ 1'b0 ;
  assign n43525 = n15922 & ~n31831 ;
  assign n43526 = ( ~n28800 & n41225 ) | ( ~n28800 & n43525 ) | ( n41225 & n43525 ) ;
  assign n43527 = n3000 & n12640 ;
  assign n43528 = n43527 ^ n16828 ^ n2448 ;
  assign n43529 = n9953 & ~n25927 ;
  assign n43530 = n24923 & n43529 ;
  assign n43531 = ( n632 & n9654 ) | ( n632 & n43530 ) | ( n9654 & n43530 ) ;
  assign n43532 = n28767 ^ n5502 ^ 1'b0 ;
  assign n43533 = n42465 | n43532 ;
  assign n43534 = n43533 ^ n9294 ^ 1'b0 ;
  assign n43535 = ( n13599 & n20588 ) | ( n13599 & ~n31972 ) | ( n20588 & ~n31972 ) ;
  assign n43536 = n43535 ^ n19065 ^ 1'b0 ;
  assign n43537 = n43455 & n43536 ;
  assign n43538 = n43537 ^ n21921 ^ 1'b0 ;
  assign n43539 = ~n30605 & n43538 ;
  assign n43543 = ( n11872 & n14077 ) | ( n11872 & n35156 ) | ( n14077 & n35156 ) ;
  assign n43541 = n18620 ^ n4907 ^ n3668 ;
  assign n43542 = n36368 & n43541 ;
  assign n43544 = n43543 ^ n43542 ^ 1'b0 ;
  assign n43545 = n7544 & n43544 ;
  assign n43546 = n8538 & n43545 ;
  assign n43540 = n15294 & ~n19047 ;
  assign n43547 = n43546 ^ n43540 ^ 1'b0 ;
  assign n43548 = n43283 ^ n17477 ^ 1'b0 ;
  assign n43549 = ~n8153 & n43548 ;
  assign n43550 = n27842 ^ n3734 ^ 1'b0 ;
  assign n43551 = n36887 ^ n15798 ^ n14764 ;
  assign n43552 = ~n12388 & n14341 ;
  assign n43553 = ( n16345 & ~n38518 ) | ( n16345 & n43552 ) | ( ~n38518 & n43552 ) ;
  assign n43554 = n25760 ^ n6049 ^ 1'b0 ;
  assign n43555 = n42302 & ~n43554 ;
  assign n43556 = n18245 | n39228 ;
  assign n43557 = n36118 ^ n29509 ^ 1'b0 ;
  assign n43558 = n25129 & n43557 ;
  assign n43559 = n28210 ^ n26714 ^ 1'b0 ;
  assign n43561 = ( n6111 & ~n15660 ) | ( n6111 & n38330 ) | ( ~n15660 & n38330 ) ;
  assign n43560 = n29598 & ~n35800 ;
  assign n43562 = n43561 ^ n43560 ^ n29414 ;
  assign n43563 = ( n1966 & n13433 ) | ( n1966 & n14314 ) | ( n13433 & n14314 ) ;
  assign n43564 = n38663 & ~n43563 ;
  assign n43565 = ~n16883 & n43247 ;
  assign n43566 = n10483 ^ n361 ^ 1'b0 ;
  assign n43567 = n8945 | n43566 ;
  assign n43568 = n3278 & n5188 ;
  assign n43569 = n43568 ^ n7860 ^ 1'b0 ;
  assign n43570 = n1706 | n24841 ;
  assign n43571 = ( n5716 & n43569 ) | ( n5716 & ~n43570 ) | ( n43569 & ~n43570 ) ;
  assign n43572 = n15831 ^ n6393 ^ 1'b0 ;
  assign n43573 = n43572 ^ n4217 ^ 1'b0 ;
  assign n43574 = n43571 & n43573 ;
  assign n43575 = n27470 ^ n18438 ^ n6369 ;
  assign n43576 = n23373 & n43575 ;
  assign n43577 = ~n757 & n43576 ;
  assign n43578 = n17189 | n43577 ;
  assign n43579 = n43578 ^ n42847 ^ 1'b0 ;
  assign n43580 = n37570 ^ n37552 ^ n24529 ;
  assign n43581 = n4132 & n6133 ;
  assign n43582 = ( n9794 & n24530 ) | ( n9794 & ~n43581 ) | ( n24530 & ~n43581 ) ;
  assign n43583 = n29321 ^ n21470 ^ 1'b0 ;
  assign n43584 = ( n3129 & n30239 ) | ( n3129 & ~n43583 ) | ( n30239 & ~n43583 ) ;
  assign n43585 = n42082 & n43584 ;
  assign n43586 = ( n9286 & ~n12168 ) | ( n9286 & n24145 ) | ( ~n12168 & n24145 ) ;
  assign n43587 = n43586 ^ n37290 ^ n15551 ;
  assign n43588 = n13535 & ~n29876 ;
  assign n43589 = ~n43587 & n43588 ;
  assign n43590 = ~n9612 & n32529 ;
  assign n43591 = n43590 ^ n13341 ^ 1'b0 ;
  assign n43592 = ~n6803 & n17754 ;
  assign n43593 = n43592 ^ n20207 ^ 1'b0 ;
  assign n43594 = n18541 ^ n16794 ^ 1'b0 ;
  assign n43595 = ~n17891 & n43594 ;
  assign n43596 = ( ~n5984 & n20100 ) | ( ~n5984 & n23573 ) | ( n20100 & n23573 ) ;
  assign n43597 = ~n4095 & n24214 ;
  assign n43598 = ~n43596 & n43597 ;
  assign n43599 = n2689 | n3632 ;
  assign n43600 = n43599 ^ n730 ^ 1'b0 ;
  assign n43601 = n43600 ^ n9566 ^ 1'b0 ;
  assign n43602 = ( n13289 & ~n17617 ) | ( n13289 & n29714 ) | ( ~n17617 & n29714 ) ;
  assign n43605 = n20763 ^ n20505 ^ n7051 ;
  assign n43603 = ~n6949 & n25445 ;
  assign n43604 = n43603 ^ n21162 ^ 1'b0 ;
  assign n43606 = n43605 ^ n43604 ^ n19290 ;
  assign n43607 = n32965 ^ n12270 ^ n3501 ;
  assign n43608 = n32412 ^ n23782 ^ 1'b0 ;
  assign n43609 = n16437 | n26813 ;
  assign n43610 = n35830 & ~n43609 ;
  assign n43611 = n11445 & ~n16548 ;
  assign n43612 = n43611 ^ n31776 ^ 1'b0 ;
  assign n43613 = ( n2522 & n9240 ) | ( n2522 & ~n21367 ) | ( n9240 & ~n21367 ) ;
  assign n43614 = n20592 ^ n3469 ^ 1'b0 ;
  assign n43615 = n3149 & ~n43614 ;
  assign n43616 = ( ~n12111 & n13005 ) | ( ~n12111 & n22559 ) | ( n13005 & n22559 ) ;
  assign n43617 = n5443 & ~n14051 ;
  assign n43618 = n43617 ^ n37677 ^ n32933 ;
  assign n43619 = ( n2218 & n4840 ) | ( n2218 & n30702 ) | ( n4840 & n30702 ) ;
  assign n43620 = n5820 ^ n573 ^ 1'b0 ;
  assign n43621 = n7304 & n27299 ;
  assign n43622 = ~n43620 & n43621 ;
  assign n43623 = n26492 ^ n25966 ^ 1'b0 ;
  assign n43624 = ~n8858 & n43623 ;
  assign n43625 = n3510 & n43624 ;
  assign n43626 = n37813 ^ n3518 ^ 1'b0 ;
  assign n43627 = n33577 & n43626 ;
  assign n43628 = ~n32936 & n42157 ;
  assign n43629 = ~n22634 & n43628 ;
  assign n43630 = n4604 & n13788 ;
  assign n43631 = ~n24094 & n43630 ;
  assign n43632 = n43631 ^ n26142 ^ 1'b0 ;
  assign n43633 = n25314 ^ n18759 ^ n12733 ;
  assign n43634 = n35527 ^ n33576 ^ n10026 ;
  assign n43635 = n13273 & n43173 ;
  assign n43636 = n4224 & ~n23771 ;
  assign n43637 = ~n10167 & n43636 ;
  assign n43638 = n11924 & n43637 ;
  assign n43639 = n13316 & ~n30989 ;
  assign n43640 = n34168 ^ n24669 ^ 1'b0 ;
  assign n43641 = n43639 | n43640 ;
  assign n43642 = n10645 & n18308 ;
  assign n43643 = ( ~n8012 & n34397 ) | ( ~n8012 & n43642 ) | ( n34397 & n43642 ) ;
  assign n43644 = n43643 ^ n10857 ^ 1'b0 ;
  assign n43645 = n38619 ^ n24765 ^ n5635 ;
  assign n43646 = n43645 ^ n39975 ^ n17779 ;
  assign n43647 = n483 & ~n11557 ;
  assign n43648 = n43647 ^ n27116 ^ n4060 ;
  assign n43649 = n40906 ^ n23920 ^ n6942 ;
  assign n43650 = n43649 ^ n18917 ^ 1'b0 ;
  assign n43651 = n28259 | n43650 ;
  assign n43652 = n6049 | n17490 ;
  assign n43653 = n11325 & ~n43652 ;
  assign n43654 = n11213 & ~n25476 ;
  assign n43655 = n43654 ^ n7170 ^ 1'b0 ;
  assign n43656 = ( n4434 & n12254 ) | ( n4434 & ~n13301 ) | ( n12254 & ~n13301 ) ;
  assign n43657 = n19263 ^ n3639 ^ 1'b0 ;
  assign n43658 = n43656 | n43657 ;
  assign n43659 = ( ~n1292 & n6538 ) | ( ~n1292 & n9401 ) | ( n6538 & n9401 ) ;
  assign n43660 = ~n4652 & n43659 ;
  assign n43661 = n39282 ^ n13270 ^ n6712 ;
  assign n43665 = n2506 & n39065 ;
  assign n43666 = ~n37505 & n43665 ;
  assign n43662 = n5702 & ~n16969 ;
  assign n43663 = ~n23573 & n43662 ;
  assign n43664 = n43663 ^ n1075 ^ 1'b0 ;
  assign n43667 = n43666 ^ n43664 ^ n13116 ;
  assign n43668 = n20536 ^ n7480 ^ 1'b0 ;
  assign n43669 = n9881 | n27933 ;
  assign n43670 = n5733 | n43669 ;
  assign n43671 = n9654 | n43670 ;
  assign n43672 = n14140 ^ n4108 ^ 1'b0 ;
  assign n43673 = n43671 & n43672 ;
  assign n43678 = ( ~n7635 & n18422 ) | ( ~n7635 & n22752 ) | ( n18422 & n22752 ) ;
  assign n43674 = n19547 & ~n26619 ;
  assign n43675 = n1270 & n43674 ;
  assign n43676 = ~n39705 & n43675 ;
  assign n43677 = ( ~n9223 & n14281 ) | ( ~n9223 & n43676 ) | ( n14281 & n43676 ) ;
  assign n43679 = n43678 ^ n43677 ^ 1'b0 ;
  assign n43680 = ~x5 & n9661 ;
  assign n43681 = n43680 ^ n34319 ^ 1'b0 ;
  assign n43682 = n5663 & n43681 ;
  assign n43683 = ~n43679 & n43682 ;
  assign n43684 = n13545 ^ n8588 ^ 1'b0 ;
  assign n43685 = n43684 ^ n9790 ^ n8634 ;
  assign n43686 = n43685 ^ n33435 ^ 1'b0 ;
  assign n43687 = ~n21619 & n33645 ;
  assign n43688 = ( n17031 & n26227 ) | ( n17031 & ~n33148 ) | ( n26227 & ~n33148 ) ;
  assign n43689 = n7786 | n14740 ;
  assign n43690 = n382 & ~n13583 ;
  assign n43691 = n27510 & n43690 ;
  assign n43692 = n43691 ^ n38990 ^ n22235 ;
  assign n43693 = n29902 ^ n25323 ^ 1'b0 ;
  assign n43694 = n40026 ^ n7020 ^ n6442 ;
  assign n43695 = n23627 & ~n28250 ;
  assign n43696 = ~n13987 & n43695 ;
  assign n43697 = ( ~n3093 & n3550 ) | ( ~n3093 & n43696 ) | ( n3550 & n43696 ) ;
  assign n43698 = ( ~n13456 & n21554 ) | ( ~n13456 & n29074 ) | ( n21554 & n29074 ) ;
  assign n43699 = n43698 ^ n20905 ^ n18825 ;
  assign n43700 = ~n18518 & n43699 ;
  assign n43701 = n15857 ^ n15595 ^ n1986 ;
  assign n43702 = n18441 | n43701 ;
  assign n43703 = ( ~n10494 & n12782 ) | ( ~n10494 & n29040 ) | ( n12782 & n29040 ) ;
  assign n43704 = ( n6895 & n15556 ) | ( n6895 & ~n43703 ) | ( n15556 & ~n43703 ) ;
  assign n43705 = ~n900 & n8913 ;
  assign n43706 = n43704 & n43705 ;
  assign n43707 = ~n11371 & n13628 ;
  assign n43708 = n43706 & n43707 ;
  assign n43709 = ( n8569 & n32770 ) | ( n8569 & n39858 ) | ( n32770 & n39858 ) ;
  assign n43710 = n3292 ^ n2571 ^ 1'b0 ;
  assign n43713 = n9139 | n11411 ;
  assign n43712 = n22439 ^ n9992 ^ 1'b0 ;
  assign n43711 = n4869 & ~n25740 ;
  assign n43714 = n43713 ^ n43712 ^ n43711 ;
  assign n43715 = n22921 ^ n7036 ^ 1'b0 ;
  assign n43716 = n7551 & n43304 ;
  assign n43717 = ~n11671 & n43716 ;
  assign n43718 = ( n10069 & ~n10579 ) | ( n10069 & n43717 ) | ( ~n10579 & n43717 ) ;
  assign n43719 = n9542 ^ n6773 ^ n6005 ;
  assign n43720 = n37538 & ~n43719 ;
  assign n43721 = n43720 ^ n27793 ^ 1'b0 ;
  assign n43722 = n13364 ^ n3126 ^ 1'b0 ;
  assign n43723 = n43721 | n43722 ;
  assign n43724 = ( n11008 & n19038 ) | ( n11008 & n19311 ) | ( n19038 & n19311 ) ;
  assign n43725 = ~n36207 & n43724 ;
  assign n43726 = n43725 ^ n7577 ^ 1'b0 ;
  assign n43727 = ( n958 & ~n12020 ) | ( n958 & n22711 ) | ( ~n12020 & n22711 ) ;
  assign n43728 = n43727 ^ n28021 ^ 1'b0 ;
  assign n43729 = n20873 | n43728 ;
  assign n43730 = n43729 ^ n8663 ^ 1'b0 ;
  assign n43731 = ( n31610 & n35507 ) | ( n31610 & n43730 ) | ( n35507 & n43730 ) ;
  assign n43732 = n43731 ^ n32911 ^ 1'b0 ;
  assign n43733 = n20008 & ~n43732 ;
  assign n43734 = n31791 & n33298 ;
  assign n43735 = n7071 & ~n20660 ;
  assign n43736 = ~n43734 & n43735 ;
  assign n43737 = n5499 & ~n8306 ;
  assign n43738 = ~n12167 & n19785 ;
  assign n43739 = n43738 ^ n7412 ^ 1'b0 ;
  assign n43740 = ( n33461 & n43737 ) | ( n33461 & ~n43739 ) | ( n43737 & ~n43739 ) ;
  assign n43741 = x81 | n43740 ;
  assign n43742 = n43741 ^ n31097 ^ 1'b0 ;
  assign n43743 = n43742 ^ n32590 ^ n9803 ;
  assign n43744 = n27242 ^ n9779 ^ n2093 ;
  assign n43745 = ~n43743 & n43744 ;
  assign n43746 = n11706 ^ n10663 ^ n7163 ;
  assign n43747 = n18484 | n43746 ;
  assign n43748 = ( ~n16301 & n31189 ) | ( ~n16301 & n35080 ) | ( n31189 & n35080 ) ;
  assign n43752 = n11013 | n25779 ;
  assign n43753 = n43752 ^ n28230 ^ 1'b0 ;
  assign n43750 = n25858 ^ n11715 ^ 1'b0 ;
  assign n43751 = n43750 ^ n27888 ^ n24744 ;
  assign n43754 = n43753 ^ n43751 ^ n29171 ;
  assign n43749 = n16626 ^ n6326 ^ n2680 ;
  assign n43755 = n43754 ^ n43749 ^ 1'b0 ;
  assign n43756 = n23950 ^ n13002 ^ n11454 ;
  assign n43757 = n22173 ^ n17856 ^ n4315 ;
  assign n43758 = n26134 & ~n43757 ;
  assign n43759 = n43758 ^ n12503 ^ 1'b0 ;
  assign n43760 = n25033 ^ n18649 ^ 1'b0 ;
  assign n43761 = n1267 | n43760 ;
  assign n43762 = n7326 & n8951 ;
  assign n43763 = n43762 ^ n26458 ^ 1'b0 ;
  assign n43764 = n30114 ^ n3156 ^ 1'b0 ;
  assign n43765 = n43763 | n43764 ;
  assign n43767 = n19005 & n34081 ;
  assign n43768 = n43767 ^ n32960 ^ n18774 ;
  assign n43766 = n20528 & n22153 ;
  assign n43769 = n43768 ^ n43766 ^ 1'b0 ;
  assign n43770 = ( n15953 & n22767 ) | ( n15953 & ~n30635 ) | ( n22767 & ~n30635 ) ;
  assign n43771 = n10137 & n22004 ;
  assign n43772 = n43771 ^ n11030 ^ 1'b0 ;
  assign n43773 = n43772 ^ n41712 ^ n21386 ;
  assign n43774 = x74 | n4465 ;
  assign n43775 = n35222 & ~n43774 ;
  assign n43777 = ~n10009 & n21500 ;
  assign n43776 = n5291 & ~n17427 ;
  assign n43778 = n43777 ^ n43776 ^ n16484 ;
  assign n43779 = n8358 | n17187 ;
  assign n43780 = n43778 | n43779 ;
  assign n43781 = ( ~n6304 & n43775 ) | ( ~n6304 & n43780 ) | ( n43775 & n43780 ) ;
  assign n43782 = n3353 & ~n11847 ;
  assign n43783 = ( n19834 & n38780 ) | ( n19834 & n43782 ) | ( n38780 & n43782 ) ;
  assign n43784 = n15520 ^ n8657 ^ 1'b0 ;
  assign n43785 = n43784 ^ n18643 ^ 1'b0 ;
  assign n43786 = ~n9432 & n43785 ;
  assign n43787 = n20100 & n43786 ;
  assign n43788 = n39117 ^ n32483 ^ n14300 ;
  assign n43789 = n43788 ^ n43050 ^ n23619 ;
  assign n43790 = ( n2087 & n19999 ) | ( n2087 & n28200 ) | ( n19999 & n28200 ) ;
  assign n43791 = n42577 ^ n14206 ^ n6121 ;
  assign n43792 = n43790 & n43791 ;
  assign n43793 = n4912 ^ n3002 ^ 1'b0 ;
  assign n43794 = n9145 & n43793 ;
  assign n43795 = n29374 ^ n7791 ^ n5416 ;
  assign n43798 = n8042 & ~n8465 ;
  assign n43799 = ~n7922 & n43798 ;
  assign n43796 = n28179 ^ n8122 ^ 1'b0 ;
  assign n43797 = n10017 & ~n43796 ;
  assign n43800 = n43799 ^ n43797 ^ n11215 ;
  assign n43801 = n12213 | n38622 ;
  assign n43802 = n5689 & ~n43801 ;
  assign n43803 = n43800 & n43802 ;
  assign n43804 = ( n38847 & n43795 ) | ( n38847 & n43803 ) | ( n43795 & n43803 ) ;
  assign n43805 = n38676 ^ n16990 ^ 1'b0 ;
  assign n43806 = n19538 & n26708 ;
  assign n43807 = n18073 & n43806 ;
  assign n43808 = n7489 & n10131 ;
  assign n43809 = n43808 ^ n23455 ^ x245 ;
  assign n43810 = n10740 & n15959 ;
  assign n43811 = n8436 & n37505 ;
  assign n43812 = n43811 ^ n5135 ^ 1'b0 ;
  assign n43813 = n43812 ^ n40380 ^ 1'b0 ;
  assign n43814 = n24224 ^ n14916 ^ n13055 ;
  assign n43815 = ( n3359 & ~n17682 ) | ( n3359 & n43814 ) | ( ~n17682 & n43814 ) ;
  assign n43816 = n4215 & n17442 ;
  assign n43817 = n43816 ^ n21579 ^ 1'b0 ;
  assign n43818 = n32472 ^ n15372 ^ n14018 ;
  assign n43819 = ~n15983 & n43818 ;
  assign n43820 = ~n25709 & n43819 ;
  assign n43821 = n12622 & ~n20766 ;
  assign n43822 = n15742 & n43821 ;
  assign n43823 = ( n3444 & n4264 ) | ( n3444 & n19461 ) | ( n4264 & n19461 ) ;
  assign n43824 = n43823 ^ n673 ^ 1'b0 ;
  assign n43825 = n23940 ^ n10160 ^ n2897 ;
  assign n43826 = ( n15998 & n25525 ) | ( n15998 & n43825 ) | ( n25525 & n43825 ) ;
  assign n43827 = n38972 ^ n11001 ^ 1'b0 ;
  assign n43828 = n43826 & n43827 ;
  assign n43829 = n18687 | n24547 ;
  assign n43830 = n43829 ^ n35426 ^ n21505 ;
  assign n43831 = ( n7216 & ~n43828 ) | ( n7216 & n43830 ) | ( ~n43828 & n43830 ) ;
  assign n43832 = n17181 & n28171 ;
  assign n43833 = ( n8620 & ~n42473 ) | ( n8620 & n43832 ) | ( ~n42473 & n43832 ) ;
  assign n43834 = n43833 ^ n12234 ^ 1'b0 ;
  assign n43835 = n9421 | n24495 ;
  assign n43836 = ( n6693 & n15986 ) | ( n6693 & ~n17726 ) | ( n15986 & ~n17726 ) ;
  assign n43837 = ~n7390 & n43836 ;
  assign n43838 = n7558 & n43837 ;
  assign n43839 = n35803 ^ n7936 ^ 1'b0 ;
  assign n43840 = n9292 | n16584 ;
  assign n43841 = n43840 ^ n8176 ^ 1'b0 ;
  assign n43842 = n43841 ^ n12168 ^ n4482 ;
  assign n43843 = n5581 & n15254 ;
  assign n43844 = n43843 ^ n25235 ^ 1'b0 ;
  assign n43845 = n14697 & ~n21976 ;
  assign n43846 = n10174 | n14522 ;
  assign n43847 = n13283 & ~n43846 ;
  assign n43848 = ( n43844 & n43845 ) | ( n43844 & ~n43847 ) | ( n43845 & ~n43847 ) ;
  assign n43849 = n7240 & n13740 ;
  assign n43850 = n33137 & ~n36422 ;
  assign n43851 = ( n4429 & n10517 ) | ( n4429 & ~n26937 ) | ( n10517 & ~n26937 ) ;
  assign n43852 = ( n10924 & n15864 ) | ( n10924 & n24655 ) | ( n15864 & n24655 ) ;
  assign n43853 = n2241 & n34686 ;
  assign n43854 = n43853 ^ n24165 ^ 1'b0 ;
  assign n43855 = n43852 | n43854 ;
  assign n43856 = n30125 ^ n6691 ^ 1'b0 ;
  assign n43857 = n15091 & n43856 ;
  assign n43858 = n37902 ^ n2027 ^ 1'b0 ;
  assign n43859 = ( n2554 & n20018 ) | ( n2554 & n43858 ) | ( n20018 & n43858 ) ;
  assign n43861 = n15590 ^ n2593 ^ n820 ;
  assign n43862 = ( n1473 & n5402 ) | ( n1473 & n43861 ) | ( n5402 & n43861 ) ;
  assign n43860 = ~n10738 & n18370 ;
  assign n43863 = n43862 ^ n43860 ^ 1'b0 ;
  assign n43864 = ( n6458 & ~n16925 ) | ( n6458 & n43863 ) | ( ~n16925 & n43863 ) ;
  assign n43865 = n3702 & ~n38250 ;
  assign n43866 = n23790 | n43865 ;
  assign n43867 = n13981 & ~n43866 ;
  assign n43868 = n1873 & ~n34694 ;
  assign n43869 = n34065 ^ n28756 ^ n26058 ;
  assign n43870 = n38873 ^ n38541 ^ 1'b0 ;
  assign n43871 = n5371 & n43870 ;
  assign n43872 = n21937 & n43871 ;
  assign n43873 = n43872 ^ n31782 ^ 1'b0 ;
  assign n43874 = n30435 ^ n9675 ^ n1672 ;
  assign n43875 = n17520 ^ n4737 ^ 1'b0 ;
  assign n43876 = ~n43874 & n43875 ;
  assign n43877 = n19980 ^ n11181 ^ 1'b0 ;
  assign n43878 = ~n9522 & n43877 ;
  assign n43879 = n11507 & n43878 ;
  assign n43880 = ( n352 & n4363 ) | ( n352 & n17820 ) | ( n4363 & n17820 ) ;
  assign n43881 = n12660 ^ n6061 ^ 1'b0 ;
  assign n43882 = n16128 & n43881 ;
  assign n43883 = n43882 ^ n37175 ^ n403 ;
  assign n43884 = n43883 ^ n13044 ^ 1'b0 ;
  assign n43885 = n21927 ^ n19234 ^ n1107 ;
  assign n43886 = n29748 ^ n15558 ^ n6665 ;
  assign n43887 = ( n9812 & n20977 ) | ( n9812 & n25765 ) | ( n20977 & n25765 ) ;
  assign n43888 = n43887 ^ n42190 ^ n2819 ;
  assign n43889 = n24599 ^ n3561 ^ 1'b0 ;
  assign n43890 = n37659 | n43889 ;
  assign n43891 = n2914 | n36850 ;
  assign n43892 = ( n18663 & ~n19972 ) | ( n18663 & n43891 ) | ( ~n19972 & n43891 ) ;
  assign n43893 = n7380 & n16148 ;
  assign n43894 = ~n23834 & n43893 ;
  assign n43895 = ~n43892 & n43894 ;
  assign n43896 = ( n6541 & n8744 ) | ( n6541 & ~n18994 ) | ( n8744 & ~n18994 ) ;
  assign n43897 = ( n552 & ~n23144 ) | ( n552 & n43896 ) | ( ~n23144 & n43896 ) ;
  assign n43898 = n21681 & n43897 ;
  assign n43899 = n3515 ^ n2497 ^ 1'b0 ;
  assign n43900 = n29409 | n43899 ;
  assign n43901 = n32893 ^ n12293 ^ 1'b0 ;
  assign n43903 = n11885 ^ n10037 ^ 1'b0 ;
  assign n43902 = n19656 ^ n7783 ^ n284 ;
  assign n43904 = n43903 ^ n43902 ^ n35497 ;
  assign n43905 = n2997 & ~n9469 ;
  assign n43906 = n36197 & n43905 ;
  assign n43907 = n43906 ^ n1560 ^ 1'b0 ;
  assign n43908 = n26385 ^ n13979 ^ n5779 ;
  assign n43909 = n7148 & n28250 ;
  assign n43912 = n28756 ^ n10440 ^ n8844 ;
  assign n43910 = n25399 & ~n31036 ;
  assign n43911 = ~n3640 & n43910 ;
  assign n43913 = n43912 ^ n43911 ^ 1'b0 ;
  assign n43914 = n20848 & ~n43031 ;
  assign n43915 = n18339 & ~n33158 ;
  assign n43916 = n9764 & ~n42392 ;
  assign n43917 = n2419 & ~n17668 ;
  assign n43918 = n43917 ^ n11144 ^ 1'b0 ;
  assign n43919 = n43918 ^ n28771 ^ n18226 ;
  assign n43920 = ( n35520 & n43916 ) | ( n35520 & ~n43919 ) | ( n43916 & ~n43919 ) ;
  assign n43921 = ( n952 & n2698 ) | ( n952 & n26608 ) | ( n2698 & n26608 ) ;
  assign n43922 = n43921 ^ n22555 ^ n16179 ;
  assign n43923 = n43922 ^ n43438 ^ n10986 ;
  assign n43924 = ~n10340 & n33967 ;
  assign n43925 = ( ~n5958 & n8136 ) | ( ~n5958 & n8513 ) | ( n8136 & n8513 ) ;
  assign n43926 = n31361 & n43925 ;
  assign n43927 = n17600 | n43926 ;
  assign n43928 = n8316 & n14256 ;
  assign n43929 = ~n38478 & n43928 ;
  assign n43930 = ( n3699 & ~n8655 ) | ( n3699 & n39548 ) | ( ~n8655 & n39548 ) ;
  assign n43931 = n41273 & n43930 ;
  assign n43932 = n13719 ^ n12177 ^ n6967 ;
  assign n43933 = n35931 ^ n11087 ^ 1'b0 ;
  assign n43934 = n30815 ^ n19201 ^ n9760 ;
  assign n43935 = ( ~n4055 & n8550 ) | ( ~n4055 & n12904 ) | ( n8550 & n12904 ) ;
  assign n43936 = n21623 ^ n18008 ^ x211 ;
  assign n43937 = n43936 ^ n9981 ^ 1'b0 ;
  assign n43938 = n9799 & n43937 ;
  assign n43939 = n43938 ^ n21035 ^ 1'b0 ;
  assign n43940 = n43897 ^ n5110 ^ 1'b0 ;
  assign n43941 = n22870 & n43940 ;
  assign n43942 = x29 & n8984 ;
  assign n43943 = n43942 ^ n21122 ^ 1'b0 ;
  assign n43944 = n11878 | n15920 ;
  assign n43945 = ( n3050 & ~n12734 ) | ( n3050 & n23857 ) | ( ~n12734 & n23857 ) ;
  assign n43946 = n43945 ^ n13323 ^ 1'b0 ;
  assign n43947 = n43946 ^ n27651 ^ n11490 ;
  assign n43948 = ( n1106 & n28104 ) | ( n1106 & ~n35496 ) | ( n28104 & ~n35496 ) ;
  assign n43949 = n43948 ^ n40460 ^ 1'b0 ;
  assign n43950 = n14483 ^ n8253 ^ 1'b0 ;
  assign n43951 = n9590 & ~n43950 ;
  assign n43952 = ~n7276 & n30474 ;
  assign n43953 = n43952 ^ n22583 ^ n14532 ;
  assign n43954 = ( n6254 & n18519 ) | ( n6254 & n25810 ) | ( n18519 & n25810 ) ;
  assign n43955 = n37571 ^ x149 ^ 1'b0 ;
  assign n43956 = n25709 & ~n43955 ;
  assign n43957 = ( n21582 & ~n29618 ) | ( n21582 & n43956 ) | ( ~n29618 & n43956 ) ;
  assign n43958 = ~x224 & n43957 ;
  assign n43959 = ( n5253 & n8711 ) | ( n5253 & n10641 ) | ( n8711 & n10641 ) ;
  assign n43960 = ~n13330 & n20079 ;
  assign n43961 = ~n43959 & n43960 ;
  assign n43962 = n30173 ^ n24121 ^ n20299 ;
  assign n43963 = n9532 ^ n8510 ^ 1'b0 ;
  assign n43964 = ~n14323 & n43963 ;
  assign n43965 = n43964 ^ n37406 ^ n10275 ;
  assign n43966 = n43965 ^ n11502 ^ 1'b0 ;
  assign n43967 = n17566 | n43966 ;
  assign n43968 = n7104 & ~n27611 ;
  assign n43969 = ~n15762 & n43968 ;
  assign n43970 = ( n26562 & ~n43967 ) | ( n26562 & n43969 ) | ( ~n43967 & n43969 ) ;
  assign n43971 = n6333 | n43970 ;
  assign n43972 = n12852 ^ n10324 ^ n4080 ;
  assign n43973 = n43972 ^ n29906 ^ n10202 ;
  assign n43974 = n27128 ^ n8239 ^ n5309 ;
  assign n43975 = ( n32616 & n38557 ) | ( n32616 & ~n43974 ) | ( n38557 & ~n43974 ) ;
  assign n43979 = ~n5261 & n34265 ;
  assign n43976 = n36844 ^ n10007 ^ 1'b0 ;
  assign n43977 = n7830 | n43976 ;
  assign n43978 = n43977 ^ n42127 ^ n3541 ;
  assign n43980 = n43979 ^ n43978 ^ n26173 ;
  assign n43981 = ~n16315 & n16931 ;
  assign n43982 = ~n22256 & n43981 ;
  assign n43983 = x129 | n8881 ;
  assign n43984 = n13500 & ~n43983 ;
  assign n43985 = ~n26270 & n43984 ;
  assign n43986 = n491 | n40433 ;
  assign n43987 = n17556 & n32148 ;
  assign n43988 = n1769 & n43987 ;
  assign n43989 = n43315 ^ n41667 ^ n28129 ;
  assign n43990 = n42231 ^ n6901 ^ 1'b0 ;
  assign n43991 = n16851 | n21127 ;
  assign n43992 = n43991 ^ n3493 ^ 1'b0 ;
  assign n43993 = ( n12677 & n43990 ) | ( n12677 & n43992 ) | ( n43990 & n43992 ) ;
  assign n43994 = n31490 ^ n21496 ^ 1'b0 ;
  assign n43995 = ~n5352 & n43994 ;
  assign n43997 = ( n8949 & n9246 ) | ( n8949 & ~n23263 ) | ( n9246 & ~n23263 ) ;
  assign n43996 = n2668 & n17096 ;
  assign n43998 = n43997 ^ n43996 ^ n12872 ;
  assign n43999 = n33532 ^ n32320 ^ 1'b0 ;
  assign n44000 = n29166 & n43999 ;
  assign n44001 = n15345 & ~n22467 ;
  assign n44002 = n7974 | n28523 ;
  assign n44003 = n41353 & ~n44002 ;
  assign n44004 = ~n14174 & n35958 ;
  assign n44005 = n6307 | n44004 ;
  assign n44006 = n26939 | n44005 ;
  assign n44007 = n21774 ^ n7783 ^ 1'b0 ;
  assign n44008 = n41054 & n44007 ;
  assign n44009 = ~n4916 & n44008 ;
  assign n44010 = n44009 ^ n8647 ^ 1'b0 ;
  assign n44011 = n33808 & n44010 ;
  assign n44012 = ( n11845 & ~n16964 ) | ( n11845 & n40058 ) | ( ~n16964 & n40058 ) ;
  assign n44013 = ( n18703 & n29939 ) | ( n18703 & n44012 ) | ( n29939 & n44012 ) ;
  assign n44014 = n29589 ^ n6959 ^ 1'b0 ;
  assign n44015 = n44014 ^ n38583 ^ n11043 ;
  assign n44016 = ( n25477 & n28230 ) | ( n25477 & n37168 ) | ( n28230 & n37168 ) ;
  assign n44017 = n6138 & ~n8605 ;
  assign n44018 = ( n8330 & n18797 ) | ( n8330 & n20326 ) | ( n18797 & n20326 ) ;
  assign n44019 = n44018 ^ n43730 ^ n7886 ;
  assign n44020 = n14232 ^ n419 ^ 1'b0 ;
  assign n44021 = n44019 | n44020 ;
  assign n44022 = n983 & n5950 ;
  assign n44023 = n32130 ^ n1635 ^ 1'b0 ;
  assign n44024 = n44022 | n44023 ;
  assign n44026 = n7406 | n31969 ;
  assign n44027 = n44026 ^ n2849 ^ 1'b0 ;
  assign n44028 = ( n2421 & ~n29447 ) | ( n2421 & n44027 ) | ( ~n29447 & n44027 ) ;
  assign n44025 = ( n10113 & ~n12051 ) | ( n10113 & n14641 ) | ( ~n12051 & n14641 ) ;
  assign n44029 = n44028 ^ n44025 ^ n32024 ;
  assign n44030 = n14667 ^ n11853 ^ 1'b0 ;
  assign n44031 = ( n22989 & n33327 ) | ( n22989 & ~n44030 ) | ( n33327 & ~n44030 ) ;
  assign n44032 = ( ~n9863 & n26695 ) | ( ~n9863 & n44031 ) | ( n26695 & n44031 ) ;
  assign n44034 = n12353 & n16266 ;
  assign n44033 = n36211 ^ n18588 ^ n6782 ;
  assign n44035 = n44034 ^ n44033 ^ 1'b0 ;
  assign n44036 = n44035 ^ n41253 ^ 1'b0 ;
  assign n44037 = n9108 ^ n8994 ^ 1'b0 ;
  assign n44038 = n18331 & n44037 ;
  assign n44039 = ( n320 & n5762 ) | ( n320 & ~n44038 ) | ( n5762 & ~n44038 ) ;
  assign n44040 = ( n25955 & n33292 ) | ( n25955 & n33705 ) | ( n33292 & n33705 ) ;
  assign n44043 = n1505 | n6671 ;
  assign n44044 = n44043 ^ n5573 ^ 1'b0 ;
  assign n44042 = n8234 | n11026 ;
  assign n44045 = n44044 ^ n44042 ^ 1'b0 ;
  assign n44041 = n30876 ^ n22193 ^ n10159 ;
  assign n44046 = n44045 ^ n44041 ^ 1'b0 ;
  assign n44047 = n33618 & ~n44046 ;
  assign n44048 = n18614 ^ n16383 ^ n5140 ;
  assign n44049 = ( ~n4863 & n7833 ) | ( ~n4863 & n9042 ) | ( n7833 & n9042 ) ;
  assign n44050 = x73 & ~n9401 ;
  assign n44051 = ~n1186 & n44050 ;
  assign n44052 = ~n44049 & n44051 ;
  assign n44053 = n44048 & ~n44052 ;
  assign n44054 = n7859 & n44053 ;
  assign n44055 = n32757 ^ n24021 ^ 1'b0 ;
  assign n44056 = x139 & ~n44055 ;
  assign n44058 = n1600 | n21488 ;
  assign n44057 = n10271 ^ n497 ^ 1'b0 ;
  assign n44059 = n44058 ^ n44057 ^ n20329 ;
  assign n44060 = n2834 & n23135 ;
  assign n44061 = n44059 & n44060 ;
  assign n44062 = n13753 ^ n6514 ^ n4285 ;
  assign n44063 = ~n15049 & n35919 ;
  assign n44064 = n20361 & n44063 ;
  assign n44065 = n44062 & ~n44064 ;
  assign n44066 = n18002 & n37832 ;
  assign n44067 = n44066 ^ n10480 ^ n10105 ;
  assign n44068 = n13621 ^ n12265 ^ 1'b0 ;
  assign n44069 = ~n38254 & n44068 ;
  assign n44070 = ( x86 & ~n7710 ) | ( x86 & n44069 ) | ( ~n7710 & n44069 ) ;
  assign n44071 = n22752 ^ n16803 ^ n327 ;
  assign n44072 = n44071 ^ n27110 ^ 1'b0 ;
  assign n44073 = n17175 | n44072 ;
  assign n44074 = n44073 ^ n10259 ^ x237 ;
  assign n44075 = ( n11339 & ~n14272 ) | ( n11339 & n44074 ) | ( ~n14272 & n44074 ) ;
  assign n44076 = n836 & n40613 ;
  assign n44077 = n18305 & n22223 ;
  assign n44078 = n44077 ^ n22162 ^ 1'b0 ;
  assign n44079 = ~n44076 & n44078 ;
  assign n44080 = n25237 ^ n3933 ^ n2890 ;
  assign n44081 = n33443 | n44080 ;
  assign n44082 = n44081 ^ n9670 ^ 1'b0 ;
  assign n44083 = n21675 | n28618 ;
  assign n44084 = n25771 & n37716 ;
  assign n44085 = ~n23184 & n44084 ;
  assign n44086 = n44085 ^ n24628 ^ 1'b0 ;
  assign n44087 = n42506 ^ n20855 ^ n13563 ;
  assign n44088 = n9414 ^ n8494 ^ 1'b0 ;
  assign n44089 = n8020 | n44088 ;
  assign n44090 = n35813 & n44089 ;
  assign n44091 = ( n9907 & n15337 ) | ( n9907 & ~n44090 ) | ( n15337 & ~n44090 ) ;
  assign n44092 = n11513 & n13406 ;
  assign n44093 = ( n782 & ~n15587 ) | ( n782 & n40128 ) | ( ~n15587 & n40128 ) ;
  assign n44094 = ( n41612 & n44092 ) | ( n41612 & n44093 ) | ( n44092 & n44093 ) ;
  assign n44095 = x167 & ~n25070 ;
  assign n44096 = n44095 ^ n29376 ^ 1'b0 ;
  assign n44097 = n17586 ^ n16989 ^ n431 ;
  assign n44098 = n44097 ^ n42577 ^ 1'b0 ;
  assign n44099 = n34849 ^ n14620 ^ n9132 ;
  assign n44100 = ( n8103 & ~n44098 ) | ( n8103 & n44099 ) | ( ~n44098 & n44099 ) ;
  assign n44101 = ~n13352 & n44100 ;
  assign n44102 = ( ~n969 & n16221 ) | ( ~n969 & n38105 ) | ( n16221 & n38105 ) ;
  assign n44103 = n25188 & ~n44102 ;
  assign n44106 = ~n15403 & n16117 ;
  assign n44107 = n44106 ^ n8463 ^ 1'b0 ;
  assign n44104 = n8148 | n32371 ;
  assign n44105 = n6282 & ~n44104 ;
  assign n44108 = n44107 ^ n44105 ^ 1'b0 ;
  assign n44109 = n1360 & n2812 ;
  assign n44110 = n44109 ^ n594 ^ 1'b0 ;
  assign n44111 = n44110 ^ n25538 ^ n5309 ;
  assign n44112 = ~n8205 & n32828 ;
  assign n44113 = n32339 ^ n1776 ^ 1'b0 ;
  assign n44119 = ~n5964 & n6511 ;
  assign n44120 = n44119 ^ x94 ^ 1'b0 ;
  assign n44121 = n19435 | n22042 ;
  assign n44122 = n44120 & ~n44121 ;
  assign n44117 = n12186 | n17013 ;
  assign n44118 = n44117 ^ n21454 ^ 1'b0 ;
  assign n44123 = n44122 ^ n44118 ^ n35614 ;
  assign n44114 = n27392 ^ n20359 ^ 1'b0 ;
  assign n44115 = ~n36868 & n44114 ;
  assign n44116 = n5822 & n44115 ;
  assign n44124 = n44123 ^ n44116 ^ 1'b0 ;
  assign n44125 = n10363 & ~n34283 ;
  assign n44126 = n44125 ^ n13653 ^ 1'b0 ;
  assign n44127 = ~n1569 & n29477 ;
  assign n44128 = n5524 | n12125 ;
  assign n44129 = n43338 & ~n44128 ;
  assign n44130 = n38951 ^ n18310 ^ n9078 ;
  assign n44131 = n44130 ^ n3472 ^ 1'b0 ;
  assign n44132 = ( n14284 & ~n16470 ) | ( n14284 & n20316 ) | ( ~n16470 & n20316 ) ;
  assign n44133 = n10722 ^ n1292 ^ 1'b0 ;
  assign n44134 = n43126 & ~n44133 ;
  assign n44135 = ( ~n1646 & n3169 ) | ( ~n1646 & n44134 ) | ( n3169 & n44134 ) ;
  assign n44136 = n5306 & ~n5397 ;
  assign n44137 = n44136 ^ n4250 ^ 1'b0 ;
  assign n44138 = n915 & ~n15838 ;
  assign n44139 = n44137 & n44138 ;
  assign n44140 = ( n16675 & ~n16703 ) | ( n16675 & n44139 ) | ( ~n16703 & n44139 ) ;
  assign n44141 = ~n570 & n16765 ;
  assign n44142 = n44141 ^ n14190 ^ 1'b0 ;
  assign n44143 = ( ~n29134 & n31622 ) | ( ~n29134 & n41632 ) | ( n31622 & n41632 ) ;
  assign n44144 = n44143 ^ n16086 ^ 1'b0 ;
  assign n44145 = n8336 & n41242 ;
  assign n44146 = n44145 ^ n36073 ^ 1'b0 ;
  assign n44147 = n23973 ^ n7143 ^ 1'b0 ;
  assign n44148 = ~n21569 & n44147 ;
  assign n44149 = ~n36793 & n44148 ;
  assign n44150 = ( ~n26832 & n31512 ) | ( ~n26832 & n33456 ) | ( n31512 & n33456 ) ;
  assign n44151 = n6240 ^ n4314 ^ 1'b0 ;
  assign n44152 = n44151 ^ n14161 ^ n6820 ;
  assign n44153 = ( ~n15413 & n35990 ) | ( ~n15413 & n44152 ) | ( n35990 & n44152 ) ;
  assign n44154 = n44153 ^ n24823 ^ n19357 ;
  assign n44156 = ~n10387 & n37730 ;
  assign n44155 = ~n2217 & n15959 ;
  assign n44157 = n44156 ^ n44155 ^ 1'b0 ;
  assign n44158 = n31728 & ~n43488 ;
  assign n44159 = n5639 & n21248 ;
  assign n44160 = ~n41963 & n44159 ;
  assign n44161 = ~n2757 & n16084 ;
  assign n44162 = n12193 & n44161 ;
  assign n44163 = n44162 ^ n6744 ^ 1'b0 ;
  assign n44164 = n1638 & ~n40247 ;
  assign n44165 = ( n394 & ~n22315 ) | ( n394 & n28787 ) | ( ~n22315 & n28787 ) ;
  assign n44166 = n1823 & n15564 ;
  assign n44167 = ~n12627 & n44166 ;
  assign n44168 = n44167 ^ n31745 ^ 1'b0 ;
  assign n44169 = n32143 & n44168 ;
  assign n44170 = ( n40064 & ~n44165 ) | ( n40064 & n44169 ) | ( ~n44165 & n44169 ) ;
  assign n44171 = ( n14370 & n17522 ) | ( n14370 & n36817 ) | ( n17522 & n36817 ) ;
  assign n44172 = n7817 ^ n7187 ^ n2128 ;
  assign n44173 = ~n16214 & n44172 ;
  assign n44174 = ~n14873 & n44173 ;
  assign n44175 = n35081 | n39535 ;
  assign n44176 = n16146 & ~n44175 ;
  assign n44177 = n12874 ^ n7353 ^ 1'b0 ;
  assign n44178 = n31960 ^ n20403 ^ 1'b0 ;
  assign n44179 = ( n21102 & n36338 ) | ( n21102 & n36534 ) | ( n36338 & n36534 ) ;
  assign n44180 = ( ~n30037 & n39199 ) | ( ~n30037 & n44179 ) | ( n39199 & n44179 ) ;
  assign n44181 = n44180 ^ n20615 ^ n11741 ;
  assign n44182 = ( ~n956 & n24603 ) | ( ~n956 & n44181 ) | ( n24603 & n44181 ) ;
  assign n44183 = n3205 ^ n3022 ^ 1'b0 ;
  assign n44184 = n10216 | n44183 ;
  assign n44185 = n14944 & ~n44184 ;
  assign n44186 = ~n27533 & n44185 ;
  assign n44187 = n44186 ^ n22766 ^ 1'b0 ;
  assign n44188 = n15521 & n44187 ;
  assign n44189 = ( n19853 & ~n24966 ) | ( n19853 & n44188 ) | ( ~n24966 & n44188 ) ;
  assign n44190 = n44189 ^ n1632 ^ 1'b0 ;
  assign n44191 = n5551 ^ n1173 ^ 1'b0 ;
  assign n44192 = n2184 & n44191 ;
  assign n44193 = n2630 ^ n1261 ^ 1'b0 ;
  assign n44194 = ( n13598 & n16518 ) | ( n13598 & ~n18361 ) | ( n16518 & ~n18361 ) ;
  assign n44195 = n44194 ^ n37195 ^ 1'b0 ;
  assign n44196 = n24069 ^ n6373 ^ 1'b0 ;
  assign n44197 = ~n22478 & n44196 ;
  assign n44198 = n8838 & n30403 ;
  assign n44199 = n44198 ^ n7619 ^ 1'b0 ;
  assign n44200 = n21636 | n26830 ;
  assign n44201 = n44199 | n44200 ;
  assign n44202 = n30868 ^ n16033 ^ n8905 ;
  assign n44203 = ( n14341 & n19688 ) | ( n14341 & ~n42572 ) | ( n19688 & ~n42572 ) ;
  assign n44204 = ( n14306 & n26692 ) | ( n14306 & ~n37195 ) | ( n26692 & ~n37195 ) ;
  assign n44205 = n44204 ^ n19018 ^ n3587 ;
  assign n44206 = n13918 & n29031 ;
  assign n44207 = n13752 & ~n21777 ;
  assign n44208 = ~n31109 & n44207 ;
  assign n44209 = ( n10461 & ~n12023 ) | ( n10461 & n40385 ) | ( ~n12023 & n40385 ) ;
  assign n44210 = ~n1720 & n30941 ;
  assign n44211 = n44209 & n44210 ;
  assign n44212 = n19981 ^ n11572 ^ 1'b0 ;
  assign n44213 = n13508 ^ n4553 ^ 1'b0 ;
  assign n44214 = n44212 | n44213 ;
  assign n44215 = n44214 ^ n23526 ^ 1'b0 ;
  assign n44216 = ( n9049 & n17243 ) | ( n9049 & ~n27382 ) | ( n17243 & ~n27382 ) ;
  assign n44217 = n20728 ^ n15645 ^ n8754 ;
  assign n44218 = ( ~n23671 & n44216 ) | ( ~n23671 & n44217 ) | ( n44216 & n44217 ) ;
  assign n44219 = n29358 ^ n20862 ^ n4160 ;
  assign n44220 = ( n20487 & n40740 ) | ( n20487 & n44219 ) | ( n40740 & n44219 ) ;
  assign n44222 = ( n514 & ~n10206 ) | ( n514 & n13148 ) | ( ~n10206 & n13148 ) ;
  assign n44221 = n8646 & ~n10492 ;
  assign n44223 = n44222 ^ n44221 ^ n18797 ;
  assign n44224 = n26406 | n33283 ;
  assign n44225 = ~n1180 & n21011 ;
  assign n44226 = n32199 & n44225 ;
  assign n44227 = n31261 ^ n15390 ^ 1'b0 ;
  assign n44229 = n16983 | n19693 ;
  assign n44230 = n44229 ^ n2823 ^ 1'b0 ;
  assign n44228 = n13045 ^ n8235 ^ 1'b0 ;
  assign n44231 = n44230 ^ n44228 ^ n40037 ;
  assign n44232 = ~n11515 & n19368 ;
  assign n44233 = n44231 & n44232 ;
  assign n44234 = n39036 ^ n10577 ^ n5585 ;
  assign n44235 = n10012 | n16964 ;
  assign n44236 = n16964 & ~n44235 ;
  assign n44237 = ( n11071 & n21490 ) | ( n11071 & ~n44236 ) | ( n21490 & ~n44236 ) ;
  assign n44238 = n41717 ^ n9469 ^ n9182 ;
  assign n44239 = n32106 ^ n1179 ^ 1'b0 ;
  assign n44240 = n3742 & n12394 ;
  assign n44241 = n44240 ^ n11213 ^ 1'b0 ;
  assign n44242 = ( n5968 & n28975 ) | ( n5968 & n44241 ) | ( n28975 & n44241 ) ;
  assign n44243 = n31883 & n44242 ;
  assign n44244 = n20757 ^ n5974 ^ 1'b0 ;
  assign n44245 = n38192 | n44244 ;
  assign n44246 = n40449 | n44245 ;
  assign n44247 = ( ~n13001 & n15088 ) | ( ~n13001 & n18522 ) | ( n15088 & n18522 ) ;
  assign n44248 = ~n12274 & n44247 ;
  assign n44249 = n44248 ^ n39828 ^ 1'b0 ;
  assign n44251 = n21049 ^ n18389 ^ 1'b0 ;
  assign n44250 = n5048 & ~n12912 ;
  assign n44252 = n44251 ^ n44250 ^ 1'b0 ;
  assign n44253 = n20831 ^ n18744 ^ 1'b0 ;
  assign n44254 = n11677 ^ n10791 ^ n7698 ;
  assign n44255 = ( n12231 & n14579 ) | ( n12231 & n21908 ) | ( n14579 & n21908 ) ;
  assign n44256 = ( n24342 & n44254 ) | ( n24342 & n44255 ) | ( n44254 & n44255 ) ;
  assign n44257 = ( n10961 & n14739 ) | ( n10961 & n38213 ) | ( n14739 & n38213 ) ;
  assign n44258 = n22919 ^ n20705 ^ 1'b0 ;
  assign n44259 = ( n19381 & n23920 ) | ( n19381 & n32057 ) | ( n23920 & n32057 ) ;
  assign n44260 = n5307 & ~n44259 ;
  assign n44261 = n8210 ^ n3208 ^ 1'b0 ;
  assign n44262 = n25252 ^ n2952 ^ 1'b0 ;
  assign n44263 = n17606 & n44262 ;
  assign n44264 = n14652 & n33421 ;
  assign n44265 = ~n44263 & n44264 ;
  assign n44266 = n5720 & ~n30382 ;
  assign n44267 = n18360 & n44266 ;
  assign n44268 = n12213 & ~n42772 ;
  assign n44269 = ~n3787 & n44268 ;
  assign n44270 = n9740 ^ n2566 ^ 1'b0 ;
  assign n44271 = ~n10819 & n22120 ;
  assign n44272 = n44270 & n44271 ;
  assign n44273 = n29205 & n36183 ;
  assign n44275 = n10065 ^ n8555 ^ n3012 ;
  assign n44274 = n28640 & ~n43591 ;
  assign n44276 = n44275 ^ n44274 ^ 1'b0 ;
  assign n44277 = ( n44272 & n44273 ) | ( n44272 & n44276 ) | ( n44273 & n44276 ) ;
  assign n44278 = n38977 ^ n22705 ^ n14769 ;
  assign n44279 = ( n2960 & ~n21807 ) | ( n2960 & n44278 ) | ( ~n21807 & n44278 ) ;
  assign n44280 = ( n9200 & ~n17800 ) | ( n9200 & n37441 ) | ( ~n17800 & n37441 ) ;
  assign n44284 = n20196 ^ n1789 ^ n1406 ;
  assign n44281 = n37373 ^ n33152 ^ 1'b0 ;
  assign n44282 = n26968 & n44281 ;
  assign n44283 = ( n14499 & n33643 ) | ( n14499 & ~n44282 ) | ( n33643 & ~n44282 ) ;
  assign n44285 = n44284 ^ n44283 ^ n2094 ;
  assign n44286 = n18397 | n26422 ;
  assign n44287 = n44286 ^ n441 ^ 1'b0 ;
  assign n44288 = n19213 ^ n5599 ^ 1'b0 ;
  assign n44289 = n16618 & n44288 ;
  assign n44290 = n10732 ^ n2821 ^ 1'b0 ;
  assign n44291 = n838 & ~n44290 ;
  assign n44292 = ~n17626 & n44291 ;
  assign n44293 = n17958 & n44292 ;
  assign n44294 = ( n8295 & ~n23397 ) | ( n8295 & n44293 ) | ( ~n23397 & n44293 ) ;
  assign n44295 = n23067 & ~n44294 ;
  assign n44296 = n27971 ^ n9510 ^ 1'b0 ;
  assign n44297 = n41139 ^ n16804 ^ n2750 ;
  assign n44298 = n44297 ^ n27097 ^ n24895 ;
  assign n44299 = n12120 & n23658 ;
  assign n44300 = n2488 & n44299 ;
  assign n44301 = ( n4077 & n32371 ) | ( n4077 & ~n44300 ) | ( n32371 & ~n44300 ) ;
  assign n44302 = n31263 ^ n773 ^ 1'b0 ;
  assign n44303 = n10415 | n44302 ;
  assign n44304 = ( ~n7526 & n15949 ) | ( ~n7526 & n21190 ) | ( n15949 & n21190 ) ;
  assign n44305 = n19113 & n32187 ;
  assign n44306 = ( n40393 & n44304 ) | ( n40393 & ~n44305 ) | ( n44304 & ~n44305 ) ;
  assign n44307 = n5225 | n8976 ;
  assign n44308 = n44307 ^ n39904 ^ 1'b0 ;
  assign n44309 = n44308 ^ n9199 ^ 1'b0 ;
  assign n44310 = ( n4510 & n32324 ) | ( n4510 & n44309 ) | ( n32324 & n44309 ) ;
  assign n44311 = ~n5954 & n17270 ;
  assign n44312 = n24595 ^ n10639 ^ n6679 ;
  assign n44313 = ( n27236 & n44311 ) | ( n27236 & ~n44312 ) | ( n44311 & ~n44312 ) ;
  assign n44314 = n9854 & n22561 ;
  assign n44315 = n16486 | n19757 ;
  assign n44316 = n44315 ^ n13873 ^ 1'b0 ;
  assign n44317 = n21547 | n44316 ;
  assign n44318 = n17394 & ~n44317 ;
  assign n44319 = n33224 ^ n12341 ^ 1'b0 ;
  assign n44320 = n30910 ^ n30028 ^ n19298 ;
  assign n44327 = ~n19056 & n26728 ;
  assign n44322 = n10466 ^ n3301 ^ n866 ;
  assign n44323 = n625 & ~n44322 ;
  assign n44324 = n9798 ^ n3222 ^ 1'b0 ;
  assign n44325 = ~n44323 & n44324 ;
  assign n44326 = ~n23142 & n44325 ;
  assign n44321 = n17218 | n44169 ;
  assign n44328 = n44327 ^ n44326 ^ n44321 ;
  assign n44329 = ( n1045 & n11507 ) | ( n1045 & ~n22575 ) | ( n11507 & ~n22575 ) ;
  assign n44330 = n12124 & ~n13689 ;
  assign n44331 = n41006 ^ n22844 ^ 1'b0 ;
  assign n44332 = n43463 & n44331 ;
  assign n44333 = n14669 | n29849 ;
  assign n44334 = n44333 ^ n25050 ^ 1'b0 ;
  assign n44335 = ~n37775 & n41391 ;
  assign n44336 = n44334 & n44335 ;
  assign n44337 = n26470 ^ n24201 ^ n16774 ;
  assign n44338 = n21880 & ~n37010 ;
  assign n44339 = n36622 ^ n24600 ^ n4591 ;
  assign n44340 = n6989 ^ n4376 ^ 1'b0 ;
  assign n44341 = n44339 & ~n44340 ;
  assign n44342 = ( n723 & n6406 ) | ( n723 & ~n7227 ) | ( n6406 & ~n7227 ) ;
  assign n44343 = n24349 & ~n44342 ;
  assign n44344 = n44343 ^ n15859 ^ 1'b0 ;
  assign n44345 = ( ~n1333 & n40508 ) | ( ~n1333 & n41485 ) | ( n40508 & n41485 ) ;
  assign n44346 = ~n1247 & n5461 ;
  assign n44347 = n12668 & n20336 ;
  assign n44348 = ( ~n36041 & n44346 ) | ( ~n36041 & n44347 ) | ( n44346 & n44347 ) ;
  assign n44349 = n6130 & n12226 ;
  assign n44350 = n44349 ^ n5533 ^ 1'b0 ;
  assign n44351 = ( n11052 & ~n14235 ) | ( n11052 & n19522 ) | ( ~n14235 & n19522 ) ;
  assign n44352 = n44350 & n44351 ;
  assign n44360 = n10090 & n13496 ;
  assign n44361 = n44360 ^ n10811 ^ 1'b0 ;
  assign n44355 = n995 & n20836 ;
  assign n44356 = n14968 ^ n14878 ^ 1'b0 ;
  assign n44357 = n16681 & ~n44356 ;
  assign n44358 = ~n4036 & n44357 ;
  assign n44359 = n44355 & n44358 ;
  assign n44362 = n44361 ^ n44359 ^ n10430 ;
  assign n44353 = ( n4978 & ~n9312 ) | ( n4978 & n20718 ) | ( ~n9312 & n20718 ) ;
  assign n44354 = n44353 ^ n38510 ^ n14959 ;
  assign n44363 = n44362 ^ n44354 ^ n4146 ;
  assign n44364 = n19818 ^ n2766 ^ 1'b0 ;
  assign n44365 = n25910 & ~n44364 ;
  assign n44366 = n42948 ^ n6596 ^ n647 ;
  assign n44367 = ( ~n7167 & n7860 ) | ( ~n7167 & n44366 ) | ( n7860 & n44366 ) ;
  assign n44368 = ( n15967 & n19428 ) | ( n15967 & ~n44367 ) | ( n19428 & ~n44367 ) ;
  assign n44369 = n15989 & ~n44368 ;
  assign n44370 = n15109 & ~n27716 ;
  assign n44371 = n44370 ^ n25225 ^ 1'b0 ;
  assign n44372 = n16043 & n32834 ;
  assign n44373 = ~n24089 & n44372 ;
  assign n44374 = ~n1410 & n32782 ;
  assign n44375 = n6708 & n44374 ;
  assign n44376 = n31148 & n44375 ;
  assign n44377 = n22512 ^ n15556 ^ n10678 ;
  assign n44378 = n5583 & n39439 ;
  assign n44379 = n44378 ^ n32375 ^ n8020 ;
  assign n44380 = n33303 & ~n41558 ;
  assign n44381 = n33643 ^ n2247 ^ 1'b0 ;
  assign n44382 = n18861 & n44381 ;
  assign n44383 = n44382 ^ n11833 ^ 1'b0 ;
  assign n44384 = n5036 ^ x254 ^ 1'b0 ;
  assign n44385 = n16120 & ~n44384 ;
  assign n44386 = n26654 & n44385 ;
  assign n44387 = n44386 ^ n39153 ^ 1'b0 ;
  assign n44388 = n39853 & n44069 ;
  assign n44389 = n44388 ^ n23072 ^ 1'b0 ;
  assign n44390 = n44389 ^ n2388 ^ 1'b0 ;
  assign n44391 = ( n3068 & n7510 ) | ( n3068 & n27589 ) | ( n7510 & n27589 ) ;
  assign n44392 = ~n8357 & n41891 ;
  assign n44393 = ( n5441 & ~n23016 ) | ( n5441 & n42039 ) | ( ~n23016 & n42039 ) ;
  assign n44394 = n15266 ^ n10719 ^ 1'b0 ;
  assign n44395 = n5655 ^ n2730 ^ 1'b0 ;
  assign n44396 = n16538 ^ n9978 ^ 1'b0 ;
  assign n44397 = ~n44395 & n44396 ;
  assign n44398 = n22943 ^ n22890 ^ 1'b0 ;
  assign n44399 = n27655 | n41623 ;
  assign n44400 = n34785 ^ n27663 ^ 1'b0 ;
  assign n44401 = n4065 & ~n44400 ;
  assign n44402 = n22840 ^ n8323 ^ 1'b0 ;
  assign n44403 = ( ~n2822 & n25579 ) | ( ~n2822 & n44402 ) | ( n25579 & n44402 ) ;
  assign n44404 = n12620 & n18364 ;
  assign n44405 = n12420 ^ n2934 ^ 1'b0 ;
  assign n44406 = n4770 | n44405 ;
  assign n44407 = n14752 ^ n9654 ^ 1'b0 ;
  assign n44408 = ~n44406 & n44407 ;
  assign n44409 = n44408 ^ n31044 ^ 1'b0 ;
  assign n44410 = n36934 ^ n18045 ^ n10472 ;
  assign n44412 = n2955 & n10811 ;
  assign n44411 = ~n9169 & n20417 ;
  assign n44413 = n44412 ^ n44411 ^ 1'b0 ;
  assign n44415 = n9381 & n34129 ;
  assign n44416 = n11702 & n44415 ;
  assign n44414 = n13428 | n14614 ;
  assign n44417 = n44416 ^ n44414 ^ 1'b0 ;
  assign n44418 = n24833 ^ x163 ^ 1'b0 ;
  assign n44419 = n11727 | n44418 ;
  assign n44422 = n17216 & ~n18627 ;
  assign n44423 = n44422 ^ n35693 ^ 1'b0 ;
  assign n44421 = n28337 ^ n8078 ^ 1'b0 ;
  assign n44424 = n44423 ^ n44421 ^ n9269 ;
  assign n44420 = n39178 ^ n36574 ^ n15653 ;
  assign n44425 = n44424 ^ n44420 ^ n10817 ;
  assign n44426 = n7220 & n15610 ;
  assign n44427 = ~n23301 & n44426 ;
  assign n44428 = ( n12653 & ~n17226 ) | ( n12653 & n44427 ) | ( ~n17226 & n44427 ) ;
  assign n44429 = ( n12333 & n18070 ) | ( n12333 & n44428 ) | ( n18070 & n44428 ) ;
  assign n44430 = n44429 ^ n33123 ^ 1'b0 ;
  assign n44431 = ( ~n3126 & n4368 ) | ( ~n3126 & n36861 ) | ( n4368 & n36861 ) ;
  assign n44432 = ( ~n4977 & n22421 ) | ( ~n4977 & n34250 ) | ( n22421 & n34250 ) ;
  assign n44433 = n15686 ^ n10270 ^ n8122 ;
  assign n44434 = n24038 | n44433 ;
  assign n44435 = n44434 ^ n37954 ^ n3896 ;
  assign n44436 = n33091 | n44435 ;
  assign n44437 = n9762 | n44436 ;
  assign n44438 = n33648 ^ n10914 ^ 1'b0 ;
  assign n44439 = n17127 & n44438 ;
  assign n44440 = ~n19828 & n44439 ;
  assign n44441 = n13160 & n24232 ;
  assign n44442 = ~n6945 & n10464 ;
  assign n44443 = ~n6586 & n44442 ;
  assign n44444 = n21023 | n44443 ;
  assign n44445 = n44444 ^ n7283 ^ 1'b0 ;
  assign n44446 = ( n16136 & n44441 ) | ( n16136 & ~n44445 ) | ( n44441 & ~n44445 ) ;
  assign n44447 = ~n1423 & n16198 ;
  assign n44448 = n44447 ^ n29431 ^ 1'b0 ;
  assign n44449 = ~n9658 & n21383 ;
  assign n44450 = ( n36589 & n44448 ) | ( n36589 & n44449 ) | ( n44448 & n44449 ) ;
  assign n44451 = ( n8430 & n17529 ) | ( n8430 & n44450 ) | ( n17529 & n44450 ) ;
  assign n44454 = n18197 ^ n864 ^ 1'b0 ;
  assign n44455 = n10670 & n44454 ;
  assign n44456 = ~n36656 & n44455 ;
  assign n44453 = n17175 ^ n6555 ^ n3958 ;
  assign n44452 = ~n20867 & n26444 ;
  assign n44457 = n44456 ^ n44453 ^ n44452 ;
  assign n44458 = n31634 ^ n20619 ^ n7819 ;
  assign n44459 = ~n5433 & n10993 ;
  assign n44460 = n44459 ^ n8634 ^ 1'b0 ;
  assign n44461 = ( n28457 & ~n30371 ) | ( n28457 & n44460 ) | ( ~n30371 & n44460 ) ;
  assign n44462 = ~n26505 & n44461 ;
  assign n44463 = n43780 ^ n18745 ^ 1'b0 ;
  assign n44464 = n12311 & ~n44463 ;
  assign n44465 = n44273 ^ n21031 ^ 1'b0 ;
  assign n44469 = ( n7119 & n13483 ) | ( n7119 & ~n15745 ) | ( n13483 & ~n15745 ) ;
  assign n44470 = n44469 ^ n20567 ^ 1'b0 ;
  assign n44466 = ( n1255 & n7272 ) | ( n1255 & ~n9211 ) | ( n7272 & ~n9211 ) ;
  assign n44467 = n40593 | n44466 ;
  assign n44468 = n2726 & ~n44467 ;
  assign n44471 = n44470 ^ n44468 ^ 1'b0 ;
  assign n44472 = n2094 & ~n6254 ;
  assign n44473 = n44472 ^ n7027 ^ n5446 ;
  assign n44474 = ( ~n5618 & n18410 ) | ( ~n5618 & n38522 ) | ( n18410 & n38522 ) ;
  assign n44475 = ~n37713 & n44474 ;
  assign n44476 = n37300 ^ n4615 ^ 1'b0 ;
  assign n44477 = n38928 ^ n25881 ^ n4813 ;
  assign n44481 = ( ~n301 & n3040 ) | ( ~n301 & n17117 ) | ( n3040 & n17117 ) ;
  assign n44480 = ~n20063 & n24487 ;
  assign n44482 = n44481 ^ n44480 ^ 1'b0 ;
  assign n44478 = n16054 ^ n14793 ^ 1'b0 ;
  assign n44479 = ( ~n18070 & n21505 ) | ( ~n18070 & n44478 ) | ( n21505 & n44478 ) ;
  assign n44483 = n44482 ^ n44479 ^ n35019 ;
  assign n44484 = ( n5360 & ~n44477 ) | ( n5360 & n44483 ) | ( ~n44477 & n44483 ) ;
  assign n44485 = n14146 ^ n8937 ^ 1'b0 ;
  assign n44486 = n1145 & ~n44485 ;
  assign n44487 = n44486 ^ n11993 ^ 1'b0 ;
  assign n44488 = ~n4688 & n44487 ;
  assign n44489 = n7254 | n21164 ;
  assign n44490 = n44489 ^ n13673 ^ 1'b0 ;
  assign n44491 = n6216 | n30381 ;
  assign n44492 = x160 & n44491 ;
  assign n44493 = n8456 & n44492 ;
  assign n44494 = n36946 ^ n31285 ^ 1'b0 ;
  assign n44495 = n44494 ^ n17511 ^ 1'b0 ;
  assign n44496 = n16163 ^ n12604 ^ n1142 ;
  assign n44497 = n20433 ^ n16085 ^ n9887 ;
  assign n44498 = ~n5063 & n31524 ;
  assign n44499 = n44498 ^ n18730 ^ 1'b0 ;
  assign n44500 = ~n19018 & n44499 ;
  assign n44501 = n3138 & ~n4051 ;
  assign n44502 = ~n31437 & n44501 ;
  assign n44503 = ( n4097 & n18839 ) | ( n4097 & n26854 ) | ( n18839 & n26854 ) ;
  assign n44504 = n29758 & ~n44503 ;
  assign n44505 = ~n9705 & n44504 ;
  assign n44506 = n11765 ^ n946 ^ 1'b0 ;
  assign n44507 = n44506 ^ n1274 ^ 1'b0 ;
  assign n44508 = n44507 ^ n25774 ^ n10731 ;
  assign n44512 = ~n9612 & n33139 ;
  assign n44513 = n15233 & ~n44512 ;
  assign n44509 = n7408 & ~n43011 ;
  assign n44510 = n44509 ^ n6216 ^ 1'b0 ;
  assign n44511 = n44510 ^ n16873 ^ 1'b0 ;
  assign n44514 = n44513 ^ n44511 ^ n10851 ;
  assign n44515 = ( n15559 & n22445 ) | ( n15559 & ~n26775 ) | ( n22445 & ~n26775 ) ;
  assign n44516 = ~n2934 & n44515 ;
  assign n44517 = n21101 ^ n5240 ^ 1'b0 ;
  assign n44518 = ~n14148 & n44517 ;
  assign n44519 = ( n11855 & ~n22581 ) | ( n11855 & n44518 ) | ( ~n22581 & n44518 ) ;
  assign n44520 = n34435 | n36970 ;
  assign n44521 = n23179 ^ n4445 ^ n1497 ;
  assign n44522 = n44521 ^ n35342 ^ n12668 ;
  assign n44523 = n445 | n1624 ;
  assign n44524 = n44522 & ~n44523 ;
  assign n44525 = n42182 ^ n32672 ^ n12872 ;
  assign n44526 = n26731 & ~n34863 ;
  assign n44527 = ( n31336 & ~n37504 ) | ( n31336 & n43669 ) | ( ~n37504 & n43669 ) ;
  assign n44528 = ( n15998 & ~n28649 ) | ( n15998 & n44527 ) | ( ~n28649 & n44527 ) ;
  assign n44529 = n1074 | n5430 ;
  assign n44530 = n44529 ^ n7201 ^ 1'b0 ;
  assign n44531 = ( ~n8405 & n24103 ) | ( ~n8405 & n27074 ) | ( n24103 & n27074 ) ;
  assign n44532 = ~n7808 & n32234 ;
  assign n44533 = ~n44531 & n44532 ;
  assign n44534 = n23512 ^ n9278 ^ 1'b0 ;
  assign n44535 = ~n6346 & n44534 ;
  assign n44536 = n29656 | n30183 ;
  assign n44537 = n26374 ^ n22189 ^ 1'b0 ;
  assign n44538 = n14049 | n44537 ;
  assign n44540 = n13648 & ~n13792 ;
  assign n44539 = n24771 ^ n14652 ^ 1'b0 ;
  assign n44541 = n44540 ^ n44539 ^ n33075 ;
  assign n44542 = n14031 & n24906 ;
  assign n44543 = n44542 ^ n14691 ^ n14226 ;
  assign n44544 = ( n6222 & n10989 ) | ( n6222 & n19363 ) | ( n10989 & n19363 ) ;
  assign n44545 = n10679 | n44544 ;
  assign n44546 = ( n4117 & n9089 ) | ( n4117 & ~n44545 ) | ( n9089 & ~n44545 ) ;
  assign n44547 = n5602 ^ n5481 ^ 1'b0 ;
  assign n44548 = n44547 ^ n12560 ^ 1'b0 ;
  assign n44549 = ~n12132 & n44548 ;
  assign n44550 = n44549 ^ n34443 ^ n22282 ;
  assign n44551 = n44550 ^ n42698 ^ n16180 ;
  assign n44552 = n44551 ^ n21823 ^ n322 ;
  assign n44553 = ~n21414 & n29591 ;
  assign n44554 = n14062 ^ n354 ^ 1'b0 ;
  assign n44555 = n13881 ^ n2820 ^ 1'b0 ;
  assign n44556 = n8493 & n44555 ;
  assign n44557 = n44556 ^ n21341 ^ n14003 ;
  assign n44558 = ~n44554 & n44557 ;
  assign n44559 = n40184 & n44558 ;
  assign n44560 = n28548 ^ n4553 ^ n4066 ;
  assign n44561 = ( n11237 & n25262 ) | ( n11237 & ~n39082 ) | ( n25262 & ~n39082 ) ;
  assign n44562 = ( n29224 & n41346 ) | ( n29224 & n42729 ) | ( n41346 & n42729 ) ;
  assign n44563 = n18531 ^ n7659 ^ 1'b0 ;
  assign n44564 = ~n7110 & n44563 ;
  assign n44565 = n3422 | n27487 ;
  assign n44566 = n11495 & ~n44565 ;
  assign n44567 = n44566 ^ n32871 ^ n5524 ;
  assign n44568 = n7754 | n8198 ;
  assign n44569 = n44567 & ~n44568 ;
  assign n44570 = n13146 & ~n44569 ;
  assign n44571 = n44570 ^ n36434 ^ 1'b0 ;
  assign n44572 = n22992 | n33162 ;
  assign n44573 = n21636 | n44572 ;
  assign n44574 = n28440 | n44573 ;
  assign n44575 = ( n13127 & n17764 ) | ( n13127 & ~n29165 ) | ( n17764 & ~n29165 ) ;
  assign n44576 = n44575 ^ n5452 ^ n4351 ;
  assign n44582 = ( n13761 & ~n18289 ) | ( n13761 & n20458 ) | ( ~n18289 & n20458 ) ;
  assign n44577 = n16499 ^ n4732 ^ 1'b0 ;
  assign n44578 = n44577 ^ n6218 ^ 1'b0 ;
  assign n44579 = n14315 & ~n14486 ;
  assign n44580 = n37199 | n44579 ;
  assign n44581 = n44578 & ~n44580 ;
  assign n44583 = n44582 ^ n44581 ^ n13020 ;
  assign n44584 = ~n13141 & n13504 ;
  assign n44585 = ( n777 & n4662 ) | ( n777 & ~n19872 ) | ( n4662 & ~n19872 ) ;
  assign n44586 = n31434 | n44585 ;
  assign n44587 = n9518 ^ n5063 ^ n1056 ;
  assign n44588 = n26478 ^ n7887 ^ 1'b0 ;
  assign n44589 = n44587 | n44588 ;
  assign n44590 = n29577 ^ n25917 ^ n16626 ;
  assign n44591 = n44590 ^ n21628 ^ 1'b0 ;
  assign n44592 = n44591 ^ n25041 ^ 1'b0 ;
  assign n44593 = n29089 & n44592 ;
  assign n44594 = n477 & n7840 ;
  assign n44595 = n44594 ^ n4889 ^ 1'b0 ;
  assign n44596 = n9978 & ~n22899 ;
  assign n44597 = ~n5500 & n18839 ;
  assign n44600 = n28229 ^ n16924 ^ n8265 ;
  assign n44601 = ~n26141 & n44600 ;
  assign n44602 = n8970 & n44601 ;
  assign n44598 = ~n6708 & n21214 ;
  assign n44599 = n36067 | n44598 ;
  assign n44603 = n44602 ^ n44599 ^ n40202 ;
  assign n44604 = n44603 ^ n5629 ^ 1'b0 ;
  assign n44605 = ~n28370 & n36791 ;
  assign n44606 = n40688 & n44605 ;
  assign n44607 = ( n44597 & n44604 ) | ( n44597 & ~n44606 ) | ( n44604 & ~n44606 ) ;
  assign n44608 = n31869 ^ n29124 ^ 1'b0 ;
  assign n44609 = ( n1671 & n2737 ) | ( n1671 & ~n6514 ) | ( n2737 & ~n6514 ) ;
  assign n44610 = n44609 ^ n15773 ^ n7867 ;
  assign n44611 = n16180 ^ n10240 ^ 1'b0 ;
  assign n44612 = n33121 & ~n44611 ;
  assign n44613 = ( n5599 & n14130 ) | ( n5599 & ~n18354 ) | ( n14130 & ~n18354 ) ;
  assign n44614 = n44613 ^ n10150 ^ 1'b0 ;
  assign n44615 = ~n21175 & n44614 ;
  assign n44616 = n15818 & n38729 ;
  assign n44617 = n24446 ^ n8041 ^ 1'b0 ;
  assign n44618 = n26645 ^ n26151 ^ 1'b0 ;
  assign n44619 = n26277 | n44618 ;
  assign n44620 = n3361 & n23572 ;
  assign n44621 = ~n2436 & n15981 ;
  assign n44622 = n11879 & n44621 ;
  assign n44623 = ( ~n25829 & n44620 ) | ( ~n25829 & n44622 ) | ( n44620 & n44622 ) ;
  assign n44624 = ( n8206 & n22527 ) | ( n8206 & ~n36139 ) | ( n22527 & ~n36139 ) ;
  assign n44625 = n9963 & n44624 ;
  assign n44626 = ( n2277 & ~n6952 ) | ( n2277 & n19981 ) | ( ~n6952 & n19981 ) ;
  assign n44627 = ( ~n26329 & n35097 ) | ( ~n26329 & n44626 ) | ( n35097 & n44626 ) ;
  assign n44628 = n44627 ^ n33644 ^ n10369 ;
  assign n44631 = n3697 | n4449 ;
  assign n44629 = ~n10873 & n40280 ;
  assign n44630 = n44629 ^ n4248 ^ 1'b0 ;
  assign n44632 = n44631 ^ n44630 ^ n8478 ;
  assign n44633 = n21284 | n43757 ;
  assign n44634 = n15764 ^ n8743 ^ 1'b0 ;
  assign n44635 = ~n3198 & n44634 ;
  assign n44636 = ~n1095 & n36545 ;
  assign n44637 = n44636 ^ n34762 ^ 1'b0 ;
  assign n44639 = n19234 ^ n15693 ^ 1'b0 ;
  assign n44640 = n44639 ^ n12609 ^ 1'b0 ;
  assign n44641 = n9118 & ~n44640 ;
  assign n44638 = ~n33402 & n37624 ;
  assign n44642 = n44641 ^ n44638 ^ 1'b0 ;
  assign n44643 = n23159 ^ n2474 ^ n1487 ;
  assign n44644 = n10559 ^ n6184 ^ n1923 ;
  assign n44645 = n23857 ^ n5823 ^ n838 ;
  assign n44646 = ~n23770 & n44645 ;
  assign n44647 = n44646 ^ n9061 ^ 1'b0 ;
  assign n44648 = ~n9578 & n39927 ;
  assign n44649 = n44648 ^ n12638 ^ n4632 ;
  assign n44650 = ~n44647 & n44649 ;
  assign n44654 = ( n1415 & n18600 ) | ( n1415 & ~n19583 ) | ( n18600 & ~n19583 ) ;
  assign n44655 = n44654 ^ n37327 ^ n26110 ;
  assign n44652 = ( ~n3044 & n4208 ) | ( ~n3044 & n4443 ) | ( n4208 & n4443 ) ;
  assign n44651 = n11708 ^ n8033 ^ n2324 ;
  assign n44653 = n44652 ^ n44651 ^ n13303 ;
  assign n44656 = n44655 ^ n44653 ^ n39906 ;
  assign n44657 = n17656 & n30379 ;
  assign n44658 = ( n19626 & ~n28772 ) | ( n19626 & n44657 ) | ( ~n28772 & n44657 ) ;
  assign n44659 = n1222 | n30641 ;
  assign n44660 = n13572 | n40620 ;
  assign n44661 = n44659 & ~n44660 ;
  assign n44662 = n12915 | n44661 ;
  assign n44663 = ( n21536 & n29371 ) | ( n21536 & ~n34262 ) | ( n29371 & ~n34262 ) ;
  assign n44664 = n44663 ^ n25354 ^ 1'b0 ;
  assign n44665 = ~n39727 & n44664 ;
  assign n44666 = n44053 ^ n16786 ^ n3840 ;
  assign n44667 = n21745 & n24763 ;
  assign n44674 = ~n8460 & n17572 ;
  assign n44675 = n44674 ^ n20453 ^ 1'b0 ;
  assign n44671 = n4473 | n7879 ;
  assign n44672 = n44671 ^ n7285 ^ 1'b0 ;
  assign n44668 = n3286 & n12984 ;
  assign n44669 = n44668 ^ x30 ^ 1'b0 ;
  assign n44670 = n24188 & ~n44669 ;
  assign n44673 = n44672 ^ n44670 ^ 1'b0 ;
  assign n44676 = n44675 ^ n44673 ^ n4108 ;
  assign n44677 = ( ~n19186 & n44667 ) | ( ~n19186 & n44676 ) | ( n44667 & n44676 ) ;
  assign n44682 = n7425 ^ n3918 ^ n2386 ;
  assign n44679 = n1181 & ~n4958 ;
  assign n44680 = ~n3076 & n44679 ;
  assign n44678 = n12902 & ~n20046 ;
  assign n44681 = n44680 ^ n44678 ^ 1'b0 ;
  assign n44683 = n44682 ^ n44681 ^ n37149 ;
  assign n44684 = n9387 & ~n42405 ;
  assign n44685 = ( n19448 & n29076 ) | ( n19448 & ~n37046 ) | ( n29076 & ~n37046 ) ;
  assign n44686 = n44685 ^ n31654 ^ 1'b0 ;
  assign n44687 = n20088 ^ n8073 ^ 1'b0 ;
  assign n44688 = ~n6624 & n44687 ;
  assign n44689 = n10793 & ~n44688 ;
  assign n44690 = ( ~n8630 & n38424 ) | ( ~n8630 & n44012 ) | ( n38424 & n44012 ) ;
  assign n44691 = n44690 ^ n38337 ^ n867 ;
  assign n44692 = n44691 ^ n9473 ^ n5306 ;
  assign n44693 = n35008 ^ n25592 ^ 1'b0 ;
  assign n44694 = ~n44692 & n44693 ;
  assign n44695 = n44694 ^ n22100 ^ n4212 ;
  assign n44696 = n32069 & ~n44695 ;
  assign n44697 = ( ~n3247 & n34301 ) | ( ~n3247 & n41754 ) | ( n34301 & n41754 ) ;
  assign n44698 = ( x76 & n3968 ) | ( x76 & n28115 ) | ( n3968 & n28115 ) ;
  assign n44699 = ( ~n590 & n29312 ) | ( ~n590 & n44698 ) | ( n29312 & n44698 ) ;
  assign n44700 = n23826 ^ n17678 ^ n5029 ;
  assign n44701 = n21924 ^ n16986 ^ n10052 ;
  assign n44702 = ( n38635 & n44700 ) | ( n38635 & ~n44701 ) | ( n44700 & ~n44701 ) ;
  assign n44703 = ( n8254 & n34041 ) | ( n8254 & ~n44702 ) | ( n34041 & ~n44702 ) ;
  assign n44704 = n8098 & ~n42816 ;
  assign n44705 = n44704 ^ n16288 ^ 1'b0 ;
  assign n44706 = n44705 ^ n3369 ^ 1'b0 ;
  assign n44707 = ~n2497 & n44706 ;
  assign n44708 = ( n6822 & ~n44600 ) | ( n6822 & n44707 ) | ( ~n44600 & n44707 ) ;
  assign n44709 = n13250 | n31215 ;
  assign n44710 = ( n5217 & n22925 ) | ( n5217 & n25217 ) | ( n22925 & n25217 ) ;
  assign n44711 = n44710 ^ n17891 ^ 1'b0 ;
  assign n44712 = n44711 ^ n17565 ^ n10125 ;
  assign n44713 = n44712 ^ n35869 ^ 1'b0 ;
  assign n44714 = n44713 ^ n3016 ^ 1'b0 ;
  assign n44715 = n43057 | n44714 ;
  assign n44717 = ( n11475 & ~n17700 ) | ( n11475 & n24743 ) | ( ~n17700 & n24743 ) ;
  assign n44716 = n14153 | n22523 ;
  assign n44718 = n44717 ^ n44716 ^ 1'b0 ;
  assign n44719 = n44718 ^ n20169 ^ 1'b0 ;
  assign n44720 = n8593 & ~n44719 ;
  assign n44721 = n20910 ^ n16958 ^ 1'b0 ;
  assign n44722 = n6502 ^ n2469 ^ n1152 ;
  assign n44723 = ( n37855 & ~n44721 ) | ( n37855 & n44722 ) | ( ~n44721 & n44722 ) ;
  assign n44724 = ( ~n8757 & n26332 ) | ( ~n8757 & n32068 ) | ( n26332 & n32068 ) ;
  assign n44725 = ( n18651 & n22313 ) | ( n18651 & n44724 ) | ( n22313 & n44724 ) ;
  assign n44726 = ( n32398 & ~n37970 ) | ( n32398 & n44725 ) | ( ~n37970 & n44725 ) ;
  assign n44727 = n13797 ^ n13535 ^ 1'b0 ;
  assign n44728 = n41474 ^ n18950 ^ 1'b0 ;
  assign n44729 = ~n31492 & n44728 ;
  assign n44730 = n39256 & n44729 ;
  assign n44731 = ~n33290 & n44730 ;
  assign n44732 = n11732 & n14156 ;
  assign n44733 = n37084 & n44732 ;
  assign n44734 = n1826 | n44733 ;
  assign n44735 = n44734 ^ n26247 ^ 1'b0 ;
  assign n44736 = n35208 | n44735 ;
  assign n44737 = n44731 & ~n44736 ;
  assign n44738 = n276 | n5166 ;
  assign n44739 = n8416 | n44738 ;
  assign n44740 = ~n17846 & n37078 ;
  assign n44741 = ~n28988 & n44740 ;
  assign n44742 = n3506 | n23704 ;
  assign n44743 = n27333 & ~n44742 ;
  assign n44744 = n8392 & n16857 ;
  assign n44745 = n44744 ^ n20818 ^ n5857 ;
  assign n44746 = ~n7263 & n43587 ;
  assign n44747 = n14530 & ~n44746 ;
  assign n44748 = n44747 ^ n12087 ^ 1'b0 ;
  assign n44749 = ( n5347 & ~n37901 ) | ( n5347 & n44748 ) | ( ~n37901 & n44748 ) ;
  assign n44750 = ( n259 & ~n2553 ) | ( n259 & n19195 ) | ( ~n2553 & n19195 ) ;
  assign n44751 = n12887 & ~n44750 ;
  assign n44752 = ( ~n2036 & n5455 ) | ( ~n2036 & n44751 ) | ( n5455 & n44751 ) ;
  assign n44753 = n20937 & ~n44752 ;
  assign n44754 = n2077 & ~n11679 ;
  assign n44755 = n18722 & n44754 ;
  assign n44756 = ~n2812 & n10585 ;
  assign n44757 = ( n23736 & ~n33493 ) | ( n23736 & n44756 ) | ( ~n33493 & n44756 ) ;
  assign n44758 = n12270 & ~n27976 ;
  assign n44759 = n44758 ^ n43713 ^ 1'b0 ;
  assign n44760 = n44759 ^ n25642 ^ 1'b0 ;
  assign n44761 = n7708 & ~n17362 ;
  assign n44762 = ~n6235 & n16761 ;
  assign n44763 = n44762 ^ n27504 ^ n7204 ;
  assign n44764 = n44763 ^ n21770 ^ n9994 ;
  assign n44765 = ~n3069 & n41375 ;
  assign n44766 = n44765 ^ n17689 ^ 1'b0 ;
  assign n44767 = ~n8700 & n44766 ;
  assign n44768 = ( ~n2941 & n17527 ) | ( ~n2941 & n44767 ) | ( n17527 & n44767 ) ;
  assign n44769 = ( ~n12419 & n16213 ) | ( ~n12419 & n44768 ) | ( n16213 & n44768 ) ;
  assign n44773 = n19731 ^ n16108 ^ n10672 ;
  assign n44770 = n34328 ^ n25070 ^ 1'b0 ;
  assign n44771 = n10010 | n44770 ;
  assign n44772 = n15614 & ~n44771 ;
  assign n44774 = n44773 ^ n44772 ^ 1'b0 ;
  assign n44775 = ( ~n42340 & n44769 ) | ( ~n42340 & n44774 ) | ( n44769 & n44774 ) ;
  assign n44777 = n28928 | n34370 ;
  assign n44776 = ~n6988 & n17273 ;
  assign n44778 = n44777 ^ n44776 ^ 1'b0 ;
  assign n44780 = ( n10563 & n14474 ) | ( n10563 & n24473 ) | ( n14474 & n24473 ) ;
  assign n44779 = n30959 ^ n15643 ^ n7586 ;
  assign n44781 = n44780 ^ n44779 ^ n5599 ;
  assign n44782 = n33790 ^ n2227 ^ 1'b0 ;
  assign n44783 = n25440 & ~n26790 ;
  assign n44784 = ( n9227 & n26504 ) | ( n9227 & ~n28757 ) | ( n26504 & ~n28757 ) ;
  assign n44785 = n19521 | n44784 ;
  assign n44786 = ~n44783 & n44785 ;
  assign n44787 = ( n30724 & ~n33318 ) | ( n30724 & n42996 ) | ( ~n33318 & n42996 ) ;
  assign n44789 = n37809 ^ n11021 ^ n8276 ;
  assign n44788 = n17276 & n31326 ;
  assign n44790 = n44789 ^ n44788 ^ 1'b0 ;
  assign n44791 = ( n4175 & n11111 ) | ( n4175 & n44790 ) | ( n11111 & n44790 ) ;
  assign n44792 = ( n31631 & n40063 ) | ( n31631 & ~n41440 ) | ( n40063 & ~n41440 ) ;
  assign n44793 = n44792 ^ n12983 ^ 1'b0 ;
  assign n44794 = ~n44791 & n44793 ;
  assign n44795 = n23472 ^ n6319 ^ n1240 ;
  assign n44796 = n25316 ^ n15937 ^ 1'b0 ;
  assign n44797 = n44795 | n44796 ;
  assign n44798 = n42767 & ~n44797 ;
  assign n44799 = n22436 ^ n9431 ^ 1'b0 ;
  assign n44800 = n9804 ^ x181 ^ 1'b0 ;
  assign n44801 = ~n10692 & n44800 ;
  assign n44802 = n41842 ^ n11196 ^ n4391 ;
  assign n44805 = n2748 | n10284 ;
  assign n44804 = n38712 ^ n12296 ^ 1'b0 ;
  assign n44803 = n1477 & n37172 ;
  assign n44806 = n44805 ^ n44804 ^ n44803 ;
  assign n44809 = ( n1915 & n3977 ) | ( n1915 & n17378 ) | ( n3977 & n17378 ) ;
  assign n44810 = n44809 ^ n16256 ^ 1'b0 ;
  assign n44807 = n1943 | n14707 ;
  assign n44808 = n18120 | n44807 ;
  assign n44811 = n44810 ^ n44808 ^ n4101 ;
  assign n44812 = n1101 & ~n40304 ;
  assign n44813 = n627 | n8438 ;
  assign n44814 = n41292 ^ n28965 ^ n1462 ;
  assign n44815 = n44814 ^ n12078 ^ 1'b0 ;
  assign n44816 = x56 & n37034 ;
  assign n44817 = n8038 & ~n28000 ;
  assign n44818 = n33827 & n44817 ;
  assign n44819 = ( ~n38127 & n38275 ) | ( ~n38127 & n42766 ) | ( n38275 & n42766 ) ;
  assign n44820 = n44819 ^ n19474 ^ 1'b0 ;
  assign n44821 = n22174 ^ n4889 ^ 1'b0 ;
  assign n44822 = ~n5196 & n8926 ;
  assign n44823 = n44822 ^ n6241 ^ 1'b0 ;
  assign n44824 = n17628 ^ n1991 ^ 1'b0 ;
  assign n44825 = n44823 & n44824 ;
  assign n44826 = n44825 ^ n23700 ^ 1'b0 ;
  assign n44827 = ( n27655 & n44821 ) | ( n27655 & n44826 ) | ( n44821 & n44826 ) ;
  assign n44828 = ~n9377 & n26043 ;
  assign n44829 = n15772 & n44828 ;
  assign n44830 = n14787 & ~n44829 ;
  assign n44831 = n23524 ^ n8878 ^ n311 ;
  assign n44832 = n25163 ^ n14609 ^ 1'b0 ;
  assign n44833 = n43757 ^ n40000 ^ 1'b0 ;
  assign n44834 = n44832 & n44833 ;
  assign n44835 = n44834 ^ n37323 ^ 1'b0 ;
  assign n44836 = n2616 & n4248 ;
  assign n44837 = n38855 & ~n44836 ;
  assign n44838 = n2777 & ~n25783 ;
  assign n44839 = ( n4851 & ~n5360 ) | ( n4851 & n44838 ) | ( ~n5360 & n44838 ) ;
  assign n44840 = n41621 ^ n5545 ^ 1'b0 ;
  assign n44841 = ( n14816 & n15207 ) | ( n14816 & ~n18596 ) | ( n15207 & ~n18596 ) ;
  assign n44842 = n44841 ^ n13341 ^ n5969 ;
  assign n44843 = ( n37923 & n44840 ) | ( n37923 & n44842 ) | ( n44840 & n44842 ) ;
  assign n44844 = n8011 ^ n6918 ^ 1'b0 ;
  assign n44845 = n44844 ^ n13450 ^ n9805 ;
  assign n44846 = ( n9825 & n36437 ) | ( n9825 & n44845 ) | ( n36437 & n44845 ) ;
  assign n44847 = ~n22065 & n28817 ;
  assign n44848 = n44847 ^ n39506 ^ 1'b0 ;
  assign n44849 = ( n6549 & n8240 ) | ( n6549 & n21471 ) | ( n8240 & n21471 ) ;
  assign n44850 = ( n9417 & ~n26172 ) | ( n9417 & n44849 ) | ( ~n26172 & n44849 ) ;
  assign n44851 = ( n2747 & ~n42864 ) | ( n2747 & n44850 ) | ( ~n42864 & n44850 ) ;
  assign n44852 = n10270 & ~n44851 ;
  assign n44853 = ~n33847 & n44852 ;
  assign n44855 = n3474 | n8844 ;
  assign n44856 = n44855 ^ n1888 ^ 1'b0 ;
  assign n44854 = ( n7725 & n12215 ) | ( n7725 & ~n34797 ) | ( n12215 & ~n34797 ) ;
  assign n44857 = n44856 ^ n44854 ^ 1'b0 ;
  assign n44858 = ( ~n1385 & n16616 ) | ( ~n1385 & n31106 ) | ( n16616 & n31106 ) ;
  assign n44859 = ( n21182 & ~n44283 ) | ( n21182 & n44858 ) | ( ~n44283 & n44858 ) ;
  assign n44860 = n29052 ^ n2412 ^ 1'b0 ;
  assign n44861 = n25783 ^ n5327 ^ n1603 ;
  assign n44862 = ( n10020 & n19664 ) | ( n10020 & ~n44861 ) | ( n19664 & ~n44861 ) ;
  assign n44864 = n8158 & n14584 ;
  assign n44865 = n3865 & n44864 ;
  assign n44863 = n23968 ^ n15967 ^ 1'b0 ;
  assign n44866 = n44865 ^ n44863 ^ n40898 ;
  assign n44867 = n20032 ^ n5928 ^ 1'b0 ;
  assign n44868 = n4624 & n28979 ;
  assign n44869 = n40185 ^ n17208 ^ 1'b0 ;
  assign n44870 = n44868 & n44869 ;
  assign n44871 = n35749 ^ n29365 ^ 1'b0 ;
  assign n44872 = n14913 ^ n12728 ^ n3509 ;
  assign n44873 = n20063 & ~n44872 ;
  assign n44874 = n44873 ^ n366 ^ 1'b0 ;
  assign n44877 = n2705 & ~n7650 ;
  assign n44875 = n13464 ^ n1582 ^ 1'b0 ;
  assign n44876 = n28761 | n44875 ;
  assign n44878 = n44877 ^ n44876 ^ n6748 ;
  assign n44879 = n31346 ^ n23296 ^ n1818 ;
  assign n44880 = n44879 ^ n36081 ^ 1'b0 ;
  assign n44881 = n1938 & ~n9359 ;
  assign n44882 = n2934 & n44881 ;
  assign n44883 = n20952 & n21696 ;
  assign n44884 = ~n36287 & n44883 ;
  assign n44885 = n24582 ^ n10206 ^ 1'b0 ;
  assign n44886 = ( n10888 & n27114 ) | ( n10888 & n41556 ) | ( n27114 & n41556 ) ;
  assign n44887 = n41101 ^ n37155 ^ 1'b0 ;
  assign n44888 = n22599 ^ n7401 ^ 1'b0 ;
  assign n44889 = ( n7414 & n30564 ) | ( n7414 & n33171 ) | ( n30564 & n33171 ) ;
  assign n44890 = ( n7160 & ~n44888 ) | ( n7160 & n44889 ) | ( ~n44888 & n44889 ) ;
  assign n44891 = n5317 & n17075 ;
  assign n44892 = n44891 ^ n22914 ^ 1'b0 ;
  assign n44893 = n25520 & n32990 ;
  assign n44894 = n44893 ^ n12893 ^ 1'b0 ;
  assign n44895 = n3548 ^ n3321 ^ 1'b0 ;
  assign n44896 = n17155 ^ n9851 ^ 1'b0 ;
  assign n44897 = n25777 & ~n44896 ;
  assign n44898 = ~n44895 & n44897 ;
  assign n44899 = n44898 ^ n11438 ^ 1'b0 ;
  assign n44900 = n13256 & ~n16863 ;
  assign n44901 = n44900 ^ n12976 ^ 1'b0 ;
  assign n44902 = n21800 ^ n5094 ^ 1'b0 ;
  assign n44903 = ~n44901 & n44902 ;
  assign n44904 = ( n21421 & n25904 ) | ( n21421 & n38689 ) | ( n25904 & n38689 ) ;
  assign n44906 = n27821 ^ n19844 ^ n680 ;
  assign n44905 = n4322 & ~n5112 ;
  assign n44907 = n44906 ^ n44905 ^ 1'b0 ;
  assign n44908 = ~n14429 & n44907 ;
  assign n44909 = ( n5244 & n5549 ) | ( n5244 & n18856 ) | ( n5549 & n18856 ) ;
  assign n44910 = n44909 ^ n34604 ^ 1'b0 ;
  assign n44911 = n23820 & n44910 ;
  assign n44912 = ( n15680 & n44908 ) | ( n15680 & n44911 ) | ( n44908 & n44911 ) ;
  assign n44913 = n10552 & ~n12386 ;
  assign n44914 = n44913 ^ n20616 ^ n19827 ;
  assign n44915 = ( n11527 & ~n26745 ) | ( n11527 & n28167 ) | ( ~n26745 & n28167 ) ;
  assign n44916 = n31906 ^ n18283 ^ n15339 ;
  assign n44917 = n8864 & n35218 ;
  assign n44918 = n5017 & n9468 ;
  assign n44919 = n44918 ^ n13305 ^ n7472 ;
  assign n44920 = n41109 ^ n13131 ^ 1'b0 ;
  assign n44921 = n11318 & ~n44920 ;
  assign n44922 = ( n6534 & n6856 ) | ( n6534 & ~n31166 ) | ( n6856 & ~n31166 ) ;
  assign n44923 = n9718 & ~n28188 ;
  assign n44924 = n44923 ^ n26233 ^ 1'b0 ;
  assign n44925 = ( n14263 & ~n27594 ) | ( n14263 & n44924 ) | ( ~n27594 & n44924 ) ;
  assign n44926 = n4471 & n41974 ;
  assign n44927 = n44926 ^ n8719 ^ x0 ;
  assign n44928 = ( n4544 & ~n4952 ) | ( n4544 & n31775 ) | ( ~n4952 & n31775 ) ;
  assign n44929 = ( n4121 & ~n14821 ) | ( n4121 & n21081 ) | ( ~n14821 & n21081 ) ;
  assign n44930 = n11319 & ~n17385 ;
  assign n44931 = n44930 ^ n9378 ^ 1'b0 ;
  assign n44932 = ~n4343 & n44931 ;
  assign n44933 = n16650 ^ n10141 ^ 1'b0 ;
  assign n44934 = n25761 & n36869 ;
  assign n44935 = ~n11795 & n44934 ;
  assign n44936 = ( n11947 & ~n27281 ) | ( n11947 & n31667 ) | ( ~n27281 & n31667 ) ;
  assign n44937 = ~n3488 & n14058 ;
  assign n44938 = ~n7465 & n30101 ;
  assign n44939 = ( n15820 & n38368 ) | ( n15820 & n44938 ) | ( n38368 & n44938 ) ;
  assign n44940 = ~n5873 & n26501 ;
  assign n44941 = ~n23015 & n44940 ;
  assign n44942 = n44941 ^ n14791 ^ 1'b0 ;
  assign n44948 = n7107 & n14425 ;
  assign n44944 = n44797 ^ n29228 ^ 1'b0 ;
  assign n44945 = n36662 ^ n20905 ^ n4001 ;
  assign n44946 = n44944 & ~n44945 ;
  assign n44947 = n10451 & n44946 ;
  assign n44949 = n44948 ^ n44947 ^ 1'b0 ;
  assign n44943 = n10199 & ~n28118 ;
  assign n44950 = n44949 ^ n44943 ^ 1'b0 ;
  assign n44951 = n29914 ^ n10002 ^ n1623 ;
  assign n44952 = n44951 ^ n13735 ^ 1'b0 ;
  assign n44953 = ~n37075 & n44952 ;
  assign n44954 = n44953 ^ n18164 ^ 1'b0 ;
  assign n44955 = n25237 ^ n7703 ^ 1'b0 ;
  assign n44958 = n21397 ^ n19984 ^ 1'b0 ;
  assign n44959 = ~n9111 & n44958 ;
  assign n44957 = n9920 & n14164 ;
  assign n44956 = ~n24382 & n36437 ;
  assign n44960 = n44959 ^ n44957 ^ n44956 ;
  assign n44961 = n32460 ^ n25293 ^ n7777 ;
  assign n44962 = n15653 ^ n7180 ^ 1'b0 ;
  assign n44963 = n30675 | n44962 ;
  assign n44964 = n18509 ^ n18100 ^ 1'b0 ;
  assign n44965 = n44963 | n44964 ;
  assign n44966 = n12596 | n18743 ;
  assign n44967 = n44965 & ~n44966 ;
  assign n44968 = ( n2160 & n32672 ) | ( n2160 & n44967 ) | ( n32672 & n44967 ) ;
  assign n44969 = ~n1850 & n39472 ;
  assign n44970 = n44969 ^ n35701 ^ n15985 ;
  assign n44971 = ( n7790 & ~n26820 ) | ( n7790 & n37789 ) | ( ~n26820 & n37789 ) ;
  assign n44972 = n44971 ^ n9856 ^ n8528 ;
  assign n44973 = n21938 ^ n16006 ^ 1'b0 ;
  assign n44974 = n44973 ^ n19905 ^ n2596 ;
  assign n44975 = n44974 ^ n4810 ^ n1353 ;
  assign n44976 = n11162 ^ n10569 ^ 1'b0 ;
  assign n44977 = n1380 & ~n44976 ;
  assign n44978 = n40341 & n44977 ;
  assign n44979 = ( ~n8446 & n21189 ) | ( ~n8446 & n44978 ) | ( n21189 & n44978 ) ;
  assign n44980 = n2904 | n6750 ;
  assign n44981 = n2646 & ~n44980 ;
  assign n44982 = n25987 ^ n17156 ^ 1'b0 ;
  assign n44983 = n4536 | n44982 ;
  assign n44984 = n5885 & ~n27640 ;
  assign n44985 = n29105 ^ n2395 ^ 1'b0 ;
  assign n44986 = n26400 | n44985 ;
  assign n44987 = n44986 ^ n680 ^ 1'b0 ;
  assign n44988 = n851 & n29376 ;
  assign n44989 = n44988 ^ n34262 ^ 1'b0 ;
  assign n44990 = n11140 | n38282 ;
  assign n44991 = ~n12093 & n12805 ;
  assign n44992 = ( n1506 & n30861 ) | ( n1506 & n44991 ) | ( n30861 & n44991 ) ;
  assign n44993 = n22891 & n27260 ;
  assign n44994 = n24861 ^ n9257 ^ 1'b0 ;
  assign n44995 = ( n7206 & n33067 ) | ( n7206 & n44994 ) | ( n33067 & n44994 ) ;
  assign n44996 = n34358 ^ n17648 ^ 1'b0 ;
  assign n44997 = n42604 & ~n44996 ;
  assign n44998 = n2152 & n18977 ;
  assign n44999 = ~n20257 & n44162 ;
  assign n45002 = n8514 ^ n3225 ^ n2444 ;
  assign n45000 = n2045 & n21350 ;
  assign n45001 = n45000 ^ n12073 ^ 1'b0 ;
  assign n45003 = n45002 ^ n45001 ^ n10398 ;
  assign n45004 = ( n34757 & n37407 ) | ( n34757 & n40240 ) | ( n37407 & n40240 ) ;
  assign n45005 = n42336 ^ n34149 ^ 1'b0 ;
  assign n45006 = n45005 ^ n33634 ^ n11008 ;
  assign n45007 = n43155 ^ n40440 ^ n5500 ;
  assign n45008 = ~n14970 & n45007 ;
  assign n45009 = n45008 ^ n23573 ^ 1'b0 ;
  assign n45010 = n30028 ^ n29849 ^ n23972 ;
  assign n45011 = n45010 ^ n11312 ^ 1'b0 ;
  assign n45012 = n35027 & n45011 ;
  assign n45013 = n13364 & n34081 ;
  assign n45014 = ( n4102 & ~n4360 ) | ( n4102 & n29520 ) | ( ~n4360 & n29520 ) ;
  assign n45015 = n36445 ^ n5447 ^ 1'b0 ;
  assign n45016 = n45014 | n45015 ;
  assign n45017 = n16378 ^ n3203 ^ 1'b0 ;
  assign n45018 = n3196 | n4412 ;
  assign n45019 = n2750 & n4540 ;
  assign n45020 = n45019 ^ n37687 ^ 1'b0 ;
  assign n45021 = ( ~n4190 & n11565 ) | ( ~n4190 & n12960 ) | ( n11565 & n12960 ) ;
  assign n45022 = n45021 ^ n4107 ^ n587 ;
  assign n45023 = n22897 ^ n14821 ^ 1'b0 ;
  assign n45024 = n9449 | n14323 ;
  assign n45025 = n45024 ^ n41454 ^ 1'b0 ;
  assign n45026 = n27705 ^ n9610 ^ 1'b0 ;
  assign n45027 = ~n7487 & n45026 ;
  assign n45028 = n45027 ^ n32494 ^ 1'b0 ;
  assign n45029 = n12313 & ~n45028 ;
  assign n45030 = n11938 & n31811 ;
  assign n45036 = n6433 & ~n21574 ;
  assign n45037 = n45036 ^ n38391 ^ 1'b0 ;
  assign n45038 = n45037 ^ n10631 ^ n1212 ;
  assign n45031 = n4796 & n25030 ;
  assign n45032 = n9413 | n45031 ;
  assign n45033 = n10983 & ~n45032 ;
  assign n45034 = n24639 & ~n45033 ;
  assign n45035 = ( n17611 & n21754 ) | ( n17611 & n45034 ) | ( n21754 & n45034 ) ;
  assign n45039 = n45038 ^ n45035 ^ 1'b0 ;
  assign n45040 = n16680 ^ n15892 ^ n13708 ;
  assign n45041 = n38697 & ~n45040 ;
  assign n45042 = n45041 ^ n12734 ^ 1'b0 ;
  assign n45043 = n45042 ^ n5347 ^ 1'b0 ;
  assign n45044 = n15120 ^ n7293 ^ n7094 ;
  assign n45045 = ( n15990 & ~n17302 ) | ( n15990 & n45044 ) | ( ~n17302 & n45044 ) ;
  assign n45046 = n3757 & ~n27480 ;
  assign n45047 = n45046 ^ n16031 ^ 1'b0 ;
  assign n45048 = n45047 ^ n26793 ^ n8165 ;
  assign n45049 = n9255 & n21499 ;
  assign n45050 = n10489 & ~n45049 ;
  assign n45051 = n17533 & n45050 ;
  assign n45052 = n299 | n44797 ;
  assign n45053 = n45051 & ~n45052 ;
  assign n45054 = n22452 ^ n14684 ^ n14302 ;
  assign n45055 = n14665 ^ n10551 ^ n5064 ;
  assign n45056 = n14079 & n45055 ;
  assign n45057 = n27788 & n45056 ;
  assign n45058 = ~n45054 & n45057 ;
  assign n45059 = n35237 ^ n17499 ^ n6781 ;
  assign n45060 = n30310 ^ n13702 ^ 1'b0 ;
  assign n45061 = n45059 & n45060 ;
  assign n45062 = n45061 ^ n41988 ^ n1863 ;
  assign n45063 = n295 & n13572 ;
  assign n45064 = ~n5664 & n45063 ;
  assign n45065 = ( n5451 & n34398 ) | ( n5451 & n45064 ) | ( n34398 & n45064 ) ;
  assign n45066 = n5683 & ~n9685 ;
  assign n45067 = n45066 ^ n37422 ^ n19114 ;
  assign n45068 = n8724 & n32828 ;
  assign n45069 = ~n12333 & n45068 ;
  assign n45070 = ( n5444 & n45067 ) | ( n5444 & n45069 ) | ( n45067 & n45069 ) ;
  assign n45071 = n12946 ^ n9851 ^ 1'b0 ;
  assign n45072 = n34294 ^ n12393 ^ 1'b0 ;
  assign n45073 = n21671 | n45072 ;
  assign n45074 = ~n37861 & n40251 ;
  assign n45075 = ~n3762 & n45074 ;
  assign n45076 = ( n3105 & ~n6570 ) | ( n3105 & n9650 ) | ( ~n6570 & n9650 ) ;
  assign n45077 = ( ~n9593 & n13422 ) | ( ~n9593 & n45076 ) | ( n13422 & n45076 ) ;
  assign n45078 = ( n2623 & n41115 ) | ( n2623 & n45077 ) | ( n41115 & n45077 ) ;
  assign n45079 = n15491 ^ n8916 ^ n279 ;
  assign n45080 = n45079 ^ n32638 ^ n4131 ;
  assign n45081 = ( n6572 & ~n13699 ) | ( n6572 & n24695 ) | ( ~n13699 & n24695 ) ;
  assign n45082 = n36565 ^ n15805 ^ n7644 ;
  assign n45083 = n42731 ^ n26795 ^ n6552 ;
  assign n45084 = n45083 ^ n44270 ^ 1'b0 ;
  assign n45085 = ~n7490 & n39049 ;
  assign n45086 = ~n14902 & n24677 ;
  assign n45087 = n45086 ^ n41899 ^ n24519 ;
  assign n45088 = n21945 & n27799 ;
  assign n45089 = n33542 ^ n2478 ^ 1'b0 ;
  assign n45090 = ( n5078 & n7518 ) | ( n5078 & ~n11325 ) | ( n7518 & ~n11325 ) ;
  assign n45091 = ( ~n9046 & n31251 ) | ( ~n9046 & n45090 ) | ( n31251 & n45090 ) ;
  assign n45092 = ( n15841 & ~n25359 ) | ( n15841 & n32112 ) | ( ~n25359 & n32112 ) ;
  assign n45093 = n32782 ^ n20739 ^ n5823 ;
  assign n45094 = n45093 ^ n41075 ^ n26196 ;
  assign n45095 = n1212 & ~n45094 ;
  assign n45096 = ~n30294 & n45095 ;
  assign n45098 = n7929 ^ n4590 ^ 1'b0 ;
  assign n45099 = n18374 | n39385 ;
  assign n45100 = n45098 & ~n45099 ;
  assign n45097 = n12538 ^ n830 ^ 1'b0 ;
  assign n45101 = n45100 ^ n45097 ^ 1'b0 ;
  assign n45102 = n24698 | n45101 ;
  assign n45103 = n3509 ^ n1567 ^ 1'b0 ;
  assign n45104 = n39864 ^ n31492 ^ 1'b0 ;
  assign n45105 = n42884 & ~n45104 ;
  assign n45106 = ( ~n13073 & n13758 ) | ( ~n13073 & n45105 ) | ( n13758 & n45105 ) ;
  assign n45111 = ( ~n10310 & n14013 ) | ( ~n10310 & n17270 ) | ( n14013 & n17270 ) ;
  assign n45107 = ~n20462 & n42852 ;
  assign n45108 = n42294 & n45107 ;
  assign n45109 = n22284 | n24292 ;
  assign n45110 = n45108 & ~n45109 ;
  assign n45112 = n45111 ^ n45110 ^ 1'b0 ;
  assign n45113 = n12015 ^ n3515 ^ n2623 ;
  assign n45114 = n30097 | n45113 ;
  assign n45115 = n1077 & ~n2280 ;
  assign n45116 = n25236 & n45115 ;
  assign n45117 = ( n17838 & ~n22377 ) | ( n17838 & n45116 ) | ( ~n22377 & n45116 ) ;
  assign n45118 = n33089 ^ n14555 ^ n6098 ;
  assign n45119 = n14403 | n23115 ;
  assign n45120 = n10202 | n45119 ;
  assign n45121 = n45120 ^ n30167 ^ n7935 ;
  assign n45122 = n15224 ^ n2499 ^ 1'b0 ;
  assign n45123 = n12577 & n45122 ;
  assign n45124 = ( n16217 & n20143 ) | ( n16217 & n45123 ) | ( n20143 & n45123 ) ;
  assign n45125 = n41826 | n45124 ;
  assign n45126 = n25082 | n41778 ;
  assign n45127 = n45126 ^ n42594 ^ 1'b0 ;
  assign n45128 = ~n1438 & n6037 ;
  assign n45129 = n45128 ^ n5242 ^ 1'b0 ;
  assign n45130 = n20071 & n45129 ;
  assign n45131 = n9668 & ~n27934 ;
  assign n45132 = ~n44230 & n45131 ;
  assign n45133 = n10131 & n45132 ;
  assign n45134 = ( n4481 & n16181 ) | ( n4481 & n38306 ) | ( n16181 & n38306 ) ;
  assign n45135 = n6786 & ~n22155 ;
  assign n45136 = ~n45134 & n45135 ;
  assign n45137 = n3404 | n9607 ;
  assign n45138 = n45137 ^ n9218 ^ 1'b0 ;
  assign n45139 = ( n35432 & ~n45136 ) | ( n35432 & n45138 ) | ( ~n45136 & n45138 ) ;
  assign n45140 = ( ~n38415 & n44359 ) | ( ~n38415 & n45139 ) | ( n44359 & n45139 ) ;
  assign n45141 = n40999 ^ n16078 ^ n14979 ;
  assign n45142 = n13379 | n26724 ;
  assign n45143 = n24036 ^ n20148 ^ n7917 ;
  assign n45144 = n16694 | n36668 ;
  assign n45146 = n14712 ^ n1839 ^ x207 ;
  assign n45145 = n3145 & ~n34406 ;
  assign n45147 = n45146 ^ n45145 ^ 1'b0 ;
  assign n45148 = n28551 ^ n18928 ^ n2359 ;
  assign n45149 = n17519 | n45148 ;
  assign n45150 = n40343 ^ n21386 ^ 1'b0 ;
  assign n45151 = n4918 & n45150 ;
  assign n45152 = ~n3161 & n45151 ;
  assign n45153 = ~n45149 & n45152 ;
  assign n45155 = n40471 ^ n36035 ^ n12460 ;
  assign n45154 = n13494 | n25425 ;
  assign n45156 = n45155 ^ n45154 ^ 1'b0 ;
  assign n45157 = n33912 ^ n24673 ^ 1'b0 ;
  assign n45158 = n37279 ^ n16602 ^ n315 ;
  assign n45159 = n44953 ^ n27257 ^ n16827 ;
  assign n45160 = n34392 ^ n21714 ^ 1'b0 ;
  assign n45161 = n45160 ^ n18420 ^ n10692 ;
  assign n45165 = n18281 ^ n9740 ^ n8174 ;
  assign n45162 = ( ~x238 & n7086 ) | ( ~x238 & n9590 ) | ( n7086 & n9590 ) ;
  assign n45163 = n45162 ^ n22377 ^ 1'b0 ;
  assign n45164 = ( n33316 & ~n33558 ) | ( n33316 & n45163 ) | ( ~n33558 & n45163 ) ;
  assign n45166 = n45165 ^ n45164 ^ n36203 ;
  assign n45167 = ( n8743 & n16191 ) | ( n8743 & n34475 ) | ( n16191 & n34475 ) ;
  assign n45168 = n27709 ^ n3515 ^ 1'b0 ;
  assign n45169 = n24206 & n33046 ;
  assign n45170 = n45169 ^ n31205 ^ 1'b0 ;
  assign n45171 = n22231 & n33522 ;
  assign n45172 = n45171 ^ n27418 ^ 1'b0 ;
  assign n45173 = n36395 | n43155 ;
  assign n45174 = n45173 ^ n2362 ^ 1'b0 ;
  assign n45175 = ( ~n3502 & n23630 ) | ( ~n3502 & n24868 ) | ( n23630 & n24868 ) ;
  assign n45176 = n26489 ^ n2985 ^ n875 ;
  assign n45177 = n2479 & ~n45176 ;
  assign n45178 = n6005 & n45177 ;
  assign n45179 = n45178 ^ n11039 ^ 1'b0 ;
  assign n45180 = ( ~n17461 & n28949 ) | ( ~n17461 & n45179 ) | ( n28949 & n45179 ) ;
  assign n45181 = n22645 ^ n19270 ^ 1'b0 ;
  assign n45182 = n3920 & n35193 ;
  assign n45183 = n21909 & n45182 ;
  assign n45184 = n45181 & ~n45183 ;
  assign n45185 = n12430 & ~n26556 ;
  assign n45186 = n11224 ^ n4199 ^ 1'b0 ;
  assign n45187 = n5084 | n45186 ;
  assign n45188 = n45187 ^ n38151 ^ n17080 ;
  assign n45189 = n6851 & n17854 ;
  assign n45190 = n28771 & n45189 ;
  assign n45191 = n37123 ^ n31723 ^ 1'b0 ;
  assign n45192 = ~n25960 & n42389 ;
  assign n45193 = n45192 ^ n1694 ^ 1'b0 ;
  assign n45194 = n43155 ^ n29063 ^ n5995 ;
  assign n45195 = n25442 & ~n25692 ;
  assign n45196 = n8161 & ~n24526 ;
  assign n45197 = n45196 ^ n7658 ^ 1'b0 ;
  assign n45198 = ( n21859 & n43155 ) | ( n21859 & ~n45197 ) | ( n43155 & ~n45197 ) ;
  assign n45199 = n14075 | n44768 ;
  assign n45200 = n700 | n20382 ;
  assign n45201 = ( ~n716 & n6767 ) | ( ~n716 & n6849 ) | ( n6767 & n6849 ) ;
  assign n45202 = n40638 ^ n5507 ^ 1'b0 ;
  assign n45203 = n45201 | n45202 ;
  assign n45204 = n38915 ^ n2561 ^ 1'b0 ;
  assign n45205 = ~n11349 & n45204 ;
  assign n45206 = ~n6216 & n45205 ;
  assign n45207 = n41450 & n45206 ;
  assign n45214 = ~n4543 & n16793 ;
  assign n45208 = n3230 & n6847 ;
  assign n45209 = n45208 ^ n19847 ^ 1'b0 ;
  assign n45210 = n2860 & n25850 ;
  assign n45211 = n33486 & n45210 ;
  assign n45212 = n45209 | n45211 ;
  assign n45213 = n9255 & ~n45212 ;
  assign n45215 = n45214 ^ n45213 ^ n20453 ;
  assign n45216 = n20476 | n30705 ;
  assign n45217 = n45216 ^ n43897 ^ 1'b0 ;
  assign n45218 = n15224 & n45217 ;
  assign n45219 = ( ~n1390 & n11067 ) | ( ~n1390 & n27996 ) | ( n11067 & n27996 ) ;
  assign n45220 = ~n10076 & n34895 ;
  assign n45221 = ( ~n25064 & n30786 ) | ( ~n25064 & n45220 ) | ( n30786 & n45220 ) ;
  assign n45222 = n29483 & ~n45221 ;
  assign n45223 = n45219 | n45222 ;
  assign n45224 = n34595 ^ n14047 ^ 1'b0 ;
  assign n45225 = n45224 ^ n14581 ^ 1'b0 ;
  assign n45226 = ~n7139 & n45225 ;
  assign n45227 = n24743 ^ n9921 ^ 1'b0 ;
  assign n45228 = n3135 | n3565 ;
  assign n45229 = n26007 | n27001 ;
  assign n45230 = n45228 | n45229 ;
  assign n45231 = ( n10772 & ~n18354 ) | ( n10772 & n45230 ) | ( ~n18354 & n45230 ) ;
  assign n45232 = ~n1412 & n45231 ;
  assign n45233 = n45232 ^ n25917 ^ 1'b0 ;
  assign n45234 = n11719 ^ n5989 ^ 1'b0 ;
  assign n45235 = n28341 | n45234 ;
  assign n45236 = n31633 ^ n3465 ^ 1'b0 ;
  assign n45237 = n12174 & ~n45236 ;
  assign n45238 = ( n21639 & n40368 ) | ( n21639 & n45237 ) | ( n40368 & n45237 ) ;
  assign n45239 = n10730 ^ n2574 ^ n1429 ;
  assign n45240 = ( n18850 & ~n25883 ) | ( n18850 & n45239 ) | ( ~n25883 & n45239 ) ;
  assign n45241 = n28861 ^ n5507 ^ 1'b0 ;
  assign n45242 = n23906 | n45241 ;
  assign n45243 = n25707 & ~n45242 ;
  assign n45244 = n25127 ^ n8094 ^ n5639 ;
  assign n45245 = n36513 ^ n5659 ^ 1'b0 ;
  assign n45246 = n23906 | n45245 ;
  assign n45249 = n14481 ^ n13953 ^ 1'b0 ;
  assign n45250 = n1966 | n45249 ;
  assign n45251 = n13743 | n45250 ;
  assign n45247 = n15342 | n23898 ;
  assign n45248 = n9965 & ~n45247 ;
  assign n45252 = n45251 ^ n45248 ^ 1'b0 ;
  assign n45253 = n45252 ^ n34518 ^ 1'b0 ;
  assign n45254 = n5039 & ~n7115 ;
  assign n45255 = n40987 ^ n10442 ^ 1'b0 ;
  assign n45256 = n6777 & n28024 ;
  assign n45257 = n45256 ^ n13708 ^ n3298 ;
  assign n45259 = n2939 ^ n993 ^ 1'b0 ;
  assign n45260 = ~n22012 & n45259 ;
  assign n45258 = ( n2179 & ~n12219 ) | ( n2179 & n26843 ) | ( ~n12219 & n26843 ) ;
  assign n45261 = n45260 ^ n45258 ^ n38285 ;
  assign n45262 = n45261 ^ n43303 ^ n1639 ;
  assign n45263 = ( n14056 & n18462 ) | ( n14056 & ~n38380 ) | ( n18462 & ~n38380 ) ;
  assign n45264 = ( n8460 & n27453 ) | ( n8460 & n45263 ) | ( n27453 & n45263 ) ;
  assign n45265 = ( ~n35274 & n35523 ) | ( ~n35274 & n45264 ) | ( n35523 & n45264 ) ;
  assign n45266 = n8660 & ~n15497 ;
  assign n45267 = n6136 & n37111 ;
  assign n45268 = n575 | n27565 ;
  assign n45269 = n41621 ^ n34579 ^ 1'b0 ;
  assign n45270 = ( n1359 & n27766 ) | ( n1359 & n45269 ) | ( n27766 & n45269 ) ;
  assign n45271 = n45270 ^ n23314 ^ n3804 ;
  assign n45272 = n5433 | n44994 ;
  assign n45273 = n14844 ^ n8034 ^ n3366 ;
  assign n45274 = n14055 & n17726 ;
  assign n45275 = n45274 ^ n22081 ^ 1'b0 ;
  assign n45276 = n3257 & ~n16244 ;
  assign n45277 = n12832 & ~n29065 ;
  assign n45278 = n11074 ^ n7729 ^ n4286 ;
  assign n45279 = n45278 ^ n19419 ^ n12454 ;
  assign n45280 = n45279 ^ n10017 ^ 1'b0 ;
  assign n45281 = ~n25286 & n45280 ;
  assign n45282 = ~n2494 & n27557 ;
  assign n45283 = n45282 ^ n17585 ^ 1'b0 ;
  assign n45284 = n4690 | n10869 ;
  assign n45285 = n45284 ^ n29473 ^ 1'b0 ;
  assign n45286 = ( n29340 & ~n45283 ) | ( n29340 & n45285 ) | ( ~n45283 & n45285 ) ;
  assign n45287 = n21537 ^ n16266 ^ n10099 ;
  assign n45289 = n5868 & n12289 ;
  assign n45290 = ~n25025 & n45289 ;
  assign n45288 = ( ~n5539 & n38593 ) | ( ~n5539 & n40885 ) | ( n38593 & n40885 ) ;
  assign n45291 = n45290 ^ n45288 ^ n9089 ;
  assign n45292 = ( n34900 & n45287 ) | ( n34900 & n45291 ) | ( n45287 & n45291 ) ;
  assign n45293 = n2836 & n4208 ;
  assign n45294 = n45293 ^ n13780 ^ 1'b0 ;
  assign n45295 = ( n27348 & n40778 ) | ( n27348 & n45294 ) | ( n40778 & n45294 ) ;
  assign n45296 = ( n6115 & n11494 ) | ( n6115 & n45295 ) | ( n11494 & n45295 ) ;
  assign n45297 = n24524 ^ n3557 ^ x35 ;
  assign n45298 = n45297 ^ n21844 ^ n8559 ;
  assign n45299 = n18485 & ~n31943 ;
  assign n45300 = n31612 ^ n18522 ^ 1'b0 ;
  assign n45301 = n9921 & n13393 ;
  assign n45302 = ~n3874 & n45301 ;
  assign n45303 = n8503 & ~n13264 ;
  assign n45304 = n1283 & n45303 ;
  assign n45305 = n45304 ^ n22382 ^ 1'b0 ;
  assign n45306 = n19218 & n45305 ;
  assign n45307 = ( n23050 & n33776 ) | ( n23050 & ~n42301 ) | ( n33776 & ~n42301 ) ;
  assign n45308 = n6258 & ~n26070 ;
  assign n45309 = ( n4150 & n14558 ) | ( n4150 & n18356 ) | ( n14558 & n18356 ) ;
  assign n45310 = n45309 ^ n13186 ^ 1'b0 ;
  assign n45311 = n16908 | n45310 ;
  assign n45312 = n9914 & ~n40683 ;
  assign n45313 = n28722 & n45312 ;
  assign n45314 = n4513 & n24582 ;
  assign n45315 = n41769 & ~n42568 ;
  assign n45316 = ~n13288 & n45315 ;
  assign n45317 = n13831 | n28328 ;
  assign n45318 = n45317 ^ n322 ^ 1'b0 ;
  assign n45319 = n45318 ^ n35218 ^ n18789 ;
  assign n45320 = ( n23243 & ~n26983 ) | ( n23243 & n31771 ) | ( ~n26983 & n31771 ) ;
  assign n45321 = ( x209 & n21185 ) | ( x209 & ~n21660 ) | ( n21185 & ~n21660 ) ;
  assign n45322 = n24312 ^ n14438 ^ n3637 ;
  assign n45323 = n45322 ^ n32503 ^ n26592 ;
  assign n45324 = n33218 ^ n28359 ^ 1'b0 ;
  assign n45325 = n14735 & n45324 ;
  assign n45326 = n45325 ^ n19606 ^ 1'b0 ;
  assign n45327 = ( ~n8563 & n11261 ) | ( ~n8563 & n19193 ) | ( n11261 & n19193 ) ;
  assign n45328 = n8117 ^ n7215 ^ n6737 ;
  assign n45329 = n39002 & ~n45328 ;
  assign n45330 = ~n6395 & n45329 ;
  assign n45331 = n3958 ^ n336 ^ 1'b0 ;
  assign n45332 = ~n8995 & n16049 ;
  assign n45333 = n18729 & n27249 ;
  assign n45334 = n23998 & ~n25765 ;
  assign n45335 = n45334 ^ n24893 ^ 1'b0 ;
  assign n45336 = ( n3279 & n18417 ) | ( n3279 & n42607 ) | ( n18417 & n42607 ) ;
  assign n45337 = ( n649 & n1125 ) | ( n649 & ~n34064 ) | ( n1125 & ~n34064 ) ;
  assign n45338 = n45337 ^ n24686 ^ n11434 ;
  assign n45339 = n22286 ^ n14832 ^ 1'b0 ;
  assign n45340 = n18021 | n45339 ;
  assign n45341 = ( ~n24690 & n40401 ) | ( ~n24690 & n45340 ) | ( n40401 & n45340 ) ;
  assign n45342 = n16390 | n17047 ;
  assign n45343 = n23024 | n31658 ;
  assign n45344 = n22451 | n45343 ;
  assign n45345 = ~n5610 & n42436 ;
  assign n45346 = n45345 ^ n18356 ^ 1'b0 ;
  assign n45347 = n45346 ^ n8461 ^ 1'b0 ;
  assign n45350 = n31619 ^ n10121 ^ n7659 ;
  assign n45348 = ( n8712 & ~n27572 ) | ( n8712 & n32462 ) | ( ~n27572 & n32462 ) ;
  assign n45349 = n10974 & ~n45348 ;
  assign n45351 = n45350 ^ n45349 ^ 1'b0 ;
  assign n45352 = ( n1468 & ~n2701 ) | ( n1468 & n45222 ) | ( ~n2701 & n45222 ) ;
  assign n45353 = n8413 ^ n749 ^ 1'b0 ;
  assign n45354 = n1358 & n45353 ;
  assign n45355 = ~n32108 & n45354 ;
  assign n45356 = ~n3369 & n25006 ;
  assign n45357 = n45356 ^ n27534 ^ n25151 ;
  assign n45358 = ~n45355 & n45357 ;
  assign n45359 = n15512 & n36412 ;
  assign n45360 = n10872 & n25302 ;
  assign n45361 = n45360 ^ n1361 ^ 1'b0 ;
  assign n45362 = ( n22259 & ~n27703 ) | ( n22259 & n40790 ) | ( ~n27703 & n40790 ) ;
  assign n45363 = ( ~n45359 & n45361 ) | ( ~n45359 & n45362 ) | ( n45361 & n45362 ) ;
  assign n45364 = n38160 ^ n27823 ^ n12746 ;
  assign n45365 = ~n10410 & n34276 ;
  assign n45366 = n2065 & ~n10095 ;
  assign n45367 = n8307 & n45366 ;
  assign n45368 = n45367 ^ n43264 ^ 1'b0 ;
  assign n45369 = ~n20625 & n45368 ;
  assign n45370 = n35503 ^ n34774 ^ 1'b0 ;
  assign n45371 = n6649 | n45370 ;
  assign n45372 = n26191 | n45371 ;
  assign n45373 = n26379 ^ n9892 ^ 1'b0 ;
  assign n45374 = n45373 ^ n22917 ^ 1'b0 ;
  assign n45375 = n8962 & n45374 ;
  assign n45376 = n36371 ^ n1658 ^ 1'b0 ;
  assign n45377 = n30249 & ~n45376 ;
  assign n45378 = n27372 ^ n10593 ^ n1826 ;
  assign n45383 = ( n9203 & n11899 ) | ( n9203 & n13616 ) | ( n11899 & n13616 ) ;
  assign n45381 = n1112 & n2251 ;
  assign n45382 = n45381 ^ n7614 ^ 1'b0 ;
  assign n45379 = ( n14872 & n21209 ) | ( n14872 & ~n24451 ) | ( n21209 & ~n24451 ) ;
  assign n45380 = n45379 ^ n31919 ^ 1'b0 ;
  assign n45384 = n45383 ^ n45382 ^ n45380 ;
  assign n45385 = n32948 ^ n23460 ^ n18253 ;
  assign n45386 = n10041 | n14703 ;
  assign n45387 = n45386 ^ n35242 ^ n3239 ;
  assign n45391 = ( n4819 & n11264 ) | ( n4819 & ~n21561 ) | ( n11264 & ~n21561 ) ;
  assign n45388 = n21502 ^ n5043 ^ 1'b0 ;
  assign n45389 = n45388 ^ n19783 ^ 1'b0 ;
  assign n45390 = n5980 | n45389 ;
  assign n45392 = n45391 ^ n45390 ^ 1'b0 ;
  assign n45393 = n25540 & n26522 ;
  assign n45394 = n45393 ^ n43132 ^ 1'b0 ;
  assign n45395 = n23234 ^ n3319 ^ n915 ;
  assign n45396 = n1088 & n4852 ;
  assign n45397 = n7099 & n45396 ;
  assign n45398 = ( n12242 & ~n43874 ) | ( n12242 & n45397 ) | ( ~n43874 & n45397 ) ;
  assign n45399 = ~n9532 & n15194 ;
  assign n45400 = n19255 ^ n5440 ^ n4832 ;
  assign n45401 = n36435 & ~n45400 ;
  assign n45402 = ( n45398 & n45399 ) | ( n45398 & ~n45401 ) | ( n45399 & ~n45401 ) ;
  assign n45403 = n37865 ^ n28173 ^ n25047 ;
  assign n45404 = n45403 ^ n36298 ^ n4570 ;
  assign n45405 = n8792 ^ n367 ^ 1'b0 ;
  assign n45406 = n18836 ^ n5009 ^ 1'b0 ;
  assign n45407 = n40640 & ~n45406 ;
  assign n45408 = n34726 ^ n19373 ^ n4388 ;
  assign n45409 = n31992 & ~n45408 ;
  assign n45410 = n45409 ^ n39572 ^ n20128 ;
  assign n45411 = ~n18520 & n29551 ;
  assign n45412 = ~n45410 & n45411 ;
  assign n45413 = n13313 & ~n24907 ;
  assign n45414 = ( n13850 & ~n44707 ) | ( n13850 & n45413 ) | ( ~n44707 & n45413 ) ;
  assign n45415 = n13330 | n45414 ;
  assign n45416 = n2744 & n3289 ;
  assign n45417 = n45416 ^ n26173 ^ 1'b0 ;
  assign n45418 = n38100 & n38775 ;
  assign n45421 = n15113 ^ n13094 ^ 1'b0 ;
  assign n45419 = ( ~n9792 & n18402 ) | ( ~n9792 & n44406 ) | ( n18402 & n44406 ) ;
  assign n45420 = n10740 | n45419 ;
  assign n45422 = n45421 ^ n45420 ^ n20862 ;
  assign n45423 = n25006 ^ n9120 ^ 1'b0 ;
  assign n45424 = n45423 ^ n40686 ^ n30359 ;
  assign n45425 = n18973 ^ n16568 ^ 1'b0 ;
  assign n45426 = n28624 & ~n44803 ;
  assign n45427 = ~n23483 & n45426 ;
  assign n45428 = n11819 ^ n851 ^ 1'b0 ;
  assign n45429 = ~n12500 & n45428 ;
  assign n45430 = n25695 & ~n45429 ;
  assign n45431 = n11075 | n25141 ;
  assign n45432 = n45431 ^ n23040 ^ 1'b0 ;
  assign n45433 = n38481 ^ n33866 ^ 1'b0 ;
  assign n45434 = n1997 | n21594 ;
  assign n45435 = n2939 & ~n45434 ;
  assign n45436 = n15174 & ~n45435 ;
  assign n45437 = ( x159 & n2229 ) | ( x159 & n12103 ) | ( n2229 & n12103 ) ;
  assign n45438 = ( n3892 & ~n31836 ) | ( n3892 & n45437 ) | ( ~n31836 & n45437 ) ;
  assign n45439 = ( ~x1 & n24433 ) | ( ~x1 & n43377 ) | ( n24433 & n43377 ) ;
  assign n45440 = n35261 ^ n25013 ^ 1'b0 ;
  assign n45441 = n45388 ^ n24620 ^ n23501 ;
  assign n45442 = n33609 | n45441 ;
  assign n45445 = n381 | n21551 ;
  assign n45446 = ( n1281 & n22338 ) | ( n1281 & ~n45445 ) | ( n22338 & ~n45445 ) ;
  assign n45444 = n10988 & ~n19446 ;
  assign n45447 = n45446 ^ n45444 ^ 1'b0 ;
  assign n45443 = n13662 | n21589 ;
  assign n45448 = n45447 ^ n45443 ^ 1'b0 ;
  assign n45449 = ~n8673 & n34446 ;
  assign n45450 = ( n9691 & n14095 ) | ( n9691 & ~n34501 ) | ( n14095 & ~n34501 ) ;
  assign n45451 = n10187 & ~n16146 ;
  assign n45452 = n45451 ^ n22353 ^ 1'b0 ;
  assign n45453 = n8320 & ~n16186 ;
  assign n45454 = ~n33246 & n45453 ;
  assign n45455 = ( n45450 & n45452 ) | ( n45450 & ~n45454 ) | ( n45452 & ~n45454 ) ;
  assign n45456 = ( n17051 & n45449 ) | ( n17051 & n45455 ) | ( n45449 & n45455 ) ;
  assign n45457 = n33618 ^ n19571 ^ n18838 ;
  assign n45458 = ~n2474 & n5542 ;
  assign n45459 = ~n4734 & n45458 ;
  assign n45460 = ( ~n17224 & n33632 ) | ( ~n17224 & n45459 ) | ( n33632 & n45459 ) ;
  assign n45462 = n18631 ^ n13812 ^ 1'b0 ;
  assign n45461 = n5639 | n12188 ;
  assign n45463 = n45462 ^ n45461 ^ 1'b0 ;
  assign n45464 = ~n17711 & n34679 ;
  assign n45465 = n31905 ^ n29976 ^ 1'b0 ;
  assign n45466 = n8884 | n25639 ;
  assign n45467 = ( ~n19238 & n27540 ) | ( ~n19238 & n29288 ) | ( n27540 & n29288 ) ;
  assign n45468 = n18810 ^ n8263 ^ 1'b0 ;
  assign n45469 = n3699 & ~n4189 ;
  assign n45470 = ~n33088 & n45469 ;
  assign n45472 = n5983 ^ n1647 ^ 1'b0 ;
  assign n45471 = ~n21238 & n24985 ;
  assign n45473 = n45472 ^ n45471 ^ 1'b0 ;
  assign n45474 = n5702 & n44739 ;
  assign n45475 = ~n45473 & n45474 ;
  assign n45476 = ( n10116 & n13590 ) | ( n10116 & ~n19951 ) | ( n13590 & ~n19951 ) ;
  assign n45477 = ( ~n4444 & n8703 ) | ( ~n4444 & n21471 ) | ( n8703 & n21471 ) ;
  assign n45478 = ( n4711 & ~n9127 ) | ( n4711 & n45477 ) | ( ~n9127 & n45477 ) ;
  assign n45479 = n21393 | n32099 ;
  assign n45480 = n43075 ^ n42096 ^ 1'b0 ;
  assign n45481 = ( n6053 & n20884 ) | ( n6053 & ~n44434 ) | ( n20884 & ~n44434 ) ;
  assign n45482 = n45481 ^ n5953 ^ n1140 ;
  assign n45483 = n8657 & n32818 ;
  assign n45484 = n45483 ^ n4351 ^ 1'b0 ;
  assign n45486 = n2028 | n25489 ;
  assign n45485 = ( n9349 & ~n11443 ) | ( n9349 & n14665 ) | ( ~n11443 & n14665 ) ;
  assign n45487 = n45486 ^ n45485 ^ n27946 ;
  assign n45488 = n45487 ^ n10663 ^ x133 ;
  assign n45489 = n45488 ^ n29000 ^ 1'b0 ;
  assign n45490 = ( n4721 & n10743 ) | ( n4721 & n20905 ) | ( n10743 & n20905 ) ;
  assign n45491 = n45490 ^ n17931 ^ 1'b0 ;
  assign n45492 = ~n26916 & n45491 ;
  assign n45493 = n45492 ^ n11312 ^ n6132 ;
  assign n45494 = n6291 & ~n34207 ;
  assign n45495 = ~n21949 & n45494 ;
  assign n45496 = n45495 ^ n33205 ^ n10072 ;
  assign n45497 = ( n15315 & ~n29197 ) | ( n15315 & n29833 ) | ( ~n29197 & n29833 ) ;
  assign n45498 = ( n3383 & n20916 ) | ( n3383 & ~n45497 ) | ( n20916 & ~n45497 ) ;
  assign n45499 = n11216 & ~n14283 ;
  assign n45500 = n45499 ^ n14991 ^ 1'b0 ;
  assign n45501 = n37290 ^ n29171 ^ 1'b0 ;
  assign n45502 = ( ~n736 & n1846 ) | ( ~n736 & n25480 ) | ( n1846 & n25480 ) ;
  assign n45503 = n12083 & n45502 ;
  assign n45504 = ~n2466 & n45503 ;
  assign n45507 = ~n13976 & n21022 ;
  assign n45508 = n45507 ^ n10844 ^ n9715 ;
  assign n45505 = n9905 & ~n11118 ;
  assign n45506 = ~n1560 & n45505 ;
  assign n45509 = n45508 ^ n45506 ^ 1'b0 ;
  assign n45510 = ~n450 & n22317 ;
  assign n45511 = n45510 ^ n44450 ^ n27523 ;
  assign n45514 = n481 | n9612 ;
  assign n45512 = n5468 ^ n1132 ^ 1'b0 ;
  assign n45513 = n45512 ^ n4459 ^ n2457 ;
  assign n45515 = n45514 ^ n45513 ^ n40740 ;
  assign n45516 = ~n28693 & n29596 ;
  assign n45517 = ~n914 & n20749 ;
  assign n45518 = n45517 ^ n8593 ^ 1'b0 ;
  assign n45519 = ~n16648 & n24641 ;
  assign n45520 = n14268 | n18520 ;
  assign n45521 = n45520 ^ n16620 ^ 1'b0 ;
  assign n45522 = n6145 & n44096 ;
  assign n45523 = n21533 & n45522 ;
  assign n45524 = n26954 ^ n17272 ^ n4807 ;
  assign n45525 = ( n15499 & ~n21438 ) | ( n15499 & n22246 ) | ( ~n21438 & n22246 ) ;
  assign n45526 = n10903 | n45525 ;
  assign n45527 = ( n1422 & n6435 ) | ( n1422 & n16683 ) | ( n6435 & n16683 ) ;
  assign n45528 = n12038 ^ n4879 ^ 1'b0 ;
  assign n45529 = ( n9040 & n17010 ) | ( n9040 & n35813 ) | ( n17010 & n35813 ) ;
  assign n45530 = n45529 ^ n17438 ^ 1'b0 ;
  assign n45531 = ( n3312 & ~n8259 ) | ( n3312 & n17275 ) | ( ~n8259 & n17275 ) ;
  assign n45532 = n42662 & ~n45531 ;
  assign n45533 = n45532 ^ n541 ^ 1'b0 ;
  assign n45534 = n30994 ^ n23698 ^ 1'b0 ;
  assign n45535 = n13499 & n45534 ;
  assign n45536 = n12715 & n45535 ;
  assign n45537 = n16709 ^ n11216 ^ n2260 ;
  assign n45538 = n1758 & ~n38006 ;
  assign n45539 = ~n44774 & n45538 ;
  assign n45540 = n29933 ^ n28520 ^ 1'b0 ;
  assign n45541 = n33743 ^ n15979 ^ 1'b0 ;
  assign n45542 = n45541 ^ n26159 ^ n10559 ;
  assign n45543 = n45542 ^ n37233 ^ 1'b0 ;
  assign n45544 = ~n18414 & n27699 ;
  assign n45545 = n30224 ^ n1037 ^ 1'b0 ;
  assign n45546 = n45545 ^ n3667 ^ n3441 ;
  assign n45547 = ~n22456 & n45546 ;
  assign n45548 = ( n6991 & n17143 ) | ( n6991 & n45547 ) | ( n17143 & n45547 ) ;
  assign n45549 = n12876 ^ n7921 ^ 1'b0 ;
  assign n45550 = n22481 & ~n45549 ;
  assign n45551 = n12997 & ~n45550 ;
  assign n45553 = ( ~n8923 & n22037 ) | ( ~n8923 & n40260 ) | ( n22037 & n40260 ) ;
  assign n45554 = n45553 ^ n23046 ^ 1'b0 ;
  assign n45552 = n1363 | n15399 ;
  assign n45555 = n45554 ^ n45552 ^ 1'b0 ;
  assign n45556 = n25078 ^ n10817 ^ 1'b0 ;
  assign n45557 = n31654 ^ n4005 ^ 1'b0 ;
  assign n45558 = n45556 & ~n45557 ;
  assign n45559 = n39194 ^ n264 ^ 1'b0 ;
  assign n45560 = n10971 & ~n11930 ;
  assign n45561 = n45560 ^ n24609 ^ 1'b0 ;
  assign n45562 = n13575 ^ n5484 ^ 1'b0 ;
  assign n45563 = n45561 | n45562 ;
  assign n45564 = n45559 & ~n45563 ;
  assign n45565 = n26208 ^ n11129 ^ 1'b0 ;
  assign n45566 = ~n12807 & n15166 ;
  assign n45567 = n11251 & n45566 ;
  assign n45568 = n45567 ^ n32961 ^ n27669 ;
  assign n45569 = n31365 ^ n22382 ^ n8739 ;
  assign n45570 = n30309 ^ n4346 ^ 1'b0 ;
  assign n45571 = n28640 & ~n45570 ;
  assign n45572 = ~n5172 & n8740 ;
  assign n45574 = ( ~n3266 & n15758 ) | ( ~n3266 & n33183 ) | ( n15758 & n33183 ) ;
  assign n45573 = n10019 | n16178 ;
  assign n45575 = n45574 ^ n45573 ^ 1'b0 ;
  assign n45576 = n5238 | n33913 ;
  assign n45577 = ( ~n1294 & n14723 ) | ( ~n1294 & n35302 ) | ( n14723 & n35302 ) ;
  assign n45578 = ~n5885 & n7999 ;
  assign n45579 = n45577 & n45578 ;
  assign n45580 = n600 & ~n45579 ;
  assign n45581 = n9787 & ~n25673 ;
  assign n45582 = ( n21344 & n39125 ) | ( n21344 & ~n45581 ) | ( n39125 & ~n45581 ) ;
  assign n45583 = n17087 ^ n1522 ^ 1'b0 ;
  assign n45584 = n1854 & n45583 ;
  assign n45585 = n22669 & ~n24802 ;
  assign n45586 = n18818 ^ n16302 ^ 1'b0 ;
  assign n45587 = ~n45585 & n45586 ;
  assign n45588 = n28308 ^ n14598 ^ 1'b0 ;
  assign n45589 = n30702 | n45588 ;
  assign n45590 = ( n791 & n21468 ) | ( n791 & n28925 ) | ( n21468 & n28925 ) ;
  assign n45591 = n421 | n45590 ;
  assign n45592 = n45591 ^ n34828 ^ 1'b0 ;
  assign n45593 = n34414 ^ n33845 ^ 1'b0 ;
  assign n45594 = ~n45389 & n45593 ;
  assign n45595 = n45097 ^ n26095 ^ n861 ;
  assign n45596 = n38951 ^ n26674 ^ n13990 ;
  assign n45597 = n12467 ^ n3469 ^ x214 ;
  assign n45598 = n4547 ^ n3868 ^ 1'b0 ;
  assign n45599 = n45598 ^ n44676 ^ n44582 ;
  assign n45600 = n16047 | n16164 ;
  assign n45601 = n45600 ^ n33585 ^ 1'b0 ;
  assign n45602 = n13999 | n45601 ;
  assign n45603 = ( n11443 & ~n15118 ) | ( n11443 & n38420 ) | ( ~n15118 & n38420 ) ;
  assign n45604 = n26528 ^ n25718 ^ n25597 ;
  assign n45605 = n21248 & ~n45604 ;
  assign n45606 = n1438 & ~n10081 ;
  assign n45607 = n9976 ^ n9790 ^ 1'b0 ;
  assign n45608 = n22065 ^ n7697 ^ 1'b0 ;
  assign n45609 = n23991 ^ n19519 ^ 1'b0 ;
  assign n45610 = n16744 | n45609 ;
  assign n45611 = n32171 ^ n22738 ^ 1'b0 ;
  assign n45612 = n4922 & n7163 ;
  assign n45613 = ( ~n14141 & n45611 ) | ( ~n14141 & n45612 ) | ( n45611 & n45612 ) ;
  assign n45614 = n39736 ^ n16327 ^ n4346 ;
  assign n45615 = n36488 ^ n3523 ^ 1'b0 ;
  assign n45621 = n8170 ^ n6785 ^ 1'b0 ;
  assign n45622 = n45621 ^ n40863 ^ n6560 ;
  assign n45618 = n3301 & ~n27700 ;
  assign n45619 = n45618 ^ n23627 ^ 1'b0 ;
  assign n45616 = n12593 ^ n3621 ^ 1'b0 ;
  assign n45617 = n27382 & ~n45616 ;
  assign n45620 = n45619 ^ n45617 ^ n11519 ;
  assign n45623 = n45622 ^ n45620 ^ n25510 ;
  assign n45624 = n23583 ^ n22234 ^ n8972 ;
  assign n45625 = n4266 | n45624 ;
  assign n45626 = ~n3935 & n30719 ;
  assign n45627 = x189 & n11572 ;
  assign n45628 = n45627 ^ n39421 ^ 1'b0 ;
  assign n45629 = n36009 ^ n18341 ^ 1'b0 ;
  assign n45630 = ( n4361 & ~n6541 ) | ( n4361 & n19453 ) | ( ~n6541 & n19453 ) ;
  assign n45631 = n45630 ^ n18199 ^ n7126 ;
  assign n45632 = n15680 ^ n7791 ^ n3721 ;
  assign n45633 = n28375 ^ n9473 ^ 1'b0 ;
  assign n45634 = ~n1590 & n45633 ;
  assign n45635 = ( n17643 & n45632 ) | ( n17643 & n45634 ) | ( n45632 & n45634 ) ;
  assign n45636 = ( n10723 & ~n23331 ) | ( n10723 & n24979 ) | ( ~n23331 & n24979 ) ;
  assign n45637 = n21906 ^ n21846 ^ 1'b0 ;
  assign n45638 = n31373 ^ n14413 ^ 1'b0 ;
  assign n45639 = n11977 & ~n45638 ;
  assign n45640 = n16067 & ~n43048 ;
  assign n45641 = ~n1566 & n45640 ;
  assign n45642 = n36683 ^ n29240 ^ n24971 ;
  assign n45643 = n45642 ^ n1981 ^ 1'b0 ;
  assign n45644 = n1539 & n45643 ;
  assign n45645 = n44984 ^ n9601 ^ 1'b0 ;
  assign n45646 = ( n3156 & ~n3186 ) | ( n3156 & n4219 ) | ( ~n3186 & n4219 ) ;
  assign n45647 = n45646 ^ n16914 ^ n4390 ;
  assign n45648 = n45647 ^ n6173 ^ n5109 ;
  assign n45649 = n23703 ^ n14942 ^ n1538 ;
  assign n45650 = n3324 & ~n41046 ;
  assign n45651 = n39342 & n45650 ;
  assign n45652 = n45649 & n45651 ;
  assign n45653 = n7217 ^ x34 ^ 1'b0 ;
  assign n45654 = n34842 ^ n28716 ^ n12255 ;
  assign n45655 = n45654 ^ n43106 ^ 1'b0 ;
  assign n45656 = n20855 ^ n14534 ^ n2628 ;
  assign n45657 = n45656 ^ n13277 ^ 1'b0 ;
  assign n45658 = n15224 & ~n45657 ;
  assign n45659 = ~n13852 & n31091 ;
  assign n45660 = n45659 ^ n35439 ^ 1'b0 ;
  assign n45661 = ( n2132 & ~n7493 ) | ( n2132 & n19813 ) | ( ~n7493 & n19813 ) ;
  assign n45662 = n32777 | n45661 ;
  assign n45663 = n45662 ^ n10492 ^ 1'b0 ;
  assign n45664 = n9723 & ~n34929 ;
  assign n45665 = n45664 ^ n14404 ^ 1'b0 ;
  assign n45666 = n16551 ^ n9824 ^ 1'b0 ;
  assign n45669 = n17981 ^ n8251 ^ 1'b0 ;
  assign n45670 = n45669 ^ n25169 ^ n1559 ;
  assign n45667 = n34608 | n45279 ;
  assign n45668 = n4546 | n45667 ;
  assign n45671 = n45670 ^ n45668 ^ 1'b0 ;
  assign n45672 = n37188 & n45671 ;
  assign n45673 = ~n14698 & n44355 ;
  assign n45674 = ( n471 & n4739 ) | ( n471 & n45673 ) | ( n4739 & n45673 ) ;
  assign n45675 = n13758 ^ n5872 ^ 1'b0 ;
  assign n45676 = n45309 & ~n45675 ;
  assign n45677 = ~n18929 & n29571 ;
  assign n45678 = ~n37424 & n45677 ;
  assign n45679 = n10557 ^ n4854 ^ 1'b0 ;
  assign n45680 = n15348 & n18100 ;
  assign n45681 = n45679 & n45680 ;
  assign n45682 = n20368 ^ n18326 ^ n12023 ;
  assign n45683 = n16116 ^ n12250 ^ 1'b0 ;
  assign n45684 = n678 & ~n11013 ;
  assign n45685 = ~n45683 & n45684 ;
  assign n45686 = n45682 & ~n45685 ;
  assign n45687 = n12267 & ~n20534 ;
  assign n45688 = ~n29296 & n45687 ;
  assign n45689 = n4142 & n42623 ;
  assign n45690 = n24995 ^ n19063 ^ 1'b0 ;
  assign n45691 = n28136 | n45690 ;
  assign n45692 = n45691 ^ n3966 ^ 1'b0 ;
  assign n45693 = n45692 ^ n21406 ^ 1'b0 ;
  assign n45694 = n1690 | n45693 ;
  assign n45695 = ~n4467 & n35724 ;
  assign n45696 = n45695 ^ x227 ^ 1'b0 ;
  assign n45697 = ( n11841 & ~n24052 ) | ( n11841 & n35794 ) | ( ~n24052 & n35794 ) ;
  assign n45698 = n3251 | n15128 ;
  assign n45699 = n45697 | n45698 ;
  assign n45700 = ( n7526 & ~n45696 ) | ( n7526 & n45699 ) | ( ~n45696 & n45699 ) ;
  assign n45701 = ~n452 & n23814 ;
  assign n45704 = n5068 & n6441 ;
  assign n45705 = n45704 ^ n4356 ^ 1'b0 ;
  assign n45706 = n45705 ^ n26455 ^ n9780 ;
  assign n45702 = n4852 & n42952 ;
  assign n45703 = n14372 & n45702 ;
  assign n45707 = n45706 ^ n45703 ^ n24370 ;
  assign n45708 = ~n4446 & n28963 ;
  assign n45709 = n6290 | n45708 ;
  assign n45710 = n39440 & ~n45709 ;
  assign n45711 = n25129 ^ n20132 ^ 1'b0 ;
  assign n45712 = ~n1080 & n45711 ;
  assign n45713 = ( ~n13264 & n20826 ) | ( ~n13264 & n26422 ) | ( n20826 & n26422 ) ;
  assign n45714 = n39982 & ~n45713 ;
  assign n45715 = n45714 ^ n10986 ^ 1'b0 ;
  assign n45716 = n44722 ^ n43485 ^ 1'b0 ;
  assign n45717 = n7745 | n33454 ;
  assign n45718 = n45717 ^ n32404 ^ 1'b0 ;
  assign n45719 = n4345 ^ n1885 ^ n1773 ;
  assign n45720 = n45719 ^ n34805 ^ 1'b0 ;
  assign n45721 = n19699 & n45720 ;
  assign n45722 = ( n14164 & n17587 ) | ( n14164 & ~n19753 ) | ( n17587 & ~n19753 ) ;
  assign n45723 = n5494 & ~n45379 ;
  assign n45724 = ~n17960 & n45723 ;
  assign n45725 = n42185 ^ n18738 ^ n5715 ;
  assign n45726 = n22210 ^ n2457 ^ 1'b0 ;
  assign n45727 = ( n34944 & ~n45725 ) | ( n34944 & n45726 ) | ( ~n45725 & n45726 ) ;
  assign n45728 = n45727 ^ n2151 ^ x109 ;
  assign n45729 = ( n3972 & ~n45724 ) | ( n3972 & n45728 ) | ( ~n45724 & n45728 ) ;
  assign n45730 = n25259 ^ n9410 ^ n1199 ;
  assign n45731 = n18054 ^ n6657 ^ n2503 ;
  assign n45732 = n13273 & n23296 ;
  assign n45733 = n45732 ^ n14782 ^ 1'b0 ;
  assign n45734 = ~n8244 & n13768 ;
  assign n45735 = n24002 ^ n16111 ^ 1'b0 ;
  assign n45736 = n40194 & ~n45735 ;
  assign n45737 = n39984 ^ n8328 ^ 1'b0 ;
  assign n45738 = n20161 & n45737 ;
  assign n45739 = n45738 ^ n11778 ^ 1'b0 ;
  assign n45742 = n5910 | n28894 ;
  assign n45743 = n45742 ^ n1910 ^ 1'b0 ;
  assign n45744 = ~n42059 & n45743 ;
  assign n45745 = ~n10468 & n45744 ;
  assign n45740 = n14380 & ~n15737 ;
  assign n45741 = n25488 & n45740 ;
  assign n45746 = n45745 ^ n45741 ^ 1'b0 ;
  assign n45747 = n20798 ^ n20727 ^ 1'b0 ;
  assign n45748 = ( n30157 & n31304 ) | ( n30157 & n45747 ) | ( n31304 & n45747 ) ;
  assign n45749 = ~n17008 & n17747 ;
  assign n45750 = ( ~n12682 & n13419 ) | ( ~n12682 & n45749 ) | ( n13419 & n45749 ) ;
  assign n45751 = n32165 & n35307 ;
  assign n45752 = n30538 ^ n11081 ^ 1'b0 ;
  assign n45753 = n8805 | n38518 ;
  assign n45754 = n38845 ^ n29940 ^ 1'b0 ;
  assign n45755 = ( n5288 & n7113 ) | ( n5288 & n10426 ) | ( n7113 & n10426 ) ;
  assign n45756 = n19634 ^ n14313 ^ n8508 ;
  assign n45757 = ( n14995 & n45755 ) | ( n14995 & ~n45756 ) | ( n45755 & ~n45756 ) ;
  assign n45758 = n45757 ^ n37499 ^ 1'b0 ;
  assign n45759 = ~n45754 & n45758 ;
  assign n45760 = ~n2468 & n7201 ;
  assign n45761 = n6680 & n45760 ;
  assign n45762 = ( n10474 & n11765 ) | ( n10474 & n45761 ) | ( n11765 & n45761 ) ;
  assign n45763 = n5233 ^ x180 ^ 1'b0 ;
  assign n45764 = n5293 ^ n5048 ^ n2399 ;
  assign n45765 = n44491 ^ n26305 ^ 1'b0 ;
  assign n45766 = n45764 & n45765 ;
  assign n45767 = n45766 ^ n9567 ^ n2035 ;
  assign n45768 = ( n8243 & n16199 ) | ( n8243 & ~n26289 ) | ( n16199 & ~n26289 ) ;
  assign n45769 = ~n2719 & n15511 ;
  assign n45770 = n44648 ^ n31938 ^ 1'b0 ;
  assign n45771 = n15605 & n31256 ;
  assign n45772 = ~n4378 & n5627 ;
  assign n45773 = n45772 ^ n42020 ^ 1'b0 ;
  assign n45774 = n4847 | n45773 ;
  assign n45775 = n3178 | n45774 ;
  assign n45776 = n12736 & ~n45775 ;
  assign n45777 = n45776 ^ n14233 ^ 1'b0 ;
  assign n45778 = ~n10599 & n45777 ;
  assign n45779 = n1749 & n5087 ;
  assign n45780 = n45779 ^ n13539 ^ 1'b0 ;
  assign n45784 = n4439 | n27100 ;
  assign n45785 = n45784 ^ n3202 ^ 1'b0 ;
  assign n45781 = x200 & n1761 ;
  assign n45782 = n45781 ^ n40591 ^ 1'b0 ;
  assign n45783 = n5729 & n45782 ;
  assign n45786 = n45785 ^ n45783 ^ n36211 ;
  assign n45787 = n5658 ^ n1192 ^ 1'b0 ;
  assign n45788 = n33647 | n45787 ;
  assign n45789 = n29634 | n45788 ;
  assign n45790 = n45789 ^ n7083 ^ 1'b0 ;
  assign n45791 = n28902 ^ n18944 ^ 1'b0 ;
  assign n45792 = ( n728 & ~n6823 ) | ( n728 & n22853 ) | ( ~n6823 & n22853 ) ;
  assign n45793 = ( ~n996 & n2919 ) | ( ~n996 & n6241 ) | ( n2919 & n6241 ) ;
  assign n45794 = n45793 ^ n18320 ^ 1'b0 ;
  assign n45795 = n45792 & ~n45794 ;
  assign n45796 = ( n3330 & n45545 ) | ( n3330 & n45795 ) | ( n45545 & n45795 ) ;
  assign n45797 = n45796 ^ n25174 ^ 1'b0 ;
  assign n45798 = n45783 ^ n26219 ^ n16043 ;
  assign n45799 = n26115 ^ n15571 ^ 1'b0 ;
  assign n45800 = n25113 & n45799 ;
  assign n45801 = n5324 ^ n3177 ^ 1'b0 ;
  assign n45802 = n45800 & ~n45801 ;
  assign n45803 = n45802 ^ n31588 ^ 1'b0 ;
  assign n45804 = ~n3468 & n34041 ;
  assign n45805 = ~n3730 & n45804 ;
  assign n45806 = n39708 ^ n7051 ^ 1'b0 ;
  assign n45807 = n39119 & n45806 ;
  assign n45808 = n17495 | n36827 ;
  assign n45809 = n30001 ^ n18744 ^ 1'b0 ;
  assign n45810 = n998 & ~n20440 ;
  assign n45811 = n45809 & n45810 ;
  assign n45812 = ( n7794 & ~n27868 ) | ( n7794 & n45811 ) | ( ~n27868 & n45811 ) ;
  assign n45813 = n17349 & n37081 ;
  assign n45814 = ~n18756 & n36662 ;
  assign n45815 = n45814 ^ n24328 ^ 1'b0 ;
  assign n45816 = n6683 | n20988 ;
  assign n45818 = n36686 ^ n20082 ^ n9411 ;
  assign n45817 = n4527 | n32705 ;
  assign n45819 = n45818 ^ n45817 ^ 1'b0 ;
  assign n45820 = n6675 | n29517 ;
  assign n45821 = n16115 ^ n3173 ^ 1'b0 ;
  assign n45822 = n7139 | n45821 ;
  assign n45823 = ( ~n742 & n6973 ) | ( ~n742 & n22058 ) | ( n6973 & n22058 ) ;
  assign n45824 = ( n7216 & ~n25476 ) | ( n7216 & n38461 ) | ( ~n25476 & n38461 ) ;
  assign n45827 = ~n1737 & n25079 ;
  assign n45828 = n7025 & n45827 ;
  assign n45825 = n2233 & n7955 ;
  assign n45826 = n45825 ^ n4352 ^ 1'b0 ;
  assign n45829 = n45828 ^ n45826 ^ n30226 ;
  assign n45830 = ( n12465 & n45824 ) | ( n12465 & n45829 ) | ( n45824 & n45829 ) ;
  assign n45831 = n19038 ^ n4907 ^ 1'b0 ;
  assign n45832 = ~n33749 & n45831 ;
  assign n45833 = n45832 ^ n45728 ^ n23628 ;
  assign n45834 = n7758 & n38647 ;
  assign n45835 = n45834 ^ n33628 ^ 1'b0 ;
  assign n45836 = n27391 ^ n4535 ^ 1'b0 ;
  assign n45837 = n45836 ^ n43185 ^ n42093 ;
  assign n45838 = n17858 | n45837 ;
  assign n45839 = n24261 | n30173 ;
  assign n45840 = n45839 ^ n20155 ^ 1'b0 ;
  assign n45841 = n45840 ^ n30049 ^ 1'b0 ;
  assign n45842 = n33210 ^ n26231 ^ 1'b0 ;
  assign n45843 = n18168 & n39485 ;
  assign n45844 = n45843 ^ n4766 ^ 1'b0 ;
  assign n45845 = ~n3535 & n24677 ;
  assign n45846 = ~n45844 & n45845 ;
  assign n45847 = n26940 ^ n4872 ^ 1'b0 ;
  assign n45848 = n1298 & ~n45847 ;
  assign n45849 = ( n37789 & n40389 ) | ( n37789 & n45848 ) | ( n40389 & n45848 ) ;
  assign n45850 = n756 & n45849 ;
  assign n45851 = ~n14847 & n45850 ;
  assign n45853 = n2789 & ~n37904 ;
  assign n45854 = n45853 ^ n6472 ^ 1'b0 ;
  assign n45855 = ( ~n2091 & n40216 ) | ( ~n2091 & n45854 ) | ( n40216 & n45854 ) ;
  assign n45852 = ( n3468 & n9030 ) | ( n3468 & ~n24432 ) | ( n9030 & ~n24432 ) ;
  assign n45856 = n45855 ^ n45852 ^ 1'b0 ;
  assign n45857 = ~n45851 & n45856 ;
  assign n45858 = ~n10216 & n42205 ;
  assign n45859 = n2109 & n45858 ;
  assign n45860 = n12227 ^ n8833 ^ 1'b0 ;
  assign n45861 = ~n20640 & n45860 ;
  assign n45862 = n45861 ^ n31053 ^ 1'b0 ;
  assign n45863 = n34971 ^ n30719 ^ n27186 ;
  assign n45864 = ~n3846 & n25635 ;
  assign n45865 = n2840 | n14013 ;
  assign n45866 = n45865 ^ n17881 ^ 1'b0 ;
  assign n45867 = ( n836 & n20355 ) | ( n836 & n45866 ) | ( n20355 & n45866 ) ;
  assign n45868 = ( ~n27908 & n40087 ) | ( ~n27908 & n45867 ) | ( n40087 & n45867 ) ;
  assign n45869 = n16008 ^ n1040 ^ 1'b0 ;
  assign n45870 = n10997 & ~n45869 ;
  assign n45871 = n8365 & n12000 ;
  assign n45872 = n45871 ^ n4124 ^ 1'b0 ;
  assign n45873 = n44576 & ~n45872 ;
  assign n45874 = n45873 ^ n29306 ^ 1'b0 ;
  assign n45875 = n17590 | n23700 ;
  assign n45876 = n45875 ^ n24619 ^ 1'b0 ;
  assign n45877 = n35643 ^ n6103 ^ 1'b0 ;
  assign n45878 = n18332 | n45877 ;
  assign n45879 = n33544 | n45878 ;
  assign n45880 = n45879 ^ n25576 ^ 1'b0 ;
  assign n45881 = n34359 & ~n45880 ;
  assign n45882 = n21849 ^ n19758 ^ 1'b0 ;
  assign n45883 = n1866 & ~n45882 ;
  assign n45884 = n32661 & ~n45883 ;
  assign n45885 = ~n4949 & n7537 ;
  assign n45886 = n11447 ^ n2351 ^ n1400 ;
  assign n45887 = ( n6331 & n12207 ) | ( n6331 & ~n35931 ) | ( n12207 & ~n35931 ) ;
  assign n45888 = n3725 | n30397 ;
  assign n45889 = n45887 | n45888 ;
  assign n45890 = ~n45886 & n45889 ;
  assign n45891 = n2710 & ~n15288 ;
  assign n45892 = n45891 ^ n2989 ^ 1'b0 ;
  assign n45894 = n19373 ^ n7198 ^ 1'b0 ;
  assign n45895 = n22781 & n33859 ;
  assign n45896 = n45895 ^ n21360 ^ 1'b0 ;
  assign n45897 = n45896 ^ n9002 ^ 1'b0 ;
  assign n45898 = n45894 & ~n45897 ;
  assign n45893 = n19923 | n23106 ;
  assign n45899 = n45898 ^ n45893 ^ 1'b0 ;
  assign n45900 = n11136 & n25666 ;
  assign n45901 = n19281 ^ n17340 ^ 1'b0 ;
  assign n45902 = n45900 & ~n45901 ;
  assign n45903 = n37422 ^ n26652 ^ 1'b0 ;
  assign n45904 = n12351 & n45903 ;
  assign n45905 = ( n23592 & ~n25985 ) | ( n23592 & n44506 ) | ( ~n25985 & n44506 ) ;
  assign n45906 = n45505 ^ n23515 ^ n17123 ;
  assign n45907 = n4364 | n11352 ;
  assign n45908 = n9943 | n45907 ;
  assign n45909 = n45908 ^ n43841 ^ n20280 ;
  assign n45910 = n45909 ^ n14336 ^ n4954 ;
  assign n45911 = ~n13815 & n34502 ;
  assign n45912 = ( ~n15850 & n17419 ) | ( ~n15850 & n45911 ) | ( n17419 & n45911 ) ;
  assign n45913 = ( n11811 & n25195 ) | ( n11811 & ~n40598 ) | ( n25195 & ~n40598 ) ;
  assign n45914 = n45913 ^ n16034 ^ n2619 ;
  assign n45917 = ( ~n2583 & n4547 ) | ( ~n2583 & n26848 ) | ( n4547 & n26848 ) ;
  assign n45915 = n20468 ^ n8517 ^ 1'b0 ;
  assign n45916 = n2282 & ~n45915 ;
  assign n45918 = n45917 ^ n45916 ^ 1'b0 ;
  assign n45919 = n30271 & n35560 ;
  assign n45920 = n3892 & n45919 ;
  assign n45921 = n15063 ^ n9643 ^ 1'b0 ;
  assign n45922 = n25167 ^ n2637 ^ n536 ;
  assign n45923 = n1118 | n45922 ;
  assign n45924 = n45923 ^ n23090 ^ 1'b0 ;
  assign n45925 = n45921 & ~n45924 ;
  assign n45927 = n37371 & n41142 ;
  assign n45928 = n1331 & n45927 ;
  assign n45926 = n1638 & n5035 ;
  assign n45929 = n45928 ^ n45926 ^ 1'b0 ;
  assign n45930 = ~n6789 & n21536 ;
  assign n45931 = n28603 ^ n16779 ^ 1'b0 ;
  assign n45932 = n7539 | n45931 ;
  assign n45933 = n4471 & n45932 ;
  assign n45934 = n11347 ^ n3294 ^ 1'b0 ;
  assign n45935 = n4769 & n45934 ;
  assign n45936 = n45935 ^ n31506 ^ n2718 ;
  assign n45937 = n9287 & n20637 ;
  assign n45939 = ~x154 & n8064 ;
  assign n45940 = n45939 ^ n12739 ^ 1'b0 ;
  assign n45938 = n17962 ^ n1597 ^ 1'b0 ;
  assign n45941 = n45940 ^ n45938 ^ n1719 ;
  assign n45942 = n29241 ^ n28979 ^ 1'b0 ;
  assign n45943 = n8704 | n45942 ;
  assign n45944 = n16371 | n45943 ;
  assign n45945 = n7499 ^ n608 ^ 1'b0 ;
  assign n45946 = n20359 | n45945 ;
  assign n45947 = n3297 ^ n2877 ^ 1'b0 ;
  assign n45948 = ~n19317 & n45947 ;
  assign n45949 = n45948 ^ n8999 ^ 1'b0 ;
  assign n45950 = n45949 ^ n27491 ^ n14863 ;
  assign n45951 = n7129 & n45950 ;
  assign n45952 = n45951 ^ n27738 ^ 1'b0 ;
  assign n45953 = n33326 ^ n25465 ^ n14675 ;
  assign n45954 = n32329 ^ n24793 ^ n16484 ;
  assign n45955 = n31831 ^ n21472 ^ 1'b0 ;
  assign n45956 = n28832 ^ n12242 ^ 1'b0 ;
  assign n45957 = n1785 | n3091 ;
  assign n45958 = ( n14829 & n45956 ) | ( n14829 & n45957 ) | ( n45956 & n45957 ) ;
  assign n45959 = n11700 ^ n10945 ^ 1'b0 ;
  assign n45960 = n7914 | n45959 ;
  assign n45961 = n45960 ^ n22621 ^ n7750 ;
  assign n45962 = n8853 ^ n7364 ^ 1'b0 ;
  assign n45963 = x55 & n45962 ;
  assign n45964 = n39612 ^ n11324 ^ 1'b0 ;
  assign n45965 = ~n11153 & n23462 ;
  assign n45966 = n45965 ^ n22141 ^ 1'b0 ;
  assign n45967 = ~n42118 & n45966 ;
  assign n45968 = n45964 & n45967 ;
  assign n45969 = n45963 | n45968 ;
  assign n45970 = n486 & n38645 ;
  assign n45971 = n16514 ^ n11252 ^ 1'b0 ;
  assign n45972 = n12766 ^ n6421 ^ n4857 ;
  assign n45973 = ( ~n10934 & n13610 ) | ( ~n10934 & n45972 ) | ( n13610 & n45972 ) ;
  assign n45974 = n11186 ^ n893 ^ 1'b0 ;
  assign n45975 = n26867 | n45974 ;
  assign n45976 = n45975 ^ n17192 ^ n6079 ;
  assign n45977 = n18339 ^ n6275 ^ 1'b0 ;
  assign n45978 = n17377 ^ n7698 ^ 1'b0 ;
  assign n45979 = n34071 & ~n45978 ;
  assign n45980 = n36244 ^ n22492 ^ 1'b0 ;
  assign n45981 = n9814 & ~n45980 ;
  assign n45982 = n7801 | n14697 ;
  assign n45983 = ( n8250 & ~n9414 ) | ( n8250 & n24248 ) | ( ~n9414 & n24248 ) ;
  assign n45984 = n17727 & n45983 ;
  assign n45985 = ~n45982 & n45984 ;
  assign n45989 = n11307 ^ n8398 ^ 1'b0 ;
  assign n45990 = ~n1168 & n45989 ;
  assign n45991 = n45990 ^ n42352 ^ n10842 ;
  assign n45986 = n10628 & ~n24698 ;
  assign n45987 = ~n11159 & n37037 ;
  assign n45988 = n45986 & n45987 ;
  assign n45992 = n45991 ^ n45988 ^ 1'b0 ;
  assign n45993 = n31866 ^ n20963 ^ 1'b0 ;
  assign n45994 = ( n13518 & n30172 ) | ( n13518 & ~n42760 ) | ( n30172 & ~n42760 ) ;
  assign n45995 = n2153 | n34875 ;
  assign n45996 = n41560 | n45995 ;
  assign n45997 = n45994 & ~n45996 ;
  assign n45998 = n29899 ^ n27083 ^ n23588 ;
  assign n45999 = n7535 & ~n19408 ;
  assign n46000 = n45999 ^ n1265 ^ 1'b0 ;
  assign n46001 = n17778 ^ n8399 ^ 1'b0 ;
  assign n46004 = x228 & n33391 ;
  assign n46002 = n8726 & n27589 ;
  assign n46003 = ~n7227 & n46002 ;
  assign n46005 = n46004 ^ n46003 ^ 1'b0 ;
  assign n46006 = n25095 ^ n21621 ^ 1'b0 ;
  assign n46007 = ~n46005 & n46006 ;
  assign n46008 = n6582 & n37980 ;
  assign n46009 = n46008 ^ n1616 ^ 1'b0 ;
  assign n46010 = n35156 ^ n18388 ^ 1'b0 ;
  assign n46011 = ~n46009 & n46010 ;
  assign n46012 = n37817 ^ n30421 ^ n7135 ;
  assign n46013 = n13635 & n46012 ;
  assign n46014 = n46013 ^ n8527 ^ x152 ;
  assign n46015 = n31198 ^ n15571 ^ n7963 ;
  assign n46016 = ~n4429 & n26044 ;
  assign n46017 = n14115 & n46016 ;
  assign n46018 = n46017 ^ n5489 ^ n1336 ;
  assign n46020 = n43605 ^ n7141 ^ 1'b0 ;
  assign n46021 = ( n9974 & n12684 ) | ( n9974 & n46020 ) | ( n12684 & n46020 ) ;
  assign n46022 = n46021 ^ n31021 ^ n11724 ;
  assign n46019 = n10079 & ~n16966 ;
  assign n46023 = n46022 ^ n46019 ^ n18899 ;
  assign n46024 = n4006 & ~n11837 ;
  assign n46025 = n46024 ^ n27456 ^ n26637 ;
  assign n46026 = n3924 & ~n9458 ;
  assign n46027 = n12155 & n46026 ;
  assign n46028 = n46027 ^ n28559 ^ 1'b0 ;
  assign n46029 = n1753 | n10575 ;
  assign n46030 = x253 | n46029 ;
  assign n46031 = n15334 ^ n4446 ^ 1'b0 ;
  assign n46032 = n46030 & ~n46031 ;
  assign n46033 = n2592 | n46032 ;
  assign n46034 = ( n7678 & ~n38699 ) | ( n7678 & n46033 ) | ( ~n38699 & n46033 ) ;
  assign n46035 = ( n6273 & ~n6560 ) | ( n6273 & n17014 ) | ( ~n6560 & n17014 ) ;
  assign n46036 = ( n8551 & ~n29121 ) | ( n8551 & n46035 ) | ( ~n29121 & n46035 ) ;
  assign n46037 = ( n22585 & ~n35426 ) | ( n22585 & n46036 ) | ( ~n35426 & n46036 ) ;
  assign n46038 = n6681 & ~n44244 ;
  assign n46039 = n43584 ^ n16858 ^ 1'b0 ;
  assign n46040 = n2411 & ~n16112 ;
  assign n46041 = n46040 ^ n20718 ^ 1'b0 ;
  assign n46042 = ~n21501 & n43887 ;
  assign n46043 = n2908 & ~n27846 ;
  assign n46044 = n46043 ^ n11704 ^ 1'b0 ;
  assign n46045 = n46044 ^ n34190 ^ n7160 ;
  assign n46046 = ( ~n14140 & n21041 ) | ( ~n14140 & n21962 ) | ( n21041 & n21962 ) ;
  assign n46047 = n46046 ^ n39641 ^ 1'b0 ;
  assign n46048 = ~n28649 & n32963 ;
  assign n46049 = n7775 ^ n2472 ^ 1'b0 ;
  assign n46050 = ~n3960 & n46049 ;
  assign n46051 = ~n30350 & n46050 ;
  assign n46052 = n8506 ^ n5739 ^ 1'b0 ;
  assign n46053 = ~n2252 & n46052 ;
  assign n46054 = n13643 & ~n46053 ;
  assign n46055 = n46054 ^ n15333 ^ 1'b0 ;
  assign n46056 = ( n3719 & n46051 ) | ( n3719 & n46055 ) | ( n46051 & n46055 ) ;
  assign n46057 = n8309 & ~n12327 ;
  assign n46058 = ~n20415 & n46057 ;
  assign n46059 = n46058 ^ n19154 ^ n10037 ;
  assign n46060 = n36887 ^ n2822 ^ 1'b0 ;
  assign n46061 = n29472 ^ n6872 ^ 1'b0 ;
  assign n46062 = ~n7555 & n46061 ;
  assign n46063 = n23116 ^ n20937 ^ 1'b0 ;
  assign n46064 = n40460 & n46063 ;
  assign n46065 = ( n11376 & ~n26562 ) | ( n11376 & n43912 ) | ( ~n26562 & n43912 ) ;
  assign n46066 = n46065 ^ n16375 ^ n9654 ;
  assign n46067 = n46066 ^ n29288 ^ n12282 ;
  assign n46068 = n42740 ^ n759 ^ 1'b0 ;
  assign n46069 = n29860 ^ n20315 ^ n14906 ;
  assign n46070 = n9142 ^ n6665 ^ 1'b0 ;
  assign n46071 = n17747 & n46070 ;
  assign n46072 = ~n6684 & n7478 ;
  assign n46073 = ~n12101 & n46072 ;
  assign n46074 = n27236 ^ n19723 ^ 1'b0 ;
  assign n46075 = ~n12953 & n46074 ;
  assign n46076 = ~n11671 & n46075 ;
  assign n46079 = ~n3675 & n6042 ;
  assign n46080 = n10780 & n46079 ;
  assign n46077 = n14491 ^ n14138 ^ 1'b0 ;
  assign n46078 = ~n32501 & n46077 ;
  assign n46081 = n46080 ^ n46078 ^ 1'b0 ;
  assign n46082 = n30224 & n46081 ;
  assign n46083 = n1697 & n13349 ;
  assign n46084 = n12285 & ~n13591 ;
  assign n46085 = n9146 | n18571 ;
  assign n46086 = n7563 & ~n46085 ;
  assign n46087 = n46086 ^ n17788 ^ n16084 ;
  assign n46088 = n41706 & ~n46087 ;
  assign n46089 = ~n46084 & n46088 ;
  assign n46090 = ( n14501 & n46083 ) | ( n14501 & ~n46089 ) | ( n46083 & ~n46089 ) ;
  assign n46093 = n18733 ^ n10543 ^ 1'b0 ;
  assign n46094 = ( n11143 & ~n22082 ) | ( n11143 & n46093 ) | ( ~n22082 & n46093 ) ;
  assign n46095 = n14517 & n20092 ;
  assign n46096 = n46095 ^ n26488 ^ 1'b0 ;
  assign n46097 = ~n19509 & n46096 ;
  assign n46098 = ~n15691 & n46097 ;
  assign n46099 = ~n46094 & n46098 ;
  assign n46091 = n3734 | n22010 ;
  assign n46092 = ~n10731 & n46091 ;
  assign n46100 = n46099 ^ n46092 ^ n38705 ;
  assign n46101 = ( n3780 & n31076 ) | ( n3780 & n33593 ) | ( n31076 & n33593 ) ;
  assign n46102 = n44009 ^ n33490 ^ n6721 ;
  assign n46103 = ~n46101 & n46102 ;
  assign n46104 = n27900 ^ n12903 ^ n12090 ;
  assign n46105 = n33557 & ~n46104 ;
  assign n46106 = ~n42897 & n46105 ;
  assign n46107 = ( ~n6780 & n9023 ) | ( ~n6780 & n27476 ) | ( n9023 & n27476 ) ;
  assign n46108 = n46107 ^ n3103 ^ 1'b0 ;
  assign n46109 = n24716 ^ n7291 ^ n1512 ;
  assign n46110 = n22032 & n46109 ;
  assign n46111 = n22524 & n35033 ;
  assign n46112 = n38666 & n46111 ;
  assign n46113 = n33808 & n46112 ;
  assign n46114 = n27243 ^ n8414 ^ 1'b0 ;
  assign n46115 = ( ~n4708 & n26883 ) | ( ~n4708 & n40898 ) | ( n26883 & n40898 ) ;
  assign n46116 = n10797 & n21042 ;
  assign n46117 = ( n3921 & n10367 ) | ( n3921 & n15020 ) | ( n10367 & n15020 ) ;
  assign n46118 = n41238 ^ n8270 ^ 1'b0 ;
  assign n46119 = n46117 & n46118 ;
  assign n46120 = ( ~n25247 & n27434 ) | ( ~n25247 & n41496 ) | ( n27434 & n41496 ) ;
  assign n46121 = n46120 ^ n12867 ^ 1'b0 ;
  assign n46122 = n40225 | n46121 ;
  assign n46123 = ( ~n10197 & n25889 ) | ( ~n10197 & n27453 ) | ( n25889 & n27453 ) ;
  assign n46124 = n35858 ^ n3771 ^ 1'b0 ;
  assign n46125 = n46123 | n46124 ;
  assign n46126 = n16878 ^ n11097 ^ n6358 ;
  assign n46127 = ( n17687 & n41494 ) | ( n17687 & n46126 ) | ( n41494 & n46126 ) ;
  assign n46128 = ( ~n3242 & n15784 ) | ( ~n3242 & n46127 ) | ( n15784 & n46127 ) ;
  assign n46129 = n4577 & n41265 ;
  assign n46130 = n46129 ^ n24639 ^ n14371 ;
  assign n46131 = n30519 ^ n15865 ^ 1'b0 ;
  assign n46140 = ~n13616 & n24336 ;
  assign n46141 = n46140 ^ x9 ^ 1'b0 ;
  assign n46138 = n35158 ^ n21868 ^ 1'b0 ;
  assign n46139 = ~n19776 & n46138 ;
  assign n46132 = n39654 ^ n23475 ^ n2117 ;
  assign n46133 = n10779 | n46132 ;
  assign n46134 = n46133 ^ n7827 ^ n1461 ;
  assign n46135 = n32619 ^ n7694 ^ 1'b0 ;
  assign n46136 = n46134 | n46135 ;
  assign n46137 = n46136 ^ n10663 ^ 1'b0 ;
  assign n46142 = n46141 ^ n46139 ^ n46137 ;
  assign n46143 = n39605 ^ n17466 ^ n4027 ;
  assign n46144 = n3330 | n33074 ;
  assign n46145 = n15240 & ~n46144 ;
  assign n46146 = n46145 ^ n33400 ^ 1'b0 ;
  assign n46147 = n33792 | n46146 ;
  assign n46148 = ~n14362 & n40282 ;
  assign n46149 = n46148 ^ n1068 ^ 1'b0 ;
  assign n46150 = n25077 & ~n43600 ;
  assign n46151 = n17130 & ~n46150 ;
  assign n46152 = n46151 ^ n21837 ^ 1'b0 ;
  assign n46153 = ( n3067 & ~n11467 ) | ( n3067 & n13039 ) | ( ~n11467 & n13039 ) ;
  assign n46154 = n2394 | n19124 ;
  assign n46155 = n21619 ^ n20353 ^ 1'b0 ;
  assign n46157 = n13819 & ~n14122 ;
  assign n46158 = n46157 ^ n27851 ^ 1'b0 ;
  assign n46156 = ~n26537 & n37799 ;
  assign n46159 = n46158 ^ n46156 ^ 1'b0 ;
  assign n46160 = n44572 ^ n17349 ^ 1'b0 ;
  assign n46161 = x11 & n46160 ;
  assign n46162 = n41645 ^ n36543 ^ n18942 ;
  assign n46169 = ~n10007 & n17234 ;
  assign n46170 = ~n2407 & n46169 ;
  assign n46171 = n1274 & n46170 ;
  assign n46164 = n7479 & n32836 ;
  assign n46165 = n5766 & n46164 ;
  assign n46166 = n46165 ^ n37190 ^ n16776 ;
  assign n46163 = n8110 & ~n22307 ;
  assign n46167 = n46166 ^ n46163 ^ 1'b0 ;
  assign n46168 = n46167 ^ n6660 ^ n5725 ;
  assign n46172 = n46171 ^ n46168 ^ n16196 ;
  assign n46173 = n2450 & ~n18942 ;
  assign n46174 = n1158 & n46173 ;
  assign n46175 = n18657 & ~n46174 ;
  assign n46176 = ( n1017 & n9904 ) | ( n1017 & n46175 ) | ( n9904 & n46175 ) ;
  assign n46178 = n17427 ^ n12180 ^ 1'b0 ;
  assign n46179 = n8868 & ~n46178 ;
  assign n46177 = ~n13789 & n18000 ;
  assign n46180 = n46179 ^ n46177 ^ n42677 ;
  assign n46181 = ( n7310 & n31383 ) | ( n7310 & ~n46180 ) | ( n31383 & ~n46180 ) ;
  assign n46183 = ( ~n5699 & n6763 ) | ( ~n5699 & n13776 ) | ( n6763 & n13776 ) ;
  assign n46182 = n5982 | n35752 ;
  assign n46184 = n46183 ^ n46182 ^ 1'b0 ;
  assign n46185 = n40782 ^ n6509 ^ 1'b0 ;
  assign n46186 = n46184 | n46185 ;
  assign n46187 = n3093 & n42318 ;
  assign n46188 = n35142 ^ n12901 ^ n464 ;
  assign n46189 = ~n16018 & n46188 ;
  assign n46190 = n46189 ^ n22360 ^ 1'b0 ;
  assign n46191 = n7394 ^ x62 ^ 1'b0 ;
  assign n46192 = n5991 & ~n27631 ;
  assign n46193 = ~n4307 & n46192 ;
  assign n46194 = n46193 ^ n24740 ^ n20617 ;
  assign n46195 = ~n21736 & n28726 ;
  assign n46196 = ~n17234 & n46195 ;
  assign n46197 = n46196 ^ n34145 ^ x199 ;
  assign n46198 = n15271 | n16690 ;
  assign n46199 = n5266 | n46198 ;
  assign n46200 = ~n24067 & n46199 ;
  assign n46201 = ( ~n17609 & n23437 ) | ( ~n17609 & n46200 ) | ( n23437 & n46200 ) ;
  assign n46202 = n869 | n9700 ;
  assign n46203 = n46202 ^ n29645 ^ 1'b0 ;
  assign n46204 = ( n2792 & ~n21508 ) | ( n2792 & n46203 ) | ( ~n21508 & n46203 ) ;
  assign n46205 = n24049 ^ n11773 ^ n10896 ;
  assign n46206 = n10540 ^ n1754 ^ 1'b0 ;
  assign n46207 = n46206 ^ n36921 ^ 1'b0 ;
  assign n46208 = n16703 & ~n46207 ;
  assign n46209 = n8020 & n31474 ;
  assign n46210 = n20617 ^ n18167 ^ 1'b0 ;
  assign n46211 = n38517 & n46210 ;
  assign n46212 = n46211 ^ n8131 ^ 1'b0 ;
  assign n46213 = n9947 & ~n46212 ;
  assign n46214 = n728 & ~n24224 ;
  assign n46215 = n46214 ^ n17403 ^ n13237 ;
  assign n46216 = n32739 ^ n27100 ^ 1'b0 ;
  assign n46217 = n2201 ^ n1255 ^ 1'b0 ;
  assign n46218 = n46217 ^ n26244 ^ n2448 ;
  assign n46219 = n32754 & n35972 ;
  assign n46220 = ( n28090 & n33067 ) | ( n28090 & ~n38882 ) | ( n33067 & ~n38882 ) ;
  assign n46221 = n46220 ^ n12428 ^ 1'b0 ;
  assign n46222 = n46219 & ~n46221 ;
  assign n46223 = n46222 ^ n20118 ^ n18331 ;
  assign n46224 = n1312 & ~n33662 ;
  assign n46225 = n46224 ^ n41242 ^ 1'b0 ;
  assign n46226 = n7237 | n9195 ;
  assign n46227 = n15835 ^ n15737 ^ 1'b0 ;
  assign n46228 = n13317 & ~n46227 ;
  assign n46229 = n12456 ^ n7167 ^ n1559 ;
  assign n46230 = n46229 ^ n5570 ^ 1'b0 ;
  assign n46231 = n46228 & ~n46230 ;
  assign n46232 = n4474 & ~n25092 ;
  assign n46233 = n26663 | n31014 ;
  assign n46234 = ~n4740 & n46233 ;
  assign n46235 = ( n7589 & n42122 ) | ( n7589 & ~n46234 ) | ( n42122 & ~n46234 ) ;
  assign n46236 = n11855 ^ n10022 ^ 1'b0 ;
  assign n46237 = ~n9132 & n46236 ;
  assign n46238 = ( n14739 & ~n42348 ) | ( n14739 & n46237 ) | ( ~n42348 & n46237 ) ;
  assign n46239 = ( n3507 & n17259 ) | ( n3507 & ~n24985 ) | ( n17259 & ~n24985 ) ;
  assign n46240 = n46239 ^ n14086 ^ n2767 ;
  assign n46241 = ~n12403 & n18886 ;
  assign n46242 = n46241 ^ n18602 ^ 1'b0 ;
  assign n46243 = n33029 ^ n1475 ^ 1'b0 ;
  assign n46244 = n16844 & n46243 ;
  assign n46245 = ~n19054 & n46244 ;
  assign n46246 = n46245 ^ n21543 ^ 1'b0 ;
  assign n46247 = n23563 | n26581 ;
  assign n46248 = n46247 ^ n8447 ^ 1'b0 ;
  assign n46249 = n23249 ^ n11737 ^ n2528 ;
  assign n46250 = n46249 ^ n25476 ^ 1'b0 ;
  assign n46251 = n25769 & n46250 ;
  assign n46252 = n9199 | n11851 ;
  assign n46253 = n1655 & ~n46252 ;
  assign n46254 = ( n12756 & n28726 ) | ( n12756 & n46253 ) | ( n28726 & n46253 ) ;
  assign n46255 = ( n46237 & n46251 ) | ( n46237 & n46254 ) | ( n46251 & n46254 ) ;
  assign n46256 = n29343 ^ n18231 ^ n9472 ;
  assign n46257 = ( n3043 & n34305 ) | ( n3043 & ~n46256 ) | ( n34305 & ~n46256 ) ;
  assign n46258 = n34995 | n46257 ;
  assign n46259 = n46258 ^ n36797 ^ n13035 ;
  assign n46260 = n31600 ^ n25319 ^ 1'b0 ;
  assign n46261 = n13702 & n19164 ;
  assign n46262 = n7415 & n46261 ;
  assign n46263 = n11034 & ~n20551 ;
  assign n46264 = ( n2638 & n46262 ) | ( n2638 & ~n46263 ) | ( n46262 & ~n46263 ) ;
  assign n46265 = n46264 ^ n18769 ^ 1'b0 ;
  assign n46266 = n3813 & ~n46265 ;
  assign n46267 = ( n2860 & n14636 ) | ( n2860 & n20556 ) | ( n14636 & n20556 ) ;
  assign n46268 = n46267 ^ n5982 ^ 1'b0 ;
  assign n46269 = n18289 & n46268 ;
  assign n46270 = ( ~n12011 & n12018 ) | ( ~n12011 & n24664 ) | ( n12018 & n24664 ) ;
  assign n46271 = n9184 | n10674 ;
  assign n46272 = n4314 | n46271 ;
  assign n46273 = n46272 ^ n42729 ^ n5292 ;
  assign n46274 = ( n19299 & n46270 ) | ( n19299 & ~n46273 ) | ( n46270 & ~n46273 ) ;
  assign n46275 = n16317 & n37987 ;
  assign n46276 = n46275 ^ n25635 ^ 1'b0 ;
  assign n46277 = n46276 ^ n34454 ^ n27350 ;
  assign n46278 = n9522 ^ n1742 ^ 1'b0 ;
  assign n46279 = ( ~n22572 & n45487 ) | ( ~n22572 & n46278 ) | ( n45487 & n46278 ) ;
  assign n46280 = n14130 ^ n4482 ^ n1863 ;
  assign n46281 = n46280 ^ n15337 ^ n12383 ;
  assign n46282 = n17935 | n19248 ;
  assign n46283 = n13997 & ~n46282 ;
  assign n46284 = ( n17827 & ~n40631 ) | ( n17827 & n46283 ) | ( ~n40631 & n46283 ) ;
  assign n46286 = ( n2411 & n7646 ) | ( n2411 & ~n11021 ) | ( n7646 & ~n11021 ) ;
  assign n46287 = ( ~n8951 & n11044 ) | ( ~n8951 & n46286 ) | ( n11044 & n46286 ) ;
  assign n46285 = n17640 | n32046 ;
  assign n46288 = n46287 ^ n46285 ^ 1'b0 ;
  assign n46289 = n39013 ^ n18490 ^ 1'b0 ;
  assign n46290 = n5183 & ~n40341 ;
  assign n46291 = n46289 & n46290 ;
  assign n46292 = n5573 & n8533 ;
  assign n46293 = n30705 & n46292 ;
  assign n46294 = n8344 & n33493 ;
  assign n46295 = n46294 ^ n10514 ^ 1'b0 ;
  assign n46296 = n27510 ^ n18760 ^ n4473 ;
  assign n46297 = n45968 ^ n25067 ^ 1'b0 ;
  assign n46298 = n46296 | n46297 ;
  assign n46299 = ( n2923 & n6420 ) | ( n2923 & n8555 ) | ( n6420 & n8555 ) ;
  assign n46300 = n37543 ^ n2020 ^ 1'b0 ;
  assign n46301 = n19456 | n46300 ;
  assign n46302 = ( ~n1006 & n17842 ) | ( ~n1006 & n46301 ) | ( n17842 & n46301 ) ;
  assign n46303 = ( n3466 & ~n11008 ) | ( n3466 & n46302 ) | ( ~n11008 & n46302 ) ;
  assign n46304 = n45682 ^ n2401 ^ 1'b0 ;
  assign n46305 = n35701 & n46304 ;
  assign n46306 = ( n40786 & ~n46303 ) | ( n40786 & n46305 ) | ( ~n46303 & n46305 ) ;
  assign n46307 = ( n7790 & n10907 ) | ( n7790 & ~n30907 ) | ( n10907 & ~n30907 ) ;
  assign n46308 = n27101 ^ n21083 ^ n2803 ;
  assign n46309 = ( n12425 & ~n37795 ) | ( n12425 & n46308 ) | ( ~n37795 & n46308 ) ;
  assign n46310 = n39288 ^ n26312 ^ 1'b0 ;
  assign n46311 = ~n9721 & n25706 ;
  assign n46312 = ~n46310 & n46311 ;
  assign n46313 = n14068 ^ n10048 ^ n4644 ;
  assign n46314 = n17479 ^ n11924 ^ 1'b0 ;
  assign n46315 = ( ~n4253 & n33533 ) | ( ~n4253 & n46314 ) | ( n33533 & n46314 ) ;
  assign n46316 = ~n26652 & n46315 ;
  assign n46317 = n46316 ^ n2045 ^ 1'b0 ;
  assign n46318 = n22823 | n46317 ;
  assign n46319 = n46313 | n46318 ;
  assign n46320 = n41712 ^ n6693 ^ 1'b0 ;
  assign n46321 = n18916 | n46320 ;
  assign n46322 = n14473 & ~n46321 ;
  assign n46323 = n44464 & n46322 ;
  assign n46324 = n36083 ^ n27933 ^ n20529 ;
  assign n46325 = n27747 ^ n10000 ^ n6679 ;
  assign n46326 = ( ~n13356 & n15798 ) | ( ~n13356 & n46325 ) | ( n15798 & n46325 ) ;
  assign n46327 = n39449 ^ n19213 ^ n1665 ;
  assign n46328 = n25628 ^ n1915 ^ 1'b0 ;
  assign n46329 = ( x14 & n388 ) | ( x14 & n8619 ) | ( n388 & n8619 ) ;
  assign n46330 = n15326 & ~n46329 ;
  assign n46331 = n9526 & n46330 ;
  assign n46332 = n46331 ^ n24948 ^ n24089 ;
  assign n46333 = n5114 | n36229 ;
  assign n46334 = n35531 ^ n24261 ^ 1'b0 ;
  assign n46335 = ( n6982 & n9377 ) | ( n6982 & n15558 ) | ( n9377 & n15558 ) ;
  assign n46336 = ~n6252 & n16247 ;
  assign n46337 = ~n44486 & n46336 ;
  assign n46338 = n46335 & n46337 ;
  assign n46339 = n17813 ^ n5238 ^ 1'b0 ;
  assign n46340 = ~n46338 & n46339 ;
  assign n46341 = n6978 & n21475 ;
  assign n46342 = ( n482 & n23704 ) | ( n482 & n46341 ) | ( n23704 & n46341 ) ;
  assign n46343 = n2092 & n15228 ;
  assign n46344 = n46343 ^ n2215 ^ 1'b0 ;
  assign n46345 = ( ~n30517 & n46342 ) | ( ~n30517 & n46344 ) | ( n46342 & n46344 ) ;
  assign n46346 = n3973 & ~n11044 ;
  assign n46347 = n45040 & n46346 ;
  assign n46348 = n33446 & ~n46347 ;
  assign n46349 = ( n4417 & n16520 ) | ( n4417 & ~n46348 ) | ( n16520 & ~n46348 ) ;
  assign n46350 = ( n13154 & ~n25884 ) | ( n13154 & n26120 ) | ( ~n25884 & n26120 ) ;
  assign n46351 = n11587 ^ n5570 ^ 1'b0 ;
  assign n46352 = n46351 ^ n32272 ^ n29946 ;
  assign n46353 = n46352 ^ n32503 ^ n5085 ;
  assign n46354 = n30805 ^ n24165 ^ n20172 ;
  assign n46355 = n13798 & n21519 ;
  assign n46356 = n46355 ^ n31431 ^ 1'b0 ;
  assign n46357 = n41988 ^ n8122 ^ 1'b0 ;
  assign n46358 = n37745 & ~n46357 ;
  assign n46359 = n46358 ^ n22135 ^ 1'b0 ;
  assign n46360 = n12053 | n45604 ;
  assign n46361 = n12755 & ~n46360 ;
  assign n46362 = n46359 & n46361 ;
  assign n46363 = n45158 ^ n16855 ^ 1'b0 ;
  assign n46364 = n4514 | n37479 ;
  assign n46365 = n46364 ^ n38127 ^ 1'b0 ;
  assign n46366 = n9624 & ~n35248 ;
  assign n46367 = ( ~n4842 & n5523 ) | ( ~n4842 & n22345 ) | ( n5523 & n22345 ) ;
  assign n46368 = n46367 ^ n26519 ^ n22538 ;
  assign n46370 = n3368 ^ n1331 ^ 1'b0 ;
  assign n46371 = n41138 & ~n46370 ;
  assign n46369 = n33502 ^ n22765 ^ n12742 ;
  assign n46372 = n46371 ^ n46369 ^ n8802 ;
  assign n46373 = n44305 ^ n15491 ^ n541 ;
  assign n46374 = n44868 ^ n26639 ^ 1'b0 ;
  assign n46376 = n17342 ^ n11490 ^ 1'b0 ;
  assign n46377 = n3488 | n46376 ;
  assign n46378 = ~n8721 & n19270 ;
  assign n46379 = n859 & n46378 ;
  assign n46380 = n46379 ^ n7473 ^ n4118 ;
  assign n46381 = n46377 & ~n46380 ;
  assign n46375 = n5442 & n43937 ;
  assign n46382 = n46381 ^ n46375 ^ 1'b0 ;
  assign n46383 = ( n14656 & ~n19708 ) | ( n14656 & n46382 ) | ( ~n19708 & n46382 ) ;
  assign n46385 = n17509 ^ n1304 ^ 1'b0 ;
  assign n46386 = n24208 & n46385 ;
  assign n46387 = n3769 & ~n46386 ;
  assign n46384 = n4455 | n5089 ;
  assign n46388 = n46387 ^ n46384 ^ 1'b0 ;
  assign n46389 = n23900 ^ n4359 ^ 1'b0 ;
  assign n46390 = ~n3658 & n27906 ;
  assign n46391 = n32162 ^ n16131 ^ n7916 ;
  assign n46392 = n5840 ^ n4255 ^ 1'b0 ;
  assign n46393 = n46391 & ~n46392 ;
  assign n46394 = n35853 ^ n16784 ^ n12606 ;
  assign n46395 = n12581 & n27453 ;
  assign n46396 = n21152 & ~n40209 ;
  assign n46397 = n851 & n24247 ;
  assign n46398 = ( ~n31972 & n37015 ) | ( ~n31972 & n46397 ) | ( n37015 & n46397 ) ;
  assign n46399 = ( n10337 & n14826 ) | ( n10337 & n36291 ) | ( n14826 & n36291 ) ;
  assign n46400 = n22668 & n28805 ;
  assign n46401 = ~n32237 & n46400 ;
  assign n46402 = x159 | n457 ;
  assign n46403 = n2730 | n16034 ;
  assign n46404 = n46403 ^ n13903 ^ 1'b0 ;
  assign n46405 = ~n9455 & n15668 ;
  assign n46406 = n28189 ^ n26753 ^ n2361 ;
  assign n46409 = ( n9647 & n15391 ) | ( n9647 & n24146 ) | ( n15391 & n24146 ) ;
  assign n46407 = n6856 & n38891 ;
  assign n46408 = n8754 | n46407 ;
  assign n46410 = n46409 ^ n46408 ^ n2003 ;
  assign n46411 = ( ~n34510 & n46406 ) | ( ~n34510 & n46410 ) | ( n46406 & n46410 ) ;
  assign n46412 = n44858 ^ n42649 ^ n24473 ;
  assign n46413 = n21048 ^ n9209 ^ 1'b0 ;
  assign n46414 = ( n21628 & n24214 ) | ( n21628 & ~n46413 ) | ( n24214 & ~n46413 ) ;
  assign n46415 = n25058 ^ n24610 ^ n21573 ;
  assign n46416 = n8361 & ~n37463 ;
  assign n46417 = ~n11307 & n28873 ;
  assign n46418 = n46417 ^ n42859 ^ 1'b0 ;
  assign n46419 = n13812 ^ n13431 ^ 1'b0 ;
  assign n46420 = n19619 & n46419 ;
  assign n46421 = ~n31433 & n46420 ;
  assign n46422 = n30624 & n45304 ;
  assign n46425 = x151 & n16167 ;
  assign n46423 = n7655 & ~n14968 ;
  assign n46424 = n46423 ^ n34768 ^ 1'b0 ;
  assign n46426 = n46425 ^ n46424 ^ n23467 ;
  assign n46427 = n21340 ^ n11431 ^ n2325 ;
  assign n46428 = n25662 ^ n13771 ^ n3641 ;
  assign n46429 = ( n7694 & ~n42816 ) | ( n7694 & n46428 ) | ( ~n42816 & n46428 ) ;
  assign n46430 = ( n6270 & n13659 ) | ( n6270 & ~n23457 ) | ( n13659 & ~n23457 ) ;
  assign n46431 = n5338 & ~n46430 ;
  assign n46432 = n25020 ^ n6543 ^ 1'b0 ;
  assign n46433 = n32574 & n46432 ;
  assign n46434 = n46433 ^ n45908 ^ n9809 ;
  assign n46435 = n27972 | n40141 ;
  assign n46436 = ( n1277 & n14080 ) | ( n1277 & ~n46435 ) | ( n14080 & ~n46435 ) ;
  assign n46437 = n46436 ^ n32519 ^ 1'b0 ;
  assign n46438 = ~n17931 & n26930 ;
  assign n46439 = n15293 & n46438 ;
  assign n46440 = n7706 & ~n11892 ;
  assign n46441 = n8699 & n46440 ;
  assign n46442 = n46441 ^ n30242 ^ 1'b0 ;
  assign n46443 = n6620 & ~n16763 ;
  assign n46444 = ~n46442 & n46443 ;
  assign n46445 = ( n3110 & ~n25662 ) | ( n3110 & n32562 ) | ( ~n25662 & n32562 ) ;
  assign n46446 = n46445 ^ n26727 ^ 1'b0 ;
  assign n46447 = n28959 ^ n24254 ^ n17119 ;
  assign n46448 = n30856 ^ n4155 ^ 1'b0 ;
  assign n46449 = ~n37323 & n46448 ;
  assign n46450 = ( n22675 & n29976 ) | ( n22675 & ~n46449 ) | ( n29976 & ~n46449 ) ;
  assign n46451 = n9175 | n22373 ;
  assign n46452 = n46451 ^ n9976 ^ 1'b0 ;
  assign n46453 = n5027 | n46452 ;
  assign n46454 = ( n11077 & ~n42096 ) | ( n11077 & n46453 ) | ( ~n42096 & n46453 ) ;
  assign n46455 = n27698 & ~n33811 ;
  assign n46456 = n20504 ^ n18563 ^ 1'b0 ;
  assign n46457 = n34022 & ~n46456 ;
  assign n46458 = n27146 & n46457 ;
  assign n46459 = n23204 & n46458 ;
  assign n46460 = ~n4212 & n41408 ;
  assign n46461 = n46460 ^ n39458 ^ 1'b0 ;
  assign n46462 = n39864 ^ n7321 ^ 1'b0 ;
  assign n46463 = n34214 & ~n46462 ;
  assign n46464 = ( n13946 & n27093 ) | ( n13946 & n31166 ) | ( n27093 & n31166 ) ;
  assign n46465 = n5343 & n10737 ;
  assign n46466 = n46465 ^ n23310 ^ 1'b0 ;
  assign n46467 = n23767 & n46466 ;
  assign n46468 = n44140 | n46467 ;
  assign n46469 = n10873 & n34566 ;
  assign n46470 = n19862 ^ n18602 ^ 1'b0 ;
  assign n46471 = n17091 & ~n46470 ;
  assign n46472 = n46471 ^ n44971 ^ 1'b0 ;
  assign n46473 = ( n6360 & n45682 ) | ( n6360 & ~n46472 ) | ( n45682 & ~n46472 ) ;
  assign n46474 = ~n30466 & n45836 ;
  assign n46475 = x187 | n40494 ;
  assign n46476 = ( n24195 & ~n44263 ) | ( n24195 & n44549 ) | ( ~n44263 & n44549 ) ;
  assign n46477 = n21778 ^ n16980 ^ n11729 ;
  assign n46478 = n18086 & n46477 ;
  assign n46479 = n13621 ^ n8201 ^ 1'b0 ;
  assign n46480 = n15433 | n46479 ;
  assign n46481 = n46480 ^ n346 ^ 1'b0 ;
  assign n46482 = ~n39276 & n46481 ;
  assign n46483 = n8192 ^ n6267 ^ n5669 ;
  assign n46484 = ~n15380 & n46483 ;
  assign n46485 = n24578 & n46484 ;
  assign n46489 = n26855 ^ n26394 ^ n2995 ;
  assign n46486 = ~n2668 & n13449 ;
  assign n46487 = ~n988 & n46486 ;
  assign n46488 = x169 | n46487 ;
  assign n46490 = n46489 ^ n46488 ^ 1'b0 ;
  assign n46491 = n24321 | n34222 ;
  assign n46493 = ~n6120 & n7907 ;
  assign n46494 = n11744 & ~n18265 ;
  assign n46495 = n12050 & n46494 ;
  assign n46496 = n46495 ^ n14588 ^ 1'b0 ;
  assign n46497 = ~n46493 & n46496 ;
  assign n46492 = n1802 & ~n16115 ;
  assign n46498 = n46497 ^ n46492 ^ 1'b0 ;
  assign n46499 = ( n2759 & ~n5473 ) | ( n2759 & n10337 ) | ( ~n5473 & n10337 ) ;
  assign n46500 = ~n44120 & n46499 ;
  assign n46501 = ( n5435 & n13457 ) | ( n5435 & n46500 ) | ( n13457 & n46500 ) ;
  assign n46502 = ~n16577 & n29499 ;
  assign n46503 = ( n8418 & n43484 ) | ( n8418 & n46502 ) | ( n43484 & n46502 ) ;
  assign n46504 = n11129 & n12291 ;
  assign n46505 = n874 & n46504 ;
  assign n46506 = ( ~n11122 & n34210 ) | ( ~n11122 & n46505 ) | ( n34210 & n46505 ) ;
  assign n46507 = n13424 & ~n31331 ;
  assign n46508 = ( n27629 & n41957 ) | ( n27629 & ~n46507 ) | ( n41957 & ~n46507 ) ;
  assign n46509 = ~n436 & n36291 ;
  assign n46510 = n46509 ^ n11439 ^ 1'b0 ;
  assign n46511 = n18968 ^ n14262 ^ 1'b0 ;
  assign n46512 = n46511 ^ n14908 ^ 1'b0 ;
  assign n46513 = n16640 & n32271 ;
  assign n46514 = n27625 | n38735 ;
  assign n46515 = n46514 ^ n28320 ^ 1'b0 ;
  assign n46516 = n544 & ~n46515 ;
  assign n46517 = ~n46513 & n46516 ;
  assign n46518 = n15510 | n41669 ;
  assign n46519 = n32867 ^ n9570 ^ n6204 ;
  assign n46520 = n21765 | n29321 ;
  assign n46521 = n46520 ^ n16811 ^ 1'b0 ;
  assign n46522 = ( n13814 & ~n32055 ) | ( n13814 & n46521 ) | ( ~n32055 & n46521 ) ;
  assign n46523 = n4982 & n16952 ;
  assign n46524 = n31662 & ~n46523 ;
  assign n46525 = n488 & ~n30765 ;
  assign n46526 = n46525 ^ n31657 ^ 1'b0 ;
  assign n46527 = n46526 ^ n5328 ^ n626 ;
  assign n46530 = n17397 ^ n2595 ^ n2191 ;
  assign n46528 = n42119 ^ n34031 ^ n436 ;
  assign n46529 = n2949 | n46528 ;
  assign n46531 = n46530 ^ n46529 ^ 1'b0 ;
  assign n46532 = n37944 ^ n23076 ^ 1'b0 ;
  assign n46533 = ( ~n3821 & n5462 ) | ( ~n3821 & n16401 ) | ( n5462 & n16401 ) ;
  assign n46534 = n24411 | n42636 ;
  assign n46535 = n13506 & ~n32160 ;
  assign n46536 = ( ~n34456 & n46534 ) | ( ~n34456 & n46535 ) | ( n46534 & n46535 ) ;
  assign n46537 = n7031 | n10425 ;
  assign n46538 = n43282 & ~n46537 ;
  assign n46539 = ( ~n16818 & n23038 ) | ( ~n16818 & n46538 ) | ( n23038 & n46538 ) ;
  assign n46540 = n27575 ^ n26912 ^ n7282 ;
  assign n46541 = ( ~n648 & n4124 ) | ( ~n648 & n46540 ) | ( n4124 & n46540 ) ;
  assign n46542 = n46541 ^ n28111 ^ n18334 ;
  assign n46543 = n26518 ^ n15164 ^ 1'b0 ;
  assign n46544 = ~n1557 & n12317 ;
  assign n46545 = n7476 & ~n18814 ;
  assign n46546 = n46544 | n46545 ;
  assign n46547 = n18173 | n46546 ;
  assign n46548 = n13032 ^ n10880 ^ 1'b0 ;
  assign n46549 = n46548 ^ n25006 ^ n7308 ;
  assign n46550 = n11681 & ~n46549 ;
  assign n46551 = ~n24479 & n46550 ;
  assign n46552 = ~n35730 & n41031 ;
  assign n46553 = n4859 & n6778 ;
  assign n46554 = ( n4190 & n28330 ) | ( n4190 & ~n40533 ) | ( n28330 & ~n40533 ) ;
  assign n46557 = ~n25151 & n25724 ;
  assign n46558 = n18294 & n46557 ;
  assign n46555 = n20526 | n42242 ;
  assign n46556 = n46555 ^ n36766 ^ 1'b0 ;
  assign n46559 = n46558 ^ n46556 ^ n40170 ;
  assign n46560 = ~n4605 & n7196 ;
  assign n46561 = n11111 | n46560 ;
  assign n46562 = n46561 ^ n2002 ^ 1'b0 ;
  assign n46563 = n46562 ^ n37603 ^ n10157 ;
  assign n46564 = ( ~n27295 & n33249 ) | ( ~n27295 & n43790 ) | ( n33249 & n43790 ) ;
  assign n46565 = ( n34413 & n46563 ) | ( n34413 & ~n46564 ) | ( n46563 & ~n46564 ) ;
  assign n46566 = n17977 ^ n13208 ^ n10797 ;
  assign n46567 = n46566 ^ n26830 ^ 1'b0 ;
  assign n46568 = n19300 | n40937 ;
  assign n46569 = n23518 & ~n46568 ;
  assign n46572 = n19373 ^ n18291 ^ n17187 ;
  assign n46570 = n24188 ^ n5313 ^ n4054 ;
  assign n46571 = ~n1943 & n46570 ;
  assign n46573 = n46572 ^ n46571 ^ 1'b0 ;
  assign n46574 = n21544 | n34560 ;
  assign n46575 = n43112 & ~n46574 ;
  assign n46576 = n38366 ^ n19790 ^ n13514 ;
  assign n46577 = n41709 ^ n33088 ^ n28555 ;
  assign n46578 = n29030 ^ n12955 ^ 1'b0 ;
  assign n46579 = ~n21967 & n46578 ;
  assign n46580 = n2941 & n7013 ;
  assign n46581 = n46580 ^ n28376 ^ 1'b0 ;
  assign n46582 = n30376 ^ n15361 ^ 1'b0 ;
  assign n46583 = n4093 & ~n46582 ;
  assign n46584 = n39921 ^ n28981 ^ 1'b0 ;
  assign n46585 = n24943 ^ n2626 ^ 1'b0 ;
  assign n46586 = ( ~n8758 & n36076 ) | ( ~n8758 & n46585 ) | ( n36076 & n46585 ) ;
  assign n46588 = n26302 ^ n18931 ^ n9766 ;
  assign n46587 = ( n5710 & ~n5912 ) | ( n5710 & n30892 ) | ( ~n5912 & n30892 ) ;
  assign n46589 = n46588 ^ n46587 ^ n43184 ;
  assign n46590 = n46586 | n46589 ;
  assign n46591 = ( n4021 & n9492 ) | ( n4021 & ~n20951 ) | ( n9492 & ~n20951 ) ;
  assign n46592 = n46591 ^ n45501 ^ 1'b0 ;
  assign n46593 = n10916 | n46592 ;
  assign n46594 = n10865 ^ n1359 ^ n1153 ;
  assign n46595 = ( ~n15811 & n20805 ) | ( ~n15811 & n46594 ) | ( n20805 & n46594 ) ;
  assign n46596 = n21378 ^ n20058 ^ 1'b0 ;
  assign n46597 = ( n2333 & n28578 ) | ( n2333 & n46596 ) | ( n28578 & n46596 ) ;
  assign n46598 = ( ~n8510 & n14195 ) | ( ~n8510 & n37435 ) | ( n14195 & n37435 ) ;
  assign n46599 = n15839 & ~n46598 ;
  assign n46600 = n46599 ^ n8245 ^ 1'b0 ;
  assign n46601 = n18527 ^ n3619 ^ 1'b0 ;
  assign n46602 = n4049 & n46601 ;
  assign n46603 = n18832 & n46602 ;
  assign n46604 = ~n8620 & n46603 ;
  assign n46605 = n44506 ^ n4587 ^ 1'b0 ;
  assign n46606 = n46604 | n46605 ;
  assign n46607 = n22063 & ~n34303 ;
  assign n46608 = n46607 ^ n2081 ^ 1'b0 ;
  assign n46609 = ~n24160 & n46608 ;
  assign n46610 = n46609 ^ n30407 ^ 1'b0 ;
  assign n46611 = n4156 & ~n13999 ;
  assign n46612 = n46611 ^ n39280 ^ 1'b0 ;
  assign n46613 = n20424 | n41110 ;
  assign n46614 = n29060 & ~n46613 ;
  assign n46615 = n44478 ^ n34938 ^ n25533 ;
  assign n46616 = ~n1995 & n5995 ;
  assign n46617 = n355 & n46616 ;
  assign n46618 = n46617 ^ n31943 ^ 1'b0 ;
  assign n46619 = ~n12943 & n21520 ;
  assign n46620 = n1097 & n46619 ;
  assign n46621 = n13776 | n46620 ;
  assign n46622 = n46621 ^ n21428 ^ n5919 ;
  assign n46623 = n8598 | n23946 ;
  assign n46624 = n27553 & ~n46623 ;
  assign n46625 = n22852 | n29465 ;
  assign n46626 = n46625 ^ n32053 ^ 1'b0 ;
  assign n46627 = ~n43685 & n46626 ;
  assign n46628 = n23488 & ~n44327 ;
  assign n46629 = n13295 ^ n8411 ^ 1'b0 ;
  assign n46630 = n10259 & ~n46629 ;
  assign n46631 = n6757 & n46630 ;
  assign n46632 = n46631 ^ n28954 ^ 1'b0 ;
  assign n46633 = ( n5871 & n15533 ) | ( n5871 & n29022 ) | ( n15533 & n29022 ) ;
  assign n46634 = n46633 ^ n22803 ^ 1'b0 ;
  assign n46635 = ( n9636 & ~n18301 ) | ( n9636 & n21707 ) | ( ~n18301 & n21707 ) ;
  assign n46636 = n46635 ^ n28541 ^ 1'b0 ;
  assign n46637 = n2869 & ~n6904 ;
  assign n46638 = n34219 & n46637 ;
  assign n46639 = n25070 ^ n12972 ^ 1'b0 ;
  assign n46640 = n46638 | n46639 ;
  assign n46641 = n1938 | n46640 ;
  assign n46642 = n14744 ^ x83 ^ 1'b0 ;
  assign n46643 = n31435 & ~n46642 ;
  assign n46644 = n14032 ^ n6533 ^ 1'b0 ;
  assign n46645 = n18854 ^ n15397 ^ 1'b0 ;
  assign n46646 = n31577 & n46645 ;
  assign n46647 = n23378 & n46646 ;
  assign n46648 = n46644 & n46647 ;
  assign n46653 = n30989 ^ n8942 ^ n6971 ;
  assign n46649 = n17960 ^ n8913 ^ n1112 ;
  assign n46650 = ~n12734 & n46649 ;
  assign n46651 = n39969 & ~n46650 ;
  assign n46652 = n1433 & n46651 ;
  assign n46654 = n46653 ^ n46652 ^ 1'b0 ;
  assign n46655 = n32194 ^ n25609 ^ 1'b0 ;
  assign n46656 = n46655 ^ n10477 ^ n10080 ;
  assign n46657 = n23962 | n46656 ;
  assign n46658 = n46657 ^ n5650 ^ 1'b0 ;
  assign n46659 = n7336 & ~n10000 ;
  assign n46660 = n6750 & n46659 ;
  assign n46661 = n35544 ^ n3535 ^ 1'b0 ;
  assign n46662 = n2503 & n46661 ;
  assign n46663 = ( ~n22216 & n46660 ) | ( ~n22216 & n46662 ) | ( n46660 & n46662 ) ;
  assign n46664 = ~n7991 & n43342 ;
  assign n46665 = ( n15673 & n30329 ) | ( n15673 & ~n31169 ) | ( n30329 & ~n31169 ) ;
  assign n46666 = n46061 ^ n19963 ^ 1'b0 ;
  assign n46667 = n14564 & ~n38775 ;
  assign n46670 = n31041 ^ n26363 ^ n10970 ;
  assign n46671 = n46670 ^ n9951 ^ 1'b0 ;
  assign n46668 = n41440 ^ n37505 ^ 1'b0 ;
  assign n46669 = n14452 & n46668 ;
  assign n46672 = n46671 ^ n46669 ^ 1'b0 ;
  assign n46673 = n15428 | n24789 ;
  assign n46674 = n30133 | n46673 ;
  assign n46675 = n2325 | n27453 ;
  assign n46676 = n46675 ^ n33998 ^ 1'b0 ;
  assign n46677 = n45887 ^ n18786 ^ n4858 ;
  assign n46678 = n46677 ^ n8474 ^ n1654 ;
  assign n46679 = ( n3608 & n4319 ) | ( n3608 & ~n17434 ) | ( n4319 & ~n17434 ) ;
  assign n46680 = n12060 & ~n38533 ;
  assign n46681 = n46680 ^ n18944 ^ n3787 ;
  assign n46682 = ( n27850 & n41017 ) | ( n27850 & ~n43656 ) | ( n41017 & ~n43656 ) ;
  assign n46683 = n8537 ^ n7049 ^ n1685 ;
  assign n46684 = n37682 ^ n16395 ^ 1'b0 ;
  assign n46685 = n46683 & n46684 ;
  assign n46686 = ~n29841 & n34001 ;
  assign n46687 = n35906 & n46686 ;
  assign n46688 = n10031 & ~n14920 ;
  assign n46689 = n46688 ^ n11181 ^ 1'b0 ;
  assign n46690 = n37168 ^ n30174 ^ n7487 ;
  assign n46691 = n46690 ^ n6716 ^ 1'b0 ;
  assign n46692 = n6705 | n42895 ;
  assign n46693 = n46692 ^ n7189 ^ n2436 ;
  assign n46694 = n2028 | n25574 ;
  assign n46695 = n29029 & n46694 ;
  assign n46696 = n12669 ^ n310 ^ 1'b0 ;
  assign n46697 = n6033 | n46696 ;
  assign n46698 = n46697 ^ n18538 ^ n2868 ;
  assign n46699 = n46698 ^ n547 ^ 1'b0 ;
  assign n46700 = n12063 ^ n11075 ^ 1'b0 ;
  assign n46701 = n3074 & ~n15389 ;
  assign n46702 = ( ~n11332 & n17066 ) | ( ~n11332 & n46233 ) | ( n17066 & n46233 ) ;
  assign n46703 = n42809 ^ n3701 ^ 1'b0 ;
  assign n46704 = ~n46702 & n46703 ;
  assign n46705 = n11720 & n37954 ;
  assign n46706 = n46705 ^ n19473 ^ 1'b0 ;
  assign n46708 = n40115 ^ n11568 ^ n5556 ;
  assign n46707 = n23637 ^ n20640 ^ 1'b0 ;
  assign n46709 = n46708 ^ n46707 ^ 1'b0 ;
  assign n46710 = n46709 ^ n6136 ^ 1'b0 ;
  assign n46711 = n20591 ^ n11750 ^ n7836 ;
  assign n46712 = ( n4461 & ~n4505 ) | ( n4461 & n46711 ) | ( ~n4505 & n46711 ) ;
  assign n46713 = n43183 ^ n19648 ^ n787 ;
  assign n46714 = n9708 ^ n6805 ^ 1'b0 ;
  assign n46715 = n46714 ^ n20765 ^ n5480 ;
  assign n46716 = n12069 & ~n14395 ;
  assign n46717 = ~n25550 & n46716 ;
  assign n46718 = n46717 ^ n42589 ^ n26043 ;
  assign n46719 = n46718 ^ n25839 ^ n3502 ;
  assign n46720 = n33878 ^ n3703 ^ 1'b0 ;
  assign n46721 = n5946 | n46720 ;
  assign n46722 = n7235 & ~n46721 ;
  assign n46723 = n46722 ^ n38091 ^ 1'b0 ;
  assign n46724 = n8586 | n33141 ;
  assign n46725 = n30796 & ~n46724 ;
  assign n46726 = ( n13061 & n32539 ) | ( n13061 & ~n45280 ) | ( n32539 & ~n45280 ) ;
  assign n46727 = n17673 ^ n17407 ^ n4739 ;
  assign n46728 = ( n7293 & n9863 ) | ( n7293 & n31480 ) | ( n9863 & n31480 ) ;
  assign n46729 = n12666 & n13623 ;
  assign n46730 = ( ~n4264 & n8762 ) | ( ~n4264 & n10885 ) | ( n8762 & n10885 ) ;
  assign n46731 = n1216 & ~n46730 ;
  assign n46732 = ( ~n9174 & n22161 ) | ( ~n9174 & n30308 ) | ( n22161 & n30308 ) ;
  assign n46733 = ( n4509 & n25561 ) | ( n4509 & ~n46732 ) | ( n25561 & ~n46732 ) ;
  assign n46734 = n30960 & ~n46733 ;
  assign n46735 = ( n1409 & n11675 ) | ( n1409 & ~n17431 ) | ( n11675 & ~n17431 ) ;
  assign n46736 = n24320 ^ n3000 ^ 1'b0 ;
  assign n46737 = ~n46735 & n46736 ;
  assign n46738 = n1889 | n11701 ;
  assign n46739 = n2071 & ~n46738 ;
  assign n46740 = n34791 ^ n6267 ^ 1'b0 ;
  assign n46741 = ~n36730 & n46740 ;
  assign n46742 = ( n16015 & ~n35502 ) | ( n16015 & n46741 ) | ( ~n35502 & n46741 ) ;
  assign n46743 = n39948 ^ n428 ^ 1'b0 ;
  assign n46744 = n46743 ^ n36070 ^ n23953 ;
  assign n46745 = ( n9812 & n10589 ) | ( n9812 & ~n15055 ) | ( n10589 & ~n15055 ) ;
  assign n46746 = n27428 ^ n13548 ^ 1'b0 ;
  assign n46747 = n3746 | n46746 ;
  assign n46748 = n33357 & ~n46747 ;
  assign n46749 = n23437 & n46748 ;
  assign n46751 = n11488 ^ n11219 ^ 1'b0 ;
  assign n46752 = n16148 & n46751 ;
  assign n46750 = n14975 | n18570 ;
  assign n46753 = n46752 ^ n46750 ^ 1'b0 ;
  assign n46754 = ( n17808 & ~n46749 ) | ( n17808 & n46753 ) | ( ~n46749 & n46753 ) ;
  assign n46755 = n9921 & n19634 ;
  assign n46756 = ~n40687 & n43812 ;
  assign n46757 = n10259 & ~n14195 ;
  assign n46758 = n46757 ^ n28203 ^ n4068 ;
  assign n46759 = n4467 | n46758 ;
  assign n46760 = n46759 ^ n8438 ^ 1'b0 ;
  assign n46761 = n16026 ^ n15304 ^ 1'b0 ;
  assign n46762 = n46761 ^ n34722 ^ 1'b0 ;
  assign n46763 = n3931 & ~n46762 ;
  assign n46767 = n32235 ^ n18773 ^ n14205 ;
  assign n46764 = n31480 ^ n15875 ^ 1'b0 ;
  assign n46765 = ~n18773 & n46764 ;
  assign n46766 = ( n3524 & n22864 ) | ( n3524 & ~n46765 ) | ( n22864 & ~n46765 ) ;
  assign n46768 = n46767 ^ n46766 ^ n1888 ;
  assign n46769 = n38703 ^ n19762 ^ n4430 ;
  assign n46770 = n46769 ^ n26414 ^ n12984 ;
  assign n46772 = n15634 ^ n9924 ^ 1'b0 ;
  assign n46773 = ~n16479 & n46772 ;
  assign n46771 = n37786 & n40583 ;
  assign n46774 = n46773 ^ n46771 ^ 1'b0 ;
  assign n46775 = n46774 ^ n6703 ^ n3794 ;
  assign n46776 = n10796 ^ n6562 ^ 1'b0 ;
  assign n46777 = ~n23027 & n46776 ;
  assign n46778 = n46777 ^ n37917 ^ 1'b0 ;
  assign n46779 = n46778 ^ n5770 ^ n1517 ;
  assign n46780 = ( ~x5 & n22306 ) | ( ~x5 & n39767 ) | ( n22306 & n39767 ) ;
  assign n46781 = ~n11285 & n44151 ;
  assign n46782 = n46781 ^ n23840 ^ 1'b0 ;
  assign n46783 = ~n19545 & n28980 ;
  assign n46784 = n17267 ^ n9690 ^ 1'b0 ;
  assign n46785 = n1406 | n46784 ;
  assign n46786 = ~n5981 & n9818 ;
  assign n46787 = ~n25886 & n33045 ;
  assign n46788 = n40172 ^ n29289 ^ n1839 ;
  assign n46789 = n46788 ^ n26016 ^ n4828 ;
  assign n46790 = n46789 ^ n12159 ^ 1'b0 ;
  assign n46791 = n46790 ^ n45879 ^ n22141 ;
  assign n46792 = n13345 | n42372 ;
  assign n46796 = n14704 | n28150 ;
  assign n46797 = n46796 ^ n46217 ^ 1'b0 ;
  assign n46793 = ~n7449 & n11139 ;
  assign n46794 = n23716 & n46793 ;
  assign n46795 = n46794 ^ n24065 ^ n368 ;
  assign n46798 = n46797 ^ n46795 ^ n14842 ;
  assign n46799 = n16283 & n40694 ;
  assign n46800 = n15975 ^ n3583 ^ n716 ;
  assign n46801 = ( ~n17862 & n33542 ) | ( ~n17862 & n46800 ) | ( n33542 & n46800 ) ;
  assign n46802 = n41786 ^ n33348 ^ n23115 ;
  assign n46803 = n24751 & n31526 ;
  assign n46804 = n41173 ^ n19656 ^ n15730 ;
  assign n46805 = n46804 ^ n12313 ^ 1'b0 ;
  assign n46806 = n15460 ^ n12414 ^ 1'b0 ;
  assign n46807 = n37849 | n46806 ;
  assign n46808 = ( n21000 & ~n24999 ) | ( n21000 & n46807 ) | ( ~n24999 & n46807 ) ;
  assign n46809 = ~n33705 & n46808 ;
  assign n46810 = n14653 | n46558 ;
  assign n46811 = n46809 & ~n46810 ;
  assign n46812 = n7733 & ~n11564 ;
  assign n46813 = ( ~n19038 & n26293 ) | ( ~n19038 & n43674 ) | ( n26293 & n43674 ) ;
  assign n46814 = n46813 ^ n4705 ^ 1'b0 ;
  assign n46815 = n37581 ^ n3375 ^ 1'b0 ;
  assign n46816 = n14614 | n42286 ;
  assign n46817 = n46816 ^ n256 ^ 1'b0 ;
  assign n46818 = n17249 ^ n11676 ^ n4549 ;
  assign n46819 = n46818 ^ n39314 ^ n17999 ;
  assign n46820 = n8893 & ~n17275 ;
  assign n46821 = n15469 & ~n46820 ;
  assign n46822 = n40331 ^ n8431 ^ 1'b0 ;
  assign n46823 = n36058 & n46822 ;
  assign n46824 = n41503 ^ n33760 ^ 1'b0 ;
  assign n46825 = n4499 | n46824 ;
  assign n46826 = ( n19030 & ~n25921 ) | ( n19030 & n46825 ) | ( ~n25921 & n46825 ) ;
  assign n46827 = n46826 ^ n20550 ^ n17399 ;
  assign n46828 = n11251 & ~n12747 ;
  assign n46829 = ~n3856 & n46828 ;
  assign n46830 = n20540 ^ n10331 ^ 1'b0 ;
  assign n46832 = n45477 ^ n17201 ^ 1'b0 ;
  assign n46833 = n24787 & ~n46832 ;
  assign n46831 = n9316 & n22206 ;
  assign n46834 = n46833 ^ n46831 ^ 1'b0 ;
  assign n46835 = n46834 ^ n38769 ^ n23941 ;
  assign n46836 = n6901 & n29359 ;
  assign n46837 = n42706 & n46836 ;
  assign n46838 = n30724 & ~n46837 ;
  assign n46839 = n46838 ^ n28461 ^ 1'b0 ;
  assign n46840 = n12409 & ~n16732 ;
  assign n46841 = n46840 ^ n19645 ^ 1'b0 ;
  assign n46842 = n26259 ^ n19553 ^ 1'b0 ;
  assign n46843 = ( n22753 & n36954 ) | ( n22753 & n46842 ) | ( n36954 & n46842 ) ;
  assign n46844 = n9239 | n46843 ;
  assign n46845 = n46841 | n46844 ;
  assign n46846 = n6075 & ~n29922 ;
  assign n46847 = n46846 ^ n41511 ^ 1'b0 ;
  assign n46851 = n1730 & n10559 ;
  assign n46852 = ~n8681 & n46851 ;
  assign n46848 = n11627 & ~n29105 ;
  assign n46849 = n32130 & n46848 ;
  assign n46850 = n46849 ^ n16663 ^ n10404 ;
  assign n46853 = n46852 ^ n46850 ^ n21551 ;
  assign n46854 = n9673 | n20471 ;
  assign n46857 = n5040 ^ n3655 ^ n1947 ;
  assign n46855 = n26956 ^ n16518 ^ n14529 ;
  assign n46856 = ( ~n28770 & n40750 ) | ( ~n28770 & n46855 ) | ( n40750 & n46855 ) ;
  assign n46858 = n46857 ^ n46856 ^ n42646 ;
  assign n46859 = n15084 | n23695 ;
  assign n46860 = n15340 & ~n46859 ;
  assign n46861 = n46860 ^ n14239 ^ 1'b0 ;
  assign n46862 = ( n18810 & n25985 ) | ( n18810 & n46861 ) | ( n25985 & n46861 ) ;
  assign n46863 = n34851 ^ n7508 ^ n3336 ;
  assign n46864 = ( n8332 & n21500 ) | ( n8332 & ~n30176 ) | ( n21500 & ~n30176 ) ;
  assign n46865 = n4461 | n46864 ;
  assign n46866 = n46863 & ~n46865 ;
  assign n46867 = n1923 & n10941 ;
  assign n46868 = n26745 ^ n22840 ^ 1'b0 ;
  assign n46869 = ~n21741 & n46868 ;
  assign n46871 = n25598 ^ n20468 ^ n2773 ;
  assign n46872 = ( ~n13642 & n38877 ) | ( ~n13642 & n46871 ) | ( n38877 & n46871 ) ;
  assign n46873 = n46872 ^ n15821 ^ 1'b0 ;
  assign n46870 = ( ~n12900 & n17836 ) | ( ~n12900 & n33547 ) | ( n17836 & n33547 ) ;
  assign n46874 = n46873 ^ n46870 ^ 1'b0 ;
  assign n46875 = n46874 ^ n22016 ^ n16743 ;
  assign n46876 = n46875 ^ n34329 ^ n7537 ;
  assign n46877 = ( n27751 & n41091 ) | ( n27751 & n42875 ) | ( n41091 & n42875 ) ;
  assign n46879 = n14704 ^ n5191 ^ 1'b0 ;
  assign n46878 = ( n874 & n5529 ) | ( n874 & n12406 ) | ( n5529 & n12406 ) ;
  assign n46880 = n46879 ^ n46878 ^ 1'b0 ;
  assign n46881 = n36078 ^ n31276 ^ 1'b0 ;
  assign n46882 = n3032 | n20252 ;
  assign n46883 = n12736 & ~n15101 ;
  assign n46884 = n46883 ^ n15443 ^ 1'b0 ;
  assign n46885 = n38605 | n46884 ;
  assign n46886 = n46885 ^ n18143 ^ 1'b0 ;
  assign n46887 = n26737 & n39599 ;
  assign n46888 = n46887 ^ n42665 ^ 1'b0 ;
  assign n46889 = n29807 ^ n11675 ^ 1'b0 ;
  assign n46890 = n1795 & n46889 ;
  assign n46891 = ~n18844 & n46890 ;
  assign n46892 = n1771 | n30720 ;
  assign n46893 = n46892 ^ n35021 ^ 1'b0 ;
  assign n46894 = n3719 & ~n13719 ;
  assign n46895 = ( ~n791 & n29039 ) | ( ~n791 & n46894 ) | ( n29039 & n46894 ) ;
  assign n46896 = n43155 ^ n27572 ^ 1'b0 ;
  assign n46897 = ( n5372 & ~n18886 ) | ( n5372 & n32089 ) | ( ~n18886 & n32089 ) ;
  assign n46898 = n18625 ^ n9890 ^ n1538 ;
  assign n46899 = ( ~n2287 & n15100 ) | ( ~n2287 & n23580 ) | ( n15100 & n23580 ) ;
  assign n46900 = n15985 | n46899 ;
  assign n46901 = n46900 ^ n11131 ^ 1'b0 ;
  assign n46902 = n19326 ^ n18700 ^ n3843 ;
  assign n46903 = n30690 & ~n46902 ;
  assign n46904 = n46901 & n46903 ;
  assign n46905 = n46898 & ~n46904 ;
  assign n46906 = n14240 & ~n30720 ;
  assign n46907 = n46906 ^ n20447 ^ 1'b0 ;
  assign n46908 = n14945 ^ n14774 ^ 1'b0 ;
  assign n46909 = n24979 & n46908 ;
  assign n46910 = ( n3214 & n12384 ) | ( n3214 & ~n18298 ) | ( n12384 & ~n18298 ) ;
  assign n46911 = n10506 | n46910 ;
  assign n46912 = n46909 | n46911 ;
  assign n46913 = n30998 ^ n15688 ^ n12886 ;
  assign n46916 = ( n8982 & ~n21445 ) | ( n8982 & n26917 ) | ( ~n21445 & n26917 ) ;
  assign n46914 = n561 & n17926 ;
  assign n46915 = ~n21423 & n46914 ;
  assign n46917 = n46916 ^ n46915 ^ 1'b0 ;
  assign n46918 = ( n16185 & ~n20351 ) | ( n16185 & n46917 ) | ( ~n20351 & n46917 ) ;
  assign n46919 = n7962 | n33347 ;
  assign n46920 = ( n2828 & n15678 ) | ( n2828 & ~n46919 ) | ( n15678 & ~n46919 ) ;
  assign n46921 = ~n1660 & n25793 ;
  assign n46922 = n46921 ^ n9855 ^ 1'b0 ;
  assign n46923 = ~n5850 & n39772 ;
  assign n46924 = n46923 ^ n34477 ^ 1'b0 ;
  assign n46925 = n29157 | n45661 ;
  assign n46926 = n46924 | n46925 ;
  assign n46927 = n46926 ^ n3699 ^ 1'b0 ;
  assign n46928 = n7551 & ~n46927 ;
  assign n46929 = ( ~n20088 & n46922 ) | ( ~n20088 & n46928 ) | ( n46922 & n46928 ) ;
  assign n46930 = n41170 ^ n38784 ^ 1'b0 ;
  assign n46931 = n1521 & ~n46930 ;
  assign n46933 = n16720 | n21625 ;
  assign n46934 = n25960 & ~n46933 ;
  assign n46932 = n33195 ^ n20413 ^ 1'b0 ;
  assign n46935 = n46934 ^ n46932 ^ 1'b0 ;
  assign n46936 = n4989 ^ n2985 ^ 1'b0 ;
  assign n46937 = n6390 & ~n15699 ;
  assign n46938 = n22321 & n46937 ;
  assign n46939 = n46938 ^ n40029 ^ 1'b0 ;
  assign n46940 = n43331 ^ n24288 ^ n4132 ;
  assign n46941 = n46940 ^ n11016 ^ 1'b0 ;
  assign n46942 = n19853 ^ n11969 ^ n8549 ;
  assign n46943 = n46942 ^ n18992 ^ n11689 ;
  assign n46944 = ( n2122 & n21945 ) | ( n2122 & ~n38615 ) | ( n21945 & ~n38615 ) ;
  assign n46948 = n15052 ^ n13824 ^ n12887 ;
  assign n46947 = ( n8179 & n12334 ) | ( n8179 & ~n26097 ) | ( n12334 & ~n26097 ) ;
  assign n46945 = ~n5223 & n16700 ;
  assign n46946 = n12460 & n46945 ;
  assign n46949 = n46948 ^ n46947 ^ n46946 ;
  assign n46950 = n46949 ^ n44724 ^ n41981 ;
  assign n46951 = x118 & n4832 ;
  assign n46952 = n46951 ^ n8854 ^ 1'b0 ;
  assign n46953 = n24284 & n35634 ;
  assign n46954 = n31410 ^ n5408 ^ 1'b0 ;
  assign n46955 = n37274 & ~n46954 ;
  assign n46956 = n46955 ^ n36467 ^ 1'b0 ;
  assign n46957 = n1114 & ~n20204 ;
  assign n46958 = n46957 ^ n38252 ^ 1'b0 ;
  assign n46959 = n39847 ^ n7073 ^ 1'b0 ;
  assign n46960 = n46959 ^ n35405 ^ n5290 ;
  assign n46961 = n46958 & ~n46960 ;
  assign n46962 = n25487 ^ n3826 ^ 1'b0 ;
  assign n46963 = ( n16110 & n17384 ) | ( n16110 & n46962 ) | ( n17384 & n46962 ) ;
  assign n46964 = n46870 ^ n40926 ^ 1'b0 ;
  assign n46965 = n46964 ^ n38149 ^ n3569 ;
  assign n46967 = n42968 ^ n11178 ^ 1'b0 ;
  assign n46966 = ( n3715 & n7460 ) | ( n3715 & n14093 ) | ( n7460 & n14093 ) ;
  assign n46968 = n46967 ^ n46966 ^ n12223 ;
  assign n46969 = n2321 & n32404 ;
  assign n46970 = n46969 ^ n9752 ^ 1'b0 ;
  assign n46971 = n2897 | n46970 ;
  assign n46972 = n32763 & ~n46971 ;
  assign n46973 = n20787 ^ n7743 ^ 1'b0 ;
  assign n46974 = n27738 & ~n46973 ;
  assign n46975 = n10463 | n35427 ;
  assign n46976 = n46974 | n46975 ;
  assign n46977 = ( n1477 & ~n2702 ) | ( n1477 & n12552 ) | ( ~n2702 & n12552 ) ;
  assign n46978 = n17874 & n46977 ;
  assign n46979 = n32195 & n46978 ;
  assign n46980 = n43304 ^ n30502 ^ n19859 ;
  assign n46981 = x218 | n46980 ;
  assign n46982 = n46728 ^ n28198 ^ n11242 ;
  assign n46983 = n45287 ^ n15112 ^ n13000 ;
  assign n46984 = ~n13704 & n46752 ;
  assign n46985 = ( n12563 & ~n27325 ) | ( n12563 & n46984 ) | ( ~n27325 & n46984 ) ;
  assign n46986 = ~n4080 & n10690 ;
  assign n46987 = ~n761 & n46986 ;
  assign n46988 = n21166 & ~n46987 ;
  assign n46989 = n5344 & n15807 ;
  assign n46990 = n21282 & ~n23055 ;
  assign n46991 = n46990 ^ n38832 ^ 1'b0 ;
  assign n46992 = ( n8760 & n15130 ) | ( n8760 & n18308 ) | ( n15130 & n18308 ) ;
  assign n46993 = n1623 & ~n25247 ;
  assign n46994 = n46993 ^ n3843 ^ 1'b0 ;
  assign n46995 = n46994 ^ n14076 ^ 1'b0 ;
  assign n46996 = n21787 & n46995 ;
  assign n46997 = n4590 & n46996 ;
  assign n46998 = ( ~n34165 & n46992 ) | ( ~n34165 & n46997 ) | ( n46992 & n46997 ) ;
  assign n46999 = n29007 ^ n9789 ^ n3147 ;
  assign n47000 = n24344 ^ n20360 ^ n8729 ;
  assign n47001 = ( n2927 & n10971 ) | ( n2927 & n26432 ) | ( n10971 & n26432 ) ;
  assign n47002 = ( n40149 & n47000 ) | ( n40149 & ~n47001 ) | ( n47000 & ~n47001 ) ;
  assign n47003 = ( ~n2206 & n10615 ) | ( ~n2206 & n25686 ) | ( n10615 & n25686 ) ;
  assign n47004 = n20839 & ~n47003 ;
  assign n47005 = ~n18070 & n47004 ;
  assign n47006 = n5693 ^ n3052 ^ 1'b0 ;
  assign n47007 = n26138 & ~n47006 ;
  assign n47008 = ~n2536 & n32544 ;
  assign n47009 = n31107 ^ n26391 ^ 1'b0 ;
  assign n47010 = n9495 & n47009 ;
  assign n47011 = n39247 ^ n4276 ^ 1'b0 ;
  assign n47012 = ( n7554 & n13400 ) | ( n7554 & n15348 ) | ( n13400 & n15348 ) ;
  assign n47013 = n47012 ^ n36860 ^ n595 ;
  assign n47014 = ( ~n461 & n11604 ) | ( ~n461 & n30366 ) | ( n11604 & n30366 ) ;
  assign n47015 = n47014 ^ n42890 ^ n34041 ;
  assign n47016 = n45554 ^ n39515 ^ 1'b0 ;
  assign n47017 = ( ~n26934 & n31871 ) | ( ~n26934 & n46175 ) | ( n31871 & n46175 ) ;
  assign n47018 = ~n4478 & n23589 ;
  assign n47019 = n25314 ^ n13118 ^ 1'b0 ;
  assign n47020 = ~n25028 & n47019 ;
  assign n47021 = ~n1345 & n16974 ;
  assign n47022 = n47021 ^ n23740 ^ 1'b0 ;
  assign n47023 = n43753 ^ n9896 ^ 1'b0 ;
  assign n47024 = n47022 & n47023 ;
  assign n47025 = ~n18617 & n24876 ;
  assign n47028 = n1336 & ~n26937 ;
  assign n47026 = ( n6014 & ~n22741 ) | ( n6014 & n26492 ) | ( ~n22741 & n26492 ) ;
  assign n47027 = n47026 ^ n2177 ^ 1'b0 ;
  assign n47029 = n47028 ^ n47027 ^ 1'b0 ;
  assign n47030 = n14319 | n16258 ;
  assign n47031 = n23454 & ~n47030 ;
  assign n47032 = n47031 ^ n40041 ^ n10186 ;
  assign n47033 = n6809 ^ n6789 ^ 1'b0 ;
  assign n47034 = n47033 ^ n22315 ^ 1'b0 ;
  assign n47035 = n25939 | n47034 ;
  assign n47036 = ( n702 & n9371 ) | ( n702 & ~n10420 ) | ( n9371 & ~n10420 ) ;
  assign n47037 = n47036 ^ n574 ^ x185 ;
  assign n47038 = ~n12536 & n47037 ;
  assign n47039 = ~n43399 & n47038 ;
  assign n47040 = n14842 ^ n6777 ^ 1'b0 ;
  assign n47041 = ~n20053 & n47040 ;
  assign n47042 = n36397 ^ n30302 ^ 1'b0 ;
  assign n47043 = ~n1850 & n47042 ;
  assign n47044 = n8859 & n34003 ;
  assign n47045 = n25105 ^ n24768 ^ n6216 ;
  assign n47046 = ( n8315 & n43970 ) | ( n8315 & n47045 ) | ( n43970 & n47045 ) ;
  assign n47047 = ( n27141 & n32951 ) | ( n27141 & ~n43514 ) | ( n32951 & ~n43514 ) ;
  assign n47048 = n15084 ^ n8405 ^ n6577 ;
  assign n47049 = n28916 ^ n8701 ^ 1'b0 ;
  assign n47050 = ( n3499 & ~n12005 ) | ( n3499 & n13375 ) | ( ~n12005 & n13375 ) ;
  assign n47051 = ( n35062 & n36178 ) | ( n35062 & n47050 ) | ( n36178 & n47050 ) ;
  assign n47052 = n3402 | n7234 ;
  assign n47053 = n47052 ^ n13197 ^ 1'b0 ;
  assign n47054 = x180 & n29873 ;
  assign n47055 = n14325 & ~n16831 ;
  assign n47056 = n34341 & n40221 ;
  assign n47057 = n47055 & ~n47056 ;
  assign n47058 = n47057 ^ n38003 ^ 1'b0 ;
  assign n47059 = ( n17256 & n19756 ) | ( n17256 & ~n43572 ) | ( n19756 & ~n43572 ) ;
  assign n47060 = ( n11708 & ~n13223 ) | ( n11708 & n34149 ) | ( ~n13223 & n34149 ) ;
  assign n47061 = n29227 ^ n28811 ^ 1'b0 ;
  assign n47062 = ~n6705 & n47061 ;
  assign n47063 = ( n24337 & n47060 ) | ( n24337 & n47062 ) | ( n47060 & n47062 ) ;
  assign n47064 = ( n4430 & ~n8352 ) | ( n4430 & n18556 ) | ( ~n8352 & n18556 ) ;
  assign n47065 = n16959 ^ n15766 ^ n5244 ;
  assign n47066 = ~n47064 & n47065 ;
  assign n47067 = n24391 & n47066 ;
  assign n47068 = n8229 ^ n2965 ^ 1'b0 ;
  assign n47069 = n47067 | n47068 ;
  assign n47070 = n24826 ^ n21947 ^ n15125 ;
  assign n47071 = n19152 ^ n15572 ^ 1'b0 ;
  assign n47072 = n47070 & n47071 ;
  assign n47073 = n47069 | n47072 ;
  assign n47074 = n10678 | n12897 ;
  assign n47075 = n1378 & ~n6825 ;
  assign n47076 = n35954 ^ n15510 ^ n8779 ;
  assign n47077 = n47076 ^ n42918 ^ 1'b0 ;
  assign n47078 = n13903 & n47077 ;
  assign n47079 = n3341 & n47078 ;
  assign n47080 = ( x9 & n27404 ) | ( x9 & n28295 ) | ( n27404 & n28295 ) ;
  assign n47081 = n47080 ^ n7533 ^ n1959 ;
  assign n47082 = n23505 ^ n7927 ^ 1'b0 ;
  assign n47083 = ( n6320 & n47081 ) | ( n6320 & ~n47082 ) | ( n47081 & ~n47082 ) ;
  assign n47084 = n41004 ^ n26211 ^ n9820 ;
  assign n47085 = n17911 & n45061 ;
  assign n47087 = n35092 ^ n27153 ^ 1'b0 ;
  assign n47086 = n38935 ^ n34059 ^ 1'b0 ;
  assign n47088 = n47087 ^ n47086 ^ n28414 ;
  assign n47089 = n24594 ^ n21963 ^ 1'b0 ;
  assign n47090 = ( n1952 & n7241 ) | ( n1952 & n30876 ) | ( n7241 & n30876 ) ;
  assign n47091 = n13364 | n31731 ;
  assign n47092 = ~n47090 & n47091 ;
  assign n47093 = n47092 ^ n17675 ^ 1'b0 ;
  assign n47094 = n333 & ~n1418 ;
  assign n47095 = n1276 & n47094 ;
  assign n47096 = n47095 ^ n3052 ^ 1'b0 ;
  assign n47097 = n13264 ^ n1884 ^ 1'b0 ;
  assign n47098 = n47096 & n47097 ;
  assign n47099 = ( n3896 & n10680 ) | ( n3896 & ~n33864 ) | ( n10680 & ~n33864 ) ;
  assign n47100 = n37929 ^ n14086 ^ 1'b0 ;
  assign n47101 = n36320 & n39748 ;
  assign n47102 = ~n11807 & n47101 ;
  assign n47103 = n15600 | n47102 ;
  assign n47104 = n25661 ^ n23817 ^ 1'b0 ;
  assign n47105 = ~n8293 & n9655 ;
  assign n47106 = ~n21049 & n47105 ;
  assign n47107 = n35926 & n36030 ;
  assign n47108 = n47107 ^ n13042 ^ 1'b0 ;
  assign n47109 = n41165 ^ n11235 ^ 1'b0 ;
  assign n47110 = ~n10553 & n47109 ;
  assign n47111 = ~n44909 & n47110 ;
  assign n47112 = ( ~n1786 & n12502 ) | ( ~n1786 & n12709 ) | ( n12502 & n12709 ) ;
  assign n47113 = ( ~n46125 & n46289 ) | ( ~n46125 & n47112 ) | ( n46289 & n47112 ) ;
  assign n47114 = n30886 ^ n25415 ^ n20952 ;
  assign n47115 = n7916 & ~n10018 ;
  assign n47116 = n47115 ^ n39587 ^ 1'b0 ;
  assign n47117 = n46315 & ~n47116 ;
  assign n47118 = ~n21619 & n32024 ;
  assign n47119 = ( n13039 & n16484 ) | ( n13039 & n24931 ) | ( n16484 & n24931 ) ;
  assign n47120 = n40020 & n47119 ;
  assign n47121 = n47120 ^ n30339 ^ 1'b0 ;
  assign n47122 = ~n15320 & n16377 ;
  assign n47123 = n47122 ^ n30082 ^ 1'b0 ;
  assign n47124 = ~n33307 & n47123 ;
  assign n47125 = n16164 & ~n17010 ;
  assign n47126 = n20647 ^ n18210 ^ 1'b0 ;
  assign n47127 = n28742 ^ n18543 ^ 1'b0 ;
  assign n47128 = n47126 & n47127 ;
  assign n47129 = n736 & n6582 ;
  assign n47130 = n47129 ^ n14652 ^ 1'b0 ;
  assign n47131 = n47130 ^ n13237 ^ 1'b0 ;
  assign n47132 = ( n46341 & ~n46435 ) | ( n46341 & n47131 ) | ( ~n46435 & n47131 ) ;
  assign n47133 = n37816 ^ n13109 ^ 1'b0 ;
  assign n47134 = n19314 & ~n47133 ;
  assign n47135 = n47134 ^ n18863 ^ 1'b0 ;
  assign n47136 = n9134 ^ n4731 ^ n3987 ;
  assign n47137 = n27700 ^ n20453 ^ n9142 ;
  assign n47138 = ( n34027 & ~n47136 ) | ( n34027 & n47137 ) | ( ~n47136 & n47137 ) ;
  assign n47139 = ( n10537 & n20936 ) | ( n10537 & ~n32642 ) | ( n20936 & ~n32642 ) ;
  assign n47140 = ( n7447 & ~n47138 ) | ( n7447 & n47139 ) | ( ~n47138 & n47139 ) ;
  assign n47141 = n11777 ^ n10698 ^ 1'b0 ;
  assign n47142 = n32005 & ~n47141 ;
  assign n47143 = n8724 & n17872 ;
  assign n47144 = ~n33493 & n47143 ;
  assign n47145 = n16064 & ~n47144 ;
  assign n47146 = n2338 ^ n1194 ^ 1'b0 ;
  assign n47147 = ~n13040 & n47146 ;
  assign n47148 = ~n2522 & n5715 ;
  assign n47149 = n47148 ^ n7474 ^ 1'b0 ;
  assign n47150 = n47149 ^ n26572 ^ n8620 ;
  assign n47151 = ( ~n11118 & n23129 ) | ( ~n11118 & n47150 ) | ( n23129 & n47150 ) ;
  assign n47152 = n47151 ^ n32286 ^ 1'b0 ;
  assign n47153 = n21523 & n46280 ;
  assign n47154 = n17340 | n24238 ;
  assign n47155 = n47154 ^ n26631 ^ 1'b0 ;
  assign n47156 = n47155 ^ n43243 ^ 1'b0 ;
  assign n47157 = n47153 | n47156 ;
  assign n47158 = ~n6437 & n39363 ;
  assign n47159 = ~n12084 & n47158 ;
  assign n47160 = n11984 ^ n6207 ^ 1'b0 ;
  assign n47161 = n12972 & ~n47160 ;
  assign n47162 = n47161 ^ n6776 ^ 1'b0 ;
  assign n47164 = n16517 ^ n6869 ^ 1'b0 ;
  assign n47165 = n47164 ^ n33844 ^ n31030 ;
  assign n47166 = n47165 ^ n5673 ^ 1'b0 ;
  assign n47163 = ~x215 & n7404 ;
  assign n47167 = n47166 ^ n47163 ^ 1'b0 ;
  assign n47168 = n25999 ^ n15224 ^ n2739 ;
  assign n47170 = ( n9130 & n23667 ) | ( n9130 & n29472 ) | ( n23667 & n29472 ) ;
  assign n47169 = n28759 & n29941 ;
  assign n47171 = n47170 ^ n47169 ^ n31141 ;
  assign n47172 = n40891 ^ n26112 ^ n7921 ;
  assign n47173 = n7021 & ~n19290 ;
  assign n47174 = ~n28639 & n47173 ;
  assign n47175 = ~n45219 & n45322 ;
  assign n47176 = n45132 & n47175 ;
  assign n47177 = n6978 | n29365 ;
  assign n47178 = n47177 ^ n6719 ^ 1'b0 ;
  assign n47179 = n32277 ^ n6904 ^ n2630 ;
  assign n47180 = ~n2836 & n47179 ;
  assign n47181 = n23786 ^ n10650 ^ 1'b0 ;
  assign n47182 = n14763 & ~n47181 ;
  assign n47183 = n8376 ^ n1764 ^ 1'b0 ;
  assign n47184 = n13660 & ~n47183 ;
  assign n47185 = ( n33487 & n47182 ) | ( n33487 & n47184 ) | ( n47182 & n47184 ) ;
  assign n47186 = n7220 & ~n29365 ;
  assign n47187 = ~n8326 & n47186 ;
  assign n47188 = ( n7714 & n40569 ) | ( n7714 & n47187 ) | ( n40569 & n47187 ) ;
  assign n47189 = n4644 ^ n1465 ^ 1'b0 ;
  assign n47190 = n7814 & n47189 ;
  assign n47191 = ( n2097 & n2423 ) | ( n2097 & n24414 ) | ( n2423 & n24414 ) ;
  assign n47192 = x106 & n44115 ;
  assign n47193 = n19657 ^ n8632 ^ 1'b0 ;
  assign n47194 = n40924 ^ n2914 ^ 1'b0 ;
  assign n47195 = n1287 & n47194 ;
  assign n47196 = n1251 & n47195 ;
  assign n47197 = n38621 ^ n4350 ^ 1'b0 ;
  assign n47198 = n47196 & n47197 ;
  assign n47200 = n1056 | n31559 ;
  assign n47201 = ( n3162 & ~n19231 ) | ( n3162 & n47200 ) | ( ~n19231 & n47200 ) ;
  assign n47199 = ( n3311 & ~n6288 ) | ( n3311 & n14768 ) | ( ~n6288 & n14768 ) ;
  assign n47202 = n47201 ^ n47199 ^ n21406 ;
  assign n47203 = ~n5770 & n47202 ;
  assign n47204 = n19995 & n47203 ;
  assign n47205 = n15623 ^ n3212 ^ 1'b0 ;
  assign n47206 = ~n43270 & n47205 ;
  assign n47207 = n41157 & ~n47206 ;
  assign n47208 = n3762 & ~n13535 ;
  assign n47209 = n12997 ^ n12590 ^ 1'b0 ;
  assign n47210 = ~n34584 & n45485 ;
  assign n47211 = n14382 ^ n7101 ^ n2853 ;
  assign n47212 = n8299 ^ n335 ^ 1'b0 ;
  assign n47213 = n15830 | n28481 ;
  assign n47214 = n47212 | n47213 ;
  assign n47215 = n7491 & n37713 ;
  assign n47216 = n11409 | n13231 ;
  assign n47217 = n9454 ^ n3584 ^ 1'b0 ;
  assign n47218 = n19381 & n47217 ;
  assign n47219 = n31563 ^ n28547 ^ n7191 ;
  assign n47220 = n23579 & n23674 ;
  assign n47221 = n47220 ^ n31023 ^ 1'b0 ;
  assign n47222 = n5645 | n30572 ;
  assign n47223 = n47221 | n47222 ;
  assign n47224 = ( n10234 & n17420 ) | ( n10234 & n47223 ) | ( n17420 & n47223 ) ;
  assign n47225 = n27463 | n30174 ;
  assign n47226 = n9820 ^ n6819 ^ 1'b0 ;
  assign n47227 = n1312 & ~n14393 ;
  assign n47228 = ( n43812 & n47226 ) | ( n43812 & n47227 ) | ( n47226 & n47227 ) ;
  assign n47229 = n16503 ^ n1986 ^ 1'b0 ;
  assign n47230 = ~n26143 & n47229 ;
  assign n47231 = n47069 ^ n12413 ^ 1'b0 ;
  assign n47232 = n25976 & n47231 ;
  assign n47233 = ~n1641 & n10524 ;
  assign n47234 = ~n5168 & n47233 ;
  assign n47235 = ( n11113 & ~n24668 ) | ( n11113 & n47234 ) | ( ~n24668 & n47234 ) ;
  assign n47236 = n20924 | n47235 ;
  assign n47237 = n19532 | n47236 ;
  assign n47238 = n33084 ^ n17216 ^ 1'b0 ;
  assign n47239 = ~n13645 & n36999 ;
  assign n47240 = ~n7920 & n47239 ;
  assign n47241 = n39168 & n42897 ;
  assign n47242 = ~n29273 & n47241 ;
  assign n47243 = n15098 ^ n11229 ^ n4357 ;
  assign n47244 = ( n26209 & n34926 ) | ( n26209 & n47243 ) | ( n34926 & n47243 ) ;
  assign n47245 = n3783 & ~n22899 ;
  assign n47246 = n47245 ^ n16504 ^ 1'b0 ;
  assign n47247 = ~n9225 & n35013 ;
  assign n47248 = ~n47246 & n47247 ;
  assign n47249 = ( n2272 & n23741 ) | ( n2272 & ~n47248 ) | ( n23741 & ~n47248 ) ;
  assign n47250 = n21635 | n38717 ;
  assign n47251 = n27037 ^ n8702 ^ 1'b0 ;
  assign n47252 = n11126 | n47251 ;
  assign n47253 = n47252 ^ n6266 ^ 1'b0 ;
  assign n47254 = n34022 & ~n47253 ;
  assign n47255 = ( ~n3759 & n23045 ) | ( ~n3759 & n33043 ) | ( n23045 & n33043 ) ;
  assign n47256 = n22968 ^ n15610 ^ 1'b0 ;
  assign n47257 = n47255 | n47256 ;
  assign n47258 = n22332 ^ n21594 ^ 1'b0 ;
  assign n47259 = n4605 & ~n20462 ;
  assign n47260 = x10 & n47259 ;
  assign n47261 = n47260 ^ n1655 ^ 1'b0 ;
  assign n47262 = n6793 | n25852 ;
  assign n47263 = n47262 ^ n36317 ^ 1'b0 ;
  assign n47264 = ~n47261 & n47263 ;
  assign n47265 = n37762 ^ n37606 ^ 1'b0 ;
  assign n47266 = ~n22394 & n24084 ;
  assign n47267 = n2628 & ~n42557 ;
  assign n47268 = ( ~n6132 & n7600 ) | ( ~n6132 & n9492 ) | ( n7600 & n9492 ) ;
  assign n47269 = ( n18582 & n22677 ) | ( n18582 & ~n44685 ) | ( n22677 & ~n44685 ) ;
  assign n47270 = n31350 ^ n17332 ^ n471 ;
  assign n47271 = n9492 & n10482 ;
  assign n47272 = ~n47270 & n47271 ;
  assign n47273 = n19518 ^ n9790 ^ 1'b0 ;
  assign n47274 = n12682 | n47273 ;
  assign n47275 = n47274 ^ n14955 ^ 1'b0 ;
  assign n47279 = n11307 | n12469 ;
  assign n47276 = n6895 & ~n40659 ;
  assign n47277 = n47276 ^ n12515 ^ 1'b0 ;
  assign n47278 = n47277 ^ n13870 ^ n12955 ;
  assign n47280 = n47279 ^ n47278 ^ n35979 ;
  assign n47281 = n32485 & ~n47280 ;
  assign n47282 = n47281 ^ n24635 ^ 1'b0 ;
  assign n47284 = n12610 | n19127 ;
  assign n47285 = n47284 ^ n8935 ^ 1'b0 ;
  assign n47286 = n47285 ^ n16369 ^ 1'b0 ;
  assign n47283 = n6660 & ~n25262 ;
  assign n47287 = n47286 ^ n47283 ^ 1'b0 ;
  assign n47288 = n44733 ^ n16156 ^ 1'b0 ;
  assign n47289 = n22925 ^ n7714 ^ n5561 ;
  assign n47290 = n45248 & ~n47289 ;
  assign n47291 = ( ~n18389 & n33012 ) | ( ~n18389 & n39928 ) | ( n33012 & n39928 ) ;
  assign n47292 = n40048 & ~n41257 ;
  assign n47297 = n9751 | n16053 ;
  assign n47298 = n38761 & ~n47297 ;
  assign n47294 = n24296 ^ n6908 ^ 1'b0 ;
  assign n47295 = n36392 & ~n47294 ;
  assign n47296 = n20717 | n47295 ;
  assign n47293 = n24508 ^ n21875 ^ 1'b0 ;
  assign n47299 = n47298 ^ n47296 ^ n47293 ;
  assign n47300 = n11301 | n12874 ;
  assign n47301 = n47300 ^ n31254 ^ 1'b0 ;
  assign n47302 = n46505 ^ n1092 ^ 1'b0 ;
  assign n47303 = n6647 & n47302 ;
  assign n47304 = n24604 ^ n16325 ^ 1'b0 ;
  assign n47305 = n39871 | n46089 ;
  assign n47306 = n47305 ^ n44973 ^ 1'b0 ;
  assign n47307 = ( n6525 & ~n31154 ) | ( n6525 & n35676 ) | ( ~n31154 & n35676 ) ;
  assign n47308 = n34350 ^ n13028 ^ 1'b0 ;
  assign n47312 = n43284 ^ n6258 ^ 1'b0 ;
  assign n47310 = n15980 ^ n12849 ^ 1'b0 ;
  assign n47311 = ~n26543 & n47310 ;
  assign n47309 = ( n11289 & ~n31633 ) | ( n11289 & n33745 ) | ( ~n31633 & n33745 ) ;
  assign n47313 = n47312 ^ n47311 ^ n47309 ;
  assign n47314 = ( n6162 & ~n26466 ) | ( n6162 & n41384 ) | ( ~n26466 & n41384 ) ;
  assign n47315 = n38386 ^ n16153 ^ 1'b0 ;
  assign n47316 = n19999 | n47315 ;
  assign n47317 = n20546 & n47316 ;
  assign n47318 = n5127 | n36837 ;
  assign n47319 = n5710 & ~n15949 ;
  assign n47320 = n7157 & n47319 ;
  assign n47321 = n26781 ^ n16557 ^ n9848 ;
  assign n47322 = ~n22148 & n47321 ;
  assign n47323 = n31347 & n47322 ;
  assign n47324 = ~n8996 & n25429 ;
  assign n47325 = ( n13502 & n27288 ) | ( n13502 & n47324 ) | ( n27288 & n47324 ) ;
  assign n47326 = n34414 ^ n18549 ^ 1'b0 ;
  assign n47327 = n31010 | n47326 ;
  assign n47328 = n47327 ^ n34093 ^ n16054 ;
  assign n47329 = ( ~n7744 & n7918 ) | ( ~n7744 & n38988 ) | ( n7918 & n38988 ) ;
  assign n47330 = n40431 ^ n25013 ^ n11049 ;
  assign n47335 = n23823 | n36647 ;
  assign n47331 = n27263 ^ n6465 ^ n2124 ;
  assign n47332 = n47331 ^ n38596 ^ n1398 ;
  assign n47333 = n9519 & ~n10173 ;
  assign n47334 = n47332 & n47333 ;
  assign n47336 = n47335 ^ n47334 ^ n24931 ;
  assign n47337 = n47065 ^ n23466 ^ 1'b0 ;
  assign n47338 = ~n12093 & n47337 ;
  assign n47339 = n1944 & n30081 ;
  assign n47340 = n35908 & n47339 ;
  assign n47341 = n9411 | n46938 ;
  assign n47342 = n40432 ^ n38228 ^ n1873 ;
  assign n47345 = n23488 ^ n23070 ^ 1'b0 ;
  assign n47346 = ~n9878 & n47345 ;
  assign n47343 = n44089 ^ n23890 ^ n6329 ;
  assign n47344 = n47343 ^ n31886 ^ n12198 ;
  assign n47347 = n47346 ^ n47344 ^ n26805 ;
  assign n47348 = ( n6681 & ~n28014 ) | ( n6681 & n33249 ) | ( ~n28014 & n33249 ) ;
  assign n47349 = n47348 ^ n33189 ^ n30591 ;
  assign n47350 = ( n9618 & n23076 ) | ( n9618 & n47349 ) | ( n23076 & n47349 ) ;
  assign n47351 = n8694 ^ n3953 ^ n2824 ;
  assign n47352 = ( n22314 & ~n27928 ) | ( n22314 & n47351 ) | ( ~n27928 & n47351 ) ;
  assign n47353 = n11597 & n47352 ;
  assign n47354 = ~n28032 & n47353 ;
  assign n47355 = ~n4763 & n7634 ;
  assign n47356 = n47355 ^ n38107 ^ 1'b0 ;
  assign n47357 = n30488 ^ n706 ^ 1'b0 ;
  assign n47358 = n12576 & n21190 ;
  assign n47359 = n47358 ^ n2191 ^ 1'b0 ;
  assign n47360 = n8045 ^ n7386 ^ 1'b0 ;
  assign n47361 = n6930 & n47360 ;
  assign n47362 = n8243 ^ n5107 ^ 1'b0 ;
  assign n47363 = n47361 & n47362 ;
  assign n47364 = ~n4679 & n47363 ;
  assign n47365 = n37020 ^ n9552 ^ 1'b0 ;
  assign n47366 = ( n27700 & n29825 ) | ( n27700 & ~n29940 ) | ( n29825 & ~n29940 ) ;
  assign n47367 = n22919 & ~n37452 ;
  assign n47368 = ~n38046 & n47367 ;
  assign n47369 = n6669 & ~n8073 ;
  assign n47370 = n47369 ^ n26725 ^ 1'b0 ;
  assign n47371 = n5930 & ~n36483 ;
  assign n47372 = ~n31588 & n47371 ;
  assign n47373 = ( n47368 & n47370 ) | ( n47368 & n47372 ) | ( n47370 & n47372 ) ;
  assign n47374 = n47373 ^ n35710 ^ n11493 ;
  assign n47375 = ~n4854 & n41203 ;
  assign n47376 = n23279 & n47375 ;
  assign n47377 = n47376 ^ n16402 ^ n11273 ;
  assign n47378 = n37493 ^ n27799 ^ n12129 ;
  assign n47379 = n47378 ^ n15304 ^ n487 ;
  assign n47380 = ~n9670 & n32257 ;
  assign n47381 = ~n4941 & n47380 ;
  assign n47382 = n22101 ^ n4386 ^ 1'b0 ;
  assign n47383 = n12560 & ~n30122 ;
  assign n47384 = ~n47382 & n47383 ;
  assign n47385 = n33763 ^ n9626 ^ 1'b0 ;
  assign n47386 = n19150 | n47385 ;
  assign n47387 = n36326 ^ n10573 ^ 1'b0 ;
  assign n47388 = ~n47386 & n47387 ;
  assign n47390 = n9136 & ~n37071 ;
  assign n47389 = n9188 | n14835 ;
  assign n47391 = n47390 ^ n47389 ^ 1'b0 ;
  assign n47392 = ( n8332 & n17068 ) | ( n8332 & n40998 ) | ( n17068 & n40998 ) ;
  assign n47393 = ~n9265 & n13206 ;
  assign n47394 = n47393 ^ n30329 ^ 1'b0 ;
  assign n47396 = ( x158 & n3579 ) | ( x158 & n16143 ) | ( n3579 & n16143 ) ;
  assign n47395 = ( n6329 & ~n13961 ) | ( n6329 & n19116 ) | ( ~n13961 & n19116 ) ;
  assign n47397 = n47396 ^ n47395 ^ n7478 ;
  assign n47398 = n45079 ^ n20640 ^ 1'b0 ;
  assign n47399 = ( n21421 & n43126 ) | ( n21421 & ~n47398 ) | ( n43126 & ~n47398 ) ;
  assign n47400 = ( n47394 & n47397 ) | ( n47394 & n47399 ) | ( n47397 & n47399 ) ;
  assign n47401 = n37700 ^ n14543 ^ 1'b0 ;
  assign n47402 = n47401 ^ n40970 ^ n17362 ;
  assign n47403 = n26060 ^ n8660 ^ 1'b0 ;
  assign n47404 = ( ~n19299 & n28408 ) | ( ~n19299 & n35944 ) | ( n28408 & n35944 ) ;
  assign n47405 = n19752 & n36693 ;
  assign n47406 = n45239 ^ n35838 ^ n7952 ;
  assign n47407 = n47406 ^ n31529 ^ 1'b0 ;
  assign n47408 = ( n8468 & ~n47405 ) | ( n8468 & n47407 ) | ( ~n47405 & n47407 ) ;
  assign n47409 = ~n4437 & n47408 ;
  assign n47410 = n26629 ^ n10098 ^ 1'b0 ;
  assign n47411 = n10791 ^ n9685 ^ 1'b0 ;
  assign n47412 = n15597 ^ n2093 ^ 1'b0 ;
  assign n47413 = n26865 & n47412 ;
  assign n47414 = ~n41460 & n47413 ;
  assign n47415 = n47411 & n47414 ;
  assign n47416 = n12638 ^ n4868 ^ 1'b0 ;
  assign n47417 = n19960 | n47416 ;
  assign n47418 = n47417 ^ n10670 ^ 1'b0 ;
  assign n47419 = ~n10057 & n21803 ;
  assign n47420 = n47419 ^ n35097 ^ 1'b0 ;
  assign n47421 = n23210 & n27016 ;
  assign n47422 = n4444 | n15921 ;
  assign n47423 = n28500 ^ n14695 ^ n10373 ;
  assign n47424 = ( ~n41503 & n44123 ) | ( ~n41503 & n47423 ) | ( n44123 & n47423 ) ;
  assign n47425 = ( n3318 & ~n17548 ) | ( n3318 & n19218 ) | ( ~n17548 & n19218 ) ;
  assign n47426 = n417 & n4813 ;
  assign n47427 = n43560 & n46881 ;
  assign n47428 = ~n47426 & n47427 ;
  assign n47429 = ~n26228 & n47150 ;
  assign n47430 = ( n4529 & n36616 ) | ( n4529 & n36620 ) | ( n36616 & n36620 ) ;
  assign n47431 = n40084 | n47430 ;
  assign n47432 = n3411 ^ n1198 ^ 1'b0 ;
  assign n47433 = n5522 | n47432 ;
  assign n47434 = n47433 ^ n2982 ^ 1'b0 ;
  assign n47435 = n16068 | n47434 ;
  assign n47436 = n27729 & ~n47435 ;
  assign n47437 = n35521 ^ n15497 ^ 1'b0 ;
  assign n47438 = ( n41239 & n46003 ) | ( n41239 & ~n47437 ) | ( n46003 & ~n47437 ) ;
  assign n47439 = ( n15301 & ~n27457 ) | ( n15301 & n37820 ) | ( ~n27457 & n37820 ) ;
  assign n47440 = n30235 & n32112 ;
  assign n47441 = n31168 & n47440 ;
  assign n47442 = n8320 | n11958 ;
  assign n47443 = n47442 ^ n40052 ^ 1'b0 ;
  assign n47444 = n28032 & ~n47443 ;
  assign n47445 = ~n31624 & n47444 ;
  assign n47446 = x234 & n21796 ;
  assign n47447 = n47446 ^ n25846 ^ 1'b0 ;
  assign n47448 = ( n4857 & n25470 ) | ( n4857 & n47372 ) | ( n25470 & n47372 ) ;
  assign n47449 = n13722 ^ n2362 ^ 1'b0 ;
  assign n47450 = n40173 ^ n29443 ^ n1171 ;
  assign n47451 = n47450 ^ n21253 ^ 1'b0 ;
  assign n47452 = n47451 ^ n26882 ^ n8307 ;
  assign n47453 = n26228 ^ n15154 ^ 1'b0 ;
  assign n47454 = n12604 & n42941 ;
  assign n47455 = ~n47453 & n47454 ;
  assign n47456 = ( ~n8180 & n39681 ) | ( ~n8180 & n47455 ) | ( n39681 & n47455 ) ;
  assign n47457 = n2697 | n10356 ;
  assign n47458 = n47457 ^ n6982 ^ 1'b0 ;
  assign n47459 = n3135 & n47458 ;
  assign n47460 = n47459 ^ n6006 ^ 1'b0 ;
  assign n47463 = n5236 | n17844 ;
  assign n47462 = n11738 & ~n18922 ;
  assign n47464 = n47463 ^ n47462 ^ 1'b0 ;
  assign n47465 = n4758 & ~n47464 ;
  assign n47466 = n44089 & n47465 ;
  assign n47461 = n22006 | n27115 ;
  assign n47467 = n47466 ^ n47461 ^ 1'b0 ;
  assign n47468 = ( n1934 & n3724 ) | ( n1934 & ~n13216 ) | ( n3724 & ~n13216 ) ;
  assign n47469 = ( ~n13163 & n13687 ) | ( ~n13163 & n47468 ) | ( n13687 & n47468 ) ;
  assign n47470 = n4639 | n47469 ;
  assign n47471 = n25349 & ~n44409 ;
  assign n47472 = ~n47470 & n47471 ;
  assign n47473 = n10238 & ~n37609 ;
  assign n47474 = ( n17997 & n31683 ) | ( n17997 & ~n38882 ) | ( n31683 & ~n38882 ) ;
  assign n47475 = ( n14613 & n21589 ) | ( n14613 & n34571 ) | ( n21589 & n34571 ) ;
  assign n47476 = n38148 ^ n18385 ^ 1'b0 ;
  assign n47478 = ( n4970 & n21855 ) | ( n4970 & n24185 ) | ( n21855 & n24185 ) ;
  assign n47479 = n47478 ^ n13244 ^ 1'b0 ;
  assign n47480 = n11143 & ~n14283 ;
  assign n47481 = n47480 ^ x218 ^ 1'b0 ;
  assign n47482 = n47479 | n47481 ;
  assign n47477 = n39070 ^ n13997 ^ 1'b0 ;
  assign n47483 = n47482 ^ n47477 ^ n38006 ;
  assign n47484 = n41610 ^ n36991 ^ n25992 ;
  assign n47488 = n7679 ^ n3600 ^ 1'b0 ;
  assign n47489 = n11604 | n47488 ;
  assign n47485 = n34805 ^ n19700 ^ 1'b0 ;
  assign n47486 = n36974 | n47485 ;
  assign n47487 = n3647 & ~n47486 ;
  assign n47490 = n47489 ^ n47487 ^ 1'b0 ;
  assign n47491 = n637 & n13657 ;
  assign n47492 = ~n1430 & n47491 ;
  assign n47493 = n7090 | n44289 ;
  assign n47494 = n38350 ^ n31298 ^ 1'b0 ;
  assign n47495 = ~n45481 & n47494 ;
  assign n47496 = n10667 | n25768 ;
  assign n47497 = n22012 & ~n47496 ;
  assign n47499 = ( n4338 & ~n33171 ) | ( n4338 & n34624 ) | ( ~n33171 & n34624 ) ;
  assign n47498 = n11889 & ~n39773 ;
  assign n47500 = n47499 ^ n47498 ^ 1'b0 ;
  assign n47501 = n47500 ^ n17196 ^ 1'b0 ;
  assign n47502 = n47501 ^ n24833 ^ n18503 ;
  assign n47503 = n12546 | n44080 ;
  assign n47504 = ( n25447 & n27140 ) | ( n25447 & ~n35149 ) | ( n27140 & ~n35149 ) ;
  assign n47505 = n36427 | n47504 ;
  assign n47506 = ~n8136 & n25995 ;
  assign n47507 = ~n43516 & n47506 ;
  assign n47508 = x183 | n11428 ;
  assign n47509 = n4389 & ~n47508 ;
  assign n47510 = n47507 & n47509 ;
  assign n47511 = n37141 ^ n27689 ^ 1'b0 ;
  assign n47512 = n24853 | n47511 ;
  assign n47513 = n3746 | n35984 ;
  assign n47514 = n47513 ^ n25648 ^ 1'b0 ;
  assign n47515 = n43995 ^ n39699 ^ 1'b0 ;
  assign n47517 = n17295 | n26781 ;
  assign n47518 = n11476 | n47517 ;
  assign n47519 = n26263 & n47518 ;
  assign n47520 = n9259 & n47519 ;
  assign n47516 = n35297 & ~n41024 ;
  assign n47521 = n47520 ^ n47516 ^ 1'b0 ;
  assign n47522 = ( n8380 & ~n26621 ) | ( n8380 & n47521 ) | ( ~n26621 & n47521 ) ;
  assign n47523 = n8419 | n18596 ;
  assign n47524 = n1475 | n2702 ;
  assign n47525 = n46758 ^ n15766 ^ n10288 ;
  assign n47526 = n9248 ^ n6333 ^ 1'b0 ;
  assign n47527 = ~n14418 & n47526 ;
  assign n47528 = ( ~n11962 & n16098 ) | ( ~n11962 & n47527 ) | ( n16098 & n47527 ) ;
  assign n47529 = ( n14073 & ~n44639 ) | ( n14073 & n47528 ) | ( ~n44639 & n47528 ) ;
  assign n47530 = ~n47525 & n47529 ;
  assign n47531 = n40814 | n47530 ;
  assign n47532 = n31049 | n47531 ;
  assign n47533 = n35081 & n35287 ;
  assign n47534 = n2961 & n28484 ;
  assign n47535 = ( ~n11677 & n21331 ) | ( ~n11677 & n27077 ) | ( n21331 & n27077 ) ;
  assign n47536 = n47535 ^ n733 ^ 1'b0 ;
  assign n47537 = n28304 & n47536 ;
  assign n47538 = n4283 | n7448 ;
  assign n47539 = n28036 ^ n27999 ^ 1'b0 ;
  assign n47540 = n28414 & n47539 ;
  assign n47541 = ( n20614 & n47538 ) | ( n20614 & ~n47540 ) | ( n47538 & ~n47540 ) ;
  assign n47542 = n7515 ^ n688 ^ 1'b0 ;
  assign n47543 = n22479 | n40444 ;
  assign n47544 = n42792 & ~n47543 ;
  assign n47545 = n47544 ^ n44125 ^ 1'b0 ;
  assign n47546 = ( n4700 & ~n15300 ) | ( n4700 & n19796 ) | ( ~n15300 & n19796 ) ;
  assign n47547 = n36334 | n45359 ;
  assign n47548 = n47547 ^ n16051 ^ 1'b0 ;
  assign n47549 = n36050 ^ n29941 ^ 1'b0 ;
  assign n47550 = n35710 ^ n24227 ^ n7555 ;
  assign n47551 = n47550 ^ n47037 ^ n24049 ;
  assign n47552 = n20894 & n25419 ;
  assign n47553 = n10840 & ~n13814 ;
  assign n47554 = n4100 & ~n47553 ;
  assign n47555 = n47554 ^ n2274 ^ 1'b0 ;
  assign n47556 = n416 | n47555 ;
  assign n47559 = n46990 ^ n4810 ^ 1'b0 ;
  assign n47557 = ~n5507 & n22035 ;
  assign n47558 = n47557 ^ n10531 ^ 1'b0 ;
  assign n47560 = n47559 ^ n47558 ^ n2582 ;
  assign n47561 = ( n17364 & n19436 ) | ( n17364 & ~n24248 ) | ( n19436 & ~n24248 ) ;
  assign n47562 = n40408 & ~n47561 ;
  assign n47563 = n47562 ^ n26262 ^ 1'b0 ;
  assign n47564 = n17898 ^ n14926 ^ 1'b0 ;
  assign n47565 = n3876 | n40889 ;
  assign n47566 = n47565 ^ n10660 ^ 1'b0 ;
  assign n47567 = n5135 | n7615 ;
  assign n47568 = n47567 ^ n21206 ^ n10127 ;
  assign n47569 = ( n24749 & n39607 ) | ( n24749 & ~n45414 ) | ( n39607 & ~n45414 ) ;
  assign n47570 = ~n2731 & n14134 ;
  assign n47571 = n37367 ^ n6216 ^ 1'b0 ;
  assign n47572 = n47570 & n47571 ;
  assign n47573 = n8085 & ~n46074 ;
  assign n47574 = n36458 ^ n31510 ^ n24097 ;
  assign n47575 = n3690 | n9615 ;
  assign n47576 = n47574 | n47575 ;
  assign n47577 = n47576 ^ n3885 ^ 1'b0 ;
  assign n47578 = n24760 & ~n34434 ;
  assign n47579 = n18934 | n47578 ;
  assign n47580 = n47579 ^ n34751 ^ 1'b0 ;
  assign n47581 = n44041 ^ n35312 ^ 1'b0 ;
  assign n47584 = ~n3918 & n6955 ;
  assign n47582 = n17875 | n33215 ;
  assign n47583 = n18242 | n47582 ;
  assign n47585 = n47584 ^ n47583 ^ n43298 ;
  assign n47586 = n12161 ^ n8810 ^ 1'b0 ;
  assign n47587 = n39451 ^ n25175 ^ 1'b0 ;
  assign n47588 = n13907 & n47587 ;
  assign n47589 = n47588 ^ n14235 ^ n11389 ;
  assign n47590 = ( n2399 & n26959 ) | ( n2399 & ~n35994 ) | ( n26959 & ~n35994 ) ;
  assign n47591 = ~n39637 & n47590 ;
  assign n47592 = ~n23314 & n37427 ;
  assign n47593 = n47592 ^ n1221 ^ 1'b0 ;
  assign n47594 = n16812 & n17461 ;
  assign n47595 = ~n11938 & n47594 ;
  assign n47596 = n6743 & ~n47595 ;
  assign n47597 = n47596 ^ n17244 ^ 1'b0 ;
  assign n47598 = n38977 ^ n35316 ^ 1'b0 ;
  assign n47599 = n26687 | n41882 ;
  assign n47600 = n20797 ^ n16854 ^ n1822 ;
  assign n47601 = n8375 & ~n47600 ;
  assign n47602 = n3460 & n5313 ;
  assign n47603 = n47602 ^ n19421 ^ n15238 ;
  assign n47604 = n47603 ^ n23378 ^ 1'b0 ;
  assign n47605 = ( ~n3787 & n18156 ) | ( ~n3787 & n20231 ) | ( n18156 & n20231 ) ;
  assign n47606 = n47605 ^ n4851 ^ 1'b0 ;
  assign n47607 = n39387 ^ n16658 ^ 1'b0 ;
  assign n47608 = n33760 & n47607 ;
  assign n47609 = n4605 & n16701 ;
  assign n47610 = n47609 ^ n8487 ^ 1'b0 ;
  assign n47612 = n42352 ^ n40179 ^ 1'b0 ;
  assign n47611 = n36686 & ~n47351 ;
  assign n47613 = n47612 ^ n47611 ^ 1'b0 ;
  assign n47614 = n33662 ^ n19262 ^ n10628 ;
  assign n47615 = n1903 | n47614 ;
  assign n47616 = n4677 & n47615 ;
  assign n47617 = n28457 ^ n18467 ^ x163 ;
  assign n47618 = n41926 ^ n4522 ^ 1'b0 ;
  assign n47619 = ( n6501 & n19674 ) | ( n6501 & n47618 ) | ( n19674 & n47618 ) ;
  assign n47620 = ( n15414 & n25155 ) | ( n15414 & ~n41749 ) | ( n25155 & ~n41749 ) ;
  assign n47621 = n47620 ^ n41393 ^ n20069 ;
  assign n47622 = ~n7889 & n27086 ;
  assign n47623 = n47478 & n47622 ;
  assign n47624 = ( n11743 & n13380 ) | ( n11743 & n34148 ) | ( n13380 & n34148 ) ;
  assign n47625 = ~n11724 & n34762 ;
  assign n47626 = ~n47624 & n47625 ;
  assign n47627 = n38666 ^ n14816 ^ 1'b0 ;
  assign n47628 = ( n11354 & n21497 ) | ( n11354 & ~n47627 ) | ( n21497 & ~n47627 ) ;
  assign n47629 = ( n8437 & n20942 ) | ( n8437 & ~n47628 ) | ( n20942 & ~n47628 ) ;
  assign n47630 = n27004 ^ n1876 ^ n333 ;
  assign n47631 = ( ~n3390 & n8403 ) | ( ~n3390 & n47630 ) | ( n8403 & n47630 ) ;
  assign n47632 = n31570 ^ n16410 ^ n13788 ;
  assign n47633 = n11590 ^ n3073 ^ 1'b0 ;
  assign n47634 = n12173 | n41327 ;
  assign n47635 = n47634 ^ n20821 ^ 1'b0 ;
  assign n47636 = ~n13859 & n24710 ;
  assign n47637 = ~n28148 & n28325 ;
  assign n47638 = n47636 & n47637 ;
  assign n47639 = n14077 ^ n11013 ^ 1'b0 ;
  assign n47640 = ~n43867 & n47639 ;
  assign n47641 = n47640 ^ n27993 ^ 1'b0 ;
  assign n47642 = n33483 ^ n12300 ^ 1'b0 ;
  assign n47643 = n756 | n47642 ;
  assign n47644 = n17219 | n42800 ;
  assign n47646 = n25338 ^ n6479 ^ 1'b0 ;
  assign n47645 = n33821 ^ n26984 ^ 1'b0 ;
  assign n47647 = n47646 ^ n47645 ^ n37779 ;
  assign n47648 = n2261 & ~n10520 ;
  assign n47649 = n47648 ^ n5102 ^ 1'b0 ;
  assign n47650 = ( n13776 & ~n14834 ) | ( n13776 & n47649 ) | ( ~n14834 & n47649 ) ;
  assign n47651 = n22855 ^ n10222 ^ n8657 ;
  assign n47652 = n47651 ^ n5239 ^ n1163 ;
  assign n47653 = ( n30431 & n36905 ) | ( n30431 & n39594 ) | ( n36905 & n39594 ) ;
  assign n47654 = ~n31808 & n35058 ;
  assign n47655 = n47654 ^ n4150 ^ 1'b0 ;
  assign n47656 = n24138 & n32148 ;
  assign n47657 = ~n18256 & n47656 ;
  assign n47658 = ( ~n4592 & n5779 ) | ( ~n4592 & n10896 ) | ( n5779 & n10896 ) ;
  assign n47659 = n25781 & n47658 ;
  assign n47660 = n44726 & n47659 ;
  assign n47661 = n4749 | n34585 ;
  assign n47662 = n47661 ^ n11706 ^ 1'b0 ;
  assign n47663 = n35215 ^ n34676 ^ n18335 ;
  assign n47664 = n1105 ^ n317 ^ 1'b0 ;
  assign n47665 = ~n11632 & n47664 ;
  assign n47666 = ( n24526 & n27429 ) | ( n24526 & n47665 ) | ( n27429 & n47665 ) ;
  assign n47667 = n21134 & n22060 ;
  assign n47668 = n2337 & ~n9106 ;
  assign n47669 = n47668 ^ n22332 ^ 1'b0 ;
  assign n47670 = ( ~n9131 & n47667 ) | ( ~n9131 & n47669 ) | ( n47667 & n47669 ) ;
  assign n47671 = ( n37301 & ~n45138 ) | ( n37301 & n47670 ) | ( ~n45138 & n47670 ) ;
  assign n47672 = n5953 & ~n9190 ;
  assign n47673 = n47672 ^ n26404 ^ 1'b0 ;
  assign n47674 = n47673 ^ n14927 ^ 1'b0 ;
  assign n47675 = ~n4310 & n7503 ;
  assign n47676 = n39834 & ~n47675 ;
  assign n47677 = n47676 ^ n18193 ^ 1'b0 ;
  assign n47679 = ( n13077 & n15091 ) | ( n13077 & n15109 ) | ( n15091 & n15109 ) ;
  assign n47678 = n4286 & n17722 ;
  assign n47680 = n47679 ^ n47678 ^ 1'b0 ;
  assign n47681 = n29777 ^ n25974 ^ 1'b0 ;
  assign n47682 = n36878 & ~n47681 ;
  assign n47683 = n1959 & ~n15007 ;
  assign n47684 = n47683 ^ n6462 ^ 1'b0 ;
  assign n47685 = n47684 ^ n39263 ^ 1'b0 ;
  assign n47686 = n39971 ^ n22847 ^ 1'b0 ;
  assign n47687 = ( n5965 & n21863 ) | ( n5965 & n47686 ) | ( n21863 & n47686 ) ;
  assign n47688 = ( n1885 & n28601 ) | ( n1885 & ~n33067 ) | ( n28601 & ~n33067 ) ;
  assign n47689 = n1098 & ~n26689 ;
  assign n47690 = n47689 ^ n2928 ^ 1'b0 ;
  assign n47692 = n16733 & ~n18197 ;
  assign n47693 = n9978 | n19290 ;
  assign n47694 = n47692 | n47693 ;
  assign n47691 = n32946 & n45385 ;
  assign n47695 = n47694 ^ n47691 ^ 1'b0 ;
  assign n47696 = n14952 | n16104 ;
  assign n47697 = n18717 & ~n34156 ;
  assign n47699 = n1570 | n15752 ;
  assign n47700 = n3218 & ~n47699 ;
  assign n47701 = ( n355 & n18349 ) | ( n355 & n47700 ) | ( n18349 & n47700 ) ;
  assign n47702 = n42341 | n47701 ;
  assign n47698 = n14594 | n31316 ;
  assign n47703 = n47702 ^ n47698 ^ 1'b0 ;
  assign n47704 = ~n14233 & n23240 ;
  assign n47705 = n47704 ^ n38653 ^ n33308 ;
  assign n47708 = n18770 & ~n25018 ;
  assign n47706 = n13056 ^ n11407 ^ 1'b0 ;
  assign n47707 = n25567 & ~n47706 ;
  assign n47709 = n47708 ^ n47707 ^ n42009 ;
  assign n47710 = ( n4223 & n13035 ) | ( n4223 & n42926 ) | ( n13035 & n42926 ) ;
  assign n47711 = n47710 ^ n3509 ^ n2087 ;
  assign n47712 = n26198 ^ n17549 ^ 1'b0 ;
  assign n47713 = n1331 | n47712 ;
  assign n47714 = n35357 | n47076 ;
  assign n47715 = ( ~n44406 & n47713 ) | ( ~n44406 & n47714 ) | ( n47713 & n47714 ) ;
  assign n47716 = n22878 ^ n7873 ^ 1'b0 ;
  assign n47717 = n26352 | n47716 ;
  assign n47718 = n6252 & n21413 ;
  assign n47719 = n1506 & ~n47718 ;
  assign n47720 = n47719 ^ n33163 ^ 1'b0 ;
  assign n47721 = n47720 ^ n3716 ^ 1'b0 ;
  assign n47722 = n32089 & ~n47721 ;
  assign n47723 = n20630 | n21654 ;
  assign n47724 = n47723 ^ n27141 ^ 1'b0 ;
  assign n47725 = n47724 ^ n38652 ^ 1'b0 ;
  assign n47726 = n1431 | n6344 ;
  assign n47727 = n38546 | n47726 ;
  assign n47728 = ( n25136 & n27621 ) | ( n25136 & n44423 ) | ( n27621 & n44423 ) ;
  assign n47729 = n13291 ^ x85 ^ 1'b0 ;
  assign n47730 = n29986 ^ n12441 ^ 1'b0 ;
  assign n47731 = ( n31226 & n47729 ) | ( n31226 & ~n47730 ) | ( n47729 & ~n47730 ) ;
  assign n47732 = ( ~n4114 & n32984 ) | ( ~n4114 & n39587 ) | ( n32984 & n39587 ) ;
  assign n47733 = n47732 ^ n8346 ^ 1'b0 ;
  assign n47734 = n23089 ^ n20316 ^ 1'b0 ;
  assign n47735 = n8645 | n26928 ;
  assign n47736 = n41745 & ~n43163 ;
  assign n47737 = n13254 & n47736 ;
  assign n47738 = ~n15663 & n44234 ;
  assign n47739 = n9225 & n47738 ;
  assign n47740 = n16734 ^ n8707 ^ 1'b0 ;
  assign n47741 = n18259 & n47740 ;
  assign n47742 = n14137 & n30809 ;
  assign n47743 = n47741 & n47742 ;
  assign n47744 = n47743 ^ n10216 ^ 1'b0 ;
  assign n47745 = n955 & n47744 ;
  assign n47746 = n47745 ^ n35617 ^ 1'b0 ;
  assign n47747 = n15081 & ~n25628 ;
  assign n47748 = ( ~n27012 & n36290 ) | ( ~n27012 & n47747 ) | ( n36290 & n47747 ) ;
  assign n47749 = n47748 ^ n5677 ^ 1'b0 ;
  assign n47750 = n47746 & n47749 ;
  assign n47751 = n23985 ^ n15681 ^ 1'b0 ;
  assign n47752 = ( ~n5689 & n18509 ) | ( ~n5689 & n25717 ) | ( n18509 & n25717 ) ;
  assign n47753 = n47752 ^ n37427 ^ n26233 ;
  assign n47754 = n10257 ^ n8450 ^ n6666 ;
  assign n47758 = n16230 ^ n3315 ^ 1'b0 ;
  assign n47759 = n6826 & n47758 ;
  assign n47755 = ~n8335 & n22613 ;
  assign n47756 = ~n11235 & n47755 ;
  assign n47757 = ( n20424 & ~n30758 ) | ( n20424 & n47756 ) | ( ~n30758 & n47756 ) ;
  assign n47760 = n47759 ^ n47757 ^ n39233 ;
  assign n47761 = ( n9446 & ~n18992 ) | ( n9446 & n21403 ) | ( ~n18992 & n21403 ) ;
  assign n47762 = n33927 ^ n3100 ^ 1'b0 ;
  assign n47763 = n10432 & ~n47762 ;
  assign n47764 = n47763 ^ n15169 ^ 1'b0 ;
  assign n47765 = n22203 & ~n47764 ;
  assign n47766 = n47765 ^ n22026 ^ n21581 ;
  assign n47767 = n45445 ^ n17676 ^ n3202 ;
  assign n47768 = n12433 ^ n8044 ^ n1035 ;
  assign n47769 = n46552 & n47768 ;
  assign n47770 = ~n47767 & n47769 ;
  assign n47771 = n12880 & ~n38963 ;
  assign n47772 = n1403 & n47771 ;
  assign n47773 = n40751 ^ n7563 ^ 1'b0 ;
  assign n47774 = n32092 ^ n11212 ^ n6575 ;
  assign n47775 = n24595 ^ n6672 ^ n4386 ;
  assign n47776 = n25850 | n47775 ;
  assign n47777 = ( n6985 & n11743 ) | ( n6985 & ~n43162 ) | ( n11743 & ~n43162 ) ;
  assign n47778 = n6742 ^ n5663 ^ 1'b0 ;
  assign n47779 = n43371 & n47778 ;
  assign n47780 = ~n9697 & n16858 ;
  assign n47781 = ~n47779 & n47780 ;
  assign n47782 = n20896 ^ n14835 ^ 1'b0 ;
  assign n47783 = n35529 & n47782 ;
  assign n47784 = n46794 ^ n39103 ^ n7049 ;
  assign n47785 = n47784 ^ n4001 ^ 1'b0 ;
  assign n47786 = n22642 ^ n21892 ^ 1'b0 ;
  assign n47787 = ~n43033 & n47786 ;
  assign n47788 = n393 & ~n5251 ;
  assign n47789 = ~n41590 & n47788 ;
  assign n47790 = n4756 ^ n4473 ^ n988 ;
  assign n47791 = n44557 & n47790 ;
  assign n47792 = n22581 ^ n12245 ^ 1'b0 ;
  assign n47793 = n47792 ^ n44398 ^ n38529 ;
  assign n47794 = n16701 & n43784 ;
  assign n47795 = ~n4054 & n47794 ;
  assign n47796 = ( n18349 & n24532 ) | ( n18349 & ~n47795 ) | ( n24532 & ~n47795 ) ;
  assign n47797 = ~n5446 & n32337 ;
  assign n47798 = n47797 ^ n2199 ^ 1'b0 ;
  assign n47799 = n47798 ^ n20050 ^ 1'b0 ;
  assign n47800 = ~n8916 & n45391 ;
  assign n47801 = n47800 ^ n25994 ^ 1'b0 ;
  assign n47802 = n34964 & ~n42585 ;
  assign n47803 = n6242 & ~n40861 ;
  assign n47804 = n47803 ^ n7201 ^ 1'b0 ;
  assign n47805 = ~n7921 & n7927 ;
  assign n47806 = n47805 ^ n5424 ^ 1'b0 ;
  assign n47807 = n19180 | n47806 ;
  assign n47808 = n46377 & ~n47807 ;
  assign n47809 = ~n24813 & n42386 ;
  assign n47810 = ~n2945 & n47809 ;
  assign n47811 = n14319 ^ n6645 ^ 1'b0 ;
  assign n47812 = ( n7294 & n10553 ) | ( n7294 & ~n37406 ) | ( n10553 & ~n37406 ) ;
  assign n47813 = ( n36625 & n47811 ) | ( n36625 & n47812 ) | ( n47811 & n47812 ) ;
  assign n47814 = n47813 ^ n35460 ^ 1'b0 ;
  assign n47815 = ( n3334 & ~n36178 ) | ( n3334 & n47814 ) | ( ~n36178 & n47814 ) ;
  assign n47816 = n33072 ^ n21629 ^ n20715 ;
  assign n47817 = n7688 & ~n35006 ;
  assign n47818 = ( ~n7790 & n32724 ) | ( ~n7790 & n47817 ) | ( n32724 & n47817 ) ;
  assign n47819 = n8235 ^ n4637 ^ 1'b0 ;
  assign n47820 = n43660 ^ n32820 ^ 1'b0 ;
  assign n47821 = n2555 & ~n47820 ;
  assign n47822 = ~n5530 & n11459 ;
  assign n47823 = n23426 & n43468 ;
  assign n47824 = n9455 ^ n3549 ^ n1646 ;
  assign n47825 = n47824 ^ n40136 ^ n31388 ;
  assign n47826 = ~n40999 & n47825 ;
  assign n47827 = n12331 & n47826 ;
  assign n47828 = ~n4652 & n39904 ;
  assign n47829 = ~n10783 & n47828 ;
  assign n47830 = n15061 & ~n47829 ;
  assign n47831 = n47830 ^ n17727 ^ 1'b0 ;
  assign n47832 = n15318 | n47831 ;
  assign n47833 = n47832 ^ n14396 ^ 1'b0 ;
  assign n47834 = n5789 | n28378 ;
  assign n47835 = n11082 & n47834 ;
  assign n47836 = n47835 ^ n20845 ^ 1'b0 ;
  assign n47837 = n47836 ^ n44895 ^ 1'b0 ;
  assign n47838 = n13312 ^ n9319 ^ 1'b0 ;
  assign n47839 = n47838 ^ n37837 ^ n11121 ;
  assign n47840 = n24952 & n47839 ;
  assign n47841 = ~n2520 & n11865 ;
  assign n47842 = ( n41664 & ~n45995 ) | ( n41664 & n47841 ) | ( ~n45995 & n47841 ) ;
  assign n47843 = n307 & ~n27050 ;
  assign n47844 = n5974 & n47843 ;
  assign n47845 = ( n22161 & n39762 ) | ( n22161 & ~n47844 ) | ( n39762 & ~n47844 ) ;
  assign n47846 = ~n33015 & n47382 ;
  assign n47847 = ~n5828 & n35915 ;
  assign n47848 = n47847 ^ n36819 ^ 1'b0 ;
  assign n47849 = ( n12517 & n15925 ) | ( n12517 & n19473 ) | ( n15925 & n19473 ) ;
  assign n47850 = n47849 ^ n44648 ^ n20356 ;
  assign n47851 = ( n6591 & ~n23700 ) | ( n6591 & n27594 ) | ( ~n23700 & n27594 ) ;
  assign n47852 = n20189 & ~n36634 ;
  assign n47853 = n40024 & n47852 ;
  assign n47854 = ( n26627 & n33201 ) | ( n26627 & ~n47853 ) | ( n33201 & ~n47853 ) ;
  assign n47855 = ( n24190 & ~n47851 ) | ( n24190 & n47854 ) | ( ~n47851 & n47854 ) ;
  assign n47856 = ( n813 & n28401 ) | ( n813 & ~n29237 ) | ( n28401 & ~n29237 ) ;
  assign n47857 = n10228 & n34988 ;
  assign n47858 = n31363 ^ n5531 ^ 1'b0 ;
  assign n47859 = ~n8433 & n16287 ;
  assign n47860 = n47859 ^ n24128 ^ 1'b0 ;
  assign n47861 = ~n22175 & n47860 ;
  assign n47862 = n10325 | n23710 ;
  assign n47863 = n26296 | n47862 ;
  assign n47864 = ( ~n4359 & n9287 ) | ( ~n4359 & n41106 ) | ( n9287 & n41106 ) ;
  assign n47865 = n47864 ^ n27372 ^ n8789 ;
  assign n47866 = ( n7978 & n12648 ) | ( n7978 & ~n14144 ) | ( n12648 & ~n14144 ) ;
  assign n47867 = n9107 & ~n32432 ;
  assign n47868 = n27674 ^ n27065 ^ 1'b0 ;
  assign n47869 = n7950 | n47868 ;
  assign n47870 = ( n10448 & n19231 ) | ( n10448 & n47869 ) | ( n19231 & n47869 ) ;
  assign n47871 = n4714 & ~n14443 ;
  assign n47872 = ( n9772 & n32015 ) | ( n9772 & ~n47871 ) | ( n32015 & ~n47871 ) ;
  assign n47873 = n11707 & n15522 ;
  assign n47874 = n8850 | n17433 ;
  assign n47875 = n47874 ^ n19441 ^ 1'b0 ;
  assign n47876 = n32879 & n47875 ;
  assign n47877 = n17689 ^ n14910 ^ 1'b0 ;
  assign n47878 = ~n24261 & n47877 ;
  assign n47879 = n16447 | n26441 ;
  assign n47880 = n47879 ^ n16005 ^ 1'b0 ;
  assign n47881 = ~n2889 & n47880 ;
  assign n47882 = n23010 & n47881 ;
  assign n47883 = n5250 | n41752 ;
  assign n47884 = n4292 & ~n28633 ;
  assign n47885 = n47884 ^ n3534 ^ 1'b0 ;
  assign n47886 = ( n3960 & ~n18424 ) | ( n3960 & n47885 ) | ( ~n18424 & n47885 ) ;
  assign n47887 = n9266 | n30901 ;
  assign n47888 = ( n774 & n22958 ) | ( n774 & ~n47887 ) | ( n22958 & ~n47887 ) ;
  assign n47889 = n534 & n1559 ;
  assign n47890 = n47889 ^ n15868 ^ 1'b0 ;
  assign n47891 = n1385 | n3894 ;
  assign n47892 = ~n10575 & n47891 ;
  assign n47893 = n42246 & n47892 ;
  assign n47894 = ( n45348 & n47890 ) | ( n45348 & ~n47893 ) | ( n47890 & ~n47893 ) ;
  assign n47895 = n11620 & n13147 ;
  assign n47896 = ~n5815 & n47895 ;
  assign n47897 = n47896 ^ n25386 ^ 1'b0 ;
  assign n47898 = n22191 & ~n47897 ;
  assign n47899 = n47898 ^ n16064 ^ n7050 ;
  assign n47900 = n47899 ^ n42030 ^ n15949 ;
  assign n47901 = n33781 ^ n19951 ^ 1'b0 ;
  assign n47902 = ( n3870 & n16895 ) | ( n3870 & ~n24243 ) | ( n16895 & ~n24243 ) ;
  assign n47903 = n47902 ^ n31960 ^ 1'b0 ;
  assign n47904 = n47901 | n47903 ;
  assign n47905 = n11747 & n28759 ;
  assign n47906 = n9252 | n26551 ;
  assign n47907 = n47906 ^ x207 ^ 1'b0 ;
  assign n47908 = n47905 & ~n47907 ;
  assign n47909 = n10080 ^ n6216 ^ 1'b0 ;
  assign n47910 = ~n16316 & n47909 ;
  assign n47911 = n11564 ^ n1961 ^ 1'b0 ;
  assign n47912 = n23343 & ~n32129 ;
  assign n47913 = n47912 ^ n42046 ^ 1'b0 ;
  assign n47914 = n47913 ^ n36977 ^ n3478 ;
  assign n47915 = n15551 ^ n7116 ^ 1'b0 ;
  assign n47916 = n20179 & n47915 ;
  assign n47917 = ~n47914 & n47916 ;
  assign n47918 = n47917 ^ n10989 ^ 1'b0 ;
  assign n47919 = n37041 ^ n34007 ^ n25695 ;
  assign n47920 = n47919 ^ n38855 ^ n2402 ;
  assign n47921 = n39467 ^ n3918 ^ 1'b0 ;
  assign n47922 = n39084 ^ n11535 ^ n10844 ;
  assign n47923 = ( ~x62 & n25156 ) | ( ~x62 & n42356 ) | ( n25156 & n42356 ) ;
  assign n47924 = n47923 ^ n10255 ^ 1'b0 ;
  assign n47925 = n12306 & n18226 ;
  assign n47926 = ~n11829 & n47925 ;
  assign n47927 = ~n20344 & n36164 ;
  assign n47928 = n20842 & n47927 ;
  assign n47929 = n28897 ^ n12953 ^ 1'b0 ;
  assign n47930 = ~n47928 & n47929 ;
  assign n47931 = n25117 ^ x102 ^ 1'b0 ;
  assign n47932 = n17925 ^ n810 ^ 1'b0 ;
  assign n47933 = ~n47931 & n47932 ;
  assign n47934 = n8258 ^ n6216 ^ 1'b0 ;
  assign n47935 = n47934 ^ n34820 ^ 1'b0 ;
  assign n47936 = n7815 | n12536 ;
  assign n47937 = n47936 ^ n9086 ^ 1'b0 ;
  assign n47938 = n9280 & n43273 ;
  assign n47939 = ( n34524 & n47937 ) | ( n34524 & ~n47938 ) | ( n47937 & ~n47938 ) ;
  assign n47940 = ( n9503 & n22623 ) | ( n9503 & n47939 ) | ( n22623 & n47939 ) ;
  assign n47941 = n1706 | n17885 ;
  assign n47942 = n47941 ^ n35448 ^ 1'b0 ;
  assign n47943 = n19113 ^ n7382 ^ n6433 ;
  assign n47944 = n47943 ^ n39338 ^ 1'b0 ;
  assign n47945 = n21865 ^ n3534 ^ 1'b0 ;
  assign n47946 = n26848 | n47945 ;
  assign n47947 = n16283 | n42923 ;
  assign n47950 = n1233 | n13924 ;
  assign n47948 = n12767 & ~n22209 ;
  assign n47949 = n47948 ^ n25784 ^ 1'b0 ;
  assign n47951 = n47950 ^ n47949 ^ n41865 ;
  assign n47952 = n21006 ^ n16181 ^ 1'b0 ;
  assign n47953 = n44071 ^ n41554 ^ n6464 ;
  assign n47954 = n7212 & ~n13633 ;
  assign n47955 = n47954 ^ n26861 ^ 1'b0 ;
  assign n47956 = n27873 ^ n3026 ^ 1'b0 ;
  assign n47957 = n44733 | n47956 ;
  assign n47959 = ~n4799 & n13241 ;
  assign n47960 = n21590 & n47959 ;
  assign n47961 = ~n10831 & n47960 ;
  assign n47958 = ( ~n12838 & n24235 ) | ( ~n12838 & n37371 ) | ( n24235 & n37371 ) ;
  assign n47962 = n47961 ^ n47958 ^ n11113 ;
  assign n47963 = ( n4844 & n11899 ) | ( n4844 & n47962 ) | ( n11899 & n47962 ) ;
  assign n47964 = n2699 ^ n2063 ^ 1'b0 ;
  assign n47965 = n25115 | n47964 ;
  assign n47966 = n47965 ^ n5102 ^ 1'b0 ;
  assign n47967 = n35149 | n42006 ;
  assign n47968 = n35096 ^ n32143 ^ 1'b0 ;
  assign n47970 = ~n5516 & n11621 ;
  assign n47969 = ~n2216 & n39727 ;
  assign n47971 = n47970 ^ n47969 ^ n7145 ;
  assign n47972 = n32418 & ~n32676 ;
  assign n47973 = ~n2968 & n23393 ;
  assign n47974 = ~n19756 & n47973 ;
  assign n47975 = ( n17186 & n26917 ) | ( n17186 & n38705 ) | ( n26917 & n38705 ) ;
  assign n47976 = n47974 & ~n47975 ;
  assign n47977 = ~n4597 & n44750 ;
  assign n47978 = n39886 & n47977 ;
  assign n47979 = ( n8531 & n13283 ) | ( n8531 & n14370 ) | ( n13283 & n14370 ) ;
  assign n47980 = n4257 & n47979 ;
  assign n47981 = n34018 & n47980 ;
  assign n47982 = n47981 ^ n26854 ^ n5481 ;
  assign n47983 = n40360 ^ n39994 ^ 1'b0 ;
  assign n47984 = n42738 | n47983 ;
  assign n47985 = n43453 & ~n47984 ;
  assign n47986 = ~n47982 & n47985 ;
  assign n47987 = n28292 & n38768 ;
  assign n47988 = n18097 ^ n13398 ^ 1'b0 ;
  assign n47989 = n23489 ^ n15213 ^ n11030 ;
  assign n47990 = ( n47987 & n47988 ) | ( n47987 & ~n47989 ) | ( n47988 & ~n47989 ) ;
  assign n47991 = ( n4567 & n14180 ) | ( n4567 & ~n25143 ) | ( n14180 & ~n25143 ) ;
  assign n47992 = n47991 ^ n30710 ^ n1438 ;
  assign n47993 = ( ~n4536 & n9799 ) | ( ~n4536 & n14922 ) | ( n9799 & n14922 ) ;
  assign n47994 = n22555 ^ n20663 ^ 1'b0 ;
  assign n47995 = ~n40187 & n47994 ;
  assign n47996 = n47995 ^ n45382 ^ n32890 ;
  assign n47997 = n41353 ^ n15969 ^ 1'b0 ;
  assign n47998 = ~n27065 & n47997 ;
  assign n47999 = n893 & ~n12278 ;
  assign n48000 = n34220 ^ n2965 ^ 1'b0 ;
  assign n48001 = ~n47999 & n48000 ;
  assign n48002 = n25013 & n48001 ;
  assign n48003 = n48002 ^ n4849 ^ 1'b0 ;
  assign n48004 = n1057 & ~n36209 ;
  assign n48005 = ~n8663 & n48004 ;
  assign n48006 = ( n11500 & n30058 ) | ( n11500 & ~n48005 ) | ( n30058 & ~n48005 ) ;
  assign n48007 = n48006 ^ n46055 ^ 1'b0 ;
  assign n48008 = ( n12596 & n41803 ) | ( n12596 & n44130 ) | ( n41803 & n44130 ) ;
  assign n48009 = n19414 ^ n15460 ^ 1'b0 ;
  assign n48010 = n3518 & n8159 ;
  assign n48011 = ( n41844 & ~n48009 ) | ( n41844 & n48010 ) | ( ~n48009 & n48010 ) ;
  assign n48012 = n25041 ^ n12300 ^ 1'b0 ;
  assign n48013 = ( ~n17186 & n29510 ) | ( ~n17186 & n48012 ) | ( n29510 & n48012 ) ;
  assign n48014 = n35288 ^ n7412 ^ 1'b0 ;
  assign n48015 = n13587 | n48014 ;
  assign n48016 = n17141 & ~n48015 ;
  assign n48017 = n11690 ^ n3209 ^ 1'b0 ;
  assign n48018 = n28305 & n48017 ;
  assign n48019 = n22366 & ~n45475 ;
  assign n48020 = ~n13396 & n48019 ;
  assign n48021 = n8754 ^ n5640 ^ 1'b0 ;
  assign n48022 = n4350 | n48021 ;
  assign n48023 = n11773 ^ n6862 ^ 1'b0 ;
  assign n48024 = n19322 & n48023 ;
  assign n48025 = ~n48022 & n48024 ;
  assign n48026 = n48025 ^ n7321 ^ n1981 ;
  assign n48027 = n22026 & ~n31621 ;
  assign n48030 = n11527 ^ n728 ^ 1'b0 ;
  assign n48031 = n341 & ~n48030 ;
  assign n48028 = n21929 & ~n22102 ;
  assign n48029 = ~n26655 & n48028 ;
  assign n48032 = n48031 ^ n48029 ^ n15153 ;
  assign n48033 = n48032 ^ n41968 ^ n29894 ;
  assign n48034 = n12996 ^ n12140 ^ 1'b0 ;
  assign n48035 = n22308 & n48034 ;
  assign n48036 = n3885 & n48035 ;
  assign n48037 = n48036 ^ n1793 ^ 1'b0 ;
  assign n48038 = n39787 & ~n43269 ;
  assign n48039 = n48038 ^ n9320 ^ 1'b0 ;
  assign n48040 = ~n8566 & n35062 ;
  assign n48041 = n4364 & n48040 ;
  assign n48042 = n43908 ^ n22961 ^ 1'b0 ;
  assign n48043 = ~n48041 & n48042 ;
  assign n48046 = n26944 ^ n1159 ^ 1'b0 ;
  assign n48044 = n2006 & n12000 ;
  assign n48045 = n26124 & n48044 ;
  assign n48047 = n48046 ^ n48045 ^ n14766 ;
  assign n48048 = ~n13518 & n16901 ;
  assign n48049 = n48048 ^ n3156 ^ 1'b0 ;
  assign n48050 = n48049 ^ n22631 ^ n18530 ;
  assign n48051 = ( n13708 & n32792 ) | ( n13708 & ~n48050 ) | ( n32792 & ~n48050 ) ;
  assign n48052 = n32466 ^ n18998 ^ 1'b0 ;
  assign n48053 = ~n9403 & n10403 ;
  assign n48054 = ~n31704 & n32043 ;
  assign n48055 = n3323 ^ n813 ^ 1'b0 ;
  assign n48056 = n6976 & n23843 ;
  assign n48057 = ~n48055 & n48056 ;
  assign n48058 = n25033 ^ n5966 ^ 1'b0 ;
  assign n48059 = ~n6899 & n25344 ;
  assign n48060 = n48059 ^ n19673 ^ 1'b0 ;
  assign n48061 = ( n28030 & n36457 ) | ( n28030 & ~n48060 ) | ( n36457 & ~n48060 ) ;
  assign n48062 = n38456 ^ n30838 ^ 1'b0 ;
  assign n48063 = n39802 ^ n15334 ^ n431 ;
  assign n48064 = n42484 ^ n39488 ^ n32032 ;
  assign n48065 = n29921 ^ n16951 ^ n5737 ;
  assign n48066 = ~n8689 & n48065 ;
  assign n48067 = x62 & n22573 ;
  assign n48068 = n21587 | n31504 ;
  assign n48069 = n48068 ^ n13991 ^ 1'b0 ;
  assign n48070 = n14320 & ~n48069 ;
  assign n48071 = ~n29439 & n48070 ;
  assign n48072 = ( ~n3517 & n5970 ) | ( ~n3517 & n20144 ) | ( n5970 & n20144 ) ;
  assign n48073 = n48072 ^ n23544 ^ n7980 ;
  assign n48074 = n48073 ^ n10995 ^ 1'b0 ;
  assign n48075 = n2337 & ~n48074 ;
  assign n48076 = n14393 ^ n2782 ^ 1'b0 ;
  assign n48077 = ~n1455 & n30688 ;
  assign n48078 = ( n15949 & n20611 ) | ( n15949 & n35232 ) | ( n20611 & n35232 ) ;
  assign n48079 = n9350 & ~n9825 ;
  assign n48080 = ( n16427 & ~n48078 ) | ( n16427 & n48079 ) | ( ~n48078 & n48079 ) ;
  assign n48081 = n28702 ^ n17004 ^ n1532 ;
  assign n48082 = ~n1919 & n20503 ;
  assign n48083 = ~n23329 & n48082 ;
  assign n48084 = n48083 ^ n2830 ^ 1'b0 ;
  assign n48085 = ( n16128 & ~n27842 ) | ( n16128 & n35355 ) | ( ~n27842 & n35355 ) ;
  assign n48086 = n48085 ^ n3413 ^ n2444 ;
  assign n48087 = n16489 ^ n3437 ^ 1'b0 ;
  assign n48088 = n43206 & n48087 ;
  assign n48089 = n12053 & n47506 ;
  assign n48090 = n48089 ^ n3872 ^ 1'b0 ;
  assign n48091 = n24394 & n48090 ;
  assign n48092 = ~n31154 & n48091 ;
  assign n48093 = n3459 | n22873 ;
  assign n48094 = n48092 & ~n48093 ;
  assign n48095 = n600 & n6460 ;
  assign n48096 = ~n11542 & n48095 ;
  assign n48097 = n40937 | n48096 ;
  assign n48098 = n48097 ^ n21683 ^ 1'b0 ;
  assign n48100 = n2310 & n24154 ;
  assign n48101 = n48100 ^ n10427 ^ 1'b0 ;
  assign n48099 = n22106 & n22190 ;
  assign n48102 = n48101 ^ n48099 ^ 1'b0 ;
  assign n48103 = n18106 & ~n48102 ;
  assign n48105 = n14704 ^ n10899 ^ 1'b0 ;
  assign n48106 = n9032 & n48105 ;
  assign n48104 = ( ~n4922 & n17391 ) | ( ~n4922 & n31666 ) | ( n17391 & n31666 ) ;
  assign n48107 = n48106 ^ n48104 ^ 1'b0 ;
  assign n48108 = n31963 ^ n24771 ^ n19868 ;
  assign n48109 = ( ~n14701 & n48107 ) | ( ~n14701 & n48108 ) | ( n48107 & n48108 ) ;
  assign n48110 = n8907 ^ n6334 ^ 1'b0 ;
  assign n48111 = n30626 | n48110 ;
  assign n48112 = n48111 ^ n28212 ^ n26088 ;
  assign n48113 = n29149 | n48112 ;
  assign n48114 = ( ~n10043 & n16693 ) | ( ~n10043 & n18994 ) | ( n16693 & n18994 ) ;
  assign n48115 = n20840 & ~n48114 ;
  assign n48116 = ~n20542 & n31637 ;
  assign n48117 = n3204 & n17065 ;
  assign n48118 = n2461 & n48117 ;
  assign n48119 = n13448 & n24296 ;
  assign n48120 = n29693 ^ n25807 ^ n16912 ;
  assign n48121 = n10245 | n48120 ;
  assign n48122 = n46958 | n48121 ;
  assign n48123 = n24441 ^ n13787 ^ 1'b0 ;
  assign n48124 = n11829 & ~n33393 ;
  assign n48125 = n48124 ^ n39893 ^ 1'b0 ;
  assign n48126 = ( n6043 & n20742 ) | ( n6043 & n23569 ) | ( n20742 & n23569 ) ;
  assign n48132 = n4779 ^ n3160 ^ 1'b0 ;
  assign n48130 = n34406 ^ n23549 ^ n4459 ;
  assign n48127 = n44322 ^ n23118 ^ 1'b0 ;
  assign n48128 = n2122 & ~n48127 ;
  assign n48129 = ( n20321 & n23973 ) | ( n20321 & ~n48128 ) | ( n23973 & ~n48128 ) ;
  assign n48131 = n48130 ^ n48129 ^ n34410 ;
  assign n48133 = n48132 ^ n48131 ^ n11982 ;
  assign n48134 = ( n16786 & ~n24966 ) | ( n16786 & n31633 ) | ( ~n24966 & n31633 ) ;
  assign n48135 = n16522 ^ n8176 ^ 1'b0 ;
  assign n48136 = n19424 ^ n7116 ^ 1'b0 ;
  assign n48137 = n48136 ^ n47901 ^ 1'b0 ;
  assign n48138 = n5735 & ~n48137 ;
  assign n48139 = n48138 ^ n38369 ^ 1'b0 ;
  assign n48140 = ~n27070 & n48139 ;
  assign n48141 = n27277 ^ n4622 ^ 1'b0 ;
  assign n48142 = n33637 | n48141 ;
  assign n48143 = n473 & ~n14148 ;
  assign n48144 = n48142 & n48143 ;
  assign n48145 = n37635 ^ n33648 ^ n17337 ;
  assign n48146 = n44722 ^ n23695 ^ 1'b0 ;
  assign n48147 = n11977 ^ n10727 ^ n832 ;
  assign n48148 = n28041 & n36564 ;
  assign n48149 = n48148 ^ n9164 ^ 1'b0 ;
  assign n48150 = ~n3245 & n12051 ;
  assign n48151 = ~n22983 & n48150 ;
  assign n48152 = n48151 ^ n19176 ^ 1'b0 ;
  assign n48153 = ~n7412 & n48152 ;
  assign n48154 = ~n48149 & n48153 ;
  assign n48155 = n48147 | n48154 ;
  assign n48156 = n25833 ^ n4101 ^ n2663 ;
  assign n48157 = ( n3127 & n11283 ) | ( n3127 & n48156 ) | ( n11283 & n48156 ) ;
  assign n48158 = ~n41007 & n48157 ;
  assign n48159 = n9585 & n27329 ;
  assign n48160 = n48159 ^ n29634 ^ 1'b0 ;
  assign n48161 = ( n4398 & n38705 ) | ( n4398 & n48160 ) | ( n38705 & n48160 ) ;
  assign n48162 = n30547 ^ n17757 ^ n1199 ;
  assign n48163 = n13227 | n22264 ;
  assign n48164 = n48163 ^ n46671 ^ 1'b0 ;
  assign n48165 = n21884 & n48164 ;
  assign n48166 = n3021 & n48165 ;
  assign n48167 = n9458 | n13461 ;
  assign n48168 = n13554 ^ n7004 ^ 1'b0 ;
  assign n48169 = ~n48167 & n48168 ;
  assign n48170 = n26489 ^ n3268 ^ 1'b0 ;
  assign n48173 = n31304 ^ n4223 ^ 1'b0 ;
  assign n48174 = ~n9434 & n48173 ;
  assign n48171 = n46511 ^ n20988 ^ 1'b0 ;
  assign n48172 = n12081 & ~n48171 ;
  assign n48175 = n48174 ^ n48172 ^ 1'b0 ;
  assign n48176 = n17428 ^ n16377 ^ 1'b0 ;
  assign n48177 = n48176 ^ n33446 ^ n14602 ;
  assign n48178 = n48177 ^ n11503 ^ 1'b0 ;
  assign n48179 = ( ~n18089 & n18695 ) | ( ~n18089 & n43825 ) | ( n18695 & n43825 ) ;
  assign n48180 = ( n11090 & n16838 ) | ( n11090 & n24781 ) | ( n16838 & n24781 ) ;
  assign n48181 = n30818 ^ n6802 ^ 1'b0 ;
  assign n48182 = ( n7139 & n19691 ) | ( n7139 & n27743 ) | ( n19691 & n27743 ) ;
  assign n48183 = ( n48180 & n48181 ) | ( n48180 & n48182 ) | ( n48181 & n48182 ) ;
  assign n48184 = n48183 ^ n29443 ^ n14691 ;
  assign n48185 = ~n27004 & n48184 ;
  assign n48186 = n36871 ^ n17807 ^ 1'b0 ;
  assign n48187 = ~n11498 & n31760 ;
  assign n48188 = n3418 & n48187 ;
  assign n48189 = n4762 | n25163 ;
  assign n48190 = n4604 | n48189 ;
  assign n48191 = n24530 | n44941 ;
  assign n48192 = n37584 & ~n48191 ;
  assign n48193 = n46347 ^ n12233 ^ 1'b0 ;
  assign n48194 = n48192 | n48193 ;
  assign n48195 = ( n3182 & n13251 ) | ( n3182 & ~n20247 ) | ( n13251 & ~n20247 ) ;
  assign n48199 = n18093 ^ n5522 ^ 1'b0 ;
  assign n48200 = n42061 & ~n48199 ;
  assign n48196 = n30785 ^ n8970 ^ 1'b0 ;
  assign n48197 = n9953 & n48196 ;
  assign n48198 = ( n8227 & n16733 ) | ( n8227 & ~n48197 ) | ( n16733 & ~n48197 ) ;
  assign n48201 = n48200 ^ n48198 ^ n40664 ;
  assign n48202 = ( n11270 & n32759 ) | ( n11270 & ~n34732 ) | ( n32759 & ~n34732 ) ;
  assign n48203 = n17812 ^ n12489 ^ 1'b0 ;
  assign n48204 = ~n2094 & n48203 ;
  assign n48205 = n22475 ^ n9169 ^ 1'b0 ;
  assign n48206 = n1360 & n3197 ;
  assign n48207 = n48206 ^ n3085 ^ 1'b0 ;
  assign n48208 = n48205 | n48207 ;
  assign n48209 = n48204 | n48208 ;
  assign n48210 = n43284 ^ n29241 ^ n14672 ;
  assign n48211 = n48210 ^ n8339 ^ 1'b0 ;
  assign n48212 = n48209 & ~n48211 ;
  assign n48213 = n31986 | n38886 ;
  assign n48214 = ( ~n2031 & n6843 ) | ( ~n2031 & n34705 ) | ( n6843 & n34705 ) ;
  assign n48215 = n48213 | n48214 ;
  assign n48216 = n33808 ^ n18268 ^ 1'b0 ;
  assign n48217 = ~n12119 & n48216 ;
  assign n48218 = n6574 | n8468 ;
  assign n48219 = n4799 & ~n48218 ;
  assign n48220 = ( n6428 & n15658 ) | ( n6428 & n39889 ) | ( n15658 & n39889 ) ;
  assign n48221 = ( n25521 & n41613 ) | ( n25521 & n42699 ) | ( n41613 & n42699 ) ;
  assign n48222 = n35692 ^ n17244 ^ n1830 ;
  assign n48223 = n11353 ^ n4187 ^ 1'b0 ;
  assign n48224 = n22651 ^ n9393 ^ 1'b0 ;
  assign n48225 = ( ~n37030 & n48223 ) | ( ~n37030 & n48224 ) | ( n48223 & n48224 ) ;
  assign n48226 = n15194 & n42740 ;
  assign n48227 = ~n24042 & n37887 ;
  assign n48228 = n48227 ^ n27654 ^ 1'b0 ;
  assign n48229 = n26288 ^ n24814 ^ 1'b0 ;
  assign n48230 = n17696 | n48229 ;
  assign n48231 = n18650 & n33777 ;
  assign n48232 = n48230 & n48231 ;
  assign n48233 = ( ~n26336 & n36791 ) | ( ~n26336 & n40017 ) | ( n36791 & n40017 ) ;
  assign n48234 = n3246 ^ x222 ^ 1'b0 ;
  assign n48235 = ~n9161 & n48234 ;
  assign n48236 = n48235 ^ n6647 ^ n2460 ;
  assign n48237 = n48236 ^ n3174 ^ 1'b0 ;
  assign n48238 = n25415 | n48237 ;
  assign n48239 = ( n5292 & ~n21090 ) | ( n5292 & n48238 ) | ( ~n21090 & n48238 ) ;
  assign n48240 = n9174 & n20713 ;
  assign n48241 = n1854 & ~n17768 ;
  assign n48242 = n22204 ^ n19687 ^ 1'b0 ;
  assign n48243 = n48241 & ~n48242 ;
  assign n48244 = n48243 ^ n36994 ^ x66 ;
  assign n48245 = n3756 & ~n18985 ;
  assign n48246 = n12222 & n48245 ;
  assign n48247 = n48246 ^ n30198 ^ 1'b0 ;
  assign n48248 = n11323 & n21166 ;
  assign n48249 = n48248 ^ n15140 ^ 1'b0 ;
  assign n48250 = n29783 | n48249 ;
  assign n48251 = n42803 | n48250 ;
  assign n48252 = n42793 ^ n21043 ^ 1'b0 ;
  assign n48253 = n48251 & ~n48252 ;
  assign n48254 = n47854 ^ n3096 ^ 1'b0 ;
  assign n48255 = ~n20867 & n48254 ;
  assign n48256 = n14368 & n39361 ;
  assign n48257 = n48256 ^ n1733 ^ 1'b0 ;
  assign n48258 = n923 & n7676 ;
  assign n48259 = n48258 ^ n1812 ^ 1'b0 ;
  assign n48262 = n7628 & ~n8603 ;
  assign n48263 = n48262 ^ n44350 ^ n8318 ;
  assign n48260 = n10862 | n27461 ;
  assign n48261 = n23962 & ~n48260 ;
  assign n48264 = n48263 ^ n48261 ^ n24115 ;
  assign n48265 = n17586 & n28726 ;
  assign n48266 = n19302 ^ n4346 ^ n1988 ;
  assign n48267 = ( n2119 & ~n19699 ) | ( n2119 & n22992 ) | ( ~n19699 & n22992 ) ;
  assign n48268 = n26911 ^ n16834 ^ 1'b0 ;
  assign n48269 = n20994 & n37643 ;
  assign n48270 = n2006 & n48269 ;
  assign n48271 = n48268 & ~n48270 ;
  assign n48272 = n16375 & ~n22218 ;
  assign n48273 = n26773 ^ n6595 ^ 1'b0 ;
  assign n48274 = n2365 & ~n48273 ;
  assign n48275 = n45800 ^ n31918 ^ 1'b0 ;
  assign n48276 = n12069 & ~n48275 ;
  assign n48277 = n20096 & n48276 ;
  assign n48278 = n48277 ^ n20870 ^ 1'b0 ;
  assign n48279 = n24700 ^ n7939 ^ 1'b0 ;
  assign n48280 = n48278 & n48279 ;
  assign n48281 = n38658 ^ n11584 ^ n8502 ;
  assign n48282 = ( n13412 & n13976 ) | ( n13412 & n30527 ) | ( n13976 & n30527 ) ;
  assign n48283 = n6175 | n39753 ;
  assign n48284 = n48283 ^ n22698 ^ 1'b0 ;
  assign n48285 = ( n12914 & n48282 ) | ( n12914 & n48284 ) | ( n48282 & n48284 ) ;
  assign n48286 = n30214 ^ n14354 ^ 1'b0 ;
  assign n48287 = ( n7172 & n28562 ) | ( n7172 & n38770 ) | ( n28562 & n38770 ) ;
  assign n48289 = ~n14607 & n25396 ;
  assign n48290 = n48289 ^ n11649 ^ 1'b0 ;
  assign n48288 = ( ~n12390 & n33015 ) | ( ~n12390 & n42797 ) | ( n33015 & n42797 ) ;
  assign n48291 = n48290 ^ n48288 ^ n5969 ;
  assign n48292 = n3739 & n26188 ;
  assign n48293 = n48292 ^ n26951 ^ 1'b0 ;
  assign n48294 = n46353 & ~n48293 ;
  assign n48295 = n18462 & n46802 ;
  assign n48296 = ~n2402 & n48295 ;
  assign n48297 = n20177 & n42577 ;
  assign n48298 = ~n29011 & n48297 ;
  assign n48299 = n28261 ^ n2834 ^ 1'b0 ;
  assign n48300 = n17896 & ~n48299 ;
  assign n48301 = n27386 ^ n24420 ^ n11183 ;
  assign n48302 = n12974 | n24174 ;
  assign n48303 = n297 & ~n48302 ;
  assign n48304 = ( ~n5369 & n22912 ) | ( ~n5369 & n48303 ) | ( n22912 & n48303 ) ;
  assign n48305 = ( n10332 & ~n34599 ) | ( n10332 & n39255 ) | ( ~n34599 & n39255 ) ;
  assign n48306 = n23963 ^ n1434 ^ 1'b0 ;
  assign n48307 = n22989 & n40977 ;
  assign n48308 = ~n686 & n46530 ;
  assign n48309 = n48308 ^ n15912 ^ 1'b0 ;
  assign n48310 = n15344 ^ n14331 ^ 1'b0 ;
  assign n48311 = ( n6340 & n19940 ) | ( n6340 & ~n48310 ) | ( n19940 & ~n48310 ) ;
  assign n48312 = n48311 ^ n24135 ^ n1939 ;
  assign n48313 = ( ~n13363 & n32820 ) | ( ~n13363 & n48312 ) | ( n32820 & n48312 ) ;
  assign n48314 = n16836 ^ n2549 ^ 1'b0 ;
  assign n48315 = n48313 & ~n48314 ;
  assign n48316 = ~n11197 & n25663 ;
  assign n48317 = n13914 & n28608 ;
  assign n48318 = n3363 & n48317 ;
  assign n48319 = ( n2444 & ~n3298 ) | ( n2444 & n32948 ) | ( ~n3298 & n32948 ) ;
  assign n48320 = n48319 ^ n38889 ^ n17516 ;
  assign n48321 = n48320 ^ n42096 ^ n1315 ;
  assign n48322 = ~n42195 & n48321 ;
  assign n48323 = n25065 ^ n18772 ^ 1'b0 ;
  assign n48324 = n28007 ^ n20236 ^ n12897 ;
  assign n48325 = n1910 | n8781 ;
  assign n48326 = n48325 ^ n13818 ^ 1'b0 ;
  assign n48327 = n48326 ^ n39210 ^ 1'b0 ;
  assign n48328 = ~n16677 & n35135 ;
  assign n48329 = n10722 & n48328 ;
  assign n48330 = ~n5324 & n13379 ;
  assign n48331 = n48329 & n48330 ;
  assign n48332 = n41978 & n48331 ;
  assign n48333 = ( n11825 & ~n13873 ) | ( n11825 & n48332 ) | ( ~n13873 & n48332 ) ;
  assign n48334 = n2229 & n4701 ;
  assign n48335 = ~n14452 & n48334 ;
  assign n48336 = n42438 ^ x104 ^ 1'b0 ;
  assign n48337 = n32718 ^ x43 ^ 1'b0 ;
  assign n48338 = n11995 & ~n48337 ;
  assign n48339 = ~n10446 & n12832 ;
  assign n48340 = n48339 ^ n33246 ^ 1'b0 ;
  assign n48346 = n9472 ^ n3204 ^ n2741 ;
  assign n48341 = ( n17294 & n20104 ) | ( n17294 & n45328 ) | ( n20104 & n45328 ) ;
  assign n48342 = n48341 ^ n13890 ^ 1'b0 ;
  assign n48343 = ( ~n36088 & n41454 ) | ( ~n36088 & n48342 ) | ( n41454 & n48342 ) ;
  assign n48344 = n336 & n48343 ;
  assign n48345 = n48344 ^ n19758 ^ 1'b0 ;
  assign n48347 = n48346 ^ n48345 ^ n14232 ;
  assign n48350 = n2583 & n15132 ;
  assign n48348 = ~n2765 & n3364 ;
  assign n48349 = ( n5233 & ~n13186 ) | ( n5233 & n48348 ) | ( ~n13186 & n48348 ) ;
  assign n48351 = n48350 ^ n48349 ^ n2548 ;
  assign n48352 = n37247 ^ n25505 ^ 1'b0 ;
  assign n48353 = ( n15578 & ~n23830 ) | ( n15578 & n30118 ) | ( ~n23830 & n30118 ) ;
  assign n48354 = n3390 | n27692 ;
  assign n48355 = n26669 | n48354 ;
  assign n48356 = n8976 | n33070 ;
  assign n48357 = n23098 & ~n48356 ;
  assign n48358 = n48357 ^ n32890 ^ 1'b0 ;
  assign n48359 = n14912 ^ n9555 ^ 1'b0 ;
  assign n48360 = n23501 & n48359 ;
  assign n48361 = ( ~n1700 & n8151 ) | ( ~n1700 & n48360 ) | ( n8151 & n48360 ) ;
  assign n48362 = n48361 ^ n8281 ^ 1'b0 ;
  assign n48363 = ~n11146 & n48362 ;
  assign n48364 = ( n504 & n2122 ) | ( n504 & ~n33377 ) | ( n2122 & ~n33377 ) ;
  assign n48365 = n6196 & n20420 ;
  assign n48366 = ~n28905 & n48365 ;
  assign n48367 = n48366 ^ n43916 ^ 1'b0 ;
  assign n48368 = n16584 | n41263 ;
  assign n48369 = n7801 | n16379 ;
  assign n48370 = ~n27252 & n48369 ;
  assign n48375 = n38666 ^ n13007 ^ 1'b0 ;
  assign n48371 = n18086 & ~n31996 ;
  assign n48372 = n48371 ^ n17838 ^ 1'b0 ;
  assign n48373 = n48372 ^ n44729 ^ x169 ;
  assign n48374 = n23572 & n48373 ;
  assign n48376 = n48375 ^ n48374 ^ 1'b0 ;
  assign n48377 = n22867 ^ n11674 ^ 1'b0 ;
  assign n48378 = n18625 & n48377 ;
  assign n48379 = ~n1148 & n36429 ;
  assign n48380 = n8813 | n8895 ;
  assign n48381 = n48380 ^ n12225 ^ n11248 ;
  assign n48382 = ~n48379 & n48381 ;
  assign n48384 = n4368 & ~n22418 ;
  assign n48383 = ~n6256 & n44633 ;
  assign n48385 = n48384 ^ n48383 ^ 1'b0 ;
  assign n48386 = ( n2276 & n7700 ) | ( n2276 & n46579 ) | ( n7700 & n46579 ) ;
  assign n48387 = n48386 ^ n16593 ^ 1'b0 ;
  assign n48390 = ( n8247 & ~n21976 ) | ( n8247 & n32768 ) | ( ~n21976 & n32768 ) ;
  assign n48391 = n26128 ^ n22397 ^ 1'b0 ;
  assign n48392 = ~n48390 & n48391 ;
  assign n48389 = n13447 ^ n715 ^ 1'b0 ;
  assign n48388 = n35251 ^ n2795 ^ 1'b0 ;
  assign n48393 = n48392 ^ n48389 ^ n48388 ;
  assign n48394 = ~n6022 & n15499 ;
  assign n48395 = n17932 ^ n11003 ^ 1'b0 ;
  assign n48396 = ~n17143 & n48395 ;
  assign n48397 = n48396 ^ n5271 ^ 1'b0 ;
  assign n48398 = n3968 | n13037 ;
  assign n48399 = ~x72 & n48398 ;
  assign n48400 = n48399 ^ n44494 ^ n14600 ;
  assign n48401 = n47405 ^ n22292 ^ 1'b0 ;
  assign n48402 = ~n1033 & n48401 ;
  assign n48403 = n48402 ^ n21715 ^ 1'b0 ;
  assign n48404 = ~n2702 & n48403 ;
  assign n48405 = n34756 ^ n21910 ^ 1'b0 ;
  assign n48406 = ( n907 & ~n11303 ) | ( n907 & n12967 ) | ( ~n11303 & n12967 ) ;
  assign n48409 = ( x204 & n4980 ) | ( x204 & n6279 ) | ( n4980 & n6279 ) ;
  assign n48408 = ( n22384 & n27342 ) | ( n22384 & n29113 ) | ( n27342 & n29113 ) ;
  assign n48407 = n38094 ^ n4632 ^ 1'b0 ;
  assign n48410 = n48409 ^ n48408 ^ n48407 ;
  assign n48411 = n34527 ^ n30220 ^ 1'b0 ;
  assign n48412 = n48410 | n48411 ;
  assign n48413 = n11896 ^ n4918 ^ 1'b0 ;
  assign n48414 = n269 & ~n48413 ;
  assign n48415 = n5933 ^ n3140 ^ n2466 ;
  assign n48416 = ( n10645 & n48414 ) | ( n10645 & ~n48415 ) | ( n48414 & ~n48415 ) ;
  assign n48417 = n48032 ^ n10546 ^ n3508 ;
  assign n48418 = n18434 ^ n5126 ^ 1'b0 ;
  assign n48419 = n20871 & n48418 ;
  assign n48420 = n48419 ^ n35156 ^ n33819 ;
  assign n48421 = n27157 ^ n2925 ^ 1'b0 ;
  assign n48422 = n7927 & n48421 ;
  assign n48423 = n48422 ^ n13972 ^ 1'b0 ;
  assign n48424 = n18738 | n48423 ;
  assign n48425 = n755 & ~n48424 ;
  assign n48426 = n48425 ^ n22206 ^ 1'b0 ;
  assign n48427 = n48426 ^ n22808 ^ n5730 ;
  assign n48428 = n25864 ^ x158 ^ 1'b0 ;
  assign n48429 = n17232 | n48428 ;
  assign n48430 = ( ~n12396 & n47527 ) | ( ~n12396 & n48429 ) | ( n47527 & n48429 ) ;
  assign n48431 = n15826 ^ n373 ^ 1'b0 ;
  assign n48432 = n13605 & n34608 ;
  assign n48433 = ( n39658 & ~n48431 ) | ( n39658 & n48432 ) | ( ~n48431 & n48432 ) ;
  assign n48434 = n48433 ^ n34543 ^ 1'b0 ;
  assign n48435 = n33378 | n37049 ;
  assign n48436 = n48435 ^ n7659 ^ 1'b0 ;
  assign n48437 = n479 & n7252 ;
  assign n48438 = ~n1052 & n48437 ;
  assign n48439 = ( ~n16541 & n33577 ) | ( ~n16541 & n48438 ) | ( n33577 & n48438 ) ;
  assign n48440 = n48439 ^ n3670 ^ 1'b0 ;
  assign n48441 = n16332 ^ n9151 ^ 1'b0 ;
  assign n48442 = n48441 ^ n23920 ^ n8800 ;
  assign n48443 = n8943 | n43522 ;
  assign n48444 = n48443 ^ n22685 ^ 1'b0 ;
  assign n48445 = n23365 & n48444 ;
  assign n48446 = ( ~n9650 & n18639 ) | ( ~n9650 & n40017 ) | ( n18639 & n40017 ) ;
  assign n48447 = n48446 ^ n11083 ^ 1'b0 ;
  assign n48448 = n4482 | n10599 ;
  assign n48449 = n48448 ^ n28402 ^ 1'b0 ;
  assign n48450 = n2382 | n48449 ;
  assign n48451 = ( n29660 & n48447 ) | ( n29660 & n48450 ) | ( n48447 & n48450 ) ;
  assign n48452 = ~n4436 & n44089 ;
  assign n48453 = n20173 & n27686 ;
  assign n48454 = n48453 ^ n41997 ^ 1'b0 ;
  assign n48455 = n9357 & n25345 ;
  assign n48456 = n48455 ^ n3666 ^ 1'b0 ;
  assign n48457 = n35575 ^ n9280 ^ 1'b0 ;
  assign n48458 = n38642 & n48457 ;
  assign n48459 = n33193 ^ n20484 ^ n4148 ;
  assign n48460 = n48459 ^ n27694 ^ 1'b0 ;
  assign n48461 = ~n13339 & n48460 ;
  assign n48462 = n33517 | n48461 ;
  assign n48463 = n39000 ^ n4825 ^ n1483 ;
  assign n48464 = n5589 | n38166 ;
  assign n48465 = n16927 & ~n48464 ;
  assign n48466 = ( n7441 & ~n36012 ) | ( n7441 & n48465 ) | ( ~n36012 & n48465 ) ;
  assign n48467 = n28643 ^ n21589 ^ n5394 ;
  assign n48468 = n48467 ^ n3844 ^ n1906 ;
  assign n48469 = ( n9553 & ~n21497 ) | ( n9553 & n48468 ) | ( ~n21497 & n48468 ) ;
  assign n48470 = n38021 ^ n25347 ^ n19259 ;
  assign n48471 = n48470 ^ n8480 ^ 1'b0 ;
  assign n48472 = n48471 ^ n8392 ^ n7980 ;
  assign n48473 = ~n10096 & n32080 ;
  assign n48474 = ~n8913 & n48473 ;
  assign n48477 = n42297 ^ n40005 ^ 1'b0 ;
  assign n48478 = ~n32488 & n48477 ;
  assign n48479 = n48478 ^ n29515 ^ 1'b0 ;
  assign n48475 = n38315 ^ n26284 ^ 1'b0 ;
  assign n48476 = n30671 | n48475 ;
  assign n48480 = n48479 ^ n48476 ^ 1'b0 ;
  assign n48481 = n25170 ^ n20538 ^ n17943 ;
  assign n48482 = n48481 ^ n45097 ^ n12399 ;
  assign n48483 = ( n12428 & n39296 ) | ( n12428 & ~n48482 ) | ( n39296 & ~n48482 ) ;
  assign n48484 = n38105 ^ n34298 ^ 1'b0 ;
  assign n48485 = ( ~n12488 & n17256 ) | ( ~n12488 & n48484 ) | ( n17256 & n48484 ) ;
  assign n48486 = n22418 ^ n16122 ^ n8045 ;
  assign n48487 = ~n11082 & n12899 ;
  assign n48488 = n32269 | n48487 ;
  assign n48489 = n44194 | n45376 ;
  assign n48490 = n19172 & n42638 ;
  assign n48491 = ( ~n6582 & n13181 ) | ( ~n6582 & n18449 ) | ( n13181 & n18449 ) ;
  assign n48492 = ( n5673 & ~n7061 ) | ( n5673 & n48491 ) | ( ~n7061 & n48491 ) ;
  assign n48493 = ( n16623 & ~n34029 ) | ( n16623 & n48492 ) | ( ~n34029 & n48492 ) ;
  assign n48494 = n34029 ^ n12311 ^ 1'b0 ;
  assign n48495 = ~n48493 & n48494 ;
  assign n48496 = n37430 ^ n4898 ^ 1'b0 ;
  assign n48497 = n23448 & n48496 ;
  assign n48498 = ( ~n809 & n2580 ) | ( ~n809 & n30101 ) | ( n2580 & n30101 ) ;
  assign n48499 = n39483 ^ n17081 ^ 1'b0 ;
  assign n48500 = ( n48497 & ~n48498 ) | ( n48497 & n48499 ) | ( ~n48498 & n48499 ) ;
  assign n48501 = n15175 ^ n2359 ^ 1'b0 ;
  assign n48502 = n48500 | n48501 ;
  assign n48503 = n9738 & n13464 ;
  assign n48504 = n48503 ^ n15156 ^ 1'b0 ;
  assign n48505 = n26115 | n48504 ;
  assign n48506 = n26768 & ~n48505 ;
  assign n48507 = n21902 & ~n29669 ;
  assign n48508 = n25226 ^ n19197 ^ n1907 ;
  assign n48509 = n48508 ^ n43696 ^ n13653 ;
  assign n48510 = n48509 ^ n1452 ^ n1051 ;
  assign n48514 = ( ~n1150 & n12304 ) | ( ~n1150 & n15422 ) | ( n12304 & n15422 ) ;
  assign n48511 = n11784 | n28152 ;
  assign n48512 = n13347 & ~n48511 ;
  assign n48513 = ( n2021 & ~n40516 ) | ( n2021 & n48512 ) | ( ~n40516 & n48512 ) ;
  assign n48515 = n48514 ^ n48513 ^ n791 ;
  assign n48516 = ( n21229 & ~n48510 ) | ( n21229 & n48515 ) | ( ~n48510 & n48515 ) ;
  assign n48517 = n44255 ^ n16117 ^ n2783 ;
  assign n48518 = ( n3247 & n28352 ) | ( n3247 & n48517 ) | ( n28352 & n48517 ) ;
  assign n48519 = ( n776 & ~n25396 ) | ( n776 & n45031 ) | ( ~n25396 & n45031 ) ;
  assign n48520 = n37464 ^ n6260 ^ 1'b0 ;
  assign n48521 = n6941 ^ n2639 ^ 1'b0 ;
  assign n48522 = n2356 ^ n1945 ^ 1'b0 ;
  assign n48523 = ~n2550 & n48522 ;
  assign n48524 = n5675 ^ n3559 ^ 1'b0 ;
  assign n48525 = n15547 & ~n48524 ;
  assign n48526 = ~n5964 & n44234 ;
  assign n48527 = n40284 & n48526 ;
  assign n48528 = n30042 & n40317 ;
  assign n48529 = n18769 ^ n10301 ^ n10027 ;
  assign n48530 = ( n9790 & n23163 ) | ( n9790 & n46560 ) | ( n23163 & n46560 ) ;
  assign n48531 = n48530 ^ n5735 ^ 1'b0 ;
  assign n48532 = n7270 & n48531 ;
  assign n48533 = n48532 ^ n29959 ^ n11532 ;
  assign n48534 = ~n6150 & n30362 ;
  assign n48535 = n2332 & ~n23684 ;
  assign n48536 = ~n30116 & n48535 ;
  assign n48537 = n48536 ^ n12719 ^ 1'b0 ;
  assign n48538 = n18116 | n48537 ;
  assign n48539 = n7679 ^ n6789 ^ 1'b0 ;
  assign n48540 = n3892 | n42200 ;
  assign n48541 = n48539 & ~n48540 ;
  assign n48542 = n36267 ^ n3653 ^ 1'b0 ;
  assign n48543 = n8490 | n15781 ;
  assign n48544 = n48543 ^ n16920 ^ n15085 ;
  assign n48545 = n48544 ^ n5436 ^ 1'b0 ;
  assign n48546 = n35555 & n48545 ;
  assign n48547 = n25392 ^ n11565 ^ n561 ;
  assign n48548 = n26443 & ~n48547 ;
  assign n48549 = n9702 & n48548 ;
  assign n48550 = ( n8764 & ~n26743 ) | ( n8764 & n48549 ) | ( ~n26743 & n48549 ) ;
  assign n48551 = n48550 ^ n4073 ^ n1832 ;
  assign n48552 = n48546 & ~n48551 ;
  assign n48553 = n22635 ^ n16167 ^ n14277 ;
  assign n48554 = n48553 ^ n13830 ^ 1'b0 ;
  assign n48555 = ( n12792 & ~n13039 ) | ( n12792 & n37860 ) | ( ~n13039 & n37860 ) ;
  assign n48556 = ( ~n10674 & n14117 ) | ( ~n10674 & n19229 ) | ( n14117 & n19229 ) ;
  assign n48557 = n48556 ^ n27962 ^ n419 ;
  assign n48558 = n10781 & n23132 ;
  assign n48559 = n21800 ^ n9894 ^ 1'b0 ;
  assign n48560 = n299 | n25104 ;
  assign n48561 = x62 | n48560 ;
  assign n48562 = n42030 ^ n1454 ^ 1'b0 ;
  assign n48563 = ( n12843 & n48561 ) | ( n12843 & ~n48562 ) | ( n48561 & ~n48562 ) ;
  assign n48564 = n37935 | n40645 ;
  assign n48565 = n48563 | n48564 ;
  assign n48566 = n1705 & ~n43691 ;
  assign n48567 = n35353 ^ n28585 ^ n13571 ;
  assign n48568 = ~n15590 & n19744 ;
  assign n48569 = n2781 & ~n48568 ;
  assign n48571 = ( n6274 & n7422 ) | ( n6274 & n45278 ) | ( n7422 & n45278 ) ;
  assign n48570 = n19645 ^ n4242 ^ x36 ;
  assign n48572 = n48571 ^ n48570 ^ n34097 ;
  assign n48573 = n29840 ^ n4675 ^ 1'b0 ;
  assign n48574 = n6611 & ~n48573 ;
  assign n48575 = n11649 & ~n37659 ;
  assign n48576 = n48575 ^ n32585 ^ 1'b0 ;
  assign n48577 = ( n2000 & n2231 ) | ( n2000 & ~n13135 ) | ( n2231 & ~n13135 ) ;
  assign n48578 = ( n2370 & n2854 ) | ( n2370 & n48577 ) | ( n2854 & n48577 ) ;
  assign n48579 = n48578 ^ n9334 ^ 1'b0 ;
  assign n48580 = n16765 ^ n10000 ^ 1'b0 ;
  assign n48581 = x94 | n36026 ;
  assign n48582 = n11984 | n43269 ;
  assign n48583 = n48581 | n48582 ;
  assign n48584 = n15699 ^ n13190 ^ 1'b0 ;
  assign n48585 = ~n7028 & n32175 ;
  assign n48586 = n29366 ^ n7878 ^ 1'b0 ;
  assign n48587 = n23295 | n48586 ;
  assign n48588 = ( n41543 & ~n48585 ) | ( n41543 & n48587 ) | ( ~n48585 & n48587 ) ;
  assign n48589 = n31993 ^ n12489 ^ 1'b0 ;
  assign n48590 = n29727 & n48589 ;
  assign n48591 = n38656 ^ n27438 ^ n10952 ;
  assign n48592 = ( ~n3750 & n10729 ) | ( ~n3750 & n48591 ) | ( n10729 & n48591 ) ;
  assign n48593 = n46274 ^ n21138 ^ 1'b0 ;
  assign n48594 = n42226 ^ n15278 ^ 1'b0 ;
  assign n48595 = n18389 ^ n3737 ^ 1'b0 ;
  assign n48596 = n20097 | n48595 ;
  assign n48597 = n34437 ^ n1312 ^ 1'b0 ;
  assign n48598 = n2255 | n48597 ;
  assign n48599 = n256 & n48598 ;
  assign n48600 = n8156 ^ n6406 ^ n2403 ;
  assign n48601 = n38180 ^ n12746 ^ 1'b0 ;
  assign n48602 = n31568 ^ n21880 ^ 1'b0 ;
  assign n48603 = ~n23161 & n48602 ;
  assign n48604 = n2745 | n40913 ;
  assign n48605 = n37100 & ~n48604 ;
  assign n48606 = n48605 ^ n6132 ^ 1'b0 ;
  assign n48607 = n22037 ^ n4064 ^ n3004 ;
  assign n48608 = ~n48606 & n48607 ;
  assign n48609 = n48608 ^ n35234 ^ n31145 ;
  assign n48610 = ( n25314 & ~n29671 ) | ( n25314 & n39101 ) | ( ~n29671 & n39101 ) ;
  assign n48611 = ( n19233 & n30107 ) | ( n19233 & ~n48610 ) | ( n30107 & ~n48610 ) ;
  assign n48612 = ( n4639 & n27732 ) | ( n4639 & ~n43018 ) | ( n27732 & ~n43018 ) ;
  assign n48613 = ( n48609 & n48611 ) | ( n48609 & n48612 ) | ( n48611 & n48612 ) ;
  assign n48614 = n48395 ^ n20963 ^ 1'b0 ;
  assign n48615 = n35502 ^ n12201 ^ n7806 ;
  assign n48616 = ( n35979 & n48614 ) | ( n35979 & ~n48615 ) | ( n48614 & ~n48615 ) ;
  assign n48617 = n9165 ^ x123 ^ 1'b0 ;
  assign n48618 = n1516 | n24494 ;
  assign n48619 = n48617 | n48618 ;
  assign n48620 = ~n28230 & n38420 ;
  assign n48621 = n32699 & n48620 ;
  assign n48622 = n48621 ^ n21044 ^ 1'b0 ;
  assign n48623 = n39787 & n48622 ;
  assign n48624 = n26725 | n27039 ;
  assign n48625 = n471 | n17690 ;
  assign n48626 = n48625 ^ n36445 ^ 1'b0 ;
  assign n48627 = n25453 | n48626 ;
  assign n48628 = n25056 ^ n13168 ^ n8500 ;
  assign n48629 = n37530 ^ n6158 ^ 1'b0 ;
  assign n48630 = n10941 & ~n48629 ;
  assign n48631 = n24052 | n48630 ;
  assign n48632 = n3550 & n47055 ;
  assign n48633 = ~n20844 & n48632 ;
  assign n48634 = n48633 ^ n31307 ^ n5714 ;
  assign n48635 = n32868 ^ n20793 ^ n2533 ;
  assign n48636 = n26058 & ~n37471 ;
  assign n48637 = ~n9247 & n47718 ;
  assign n48638 = n4414 & n13203 ;
  assign n48639 = ~n47834 & n48638 ;
  assign n48640 = n27800 & n30854 ;
  assign n48641 = n6339 | n27808 ;
  assign n48642 = n48641 ^ n23016 ^ 1'b0 ;
  assign n48643 = n15798 ^ n4410 ^ n2492 ;
  assign n48644 = n48643 ^ n22102 ^ 1'b0 ;
  assign n48645 = n31587 | n48644 ;
  assign n48646 = n18521 | n46743 ;
  assign n48647 = ( n4488 & n16873 ) | ( n4488 & ~n47558 ) | ( n16873 & ~n47558 ) ;
  assign n48653 = n6785 & ~n12801 ;
  assign n48654 = n5289 & n48653 ;
  assign n48655 = n48654 ^ n11389 ^ 1'b0 ;
  assign n48651 = ( n10502 & n10834 ) | ( n10502 & n41253 ) | ( n10834 & n41253 ) ;
  assign n48648 = n8295 ^ n7651 ^ n6823 ;
  assign n48649 = n48648 ^ n40058 ^ n7042 ;
  assign n48650 = n38692 | n48649 ;
  assign n48652 = n48651 ^ n48650 ^ 1'b0 ;
  assign n48656 = n48655 ^ n48652 ^ n6181 ;
  assign n48657 = n22121 | n38382 ;
  assign n48665 = n14577 & ~n16904 ;
  assign n48666 = n48665 ^ n33454 ^ 1'b0 ;
  assign n48664 = ( n12658 & n20437 ) | ( n12658 & ~n20454 ) | ( n20437 & ~n20454 ) ;
  assign n48667 = n48666 ^ n48664 ^ n5618 ;
  assign n48661 = n7228 | n8438 ;
  assign n48662 = n48661 ^ n6344 ^ 1'b0 ;
  assign n48658 = n21742 ^ n18796 ^ 1'b0 ;
  assign n48659 = n20204 | n48658 ;
  assign n48660 = n6869 & ~n48659 ;
  assign n48663 = n48662 ^ n48660 ^ n12496 ;
  assign n48668 = n48667 ^ n48663 ^ 1'b0 ;
  assign n48669 = n5064 & n39903 ;
  assign n48670 = ~n26962 & n48669 ;
  assign n48671 = n48670 ^ n27832 ^ 1'b0 ;
  assign n48672 = n23055 ^ n16895 ^ 1'b0 ;
  assign n48673 = n27457 & ~n48672 ;
  assign n48674 = n48673 ^ n39165 ^ 1'b0 ;
  assign n48675 = n15736 ^ n5112 ^ 1'b0 ;
  assign n48676 = ~n5042 & n48675 ;
  assign n48677 = x102 & n27288 ;
  assign n48678 = ~n5458 & n48677 ;
  assign n48679 = ( n5381 & ~n22214 ) | ( n5381 & n45761 ) | ( ~n22214 & n45761 ) ;
  assign n48680 = n47614 ^ n26220 ^ n8034 ;
  assign n48681 = n27238 & ~n33079 ;
  assign n48682 = n3187 | n29745 ;
  assign n48683 = n7022 ^ n6085 ^ 1'b0 ;
  assign n48684 = ~n33775 & n48683 ;
  assign n48685 = n48684 ^ n16729 ^ 1'b0 ;
  assign n48686 = ~n48682 & n48685 ;
  assign n48687 = n14516 & n40459 ;
  assign n48688 = n14445 & n48687 ;
  assign n48689 = n45917 ^ n7864 ^ 1'b0 ;
  assign n48690 = n48688 | n48689 ;
  assign n48691 = ( n10394 & n23812 ) | ( n10394 & ~n45429 ) | ( n23812 & ~n45429 ) ;
  assign n48692 = n10971 & ~n32935 ;
  assign n48693 = n48692 ^ n16960 ^ 1'b0 ;
  assign n48694 = ( n20982 & n48691 ) | ( n20982 & n48693 ) | ( n48691 & n48693 ) ;
  assign n48695 = ( n10617 & n38596 ) | ( n10617 & ~n48694 ) | ( n38596 & ~n48694 ) ;
  assign n48696 = n48695 ^ n30721 ^ 1'b0 ;
  assign n48697 = n5760 ^ n2286 ^ 1'b0 ;
  assign n48698 = ~n3788 & n48697 ;
  assign n48701 = ( n774 & n980 ) | ( n774 & ~n13337 ) | ( n980 & ~n13337 ) ;
  assign n48699 = ~n17385 & n31813 ;
  assign n48700 = n48699 ^ n1705 ^ 1'b0 ;
  assign n48702 = n48701 ^ n48700 ^ 1'b0 ;
  assign n48703 = n48698 & ~n48702 ;
  assign n48704 = ( n26672 & ~n43698 ) | ( n26672 & n48703 ) | ( ~n43698 & n48703 ) ;
  assign n48705 = ( ~n13659 & n19900 ) | ( ~n13659 & n31728 ) | ( n19900 & n31728 ) ;
  assign n48706 = ~n18365 & n24009 ;
  assign n48707 = n48706 ^ n2329 ^ 1'b0 ;
  assign n48708 = n48707 ^ n24725 ^ n22934 ;
  assign n48709 = ( n9718 & ~n31571 ) | ( n9718 & n46563 ) | ( ~n31571 & n46563 ) ;
  assign n48710 = n48709 ^ n2221 ^ n857 ;
  assign n48711 = n12841 | n21808 ;
  assign n48712 = ( ~n6791 & n22470 ) | ( ~n6791 & n42050 ) | ( n22470 & n42050 ) ;
  assign n48713 = n11427 & ~n48712 ;
  assign n48714 = n1773 | n16709 ;
  assign n48715 = n48714 ^ n17186 ^ 1'b0 ;
  assign n48716 = n33618 ^ n6283 ^ 1'b0 ;
  assign n48717 = n9146 & n48716 ;
  assign n48718 = n40782 ^ n21159 ^ 1'b0 ;
  assign n48719 = n9260 | n26121 ;
  assign n48720 = n48719 ^ n21046 ^ 1'b0 ;
  assign n48721 = n48720 ^ n10434 ^ n6514 ;
  assign n48723 = ~n10536 & n13433 ;
  assign n48722 = n41190 ^ n30976 ^ n5737 ;
  assign n48724 = n48723 ^ n48722 ^ n11166 ;
  assign n48725 = n42423 ^ n11106 ^ 1'b0 ;
  assign n48726 = n13073 ^ n12849 ^ n1611 ;
  assign n48727 = n6809 ^ n3887 ^ n2606 ;
  assign n48728 = n48727 ^ n37956 ^ n19644 ;
  assign n48729 = ~n10212 & n19634 ;
  assign n48730 = ~n48728 & n48729 ;
  assign n48731 = n43032 ^ n3958 ^ 1'b0 ;
  assign n48732 = n12739 ^ n2240 ^ 1'b0 ;
  assign n48733 = n30022 | n48732 ;
  assign n48734 = n11058 ^ n6866 ^ n5229 ;
  assign n48735 = n48734 ^ n18682 ^ n11138 ;
  assign n48736 = n48735 ^ n35701 ^ 1'b0 ;
  assign n48737 = n35234 ^ n13536 ^ n10150 ;
  assign n48738 = ( n7602 & n10108 ) | ( n7602 & ~n23321 ) | ( n10108 & ~n23321 ) ;
  assign n48739 = n29263 ^ n28613 ^ 1'b0 ;
  assign n48740 = ( n1582 & ~n33308 ) | ( n1582 & n48739 ) | ( ~n33308 & n48739 ) ;
  assign n48741 = ( n42328 & n48738 ) | ( n42328 & n48740 ) | ( n48738 & n48740 ) ;
  assign n48742 = n43122 ^ n26397 ^ 1'b0 ;
  assign n48743 = n48742 ^ n15741 ^ n13480 ;
  assign n48744 = ~n2336 & n16698 ;
  assign n48745 = n48744 ^ n5848 ^ n3226 ;
  assign n48746 = n23313 ^ n4904 ^ n3366 ;
  assign n48747 = n34454 | n48746 ;
  assign n48748 = n19300 | n21904 ;
  assign n48749 = n48748 ^ n37123 ^ 1'b0 ;
  assign n48750 = n26477 & ~n48749 ;
  assign n48751 = n7850 & n20380 ;
  assign n48752 = n41588 ^ n21914 ^ n14141 ;
  assign n48753 = n48752 ^ n16776 ^ 1'b0 ;
  assign n48754 = n31009 ^ n855 ^ 1'b0 ;
  assign n48755 = n22690 ^ n394 ^ 1'b0 ;
  assign n48756 = ( n13424 & ~n22125 ) | ( n13424 & n36009 ) | ( ~n22125 & n36009 ) ;
  assign n48757 = n8844 | n16843 ;
  assign n48758 = n48757 ^ n32337 ^ 1'b0 ;
  assign n48759 = ( ~n12726 & n18421 ) | ( ~n12726 & n48758 ) | ( n18421 & n48758 ) ;
  assign n48760 = ( ~n1059 & n36693 ) | ( ~n1059 & n38800 ) | ( n36693 & n38800 ) ;
  assign n48761 = ~n11992 & n31905 ;
  assign n48762 = n23324 ^ n19914 ^ 1'b0 ;
  assign n48763 = n41950 ^ n18340 ^ n4550 ;
  assign n48764 = n13303 & n48763 ;
  assign n48765 = n17954 ^ n6856 ^ 1'b0 ;
  assign n48766 = x5 & n48765 ;
  assign n48767 = n48766 ^ n2668 ^ 1'b0 ;
  assign n48768 = ( n4739 & n8063 ) | ( n4739 & ~n18796 ) | ( n8063 & ~n18796 ) ;
  assign n48769 = ( ~n8006 & n25408 ) | ( ~n8006 & n28658 ) | ( n25408 & n28658 ) ;
  assign n48770 = n48769 ^ n1543 ^ 1'b0 ;
  assign n48771 = n44284 & n48770 ;
  assign n48772 = n23484 ^ n10811 ^ n9078 ;
  assign n48773 = n1192 & n48772 ;
  assign n48774 = ( n2324 & ~n8939 ) | ( n2324 & n30781 ) | ( ~n8939 & n30781 ) ;
  assign n48775 = n48774 ^ n37870 ^ x168 ;
  assign n48776 = n6689 | n37654 ;
  assign n48777 = n17125 | n48776 ;
  assign n48781 = n39467 ^ n20438 ^ 1'b0 ;
  assign n48778 = n48138 ^ n3546 ^ 1'b0 ;
  assign n48779 = n8584 | n48778 ;
  assign n48780 = n48779 ^ n23207 ^ n7568 ;
  assign n48782 = n48781 ^ n48780 ^ n9595 ;
  assign n48783 = n48782 ^ n30652 ^ n18314 ;
  assign n48784 = n10264 ^ n6464 ^ 1'b0 ;
  assign n48785 = n3643 | n9931 ;
  assign n48786 = n22224 ^ n18839 ^ n7862 ;
  assign n48787 = n10791 & ~n48786 ;
  assign n48788 = ~n7128 & n48787 ;
  assign n48790 = ~n12345 & n36468 ;
  assign n48791 = ~n13332 & n48790 ;
  assign n48792 = n13910 ^ n4052 ^ 1'b0 ;
  assign n48793 = n13967 | n48792 ;
  assign n48794 = ~n48791 & n48793 ;
  assign n48789 = n14539 & n27457 ;
  assign n48795 = n48794 ^ n48789 ^ 1'b0 ;
  assign n48798 = n8125 & ~n15562 ;
  assign n48799 = n48798 ^ n15644 ^ n9267 ;
  assign n48796 = n5136 & n16338 ;
  assign n48797 = n48796 ^ n10898 ^ 1'b0 ;
  assign n48800 = n48799 ^ n48797 ^ 1'b0 ;
  assign n48801 = n27054 ^ n10672 ^ n543 ;
  assign n48802 = n12763 & ~n42456 ;
  assign n48803 = n34912 & n48802 ;
  assign n48804 = n48803 ^ n19005 ^ 1'b0 ;
  assign n48805 = ( n1805 & ~n48801 ) | ( n1805 & n48804 ) | ( ~n48801 & n48804 ) ;
  assign n48806 = ( n11013 & n24088 ) | ( n11013 & n41247 ) | ( n24088 & n41247 ) ;
  assign n48807 = ( ~n11298 & n15378 ) | ( ~n11298 & n21247 ) | ( n15378 & n21247 ) ;
  assign n48808 = n15548 | n34825 ;
  assign n48809 = n31860 | n48808 ;
  assign n48810 = n48809 ^ n25622 ^ 1'b0 ;
  assign n48811 = n45964 ^ n5601 ^ 1'b0 ;
  assign n48812 = n48811 ^ n20016 ^ 1'b0 ;
  assign n48813 = ( ~n48807 & n48810 ) | ( ~n48807 & n48812 ) | ( n48810 & n48812 ) ;
  assign n48816 = n4453 & n4706 ;
  assign n48817 = n26587 & n48816 ;
  assign n48814 = ~n3802 & n13582 ;
  assign n48815 = n48814 ^ n20727 ^ 1'b0 ;
  assign n48818 = n48817 ^ n48815 ^ n40740 ;
  assign n48819 = ~n9816 & n28565 ;
  assign n48820 = n43269 & n48819 ;
  assign n48821 = ( n2820 & n3044 ) | ( n2820 & n26478 ) | ( n3044 & n26478 ) ;
  assign n48822 = n48821 ^ n26731 ^ n17682 ;
  assign n48823 = ~n26416 & n35015 ;
  assign n48824 = ~n48822 & n48823 ;
  assign n48825 = n9534 & n22277 ;
  assign n48826 = n48825 ^ n16620 ^ 1'b0 ;
  assign n48827 = x88 | n11349 ;
  assign n48828 = n1099 & ~n6829 ;
  assign n48829 = n22594 & n48828 ;
  assign n48830 = n19793 ^ n12267 ^ 1'b0 ;
  assign n48831 = n30361 & ~n48830 ;
  assign n48834 = ( n6994 & ~n37544 ) | ( n6994 & n37690 ) | ( ~n37544 & n37690 ) ;
  assign n48835 = n47527 ^ n25323 ^ 1'b0 ;
  assign n48836 = ~n48834 & n48835 ;
  assign n48837 = n48836 ^ n7644 ^ 1'b0 ;
  assign n48832 = ~n5975 & n24381 ;
  assign n48833 = ~n30741 & n48832 ;
  assign n48838 = n48837 ^ n48833 ^ 1'b0 ;
  assign n48839 = n48838 ^ n7084 ^ n4005 ;
  assign n48840 = n11357 ^ n520 ^ 1'b0 ;
  assign n48841 = n20871 & n48840 ;
  assign n48842 = n9162 ^ x170 ^ 1'b0 ;
  assign n48843 = ~n2781 & n48842 ;
  assign n48844 = n17419 & n37938 ;
  assign n48845 = n48844 ^ n4577 ^ 1'b0 ;
  assign n48846 = n48843 & ~n48845 ;
  assign n48847 = n19157 | n24029 ;
  assign n48848 = n650 | n48847 ;
  assign n48849 = ~n11832 & n27256 ;
  assign n48850 = n7555 | n10577 ;
  assign n48851 = n1710 & n48850 ;
  assign n48852 = ~n48849 & n48851 ;
  assign n48853 = n11744 & ~n25966 ;
  assign n48854 = n6634 & n48853 ;
  assign n48855 = ( n2782 & n11339 ) | ( n2782 & ~n46651 ) | ( n11339 & ~n46651 ) ;
  assign n48856 = ( n7104 & ~n8655 ) | ( n7104 & n26485 ) | ( ~n8655 & n26485 ) ;
  assign n48857 = n25003 ^ n21787 ^ n2889 ;
  assign n48858 = ( n5838 & n20942 ) | ( n5838 & ~n48857 ) | ( n20942 & ~n48857 ) ;
  assign n48859 = n33115 ^ n26688 ^ n18470 ;
  assign n48860 = n48859 ^ n38616 ^ n16489 ;
  assign n48861 = n13330 | n13721 ;
  assign n48862 = n48861 ^ n6624 ^ 1'b0 ;
  assign n48863 = n4963 & n19282 ;
  assign n48864 = ~n45205 & n48863 ;
  assign n48865 = n5869 & n38487 ;
  assign n48866 = n48865 ^ n18513 ^ 1'b0 ;
  assign n48867 = ~n37155 & n48866 ;
  assign n48868 = ( ~n4629 & n7597 ) | ( ~n4629 & n15017 ) | ( n7597 & n15017 ) ;
  assign n48869 = n2369 | n48868 ;
  assign n48870 = n48869 ^ n44585 ^ 1'b0 ;
  assign n48871 = n13382 | n20683 ;
  assign n48872 = n14268 ^ n5829 ^ 1'b0 ;
  assign n48873 = n1488 | n48872 ;
  assign n48874 = n44906 ^ n17414 ^ n2497 ;
  assign n48879 = n20193 ^ n8776 ^ 1'b0 ;
  assign n48880 = n28014 | n48879 ;
  assign n48875 = n7232 ^ n747 ^ 1'b0 ;
  assign n48876 = n7596 & ~n48875 ;
  assign n48877 = ~n20614 & n43833 ;
  assign n48878 = ~n48876 & n48877 ;
  assign n48881 = n48880 ^ n48878 ^ n23909 ;
  assign n48882 = ~n32969 & n33015 ;
  assign n48883 = n47144 ^ n43530 ^ n15543 ;
  assign n48884 = n48883 ^ n18302 ^ n3035 ;
  assign n48885 = n7473 & ~n45852 ;
  assign n48886 = n48568 ^ n22115 ^ n13436 ;
  assign n48887 = n5751 & n28542 ;
  assign n48888 = n48887 ^ n2533 ^ 1'b0 ;
  assign n48889 = n4794 & n48888 ;
  assign n48890 = n44515 ^ n33734 ^ 1'b0 ;
  assign n48891 = ( n1928 & n24434 ) | ( n1928 & ~n47686 ) | ( n24434 & ~n47686 ) ;
  assign n48892 = n48891 ^ n43232 ^ n18243 ;
  assign n48898 = n4177 & n23332 ;
  assign n48895 = n10438 & n11658 ;
  assign n48896 = n48895 ^ n6107 ^ 1'b0 ;
  assign n48894 = n5064 & ~n24450 ;
  assign n48897 = n48896 ^ n48894 ^ 1'b0 ;
  assign n48893 = ( ~n6370 & n14418 ) | ( ~n6370 & n28538 ) | ( n14418 & n28538 ) ;
  assign n48899 = n48898 ^ n48897 ^ n48893 ;
  assign n48900 = n4837 | n8169 ;
  assign n48901 = n2705 | n48900 ;
  assign n48902 = n48901 ^ n27910 ^ 1'b0 ;
  assign n48903 = n2883 | n21329 ;
  assign n48904 = n48903 ^ n41932 ^ n11440 ;
  assign n48905 = n6203 | n48904 ;
  assign n48906 = n37384 ^ n33435 ^ 1'b0 ;
  assign n48907 = n31639 ^ n20840 ^ 1'b0 ;
  assign n48908 = ~n21856 & n48907 ;
  assign n48909 = n29807 ^ n20810 ^ 1'b0 ;
  assign n48910 = ~n1278 & n48909 ;
  assign n48911 = n16075 & ~n46341 ;
  assign n48912 = n35330 & n48911 ;
  assign n48913 = n12782 ^ n10650 ^ n9687 ;
  assign n48914 = n48912 & ~n48913 ;
  assign n48915 = n48914 ^ n8969 ^ n1393 ;
  assign n48916 = n11150 | n17920 ;
  assign n48917 = n48916 ^ n19860 ^ 1'b0 ;
  assign n48918 = ( n6865 & n25178 ) | ( n6865 & n48917 ) | ( n25178 & n48917 ) ;
  assign n48919 = ( n8510 & n15391 ) | ( n8510 & n47386 ) | ( n15391 & n47386 ) ;
  assign n48920 = n33662 ^ n15087 ^ 1'b0 ;
  assign n48921 = n13007 & ~n48920 ;
  assign n48922 = n48921 ^ n27248 ^ n15820 ;
  assign n48925 = n44452 ^ n6414 ^ 1'b0 ;
  assign n48923 = n48311 ^ n20321 ^ 1'b0 ;
  assign n48924 = n1975 & ~n48923 ;
  assign n48926 = n48925 ^ n48924 ^ n36626 ;
  assign n48927 = ~n4030 & n5208 ;
  assign n48928 = n31334 & n48927 ;
  assign n48929 = n7354 | n48928 ;
  assign n48930 = n48929 ^ n37564 ^ 1'b0 ;
  assign n48931 = n3577 | n28551 ;
  assign n48932 = n2213 | n48931 ;
  assign n48933 = n34081 | n48932 ;
  assign n48934 = n12223 & n48933 ;
  assign n48935 = n48934 ^ n24084 ^ 1'b0 ;
  assign n48936 = n21049 & n29300 ;
  assign n48937 = n48936 ^ n29930 ^ 1'b0 ;
  assign n48938 = ~n23644 & n35588 ;
  assign n48939 = n5416 & n12905 ;
  assign n48940 = n48939 ^ n19940 ^ 1'b0 ;
  assign n48941 = n22498 ^ n19210 ^ 1'b0 ;
  assign n48942 = ~n2602 & n4612 ;
  assign n48943 = n48942 ^ n43018 ^ n30543 ;
  assign n48944 = n13449 ^ n11019 ^ n3171 ;
  assign n48945 = ( n18222 & n22326 ) | ( n18222 & ~n48944 ) | ( n22326 & ~n48944 ) ;
  assign n48946 = ( n7941 & n9145 ) | ( n7941 & ~n23181 ) | ( n9145 & ~n23181 ) ;
  assign n48947 = n48946 ^ n20015 ^ n18841 ;
  assign n48950 = n10890 ^ n1930 ^ 1'b0 ;
  assign n48951 = n10159 | n48950 ;
  assign n48952 = n48951 ^ n8354 ^ n8156 ;
  assign n48948 = ~n4617 & n17783 ;
  assign n48949 = n48948 ^ n17836 ^ 1'b0 ;
  assign n48953 = n48952 ^ n48949 ^ n31252 ;
  assign n48954 = ( n7722 & n22478 ) | ( n7722 & n34904 ) | ( n22478 & n34904 ) ;
  assign n48955 = ~n543 & n48954 ;
  assign n48956 = ~n39452 & n48955 ;
  assign n48957 = n3666 ^ n1738 ^ 1'b0 ;
  assign n48958 = n19231 ^ n4360 ^ 1'b0 ;
  assign n48959 = ~n17279 & n25859 ;
  assign n48960 = n11641 & n48959 ;
  assign n48961 = ~n7974 & n39605 ;
  assign n48962 = n48961 ^ n28087 ^ 1'b0 ;
  assign n48965 = n12381 & n32098 ;
  assign n48963 = ( n2368 & n14900 ) | ( n2368 & n43701 ) | ( n14900 & n43701 ) ;
  assign n48964 = n48963 ^ n15269 ^ n4809 ;
  assign n48966 = n48965 ^ n48964 ^ n36849 ;
  assign n48967 = ( ~n28003 & n37733 ) | ( ~n28003 & n48966 ) | ( n37733 & n48966 ) ;
  assign n48968 = n34730 ^ n12437 ^ 1'b0 ;
  assign n48969 = ( n1690 & ~n3410 ) | ( n1690 & n48968 ) | ( ~n3410 & n48968 ) ;
  assign n48970 = ( n759 & n27238 ) | ( n759 & n48969 ) | ( n27238 & n48969 ) ;
  assign n48971 = n29084 ^ n21059 ^ n19253 ;
  assign n48972 = n31337 ^ n17186 ^ n9363 ;
  assign n48973 = ( n3482 & n21570 ) | ( n3482 & ~n34811 ) | ( n21570 & ~n34811 ) ;
  assign n48974 = n48973 ^ x188 ^ 1'b0 ;
  assign n48975 = n24054 | n48974 ;
  assign n48976 = ( n540 & n6628 ) | ( n540 & n18763 ) | ( n6628 & n18763 ) ;
  assign n48977 = n48976 ^ n14106 ^ 1'b0 ;
  assign n48978 = n21856 | n48977 ;
  assign n48979 = n12347 & ~n33565 ;
  assign n48980 = n48979 ^ n1723 ^ 1'b0 ;
  assign n48981 = n32199 ^ n27288 ^ n17208 ;
  assign n48982 = n12519 | n21611 ;
  assign n48983 = n48982 ^ n34302 ^ n12320 ;
  assign n48984 = n10848 & n24322 ;
  assign n48985 = n48984 ^ n47274 ^ n9429 ;
  assign n48986 = ( n17208 & n38800 ) | ( n17208 & n43330 ) | ( n38800 & n43330 ) ;
  assign n48987 = n10926 ^ n5344 ^ 1'b0 ;
  assign n48988 = n11357 & n48987 ;
  assign n48989 = ( n2329 & n16547 ) | ( n2329 & ~n48988 ) | ( n16547 & ~n48988 ) ;
  assign n48991 = n7714 & n15870 ;
  assign n48992 = n28873 & n48991 ;
  assign n48990 = ( n2031 & n40496 ) | ( n2031 & n41128 ) | ( n40496 & n41128 ) ;
  assign n48993 = n48992 ^ n48990 ^ n24397 ;
  assign n48994 = n46328 ^ n35081 ^ 1'b0 ;
  assign n48995 = n38563 ^ n23371 ^ 1'b0 ;
  assign n48996 = n26390 & n48995 ;
  assign n48997 = n13121 ^ n8869 ^ 1'b0 ;
  assign n48998 = n31344 & n48997 ;
  assign n48999 = ~n6199 & n48998 ;
  assign n49000 = n1986 & n48999 ;
  assign n49001 = n9829 | n23817 ;
  assign n49002 = n46490 ^ n27764 ^ 1'b0 ;
  assign n49003 = ~n40620 & n49002 ;
  assign n49004 = ~n18678 & n26379 ;
  assign n49005 = ( n1099 & n25385 ) | ( n1099 & ~n49004 ) | ( n25385 & ~n49004 ) ;
  assign n49006 = ( n5680 & ~n25514 ) | ( n5680 & n47423 ) | ( ~n25514 & n47423 ) ;
  assign n49007 = n26802 & ~n33239 ;
  assign n49008 = n25247 ^ n22291 ^ 1'b0 ;
  assign n49009 = n2333 & ~n49008 ;
  assign n49010 = n49009 ^ n14628 ^ 1'b0 ;
  assign n49011 = n18936 & n31533 ;
  assign n49012 = ( n14183 & n29868 ) | ( n14183 & n49011 ) | ( n29868 & n49011 ) ;
  assign n49013 = n17640 ^ n1888 ^ 1'b0 ;
  assign n49014 = n22548 & n49013 ;
  assign n49015 = n25477 & ~n49014 ;
  assign n49016 = ~n41882 & n49015 ;
  assign n49017 = n15957 ^ n15058 ^ n3301 ;
  assign n49018 = n15058 | n49017 ;
  assign n49019 = n49016 & ~n49018 ;
  assign n49020 = n2861 & ~n3034 ;
  assign n49021 = n49020 ^ n42607 ^ 1'b0 ;
  assign n49022 = ~n5937 & n32283 ;
  assign n49023 = ( n2545 & n8593 ) | ( n2545 & ~n30679 ) | ( n8593 & ~n30679 ) ;
  assign n49024 = n32425 & n49023 ;
  assign n49025 = ( n25242 & n25777 ) | ( n25242 & n30962 ) | ( n25777 & n30962 ) ;
  assign n49026 = n7897 & ~n15288 ;
  assign n49027 = n49026 ^ n1283 ^ 1'b0 ;
  assign n49028 = n49027 ^ n21687 ^ 1'b0 ;
  assign n49029 = n6129 | n42707 ;
  assign n49030 = n6267 | n20210 ;
  assign n49031 = n49030 ^ n5408 ^ 1'b0 ;
  assign n49032 = n15594 ^ n15244 ^ n3197 ;
  assign n49033 = ~n9251 & n31202 ;
  assign n49034 = ~n14575 & n49033 ;
  assign n49035 = n310 & ~n49034 ;
  assign n49036 = n49032 & n49035 ;
  assign n49037 = n16659 ^ n10098 ^ 1'b0 ;
  assign n49038 = ~n40530 & n49037 ;
  assign n49039 = n6740 & ~n11150 ;
  assign n49040 = n49039 ^ n10606 ^ 1'b0 ;
  assign n49041 = ( n1599 & ~n4562 ) | ( n1599 & n49040 ) | ( ~n4562 & n49040 ) ;
  assign n49042 = n5568 ^ n1662 ^ 1'b0 ;
  assign n49043 = n49042 ^ n31524 ^ n7136 ;
  assign n49044 = ( n36097 & n45187 ) | ( n36097 & ~n49043 ) | ( n45187 & ~n49043 ) ;
  assign n49045 = n40990 ^ n12287 ^ n10026 ;
  assign n49046 = n1877 & ~n24863 ;
  assign n49047 = n49046 ^ n34074 ^ 1'b0 ;
  assign n49048 = n38972 | n49047 ;
  assign n49049 = n11782 ^ n3375 ^ 1'b0 ;
  assign n49050 = n26898 & n49049 ;
  assign n49051 = n16620 & n23146 ;
  assign n49052 = n46331 & n49051 ;
  assign n49053 = n32177 ^ n31337 ^ n7143 ;
  assign n49054 = ~n7110 & n23422 ;
  assign n49055 = ~n36537 & n49054 ;
  assign n49056 = n49055 ^ x235 ^ 1'b0 ;
  assign n49057 = ( n1887 & n35232 ) | ( n1887 & ~n47166 ) | ( n35232 & ~n47166 ) ;
  assign n49061 = n2261 & ~n21490 ;
  assign n49058 = ( x172 & n3998 ) | ( x172 & n17981 ) | ( n3998 & n17981 ) ;
  assign n49059 = ~n24401 & n49058 ;
  assign n49060 = ~n24505 & n49059 ;
  assign n49062 = n49061 ^ n49060 ^ n41045 ;
  assign n49063 = n7515 & ~n19886 ;
  assign n49064 = ~n18052 & n49063 ;
  assign n49065 = n9291 & ~n30864 ;
  assign n49066 = ~n2504 & n49065 ;
  assign n49067 = n37438 & n44153 ;
  assign n49068 = ~n5633 & n27236 ;
  assign n49069 = n49068 ^ n13549 ^ 1'b0 ;
  assign n49070 = n25117 & ~n49069 ;
  assign n49071 = ~n49067 & n49070 ;
  assign n49072 = n41586 ^ n25598 ^ n744 ;
  assign n49073 = n7422 & ~n26488 ;
  assign n49074 = n27401 ^ n26860 ^ 1'b0 ;
  assign n49075 = n7551 & ~n49074 ;
  assign n49076 = n17170 | n23402 ;
  assign n49077 = n49076 ^ n19467 ^ 1'b0 ;
  assign n49078 = ( n34351 & n49075 ) | ( n34351 & n49077 ) | ( n49075 & n49077 ) ;
  assign n49079 = n15528 & ~n22216 ;
  assign n49080 = n49079 ^ n18361 ^ 1'b0 ;
  assign n49081 = ( ~n3913 & n13262 ) | ( ~n3913 & n49080 ) | ( n13262 & n49080 ) ;
  assign n49082 = ~n45217 & n49081 ;
  assign n49083 = n47583 ^ n12900 ^ 1'b0 ;
  assign n49084 = n44648 ^ n9825 ^ 1'b0 ;
  assign n49085 = ~n18441 & n49084 ;
  assign n49086 = n8087 & ~n14846 ;
  assign n49087 = n49086 ^ n23018 ^ 1'b0 ;
  assign n49088 = n28451 & ~n38807 ;
  assign n49089 = n11878 & ~n25474 ;
  assign n49090 = n6384 & n49089 ;
  assign n49091 = n24538 ^ n15975 ^ n5291 ;
  assign n49092 = n28244 ^ n21787 ^ 1'b0 ;
  assign n49093 = n18255 ^ n17381 ^ 1'b0 ;
  assign n49094 = n32828 ^ n2553 ^ 1'b0 ;
  assign n49095 = n49094 ^ n40620 ^ n34892 ;
  assign n49096 = ~n11631 & n21453 ;
  assign n49097 = ( n24161 & ~n38760 ) | ( n24161 & n49096 ) | ( ~n38760 & n49096 ) ;
  assign n49098 = n38517 ^ n21761 ^ 1'b0 ;
  assign n49099 = n4157 | n49098 ;
  assign n49100 = n49099 ^ n15476 ^ n5141 ;
  assign n49101 = n49100 ^ n16852 ^ 1'b0 ;
  assign n49102 = ( ~n17863 & n32303 ) | ( ~n17863 & n41709 ) | ( n32303 & n41709 ) ;
  assign n49103 = n49102 ^ n30037 ^ 1'b0 ;
  assign n49104 = n45487 ^ n41393 ^ n14462 ;
  assign n49105 = n49103 | n49104 ;
  assign n49106 = n7134 & n41277 ;
  assign n49107 = ( n3296 & n12430 ) | ( n3296 & n42336 ) | ( n12430 & n42336 ) ;
  assign n49108 = n49107 ^ n44792 ^ 1'b0 ;
  assign n49109 = n33425 & ~n45932 ;
  assign n49110 = ( n3791 & ~n3803 ) | ( n3791 & n12050 ) | ( ~n3803 & n12050 ) ;
  assign n49113 = n31727 ^ n13664 ^ n11781 ;
  assign n49111 = n19775 ^ n3503 ^ 1'b0 ;
  assign n49112 = n49111 ^ n30510 ^ n20683 ;
  assign n49114 = n49113 ^ n49112 ^ n47869 ;
  assign n49115 = n15017 & ~n23103 ;
  assign n49116 = n49115 ^ n25597 ^ 1'b0 ;
  assign n49117 = ( x215 & ~n8947 ) | ( x215 & n49116 ) | ( ~n8947 & n49116 ) ;
  assign n49118 = ~n4472 & n16018 ;
  assign n49119 = ( n9666 & n36990 ) | ( n9666 & n49118 ) | ( n36990 & n49118 ) ;
  assign n49120 = n17888 & ~n49119 ;
  assign n49121 = n27633 & ~n49120 ;
  assign n49122 = n49121 ^ n48223 ^ 1'b0 ;
  assign n49123 = n4361 ^ n992 ^ 1'b0 ;
  assign n49124 = n46334 ^ n35740 ^ n24735 ;
  assign n49125 = ( n10671 & ~n12317 ) | ( n10671 & n47362 ) | ( ~n12317 & n47362 ) ;
  assign n49127 = n13720 ^ n5214 ^ 1'b0 ;
  assign n49128 = ~n14395 & n49127 ;
  assign n49129 = n10066 & ~n34519 ;
  assign n49130 = ~n49128 & n49129 ;
  assign n49126 = ( ~n28528 & n29534 ) | ( ~n28528 & n37193 ) | ( n29534 & n37193 ) ;
  assign n49131 = n49130 ^ n49126 ^ 1'b0 ;
  assign n49132 = ( n3923 & n13242 ) | ( n3923 & ~n13568 ) | ( n13242 & ~n13568 ) ;
  assign n49133 = n5395 | n47015 ;
  assign n49134 = n640 & ~n24810 ;
  assign n49135 = n49134 ^ n27984 ^ 1'b0 ;
  assign n49136 = ~n9270 & n38337 ;
  assign n49137 = n3594 & ~n22592 ;
  assign n49138 = n11670 & n49137 ;
  assign n49139 = n41143 ^ n25096 ^ n23346 ;
  assign n49140 = n49139 ^ n22617 ^ 1'b0 ;
  assign n49142 = n34432 ^ n33832 ^ n26276 ;
  assign n49141 = n7944 | n42751 ;
  assign n49143 = n49142 ^ n49141 ^ 1'b0 ;
  assign n49144 = ( n14051 & n30987 ) | ( n14051 & ~n49143 ) | ( n30987 & ~n49143 ) ;
  assign n49145 = n37183 ^ n8805 ^ n3764 ;
  assign n49146 = n49145 ^ n23076 ^ n16377 ;
  assign n49147 = n24109 | n31788 ;
  assign n49148 = n49147 ^ n19391 ^ n3066 ;
  assign n49149 = n13101 ^ x20 ^ 1'b0 ;
  assign n49150 = n7466 & ~n49149 ;
  assign n49151 = ~n23749 & n49150 ;
  assign n49152 = n2107 & n18703 ;
  assign n49153 = ( ~n31167 & n49151 ) | ( ~n31167 & n49152 ) | ( n49151 & n49152 ) ;
  assign n49154 = n35122 ^ n20257 ^ 1'b0 ;
  assign n49155 = n6042 & n49154 ;
  assign n49156 = ( n15228 & n35908 ) | ( n15228 & n49155 ) | ( n35908 & n49155 ) ;
  assign n49157 = n22732 ^ n11366 ^ 1'b0 ;
  assign n49158 = n6729 | n49157 ;
  assign n49159 = ( ~n1548 & n17652 ) | ( ~n1548 & n38915 ) | ( n17652 & n38915 ) ;
  assign n49160 = ( n20047 & n37580 ) | ( n20047 & ~n49159 ) | ( n37580 & ~n49159 ) ;
  assign n49161 = ~n10386 & n49160 ;
  assign n49162 = ~n17453 & n20289 ;
  assign n49163 = n9690 ^ n4924 ^ 1'b0 ;
  assign n49170 = n37312 ^ n1873 ^ 1'b0 ;
  assign n49171 = n28010 & ~n49170 ;
  assign n49164 = n16101 ^ n11656 ^ n4479 ;
  assign n49165 = ~n27386 & n49164 ;
  assign n49166 = ~n22004 & n49165 ;
  assign n49167 = ( ~n5304 & n22938 ) | ( ~n5304 & n33425 ) | ( n22938 & n33425 ) ;
  assign n49168 = n22263 | n49167 ;
  assign n49169 = n49166 & ~n49168 ;
  assign n49172 = n49171 ^ n49169 ^ n29511 ;
  assign n49173 = ( n7726 & ~n17892 ) | ( n7726 & n49172 ) | ( ~n17892 & n49172 ) ;
  assign n49174 = ( n21198 & n37987 ) | ( n21198 & n39612 ) | ( n37987 & n39612 ) ;
  assign n49175 = n10233 & ~n12558 ;
  assign n49176 = ( n2925 & n4921 ) | ( n2925 & n10829 ) | ( n4921 & n10829 ) ;
  assign n49177 = ~n5185 & n5631 ;
  assign n49178 = ~n28933 & n49177 ;
  assign n49179 = n1056 | n4242 ;
  assign n49180 = n49178 & ~n49179 ;
  assign n49181 = n382 & ~n49180 ;
  assign n49182 = n49181 ^ n16599 ^ 1'b0 ;
  assign n49183 = ( n2428 & n49176 ) | ( n2428 & n49182 ) | ( n49176 & n49182 ) ;
  assign n49184 = n20948 ^ n17122 ^ n419 ;
  assign n49185 = n42190 ^ n27206 ^ 1'b0 ;
  assign n49186 = ~n2130 & n49185 ;
  assign n49187 = ( ~n2832 & n5281 ) | ( ~n2832 & n49186 ) | ( n5281 & n49186 ) ;
  assign n49188 = ( ~n41420 & n49184 ) | ( ~n41420 & n49187 ) | ( n49184 & n49187 ) ;
  assign n49189 = n3229 ^ n2475 ^ 1'b0 ;
  assign n49190 = n49189 ^ n1218 ^ 1'b0 ;
  assign n49191 = n26020 & n49190 ;
  assign n49192 = n22923 ^ n12672 ^ n12588 ;
  assign n49193 = n15359 & ~n49192 ;
  assign n49194 = n24522 ^ n6362 ^ 1'b0 ;
  assign n49195 = n26319 | n49194 ;
  assign n49196 = n3393 & ~n28034 ;
  assign n49197 = n12527 & ~n35729 ;
  assign n49198 = ~n6186 & n49197 ;
  assign n49199 = n36697 & n49198 ;
  assign n49200 = n28238 | n44254 ;
  assign n49201 = n49200 ^ n16873 ^ 1'b0 ;
  assign n49202 = ( ~n32267 & n41820 ) | ( ~n32267 & n49201 ) | ( n41820 & n49201 ) ;
  assign n49203 = ( n8670 & n48345 ) | ( n8670 & ~n48624 ) | ( n48345 & ~n48624 ) ;
  assign n49205 = n6238 | n25576 ;
  assign n49204 = n12617 & n23536 ;
  assign n49206 = n49205 ^ n49204 ^ 1'b0 ;
  assign n49207 = ~n8027 & n41891 ;
  assign n49208 = ~n38734 & n49207 ;
  assign n49209 = n49208 ^ n46627 ^ 1'b0 ;
  assign n49210 = n44510 & ~n49209 ;
  assign n49214 = n24889 ^ n14288 ^ n12282 ;
  assign n49213 = n34566 ^ n16077 ^ 1'b0 ;
  assign n49211 = n35467 ^ n18389 ^ 1'b0 ;
  assign n49212 = ~n24595 & n49211 ;
  assign n49215 = n49214 ^ n49213 ^ n49212 ;
  assign n49216 = ~n42557 & n49215 ;
  assign n49217 = n49216 ^ n19445 ^ 1'b0 ;
  assign n49218 = n36085 ^ n17524 ^ n3413 ;
  assign n49219 = ( n5658 & n30758 ) | ( n5658 & ~n49218 ) | ( n30758 & ~n49218 ) ;
  assign n49220 = ( ~n6851 & n41944 ) | ( ~n6851 & n49219 ) | ( n41944 & n49219 ) ;
  assign n49221 = n13942 ^ n4208 ^ 1'b0 ;
  assign n49222 = n43979 ^ n38194 ^ 1'b0 ;
  assign n49223 = n35794 & ~n49222 ;
  assign n49224 = n49223 ^ n12233 ^ 1'b0 ;
  assign n49225 = ~n6512 & n49224 ;
  assign n49226 = n46407 ^ n24439 ^ n5461 ;
  assign n49227 = n6216 & n49226 ;
  assign n49228 = n34265 | n49227 ;
  assign n49229 = n2735 & ~n49228 ;
  assign n49230 = ( n5474 & n25432 ) | ( n5474 & ~n49229 ) | ( n25432 & ~n49229 ) ;
  assign n49231 = n44833 ^ n703 ^ 1'b0 ;
  assign n49232 = n14288 & n49231 ;
  assign n49233 = ~n5300 & n14558 ;
  assign n49234 = n49233 ^ n40935 ^ n18683 ;
  assign n49235 = ( n2684 & n12363 ) | ( n2684 & n41148 ) | ( n12363 & n41148 ) ;
  assign n49236 = n49235 ^ n20661 ^ 1'b0 ;
  assign n49237 = n49234 & n49236 ;
  assign n49238 = n5641 | n26114 ;
  assign n49239 = n49238 ^ n35479 ^ 1'b0 ;
  assign n49240 = n36318 ^ n35382 ^ n6369 ;
  assign n49241 = n9211 & n49240 ;
  assign n49242 = n35395 & n49241 ;
  assign n49243 = n22014 & n33391 ;
  assign n49244 = n33115 ^ n8226 ^ 1'b0 ;
  assign n49245 = n49244 ^ n31804 ^ n24551 ;
  assign n49246 = ( ~n2845 & n31505 ) | ( ~n2845 & n43234 ) | ( n31505 & n43234 ) ;
  assign n49247 = n42996 ^ n39848 ^ n10334 ;
  assign n49248 = n406 & ~n35617 ;
  assign n49249 = ~n2247 & n49248 ;
  assign n49250 = ( n12794 & n16401 ) | ( n12794 & n49249 ) | ( n16401 & n49249 ) ;
  assign n49251 = n12830 ^ n10816 ^ 1'b0 ;
  assign n49252 = n33443 ^ n17420 ^ n8282 ;
  assign n49253 = ( n6568 & ~n27691 ) | ( n6568 & n48543 ) | ( ~n27691 & n48543 ) ;
  assign n49254 = n10324 | n11507 ;
  assign n49255 = n49253 | n49254 ;
  assign n49256 = n23258 & n35674 ;
  assign n49257 = n12076 & n49256 ;
  assign n49258 = n19261 ^ n15185 ^ n2211 ;
  assign n49259 = n21952 & ~n47352 ;
  assign n49260 = n10908 & n49259 ;
  assign n49261 = n49258 & n49260 ;
  assign n49265 = n18304 ^ n15453 ^ 1'b0 ;
  assign n49263 = n12394 ^ n550 ^ 1'b0 ;
  assign n49264 = n26171 & ~n49263 ;
  assign n49262 = ( ~n4450 & n10873 ) | ( ~n4450 & n14546 ) | ( n10873 & n14546 ) ;
  assign n49266 = n49265 ^ n49264 ^ n49262 ;
  assign n49267 = ( ~n27792 & n36103 ) | ( ~n27792 & n44795 ) | ( n36103 & n44795 ) ;
  assign n49268 = ( ~n26289 & n35133 ) | ( ~n26289 & n39314 ) | ( n35133 & n39314 ) ;
  assign n49269 = n49268 ^ n22829 ^ n949 ;
  assign n49270 = n49269 ^ n44494 ^ n37559 ;
  assign n49271 = n23212 ^ n16114 ^ n15466 ;
  assign n49272 = ~n4636 & n19895 ;
  assign n49273 = ( n4810 & ~n5482 ) | ( n4810 & n24048 ) | ( ~n5482 & n24048 ) ;
  assign n49274 = n20477 & n49273 ;
  assign n49276 = ~n3809 & n27157 ;
  assign n49277 = n23661 & n49276 ;
  assign n49275 = ~n11623 & n32951 ;
  assign n49278 = n49277 ^ n49275 ^ 1'b0 ;
  assign n49279 = n23590 | n29133 ;
  assign n49280 = n49279 ^ n38830 ^ 1'b0 ;
  assign n49281 = n17593 ^ n13766 ^ 1'b0 ;
  assign n49282 = n3775 | n49281 ;
  assign n49283 = n49282 ^ n48734 ^ 1'b0 ;
  assign n49284 = n49283 ^ n14973 ^ 1'b0 ;
  assign n49285 = n17106 | n49284 ;
  assign n49286 = n4730 | n30002 ;
  assign n49287 = n49286 ^ n39335 ^ 1'b0 ;
  assign n49288 = ( n3478 & ~n7408 ) | ( n3478 & n11149 ) | ( ~n7408 & n11149 ) ;
  assign n49289 = n25908 & n49288 ;
  assign n49290 = ( n4577 & n15085 ) | ( n4577 & n29501 ) | ( n15085 & n29501 ) ;
  assign n49291 = n36622 ^ n12532 ^ 1'b0 ;
  assign n49292 = n49291 ^ n17438 ^ 1'b0 ;
  assign n49293 = n49290 & ~n49292 ;
  assign n49294 = n25334 ^ n802 ^ 1'b0 ;
  assign n49295 = ~n22623 & n49294 ;
  assign n49296 = n43438 & n49295 ;
  assign n49297 = ( n22564 & n49293 ) | ( n22564 & n49296 ) | ( n49293 & n49296 ) ;
  assign n49299 = n5242 | n19257 ;
  assign n49300 = n49299 ^ n10956 ^ 1'b0 ;
  assign n49298 = n17888 ^ n10400 ^ n8472 ;
  assign n49301 = n49300 ^ n49298 ^ n2629 ;
  assign n49302 = ~n19132 & n37959 ;
  assign n49303 = n42904 ^ n8923 ^ 1'b0 ;
  assign n49304 = n1543 & ~n49303 ;
  assign n49305 = n19816 ^ n7639 ^ 1'b0 ;
  assign n49306 = ~n13252 & n49305 ;
  assign n49307 = n11005 & ~n21568 ;
  assign n49308 = n49307 ^ n45116 ^ 1'b0 ;
  assign n49309 = n3395 & n11345 ;
  assign n49310 = n49309 ^ n36031 ^ 1'b0 ;
  assign n49311 = n9455 | n49310 ;
  assign n49312 = n1758 & ~n39117 ;
  assign n49313 = n49312 ^ n30384 ^ 1'b0 ;
  assign n49314 = ( n15534 & ~n47086 ) | ( n15534 & n49313 ) | ( ~n47086 & n49313 ) ;
  assign n49315 = n37603 ^ n1776 ^ 1'b0 ;
  assign n49316 = n49315 ^ n44821 ^ n2488 ;
  assign n49317 = n31357 ^ n27682 ^ n1629 ;
  assign n49318 = n6662 ^ n1398 ^ n598 ;
  assign n49319 = n12372 ^ n5533 ^ 1'b0 ;
  assign n49320 = n2295 & ~n24941 ;
  assign n49321 = n49320 ^ n27402 ^ 1'b0 ;
  assign n49322 = n4043 & n47070 ;
  assign n49323 = ~n27471 & n49322 ;
  assign n49325 = ~n6097 & n19438 ;
  assign n49324 = n1789 | n8716 ;
  assign n49326 = n49325 ^ n49324 ^ 1'b0 ;
  assign n49327 = n40267 ^ n25175 ^ 1'b0 ;
  assign n49328 = ( n15973 & n39600 ) | ( n15973 & n49327 ) | ( n39600 & n49327 ) ;
  assign n49329 = n26390 ^ n19107 ^ n3365 ;
  assign n49330 = n47095 ^ x206 ^ 1'b0 ;
  assign n49331 = n6000 & ~n49330 ;
  assign n49332 = ( n9758 & ~n44357 ) | ( n9758 & n49331 ) | ( ~n44357 & n49331 ) ;
  assign n49333 = ~n9366 & n11303 ;
  assign n49334 = n23216 & ~n49333 ;
  assign n49335 = ~n43734 & n49334 ;
  assign n49336 = n4564 | n5112 ;
  assign n49337 = n16336 & ~n49336 ;
  assign n49338 = n49337 ^ n3041 ^ 1'b0 ;
  assign n49339 = n37233 & n42881 ;
  assign n49340 = n49339 ^ n36302 ^ 1'b0 ;
  assign n49342 = n14107 ^ n4227 ^ 1'b0 ;
  assign n49341 = ~n10934 & n30240 ;
  assign n49343 = n49342 ^ n49341 ^ 1'b0 ;
  assign n49344 = ( n1656 & n39891 ) | ( n1656 & ~n49343 ) | ( n39891 & ~n49343 ) ;
  assign n49345 = n38533 ^ n30103 ^ n7653 ;
  assign n49346 = n10954 ^ n6492 ^ 1'b0 ;
  assign n49347 = n38628 ^ n23630 ^ 1'b0 ;
  assign n49348 = ( n24087 & n49346 ) | ( n24087 & n49347 ) | ( n49346 & n49347 ) ;
  assign n49349 = n47584 ^ n9738 ^ n8458 ;
  assign n49350 = ( ~n21105 & n36532 ) | ( ~n21105 & n49349 ) | ( n36532 & n49349 ) ;
  assign n49351 = ( n9349 & n19857 ) | ( n9349 & n34867 ) | ( n19857 & n34867 ) ;
  assign n49352 = n2112 | n18723 ;
  assign n49353 = n49351 & ~n49352 ;
  assign n49354 = n33647 | n40259 ;
  assign n49355 = n49353 & ~n49354 ;
  assign n49356 = n40075 & n42157 ;
  assign n49357 = n22901 | n46391 ;
  assign n49358 = n2386 & ~n17885 ;
  assign n49359 = n37645 & n49358 ;
  assign n49360 = ~n32319 & n36851 ;
  assign n49362 = n7000 & ~n14095 ;
  assign n49361 = ~n7296 & n22966 ;
  assign n49363 = n49362 ^ n49361 ^ 1'b0 ;
  assign n49364 = n49363 ^ n34510 ^ 1'b0 ;
  assign n49365 = n36977 ^ n19266 ^ 1'b0 ;
  assign n49366 = ( ~n430 & n3844 ) | ( ~n430 & n6869 ) | ( n3844 & n6869 ) ;
  assign n49367 = ( n25388 & n35447 ) | ( n25388 & ~n49366 ) | ( n35447 & ~n49366 ) ;
  assign n49368 = n3147 & ~n20026 ;
  assign n49369 = n41190 ^ n16727 ^ 1'b0 ;
  assign n49370 = ( ~n28175 & n38755 ) | ( ~n28175 & n49369 ) | ( n38755 & n49369 ) ;
  assign n49371 = n9480 & ~n49370 ;
  assign n49372 = n8438 & n49371 ;
  assign n49373 = n19504 & ~n48065 ;
  assign n49374 = ( n6408 & ~n15456 ) | ( n6408 & n20948 ) | ( ~n15456 & n20948 ) ;
  assign n49375 = n49374 ^ n7489 ^ 1'b0 ;
  assign n49376 = n25662 ^ n10783 ^ 1'b0 ;
  assign n49377 = n4198 & n49376 ;
  assign n49378 = ( n6431 & ~n10985 ) | ( n6431 & n32513 ) | ( ~n10985 & n32513 ) ;
  assign n49380 = ( n1773 & n2104 ) | ( n1773 & ~n15990 ) | ( n2104 & ~n15990 ) ;
  assign n49379 = n32416 & ~n39315 ;
  assign n49381 = n49380 ^ n49379 ^ 1'b0 ;
  assign n49382 = ~n29329 & n41923 ;
  assign n49383 = n44062 & n49382 ;
  assign n49384 = n8580 & ~n42175 ;
  assign n49385 = n21742 & n24966 ;
  assign n49389 = ~n3043 & n25557 ;
  assign n49390 = n5387 & ~n27276 ;
  assign n49391 = ~n49389 & n49390 ;
  assign n49386 = n8686 & ~n8832 ;
  assign n49387 = n49386 ^ n11437 ^ 1'b0 ;
  assign n49388 = n49387 ^ n38097 ^ n19077 ;
  assign n49392 = n49391 ^ n49388 ^ n9186 ;
  assign n49393 = n27832 ^ n5344 ^ 1'b0 ;
  assign n49394 = n49393 ^ n44808 ^ n29018 ;
  assign n49395 = n18842 ^ n17407 ^ n6835 ;
  assign n49396 = n49395 ^ n48160 ^ n46036 ;
  assign n49397 = n36345 ^ n32787 ^ 1'b0 ;
  assign n49398 = n33075 | n49397 ;
  assign n49399 = ( ~n30241 & n31975 ) | ( ~n30241 & n49398 ) | ( n31975 & n49398 ) ;
  assign n49400 = n46267 ^ n29708 ^ 1'b0 ;
  assign n49401 = n49400 ^ n37874 ^ n14571 ;
  assign n49402 = n9262 | n43040 ;
  assign n49403 = n4283 | n25044 ;
  assign n49404 = n419 | n29756 ;
  assign n49405 = n49404 ^ n3516 ^ 1'b0 ;
  assign n49406 = n10936 ^ n5803 ^ n5715 ;
  assign n49407 = n10012 ^ n6336 ^ 1'b0 ;
  assign n49408 = n49406 & ~n49407 ;
  assign n49409 = ~n33733 & n37144 ;
  assign n49410 = ~n27496 & n49409 ;
  assign n49411 = n4119 & ~n15730 ;
  assign n49412 = ~n1617 & n34332 ;
  assign n49413 = ~n49411 & n49412 ;
  assign n49414 = n14873 ^ n7238 ^ 1'b0 ;
  assign n49415 = ( ~n2089 & n2267 ) | ( ~n2089 & n49414 ) | ( n2267 & n49414 ) ;
  assign n49416 = n49415 ^ n20437 ^ n1273 ;
  assign n49417 = n49413 | n49416 ;
  assign n49418 = n20613 ^ n9876 ^ n6964 ;
  assign n49419 = ( n2149 & n4941 ) | ( n2149 & n49418 ) | ( n4941 & n49418 ) ;
  assign n49420 = ( n14365 & ~n19095 ) | ( n14365 & n22613 ) | ( ~n19095 & n22613 ) ;
  assign n49421 = n18761 ^ n10761 ^ n6320 ;
  assign n49422 = n49421 ^ n28166 ^ 1'b0 ;
  assign n49423 = n18104 & n49422 ;
  assign n49424 = ~n32044 & n49423 ;
  assign n49425 = n8847 & ~n40567 ;
  assign n49426 = ~n18707 & n49425 ;
  assign n49427 = n49426 ^ n40247 ^ 1'b0 ;
  assign n49428 = n17216 ^ n11149 ^ 1'b0 ;
  assign n49429 = ~n10657 & n49428 ;
  assign n49430 = n49429 ^ n46342 ^ 1'b0 ;
  assign n49431 = ~n24712 & n40445 ;
  assign n49432 = n49430 & n49431 ;
  assign n49433 = n7339 | n10699 ;
  assign n49434 = n49433 ^ n20269 ^ 1'b0 ;
  assign n49435 = n27312 | n48811 ;
  assign n49436 = n49435 ^ n32033 ^ 1'b0 ;
  assign n49437 = ~n10930 & n11061 ;
  assign n49438 = n49437 ^ n39168 ^ n14320 ;
  assign n49439 = n31406 ^ n8468 ^ 1'b0 ;
  assign n49440 = n9699 & ~n49439 ;
  assign n49441 = ~n10481 & n20343 ;
  assign n49442 = ~n49440 & n49441 ;
  assign n49443 = n49442 ^ n18550 ^ 1'b0 ;
  assign n49444 = n7471 ^ n3144 ^ 1'b0 ;
  assign n49445 = ( n5585 & n40677 ) | ( n5585 & n43799 ) | ( n40677 & n43799 ) ;
  assign n49446 = n49445 ^ n7201 ^ n2175 ;
  assign n49447 = n49446 ^ n23761 ^ 1'b0 ;
  assign n49448 = n45140 ^ n20911 ^ 1'b0 ;
  assign n49449 = ~n16170 & n49448 ;
  assign n49450 = n20168 ^ n731 ^ 1'b0 ;
  assign n49451 = ~n41541 & n49450 ;
  assign n49453 = n17015 ^ n12498 ^ 1'b0 ;
  assign n49454 = n41497 & ~n49453 ;
  assign n49452 = n13263 | n30749 ;
  assign n49455 = n49454 ^ n49452 ^ 1'b0 ;
  assign n49456 = n3466 & ~n47516 ;
  assign n49457 = ~n20208 & n49456 ;
  assign n49458 = n8817 & ~n46656 ;
  assign n49459 = n10780 & n49458 ;
  assign n49460 = ( n10479 & ~n24789 ) | ( n10479 & n49459 ) | ( ~n24789 & n49459 ) ;
  assign n49461 = ( n10725 & ~n15632 ) | ( n10725 & n38513 ) | ( ~n15632 & n38513 ) ;
  assign n49462 = ~n10420 & n14265 ;
  assign n49463 = ( ~n10134 & n21598 ) | ( ~n10134 & n49462 ) | ( n21598 & n49462 ) ;
  assign n49464 = n15768 ^ n7801 ^ 1'b0 ;
  assign n49465 = n28716 & n49464 ;
  assign n49466 = n31916 ^ n27631 ^ n15743 ;
  assign n49467 = n426 & ~n49466 ;
  assign n49468 = ~n1086 & n49467 ;
  assign n49469 = ( ~n1726 & n45670 ) | ( ~n1726 & n49468 ) | ( n45670 & n49468 ) ;
  assign n49470 = n31442 ^ n12124 ^ 1'b0 ;
  assign n49471 = n28596 ^ n4624 ^ 1'b0 ;
  assign n49472 = n49470 & n49471 ;
  assign n49474 = n25600 ^ n18402 ^ n16340 ;
  assign n49475 = n25685 | n49474 ;
  assign n49473 = n18070 & ~n42325 ;
  assign n49476 = n49475 ^ n49473 ^ 1'b0 ;
  assign n49477 = n16561 & n31433 ;
  assign n49478 = ~n7308 & n21116 ;
  assign n49479 = ~n8766 & n49478 ;
  assign n49480 = n4819 & n9154 ;
  assign n49481 = n49480 ^ n17872 ^ 1'b0 ;
  assign n49482 = ( n18085 & n29825 ) | ( n18085 & n49481 ) | ( n29825 & n49481 ) ;
  assign n49483 = ~n15273 & n43818 ;
  assign n49484 = n38464 ^ n14685 ^ n12891 ;
  assign n49485 = n40499 ^ n30944 ^ 1'b0 ;
  assign n49486 = n31224 ^ n25821 ^ n15660 ;
  assign n49487 = n2175 & n6502 ;
  assign n49488 = n19381 ^ n7959 ^ 1'b0 ;
  assign n49489 = n11831 & n49488 ;
  assign n49490 = ~n6637 & n18861 ;
  assign n49491 = n49490 ^ n2630 ^ 1'b0 ;
  assign n49492 = ( n9258 & ~n29973 ) | ( n9258 & n45622 ) | ( ~n29973 & n45622 ) ;
  assign n49493 = n32375 ^ n22431 ^ n14174 ;
  assign n49494 = n19105 & ~n23420 ;
  assign n49495 = ( n12101 & n48510 ) | ( n12101 & ~n49494 ) | ( n48510 & ~n49494 ) ;
  assign n49496 = n42380 ^ n14858 ^ n4982 ;
  assign n49497 = n3699 & ~n31926 ;
  assign n49498 = n49497 ^ n10120 ^ 1'b0 ;
  assign n49502 = ( ~n13141 & n17779 ) | ( ~n13141 & n33137 ) | ( n17779 & n33137 ) ;
  assign n49499 = n38825 ^ n19993 ^ 1'b0 ;
  assign n49500 = n49499 ^ n46525 ^ n28437 ;
  assign n49501 = ~n7767 & n49500 ;
  assign n49503 = n49502 ^ n49501 ^ 1'b0 ;
  assign n49504 = n19855 & ~n20595 ;
  assign n49505 = n4004 & ~n15305 ;
  assign n49506 = n49505 ^ n20460 ^ 1'b0 ;
  assign n49508 = n25148 ^ n19795 ^ 1'b0 ;
  assign n49509 = n21825 | n49508 ;
  assign n49510 = n11517 & n49509 ;
  assign n49507 = n6553 & n49259 ;
  assign n49511 = n49510 ^ n49507 ^ 1'b0 ;
  assign n49512 = n44045 ^ n33971 ^ 1'b0 ;
  assign n49513 = ( n39152 & n49511 ) | ( n39152 & ~n49512 ) | ( n49511 & ~n49512 ) ;
  assign n49514 = n44832 ^ n41761 ^ 1'b0 ;
  assign n49515 = ( n8222 & n8964 ) | ( n8222 & n15304 ) | ( n8964 & n15304 ) ;
  assign n49516 = ( n19544 & n35652 ) | ( n19544 & ~n44513 ) | ( n35652 & ~n44513 ) ;
  assign n49517 = n19154 ^ n865 ^ 1'b0 ;
  assign n49518 = n25531 | n49517 ;
  assign n49519 = n24311 & ~n40875 ;
  assign n49520 = n4783 & n21527 ;
  assign n49521 = ~n14712 & n49520 ;
  assign n49522 = n49521 ^ n28006 ^ n18903 ;
  assign n49523 = n41074 ^ n29175 ^ 1'b0 ;
  assign n49524 = ~n10466 & n49523 ;
  assign n49525 = n49524 ^ n42862 ^ 1'b0 ;
  assign n49526 = n16001 ^ n10363 ^ n866 ;
  assign n49528 = n2158 ^ n1586 ^ 1'b0 ;
  assign n49529 = n2068 & ~n49528 ;
  assign n49527 = n4187 & n24662 ;
  assign n49530 = n49529 ^ n49527 ^ 1'b0 ;
  assign n49531 = n42613 ^ n37160 ^ n31975 ;
  assign n49532 = ~n24999 & n39401 ;
  assign n49533 = n17400 | n49532 ;
  assign n49534 = n33130 & ~n49533 ;
  assign n49535 = n30366 ^ n23668 ^ 1'b0 ;
  assign n49536 = n47090 | n49535 ;
  assign n49537 = n49536 ^ n48180 ^ 1'b0 ;
  assign n49540 = n5226 & ~n33977 ;
  assign n49541 = n49540 ^ n8910 ^ 1'b0 ;
  assign n49538 = n682 | n5470 ;
  assign n49539 = n48092 | n49538 ;
  assign n49542 = n49541 ^ n49539 ^ 1'b0 ;
  assign n49543 = ~n12891 & n49542 ;
  assign n49544 = n19598 ^ n3430 ^ n870 ;
  assign n49545 = ( n4185 & n19236 ) | ( n4185 & ~n41295 ) | ( n19236 & ~n41295 ) ;
  assign n49546 = n42389 ^ n8435 ^ 1'b0 ;
  assign n49547 = n29437 ^ n17103 ^ n2301 ;
  assign n49548 = ~n1754 & n49547 ;
  assign n49549 = n49548 ^ n31359 ^ 1'b0 ;
  assign n49550 = ( n13960 & n49546 ) | ( n13960 & n49549 ) | ( n49546 & n49549 ) ;
  assign n49551 = n49550 ^ n23146 ^ n7282 ;
  assign n49552 = n13582 ^ n11508 ^ 1'b0 ;
  assign n49553 = ( n11837 & n29176 ) | ( n11837 & n35330 ) | ( n29176 & n35330 ) ;
  assign n49554 = n17230 | n49553 ;
  assign n49555 = n35870 & ~n49554 ;
  assign n49556 = n6132 & n14120 ;
  assign n49557 = n49555 & n49556 ;
  assign n49558 = n37971 | n38206 ;
  assign n49559 = n49558 ^ n15943 ^ 1'b0 ;
  assign n49560 = n1338 & n34786 ;
  assign n49561 = n49560 ^ n41537 ^ 1'b0 ;
  assign n49562 = ( n6952 & n19363 ) | ( n6952 & ~n30808 ) | ( n19363 & ~n30808 ) ;
  assign n49563 = ( n15649 & ~n21069 ) | ( n15649 & n41954 ) | ( ~n21069 & n41954 ) ;
  assign n49564 = n6388 ^ n4240 ^ 1'b0 ;
  assign n49565 = ( n19073 & ~n23285 ) | ( n19073 & n49564 ) | ( ~n23285 & n49564 ) ;
  assign n49566 = n1359 | n49565 ;
  assign n49567 = n9874 & n10772 ;
  assign n49568 = ~n25538 & n49567 ;
  assign n49569 = n49568 ^ n26798 ^ 1'b0 ;
  assign n49570 = n37318 ^ n26388 ^ n5389 ;
  assign n49571 = n10287 | n32171 ;
  assign n49572 = n28538 | n49571 ;
  assign n49575 = n22285 ^ n963 ^ 1'b0 ;
  assign n49573 = n18371 ^ n1535 ^ x182 ;
  assign n49574 = ( ~n15678 & n20031 ) | ( ~n15678 & n49573 ) | ( n20031 & n49573 ) ;
  assign n49576 = n49575 ^ n49574 ^ n2908 ;
  assign n49577 = n49576 ^ n38658 ^ 1'b0 ;
  assign n49578 = n37898 & ~n49577 ;
  assign n49579 = n20253 ^ n8497 ^ 1'b0 ;
  assign n49580 = ~n13638 & n49579 ;
  assign n49581 = n46273 ^ n32211 ^ n7135 ;
  assign n49582 = n1674 | n6823 ;
  assign n49583 = n49581 | n49582 ;
  assign n49584 = ~n9899 & n32090 ;
  assign n49585 = n49584 ^ n11136 ^ 1'b0 ;
  assign n49586 = n36437 ^ n16406 ^ n11434 ;
  assign n49587 = ~n2684 & n14632 ;
  assign n49588 = n14518 & ~n49587 ;
  assign n49589 = n23731 & n35664 ;
  assign n49590 = ( ~n3754 & n16906 ) | ( ~n3754 & n22563 ) | ( n16906 & n22563 ) ;
  assign n49591 = n49590 ^ n11606 ^ n5730 ;
  assign n49593 = n23084 & ~n46150 ;
  assign n49594 = n1806 & n46958 ;
  assign n49595 = n49593 & n49594 ;
  assign n49592 = ( n11513 & n19458 ) | ( n11513 & ~n24284 ) | ( n19458 & ~n24284 ) ;
  assign n49596 = n49595 ^ n49592 ^ n31097 ;
  assign n49597 = n21389 & n24326 ;
  assign n49598 = n49597 ^ n6492 ^ 1'b0 ;
  assign n49599 = ( ~n9540 & n49596 ) | ( ~n9540 & n49598 ) | ( n49596 & n49598 ) ;
  assign n49600 = ~n12236 & n14873 ;
  assign n49601 = n4214 & n49600 ;
  assign n49602 = n29553 & ~n49601 ;
  assign n49603 = ~n19684 & n49602 ;
  assign n49604 = n49603 ^ n27880 ^ 1'b0 ;
  assign n49605 = n8250 & n15528 ;
  assign n49606 = n49605 ^ n21340 ^ 1'b0 ;
  assign n49607 = n43109 ^ n6844 ^ 1'b0 ;
  assign n49608 = n49606 & n49607 ;
  assign n49609 = n36150 & n49608 ;
  assign n49610 = ~n17823 & n49609 ;
  assign n49611 = n8500 | n26732 ;
  assign n49612 = ~n925 & n2408 ;
  assign n49613 = n8828 & n49612 ;
  assign n49614 = ~n19306 & n49613 ;
  assign n49615 = n26761 ^ n26703 ^ 1'b0 ;
  assign n49616 = n49614 | n49615 ;
  assign n49617 = n22397 ^ n6379 ^ n2858 ;
  assign n49618 = n33486 ^ n11418 ^ 1'b0 ;
  assign n49619 = n14293 & ~n49618 ;
  assign n49620 = n49619 ^ n43162 ^ n13778 ;
  assign n49621 = ( n10265 & n18073 ) | ( n10265 & ~n26648 ) | ( n18073 & ~n26648 ) ;
  assign n49622 = n49621 ^ n24844 ^ n5089 ;
  assign n49623 = ~n15440 & n19803 ;
  assign n49624 = n49623 ^ n9211 ^ 1'b0 ;
  assign n49625 = n11564 & n23645 ;
  assign n49626 = n6417 | n16472 ;
  assign n49627 = n49626 ^ n17747 ^ 1'b0 ;
  assign n49628 = n44547 ^ n25627 ^ n6235 ;
  assign n49629 = n40319 & n49628 ;
  assign n49630 = n6047 ^ n5671 ^ 1'b0 ;
  assign n49631 = n8350 | n27616 ;
  assign n49632 = n6202 & ~n49631 ;
  assign n49633 = n5924 | n15727 ;
  assign n49634 = n49633 ^ n32768 ^ 1'b0 ;
  assign n49635 = n49634 ^ n8220 ^ 1'b0 ;
  assign n49636 = n16892 & ~n49635 ;
  assign n49637 = n49636 ^ n15797 ^ 1'b0 ;
  assign n49638 = ( ~n1850 & n29937 ) | ( ~n1850 & n31124 ) | ( n29937 & n31124 ) ;
  assign n49639 = n49638 ^ n37208 ^ 1'b0 ;
  assign n49640 = n16675 & n39663 ;
  assign n49641 = ( ~n6476 & n8811 ) | ( ~n6476 & n16603 ) | ( n8811 & n16603 ) ;
  assign n49642 = n30229 | n41270 ;
  assign n49643 = n1427 & ~n2349 ;
  assign n49644 = n49643 ^ n23704 ^ 1'b0 ;
  assign n49645 = n38448 ^ n7218 ^ 1'b0 ;
  assign n49646 = n28500 ^ n470 ^ 1'b0 ;
  assign n49647 = n49645 & n49646 ;
  assign n49648 = ( n2110 & n2175 ) | ( n2110 & n7024 ) | ( n2175 & n7024 ) ;
  assign n49649 = n49648 ^ n42887 ^ 1'b0 ;
  assign n49650 = ~n31753 & n49649 ;
  assign n49653 = n8698 ^ n5479 ^ 1'b0 ;
  assign n49652 = ( n11614 & ~n14737 ) | ( n11614 & n22621 ) | ( ~n14737 & n22621 ) ;
  assign n49651 = ( ~n2463 & n40743 ) | ( ~n2463 & n42249 ) | ( n40743 & n42249 ) ;
  assign n49654 = n49653 ^ n49652 ^ n49651 ;
  assign n49655 = n45485 ^ n16075 ^ n8108 ;
  assign n49656 = n7176 | n20791 ;
  assign n49657 = n49656 ^ n22308 ^ 1'b0 ;
  assign n49658 = n31089 ^ n8739 ^ 1'b0 ;
  assign n49659 = ~n13764 & n49658 ;
  assign n49660 = n20192 & n30393 ;
  assign n49661 = n49660 ^ n4224 ^ 1'b0 ;
  assign n49662 = n14755 ^ n9580 ^ 1'b0 ;
  assign n49663 = ~n13804 & n49662 ;
  assign n49664 = ( n33347 & ~n36843 ) | ( n33347 & n49663 ) | ( ~n36843 & n49663 ) ;
  assign n49667 = n33180 ^ n27707 ^ 1'b0 ;
  assign n49665 = ( n1913 & ~n2659 ) | ( n1913 & n4550 ) | ( ~n2659 & n4550 ) ;
  assign n49666 = n49665 ^ n48005 ^ 1'b0 ;
  assign n49668 = n49667 ^ n49666 ^ n2464 ;
  assign n49669 = ( n5815 & n25114 ) | ( n5815 & n37082 ) | ( n25114 & n37082 ) ;
  assign n49670 = ~n25252 & n43301 ;
  assign n49671 = n35490 ^ n12677 ^ 1'b0 ;
  assign n49672 = n7551 | n14314 ;
  assign n49673 = n49671 & ~n49672 ;
  assign n49674 = n45021 ^ n751 ^ 1'b0 ;
  assign n49675 = n32033 & ~n49674 ;
  assign n49676 = n21317 ^ n12142 ^ n7732 ;
  assign n49677 = n1044 & ~n49676 ;
  assign n49678 = ~n11696 & n18786 ;
  assign n49679 = n14603 & n49678 ;
  assign n49680 = n18729 | n49679 ;
  assign n49681 = ( ~n14624 & n35158 ) | ( ~n14624 & n49680 ) | ( n35158 & n49680 ) ;
  assign n49682 = n3511 & ~n10834 ;
  assign n49683 = n15433 | n49682 ;
  assign n49684 = n37647 ^ n34794 ^ n26612 ;
  assign n49685 = n33707 & ~n34018 ;
  assign n49686 = n10185 ^ n326 ^ 1'b0 ;
  assign n49687 = ( ~n1352 & n11508 ) | ( ~n1352 & n24551 ) | ( n11508 & n24551 ) ;
  assign n49688 = n49687 ^ n25549 ^ n18976 ;
  assign n49689 = ~n49686 & n49688 ;
  assign n49690 = n26687 ^ n16186 ^ 1'b0 ;
  assign n49691 = n49689 & n49690 ;
  assign n49692 = ( ~n6714 & n8405 ) | ( ~n6714 & n9109 ) | ( n8405 & n9109 ) ;
  assign n49693 = n3369 & n9625 ;
  assign n49694 = n49693 ^ n545 ^ 1'b0 ;
  assign n49695 = n49694 ^ n2893 ^ n1971 ;
  assign n49696 = n22270 ^ n5755 ^ 1'b0 ;
  assign n49697 = n23780 | n49696 ;
  assign n49698 = ( n15115 & n18748 ) | ( n15115 & ~n49697 ) | ( n18748 & ~n49697 ) ;
  assign n49699 = ( ~n7844 & n15603 ) | ( ~n7844 & n21252 ) | ( n15603 & n21252 ) ;
  assign n49700 = ( ~n18005 & n33792 ) | ( ~n18005 & n49699 ) | ( n33792 & n49699 ) ;
  assign n49701 = n24262 ^ n23493 ^ 1'b0 ;
  assign n49702 = n2682 & n49701 ;
  assign n49703 = n14808 ^ n2691 ^ 1'b0 ;
  assign n49704 = ~n35836 & n49703 ;
  assign n49705 = ( n40171 & n49702 ) | ( n40171 & ~n49704 ) | ( n49702 & ~n49704 ) ;
  assign n49706 = n388 | n28051 ;
  assign n49707 = n49706 ^ x193 ^ 1'b0 ;
  assign n49708 = n3962 & ~n33479 ;
  assign n49709 = ~n49707 & n49708 ;
  assign n49710 = n1630 | n3656 ;
  assign n49711 = n17910 & ~n49710 ;
  assign n49712 = n13929 | n17578 ;
  assign n49713 = n49712 ^ n15646 ^ 1'b0 ;
  assign n49714 = ( ~n17807 & n44022 ) | ( ~n17807 & n49713 ) | ( n44022 & n49713 ) ;
  assign n49715 = n44821 & ~n49714 ;
  assign n49716 = n49715 ^ n10038 ^ 1'b0 ;
  assign n49717 = ( n3782 & ~n10575 ) | ( n3782 & n12761 ) | ( ~n10575 & n12761 ) ;
  assign n49718 = ~n32037 & n49717 ;
  assign n49719 = n20550 & n49718 ;
  assign n49720 = n34995 ^ n12480 ^ 1'b0 ;
  assign n49721 = ~n10036 & n26394 ;
  assign n49722 = n49721 ^ n10577 ^ n9195 ;
  assign n49724 = ~n12728 & n25590 ;
  assign n49725 = ~n32618 & n49724 ;
  assign n49726 = n49725 ^ n29618 ^ n25805 ;
  assign n49723 = n21011 ^ n17910 ^ n13497 ;
  assign n49727 = n49726 ^ n49723 ^ n10552 ;
  assign n49728 = ~n9164 & n47255 ;
  assign n49729 = n15111 & n21687 ;
  assign n49730 = ~n9886 & n49729 ;
  assign n49731 = n36978 ^ n30096 ^ n6164 ;
  assign n49732 = n49638 ^ n44985 ^ 1'b0 ;
  assign n49733 = n1655 | n49732 ;
  assign n49734 = ( n40184 & n49731 ) | ( n40184 & ~n49733 ) | ( n49731 & ~n49733 ) ;
  assign n49735 = n45139 ^ n31896 ^ 1'b0 ;
  assign n49736 = n49734 & ~n49735 ;
  assign n49737 = n11334 | n13468 ;
  assign n49738 = n11631 ^ n7143 ^ x83 ;
  assign n49739 = ( n883 & n11174 ) | ( n883 & n46540 ) | ( n11174 & n46540 ) ;
  assign n49740 = n49739 ^ n31520 ^ n27616 ;
  assign n49741 = n49740 ^ n10955 ^ n7406 ;
  assign n49742 = ( n34265 & n39452 ) | ( n34265 & ~n46940 ) | ( n39452 & ~n46940 ) ;
  assign n49743 = n6539 | n10730 ;
  assign n49744 = n49743 ^ n6437 ^ 1'b0 ;
  assign n49745 = n11414 & ~n12493 ;
  assign n49746 = ( ~n838 & n49744 ) | ( ~n838 & n49745 ) | ( n49744 & n49745 ) ;
  assign n49747 = n32219 ^ n22855 ^ n11111 ;
  assign n49748 = n5554 | n9131 ;
  assign n49749 = n25809 & ~n49748 ;
  assign n49750 = ~n49747 & n49749 ;
  assign n49751 = n1646 & n40029 ;
  assign n49752 = n49751 ^ n8705 ^ 1'b0 ;
  assign n49753 = n15323 | n49752 ;
  assign n49754 = n17470 | n18343 ;
  assign n49760 = n43034 ^ n1709 ^ 1'b0 ;
  assign n49761 = n17922 & ~n49760 ;
  assign n49756 = n1616 & n2718 ;
  assign n49755 = n830 & ~n4190 ;
  assign n49757 = n49756 ^ n49755 ^ 1'b0 ;
  assign n49758 = n18208 ^ n10300 ^ 1'b0 ;
  assign n49759 = n49757 & ~n49758 ;
  assign n49762 = n49761 ^ n49759 ^ 1'b0 ;
  assign n49763 = ~n43721 & n49762 ;
  assign n49764 = ( n33148 & n47413 ) | ( n33148 & ~n47713 ) | ( n47413 & ~n47713 ) ;
  assign n49766 = n39954 ^ n9465 ^ 1'b0 ;
  assign n49765 = ~n1303 & n21629 ;
  assign n49767 = n49766 ^ n49765 ^ 1'b0 ;
  assign n49768 = n49767 ^ n39953 ^ 1'b0 ;
  assign n49769 = n42997 ^ n2325 ^ n662 ;
  assign n49770 = ( x156 & n28589 ) | ( x156 & n45525 ) | ( n28589 & n45525 ) ;
  assign n49771 = n11664 & ~n26654 ;
  assign n49772 = ~n41115 & n49771 ;
  assign n49773 = n2213 & n4137 ;
  assign n49774 = n8823 & ~n35425 ;
  assign n49775 = n49773 & n49774 ;
  assign n49776 = n3094 & ~n28492 ;
  assign n49777 = n49776 ^ n6740 ^ 1'b0 ;
  assign n49778 = n43858 ^ n34841 ^ n6958 ;
  assign n49779 = n49778 ^ n23628 ^ n15608 ;
  assign n49780 = n23258 ^ n1380 ^ 1'b0 ;
  assign n49781 = n38960 ^ n29643 ^ n21999 ;
  assign n49785 = n31785 ^ n9501 ^ 1'b0 ;
  assign n49786 = n18978 | n49785 ;
  assign n49787 = n22169 | n49786 ;
  assign n49788 = n18596 & ~n49787 ;
  assign n49782 = n8399 ^ n1372 ^ 1'b0 ;
  assign n49783 = n4851 & n49782 ;
  assign n49784 = ( ~n4090 & n19461 ) | ( ~n4090 & n49783 ) | ( n19461 & n49783 ) ;
  assign n49789 = n49788 ^ n49784 ^ n34642 ;
  assign n49790 = n49304 ^ n14618 ^ 1'b0 ;
  assign n49791 = n36487 | n49790 ;
  assign n49792 = n19069 ^ n10308 ^ 1'b0 ;
  assign n49793 = n3087 & n49792 ;
  assign n49794 = n1827 ^ n482 ^ 1'b0 ;
  assign n49795 = ( n16072 & n21784 ) | ( n16072 & ~n22353 ) | ( n21784 & ~n22353 ) ;
  assign n49796 = x212 & ~n4528 ;
  assign n49797 = n49796 ^ n5989 ^ 1'b0 ;
  assign n49798 = ( n15506 & ~n43078 ) | ( n15506 & n49797 ) | ( ~n43078 & n49797 ) ;
  assign n49799 = ~n14552 & n49798 ;
  assign n49800 = ~n24931 & n49799 ;
  assign n49801 = n49800 ^ n24759 ^ 1'b0 ;
  assign n49802 = n34764 & ~n49801 ;
  assign n49803 = n16804 ^ n7642 ^ n1261 ;
  assign n49804 = n49802 & n49803 ;
  assign n49805 = n49804 ^ n43948 ^ 1'b0 ;
  assign n49806 = n47386 ^ n26283 ^ n974 ;
  assign n49807 = ( x72 & ~n8306 ) | ( x72 & n10990 ) | ( ~n8306 & n10990 ) ;
  assign n49808 = n32791 ^ n13605 ^ n3852 ;
  assign n49809 = ( n8939 & n46820 ) | ( n8939 & ~n49808 ) | ( n46820 & ~n49808 ) ;
  assign n49810 = n3688 | n49809 ;
  assign n49811 = n15564 | n49810 ;
  assign n49812 = n49811 ^ n45829 ^ n8745 ;
  assign n49813 = n36267 ^ n24697 ^ 1'b0 ;
  assign n49814 = n1134 & n49813 ;
  assign n49815 = n17291 & ~n36969 ;
  assign n49816 = n49815 ^ n19824 ^ 1'b0 ;
  assign n49817 = n20503 & n25662 ;
  assign n49818 = ( n9795 & ~n12692 ) | ( n9795 & n35298 ) | ( ~n12692 & n35298 ) ;
  assign n49819 = n49818 ^ n18596 ^ 1'b0 ;
  assign n49820 = ( ~n10543 & n44050 ) | ( ~n10543 & n48547 ) | ( n44050 & n48547 ) ;
  assign n49821 = n22045 ^ n14428 ^ 1'b0 ;
  assign n49822 = n17981 & ~n49821 ;
  assign n49823 = n49822 ^ n14931 ^ 1'b0 ;
  assign n49824 = n30309 ^ n19763 ^ n10030 ;
  assign n49825 = n9539 | n29171 ;
  assign n49829 = n15119 | n32724 ;
  assign n49826 = n17425 | n23027 ;
  assign n49827 = n38221 & ~n49826 ;
  assign n49828 = n6973 & ~n49827 ;
  assign n49830 = n49829 ^ n49828 ^ 1'b0 ;
  assign n49831 = ~n24217 & n49274 ;
  assign n49832 = n17218 & n49831 ;
  assign n49833 = x9 & n43743 ;
  assign n49834 = n49833 ^ n28388 ^ 1'b0 ;
  assign n49835 = ~n4369 & n23659 ;
  assign n49836 = n36870 & n49835 ;
  assign n49837 = n49836 ^ n37732 ^ 1'b0 ;
  assign n49838 = n29036 ^ n8772 ^ n4793 ;
  assign n49839 = n15448 ^ n6826 ^ 1'b0 ;
  assign n49840 = n10480 | n49839 ;
  assign n49843 = n8279 & n18652 ;
  assign n49841 = ( ~n4684 & n8448 ) | ( ~n4684 & n14891 ) | ( n8448 & n14891 ) ;
  assign n49842 = n49841 ^ n39603 ^ n9697 ;
  assign n49844 = n49843 ^ n49842 ^ n13601 ;
  assign n49845 = n38424 ^ n21160 ^ 1'b0 ;
  assign n49846 = n2443 & ~n49845 ;
  assign n49847 = ( ~n12925 & n24006 ) | ( ~n12925 & n49846 ) | ( n24006 & n49846 ) ;
  assign n49848 = n1559 & ~n24128 ;
  assign n49849 = n49847 & n49848 ;
  assign n49850 = ~n1064 & n7934 ;
  assign n49851 = ( ~x238 & n21389 ) | ( ~x238 & n34861 ) | ( n21389 & n34861 ) ;
  assign n49852 = ( ~n13684 & n28904 ) | ( ~n13684 & n29994 ) | ( n28904 & n29994 ) ;
  assign n49853 = n3504 & ~n49852 ;
  assign n49854 = ~n15975 & n49853 ;
  assign n49855 = ( n27468 & n40776 ) | ( n27468 & n49854 ) | ( n40776 & n49854 ) ;
  assign n49856 = ( ~n8346 & n19030 ) | ( ~n8346 & n49855 ) | ( n19030 & n49855 ) ;
  assign n49857 = n39103 ^ n33561 ^ 1'b0 ;
  assign n49858 = n32893 ^ n18438 ^ 1'b0 ;
  assign n49859 = n20847 & ~n49858 ;
  assign n49860 = n49859 ^ n19073 ^ n774 ;
  assign n49861 = n7123 & ~n17544 ;
  assign n49862 = n49861 ^ n18568 ^ 1'b0 ;
  assign n49868 = n29660 ^ n26412 ^ n4562 ;
  assign n49864 = n7039 & ~n24968 ;
  assign n49865 = n16686 ^ n8084 ^ 1'b0 ;
  assign n49866 = ~n49864 & n49865 ;
  assign n49867 = n8497 & n49866 ;
  assign n49869 = n49868 ^ n49867 ^ 1'b0 ;
  assign n49863 = ~n11607 & n17408 ;
  assign n49870 = n49869 ^ n49863 ^ 1'b0 ;
  assign n49871 = n15614 & ~n43799 ;
  assign n49872 = n49871 ^ n49843 ^ 1'b0 ;
  assign n49873 = n4445 & ~n12242 ;
  assign n49874 = n15154 & ~n36535 ;
  assign n49875 = ~n32681 & n44705 ;
  assign n49876 = n49875 ^ n21198 ^ 1'b0 ;
  assign n49877 = n5855 | n32734 ;
  assign n49878 = n49876 & ~n49877 ;
  assign n49879 = ( n1336 & n2291 ) | ( n1336 & n49878 ) | ( n2291 & n49878 ) ;
  assign n49880 = n27799 ^ n21727 ^ n16650 ;
  assign n49881 = ( n23703 & n27627 ) | ( n23703 & ~n48172 ) | ( n27627 & ~n48172 ) ;
  assign n49882 = n3093 ^ n464 ^ 1'b0 ;
  assign n49883 = n24519 | n49882 ;
  assign n49884 = ( ~n8380 & n10667 ) | ( ~n8380 & n49883 ) | ( n10667 & n49883 ) ;
  assign n49885 = n38848 ^ n11897 ^ 1'b0 ;
  assign n49886 = n38811 ^ n21254 ^ 1'b0 ;
  assign n49887 = n49885 & ~n49886 ;
  assign n49888 = n2798 & ~n37370 ;
  assign n49889 = n6332 & n14237 ;
  assign n49890 = n49889 ^ n7897 ^ 1'b0 ;
  assign n49891 = n34113 | n49890 ;
  assign n49892 = n49891 ^ n32688 ^ 1'b0 ;
  assign n49893 = n2642 & ~n24594 ;
  assign n49894 = n49893 ^ n18061 ^ n9769 ;
  assign n49895 = ( n16677 & ~n18341 ) | ( n16677 & n45785 ) | ( ~n18341 & n45785 ) ;
  assign n49896 = ~n20493 & n35729 ;
  assign n49897 = n4807 | n38778 ;
  assign n49898 = ( n4441 & n49896 ) | ( n4441 & ~n49897 ) | ( n49896 & ~n49897 ) ;
  assign n49899 = ( n6107 & n8910 ) | ( n6107 & ~n25894 ) | ( n8910 & ~n25894 ) ;
  assign n49900 = ~n33411 & n42508 ;
  assign n49901 = n7886 | n26166 ;
  assign n49902 = n49901 ^ n9161 ^ 1'b0 ;
  assign n49903 = ( ~n3446 & n3792 ) | ( ~n3446 & n4832 ) | ( n3792 & n4832 ) ;
  assign n49904 = n49227 | n49903 ;
  assign n49905 = n14047 | n20253 ;
  assign n49906 = n4989 ^ n334 ^ 1'b0 ;
  assign n49907 = n1819 & n49906 ;
  assign n49908 = n24246 | n49907 ;
  assign n49909 = ( n8515 & n27488 ) | ( n8515 & ~n49908 ) | ( n27488 & ~n49908 ) ;
  assign n49910 = n10998 & n39583 ;
  assign n49911 = ( n782 & ~n11496 ) | ( n782 & n25675 ) | ( ~n11496 & n25675 ) ;
  assign n49912 = ( ~n4959 & n28284 ) | ( ~n4959 & n49911 ) | ( n28284 & n49911 ) ;
  assign n49913 = n26792 ^ n17273 ^ n16764 ;
  assign n49914 = x34 | n36029 ;
  assign n49915 = n20759 & n49914 ;
  assign n49916 = ~n49913 & n49915 ;
  assign n49917 = n1977 | n6397 ;
  assign n49918 = n49917 ^ n45577 ^ 1'b0 ;
  assign n49919 = n8598 | n10995 ;
  assign n49920 = n49919 ^ n3149 ^ 1'b0 ;
  assign n49929 = n5864 & n24198 ;
  assign n49925 = n17604 & ~n24288 ;
  assign n49926 = n9951 & n49925 ;
  assign n49923 = ~n31295 & n34301 ;
  assign n49924 = n49923 ^ n13213 ^ n2026 ;
  assign n49927 = n49926 ^ n49924 ^ n4893 ;
  assign n49928 = ( n22190 & n31504 ) | ( n22190 & ~n49927 ) | ( n31504 & ~n49927 ) ;
  assign n49930 = n49929 ^ n49928 ^ n17362 ;
  assign n49921 = n17737 & n32791 ;
  assign n49922 = n49921 ^ n7566 ^ 1'b0 ;
  assign n49931 = n49930 ^ n49922 ^ 1'b0 ;
  assign n49932 = n16580 & n49931 ;
  assign n49933 = n2682 & n5173 ;
  assign n49934 = ~n15625 & n49933 ;
  assign n49935 = n21529 | n49934 ;
  assign n49936 = n44789 ^ n11775 ^ 1'b0 ;
  assign n49937 = ~n20759 & n33461 ;
  assign n49938 = n49937 ^ n49149 ^ n18443 ;
  assign n49939 = n1145 & n38979 ;
  assign n49940 = n39437 ^ n37720 ^ n13420 ;
  assign n49941 = n45373 ^ n34049 ^ 1'b0 ;
  assign n49942 = n13920 ^ n12421 ^ 1'b0 ;
  assign n49943 = n3297 | n49942 ;
  assign n49944 = n9882 & ~n49943 ;
  assign n49945 = n39449 ^ n13151 ^ 1'b0 ;
  assign n49946 = n17611 & n49945 ;
  assign n49947 = ( ~n20889 & n23590 ) | ( ~n20889 & n43679 ) | ( n23590 & n43679 ) ;
  assign n49948 = n49947 ^ n37344 ^ n13757 ;
  assign n49949 = n13365 & ~n48357 ;
  assign n49950 = n49949 ^ n38020 ^ 1'b0 ;
  assign n49951 = n49950 ^ n30643 ^ n19868 ;
  assign n49952 = n49951 ^ n22820 ^ n6441 ;
  assign n49955 = n27186 ^ n22269 ^ n11727 ;
  assign n49953 = ~n8282 & n38580 ;
  assign n49954 = n49953 ^ n29563 ^ 1'b0 ;
  assign n49956 = n49955 ^ n49954 ^ n13976 ;
  assign n49957 = n38038 ^ n31270 ^ n9825 ;
  assign n49958 = n2325 ^ x56 ^ 1'b0 ;
  assign n49959 = n14008 | n49958 ;
  assign n49960 = ( n7924 & n16730 ) | ( n7924 & ~n36680 ) | ( n16730 & ~n36680 ) ;
  assign n49961 = ~n34279 & n49960 ;
  assign n49962 = n23837 & n49961 ;
  assign n49963 = ( n7744 & n24490 ) | ( n7744 & n29432 ) | ( n24490 & n29432 ) ;
  assign n49964 = ( n14373 & n22725 ) | ( n14373 & n33506 ) | ( n22725 & n33506 ) ;
  assign n49965 = n15341 & ~n39248 ;
  assign n49966 = ( n23372 & n49964 ) | ( n23372 & n49965 ) | ( n49964 & n49965 ) ;
  assign n49967 = ( n6773 & n10456 ) | ( n6773 & ~n36164 ) | ( n10456 & ~n36164 ) ;
  assign n49968 = n21014 ^ n3107 ^ 1'b0 ;
  assign n49969 = ~n48246 & n49968 ;
  assign n49970 = n40384 ^ n14765 ^ 1'b0 ;
  assign n49971 = n23611 | n49970 ;
  assign n49972 = n19583 | n30319 ;
  assign n49973 = n14906 | n49972 ;
  assign n49974 = n49973 ^ n34734 ^ n33689 ;
  assign n49975 = n9936 ^ n7375 ^ 1'b0 ;
  assign n49976 = ( x248 & n35049 ) | ( x248 & n35883 ) | ( n35049 & n35883 ) ;
  assign n49977 = n24922 ^ n4952 ^ 1'b0 ;
  assign n49978 = n13386 & n49977 ;
  assign n49979 = ~n1449 & n49978 ;
  assign n49980 = n23192 ^ n18793 ^ 1'b0 ;
  assign n49981 = n41322 | n49980 ;
  assign n49982 = ~n31838 & n34382 ;
  assign n49983 = n49982 ^ n25178 ^ 1'b0 ;
  assign n49984 = ~n14569 & n38708 ;
  assign n49985 = ~n49983 & n49984 ;
  assign n49986 = n22765 & n25020 ;
  assign n49988 = n12959 ^ n9825 ^ 1'b0 ;
  assign n49989 = n14022 & n49988 ;
  assign n49987 = ~n8999 & n17294 ;
  assign n49990 = n49989 ^ n49987 ^ n25237 ;
  assign n49991 = ( n11188 & n15583 ) | ( n11188 & n49990 ) | ( n15583 & n49990 ) ;
  assign n49992 = n12179 & ~n46109 ;
  assign n49993 = ~n12761 & n31869 ;
  assign n49994 = n23010 & n49993 ;
  assign n49995 = n49994 ^ n44151 ^ n28728 ;
  assign n49996 = n9704 & ~n38136 ;
  assign n49997 = n17165 & n19663 ;
  assign n49998 = n49997 ^ n4803 ^ 1'b0 ;
  assign n49999 = ( n6796 & ~n15710 ) | ( n6796 & n46558 ) | ( ~n15710 & n46558 ) ;
  assign n50000 = n38652 | n44080 ;
  assign n50001 = n49999 & ~n50000 ;
  assign n50002 = n28286 ^ n5709 ^ 1'b0 ;
  assign n50013 = n22607 ^ n8689 ^ 1'b0 ;
  assign n50014 = n50013 ^ n24361 ^ n6035 ;
  assign n50009 = n26173 ^ n21816 ^ 1'b0 ;
  assign n50010 = ~n47234 & n50009 ;
  assign n50011 = n50010 ^ n16438 ^ 1'b0 ;
  assign n50012 = ~n1832 & n50011 ;
  assign n50015 = n50014 ^ n50012 ^ n21852 ;
  assign n50004 = n29732 & n37898 ;
  assign n50005 = n1124 & n50004 ;
  assign n50003 = n9618 | n33128 ;
  assign n50006 = n50005 ^ n50003 ^ 1'b0 ;
  assign n50007 = n50006 ^ n22035 ^ 1'b0 ;
  assign n50008 = n41450 | n50007 ;
  assign n50016 = n50015 ^ n50008 ^ n45800 ;
  assign n50017 = n46572 ^ n12194 ^ n4542 ;
  assign n50018 = n12988 | n46948 ;
  assign n50019 = n50018 ^ n17592 ^ 1'b0 ;
  assign n50020 = n50019 ^ n7554 ^ 1'b0 ;
  assign n50021 = n19229 | n50020 ;
  assign n50022 = n50021 ^ n32642 ^ n6960 ;
  assign n50023 = n5559 & ~n34121 ;
  assign n50024 = n2205 | n50023 ;
  assign n50025 = n18924 & ~n50024 ;
  assign n50026 = ( ~n37647 & n47752 ) | ( ~n37647 & n50025 ) | ( n47752 & n50025 ) ;
  assign n50027 = n4168 & n10127 ;
  assign n50028 = ~n41023 & n50027 ;
  assign n50029 = n50028 ^ n8741 ^ 1'b0 ;
  assign n50030 = n21565 & n50029 ;
  assign n50031 = ( n3788 & ~n17725 ) | ( n3788 & n50030 ) | ( ~n17725 & n50030 ) ;
  assign n50032 = n5413 | n21619 ;
  assign n50033 = n24179 | n50032 ;
  assign n50034 = n13689 ^ n4068 ^ 1'b0 ;
  assign n50035 = n19778 & n50034 ;
  assign n50036 = n48152 ^ n1493 ^ n791 ;
  assign n50037 = n32326 & ~n50036 ;
  assign n50038 = ~n26357 & n27603 ;
  assign n50039 = n50038 ^ n48041 ^ 1'b0 ;
  assign n50040 = n9114 | n34291 ;
  assign n50041 = n50040 ^ n23264 ^ 1'b0 ;
  assign n50042 = ( n11976 & ~n23982 ) | ( n11976 & n47649 ) | ( ~n23982 & n47649 ) ;
  assign n50043 = n50042 ^ n28106 ^ n21265 ;
  assign n50044 = ~n31129 & n47437 ;
  assign n50045 = n50044 ^ n49111 ^ 1'b0 ;
  assign n50046 = n36520 ^ n15406 ^ n10686 ;
  assign n50047 = n47453 ^ n19855 ^ n16294 ;
  assign n50048 = n29769 ^ n3579 ^ 1'b0 ;
  assign n50049 = ~n32985 & n50048 ;
  assign n50050 = ~n28252 & n38089 ;
  assign n50051 = n50050 ^ n9043 ^ 1'b0 ;
  assign n50052 = n39612 | n43209 ;
  assign n50053 = n40520 ^ n36178 ^ n30348 ;
  assign n50054 = ( n15764 & n33634 ) | ( n15764 & n35869 ) | ( n33634 & n35869 ) ;
  assign n50055 = n13512 & ~n15820 ;
  assign n50056 = ~n3085 & n50055 ;
  assign n50057 = ( n19743 & n50054 ) | ( n19743 & ~n50056 ) | ( n50054 & ~n50056 ) ;
  assign n50058 = ( ~n13795 & n26919 ) | ( ~n13795 & n50057 ) | ( n26919 & n50057 ) ;
  assign n50059 = n23581 ^ n10351 ^ n4893 ;
  assign n50060 = n50059 ^ n10917 ^ n10599 ;
  assign n50061 = n14318 ^ n7230 ^ n5860 ;
  assign n50062 = n46743 ^ n14439 ^ 1'b0 ;
  assign n50063 = ~n21479 & n50062 ;
  assign n50064 = n50061 & ~n50063 ;
  assign n50065 = n26699 ^ n9632 ^ 1'b0 ;
  assign n50066 = n37290 ^ n20448 ^ n12933 ;
  assign n50067 = n14091 & ~n15202 ;
  assign n50068 = ~n24254 & n50067 ;
  assign n50069 = n50066 & n50068 ;
  assign n50070 = n21030 & n22196 ;
  assign n50071 = n38356 ^ n17743 ^ n2113 ;
  assign n50072 = n38635 ^ n3930 ^ 1'b0 ;
  assign n50073 = n50072 ^ n12579 ^ n8591 ;
  assign n50074 = n50073 ^ n10963 ^ 1'b0 ;
  assign n50075 = ~n50071 & n50074 ;
  assign n50076 = n16786 ^ n8249 ^ n4147 ;
  assign n50077 = n841 | n2865 ;
  assign n50078 = ( ~n33372 & n50076 ) | ( ~n33372 & n50077 ) | ( n50076 & n50077 ) ;
  assign n50079 = n40420 ^ n11227 ^ n9141 ;
  assign n50080 = n10621 | n14276 ;
  assign n50081 = n25707 ^ n15989 ^ n757 ;
  assign n50082 = n50081 ^ n23391 ^ 1'b0 ;
  assign n50083 = n15320 & n50082 ;
  assign n50084 = n10126 & ~n37750 ;
  assign n50085 = n50084 ^ n27335 ^ 1'b0 ;
  assign n50086 = n15842 & ~n29498 ;
  assign n50087 = ~n30126 & n49978 ;
  assign n50088 = n21609 ^ n7410 ^ 1'b0 ;
  assign n50089 = ~n19775 & n50088 ;
  assign n50090 = ( n39098 & ~n49331 ) | ( n39098 & n50089 ) | ( ~n49331 & n50089 ) ;
  assign n50091 = n3565 & n19911 ;
  assign n50092 = n31888 ^ n16148 ^ 1'b0 ;
  assign n50093 = n50092 ^ n48461 ^ n47050 ;
  assign n50094 = ( n10002 & ~n14866 ) | ( n10002 & n21059 ) | ( ~n14866 & n21059 ) ;
  assign n50095 = n18768 ^ n1317 ^ 1'b0 ;
  assign n50096 = n32879 | n50095 ;
  assign n50097 = ~n15247 & n27445 ;
  assign n50098 = n44355 ^ n21288 ^ 1'b0 ;
  assign n50099 = n50098 ^ n11891 ^ n5380 ;
  assign n50100 = n50099 ^ n25541 ^ n16598 ;
  assign n50101 = n5153 & n10511 ;
  assign n50102 = n50101 ^ n30149 ^ 1'b0 ;
  assign n50103 = n27302 | n45219 ;
  assign n50104 = n50103 ^ n6589 ^ 1'b0 ;
  assign n50105 = ( n37802 & n50102 ) | ( n37802 & ~n50104 ) | ( n50102 & ~n50104 ) ;
  assign n50106 = n15142 ^ n14924 ^ 1'b0 ;
  assign n50107 = n48504 ^ n21476 ^ n5568 ;
  assign n50108 = n30058 ^ n10427 ^ 1'b0 ;
  assign n50109 = n50108 ^ n39197 ^ n26114 ;
  assign n50110 = n47768 ^ n8422 ^ 1'b0 ;
  assign n50111 = n45429 & n50110 ;
  assign n50112 = n5499 & ~n32593 ;
  assign n50113 = n27004 ^ n23194 ^ 1'b0 ;
  assign n50114 = ~n37090 & n50113 ;
  assign n50115 = n5372 & n28401 ;
  assign n50116 = n42867 & n50115 ;
  assign n50121 = n14446 & n22566 ;
  assign n50122 = ~n22566 & n50121 ;
  assign n50117 = n1928 & n2333 ;
  assign n50118 = ~n1928 & n50117 ;
  assign n50119 = n50118 ^ n2812 ^ n604 ;
  assign n50120 = n50119 ^ n9180 ^ n466 ;
  assign n50123 = n50122 ^ n50120 ^ n15373 ;
  assign n50124 = n32130 ^ n30624 ^ n1450 ;
  assign n50127 = n34462 ^ n3763 ^ 1'b0 ;
  assign n50128 = n17810 & n50127 ;
  assign n50125 = n18579 ^ n14601 ^ 1'b0 ;
  assign n50126 = n32150 & n50125 ;
  assign n50129 = n50128 ^ n50126 ^ n27539 ;
  assign n50130 = n44591 ^ n22923 ^ n6218 ;
  assign n50131 = n45828 ^ n29621 ^ n9959 ;
  assign n50132 = n46117 ^ n25431 ^ 1'b0 ;
  assign n50133 = ~n10572 & n50132 ;
  assign n50134 = ( n22018 & n23344 ) | ( n22018 & ~n50133 ) | ( n23344 & ~n50133 ) ;
  assign n50135 = ~n33977 & n48515 ;
  assign n50136 = n37932 & n50135 ;
  assign n50137 = n14813 & n36662 ;
  assign n50138 = n50137 ^ n22173 ^ 1'b0 ;
  assign n50139 = n45543 ^ n16064 ^ 1'b0 ;
  assign n50140 = n1482 & n50139 ;
  assign n50141 = n18005 ^ n11787 ^ n9762 ;
  assign n50142 = n13590 & ~n50141 ;
  assign n50143 = n23497 ^ n13115 ^ 1'b0 ;
  assign n50144 = n4052 & ~n50143 ;
  assign n50145 = ( n14586 & n34595 ) | ( n14586 & n48666 ) | ( n34595 & n48666 ) ;
  assign n50146 = n11357 ^ n10406 ^ n434 ;
  assign n50147 = n48174 & n50146 ;
  assign n50148 = n50147 ^ n32693 ^ n19218 ;
  assign n50149 = ~n13137 & n46765 ;
  assign n50150 = ~n9551 & n50149 ;
  assign n50151 = n50150 ^ n28403 ^ 1'b0 ;
  assign n50152 = n27059 ^ n11132 ^ 1'b0 ;
  assign n50153 = n50152 ^ n5481 ^ x112 ;
  assign n50155 = ( ~n2315 & n12904 ) | ( ~n2315 & n18695 ) | ( n12904 & n18695 ) ;
  assign n50154 = ( n492 & ~n39740 ) | ( n492 & n49227 ) | ( ~n39740 & n49227 ) ;
  assign n50156 = n50155 ^ n50154 ^ n3668 ;
  assign n50157 = n18682 & ~n50156 ;
  assign n50158 = ( n12051 & n24117 ) | ( n12051 & n50157 ) | ( n24117 & n50157 ) ;
  assign n50159 = n29326 ^ n23101 ^ n10930 ;
  assign n50160 = ~n5012 & n50159 ;
  assign n50161 = ( n6798 & n8924 ) | ( n6798 & n21264 ) | ( n8924 & n21264 ) ;
  assign n50162 = n50161 ^ n5291 ^ 1'b0 ;
  assign n50163 = n45783 & ~n50162 ;
  assign n50164 = n20659 & n24242 ;
  assign n50165 = n50164 ^ n14803 ^ 1'b0 ;
  assign n50166 = n24996 ^ n8070 ^ 1'b0 ;
  assign n50167 = n50165 & n50166 ;
  assign n50168 = ~n23012 & n29008 ;
  assign n50169 = ( n12724 & n14902 ) | ( n12724 & ~n20196 ) | ( n14902 & ~n20196 ) ;
  assign n50170 = n50169 ^ n29105 ^ 1'b0 ;
  assign n50171 = ( n11089 & ~n17359 ) | ( n11089 & n50170 ) | ( ~n17359 & n50170 ) ;
  assign n50172 = n2700 & ~n13597 ;
  assign n50173 = n5981 & n50172 ;
  assign n50174 = n50173 ^ n19007 ^ n2220 ;
  assign n50175 = n50174 ^ n48779 ^ n14450 ;
  assign n50180 = ~n13116 & n27264 ;
  assign n50176 = n44756 ^ n30764 ^ 1'b0 ;
  assign n50177 = n3591 | n50176 ;
  assign n50178 = n50177 ^ n11897 ^ 1'b0 ;
  assign n50179 = n38065 | n50178 ;
  assign n50181 = n50180 ^ n50179 ^ 1'b0 ;
  assign n50182 = n43033 ^ n21094 ^ 1'b0 ;
  assign n50183 = n29077 & ~n50182 ;
  assign n50184 = n32693 & n35575 ;
  assign n50186 = n6282 | n13272 ;
  assign n50185 = n31018 | n35357 ;
  assign n50187 = n50186 ^ n50185 ^ 1'b0 ;
  assign n50188 = n1276 | n36020 ;
  assign n50189 = n50188 ^ n35582 ^ 1'b0 ;
  assign n50190 = n1655 | n6476 ;
  assign n50191 = n50190 ^ n1801 ^ 1'b0 ;
  assign n50192 = n50191 ^ n32948 ^ 1'b0 ;
  assign n50193 = n50192 ^ n35713 ^ n25557 ;
  assign n50194 = n4793 ^ n2013 ^ 1'b0 ;
  assign n50195 = n10184 | n50194 ;
  assign n50196 = ( n9365 & n35972 ) | ( n9365 & ~n50195 ) | ( n35972 & ~n50195 ) ;
  assign n50197 = ( ~n8908 & n13683 ) | ( ~n8908 & n28003 ) | ( n13683 & n28003 ) ;
  assign n50198 = n48241 ^ n18057 ^ n12771 ;
  assign n50199 = n25138 ^ n25043 ^ n389 ;
  assign n50200 = ~n1475 & n50199 ;
  assign n50201 = n26438 & n35476 ;
  assign n50202 = n39022 ^ n30438 ^ 1'b0 ;
  assign n50203 = n8769 | n50202 ;
  assign n50204 = n7527 & ~n11999 ;
  assign n50205 = n50203 & n50204 ;
  assign n50206 = n44700 ^ n14206 ^ n2916 ;
  assign n50207 = n13621 | n50206 ;
  assign n50208 = n50205 & ~n50207 ;
  assign n50209 = n50208 ^ n5523 ^ 1'b0 ;
  assign n50210 = n50209 ^ n27350 ^ 1'b0 ;
  assign n50211 = ~n12935 & n30248 ;
  assign n50212 = n50211 ^ n19565 ^ 1'b0 ;
  assign n50213 = ~n23210 & n48606 ;
  assign n50214 = n8595 & n33717 ;
  assign n50215 = ~n38597 & n50214 ;
  assign n50216 = ~n13967 & n37673 ;
  assign n50217 = n7505 & ~n24446 ;
  assign n50218 = ( ~n11614 & n21907 ) | ( ~n11614 & n50217 ) | ( n21907 & n50217 ) ;
  assign n50219 = ( n20222 & ~n46732 ) | ( n20222 & n50218 ) | ( ~n46732 & n50218 ) ;
  assign n50220 = n4046 | n33962 ;
  assign n50221 = ( n40308 & n50219 ) | ( n40308 & n50220 ) | ( n50219 & n50220 ) ;
  assign n50222 = n19740 ^ n9109 ^ 1'b0 ;
  assign n50223 = ~n2383 & n44486 ;
  assign n50224 = n4095 & n50223 ;
  assign n50225 = n2260 & ~n40185 ;
  assign n50226 = ~n50224 & n50225 ;
  assign n50227 = ~n3376 & n4678 ;
  assign n50228 = n36078 ^ n2917 ^ 1'b0 ;
  assign n50229 = ~n27872 & n50228 ;
  assign n50230 = n392 & ~n6333 ;
  assign n50231 = n10356 & ~n15945 ;
  assign n50232 = n6387 | n15334 ;
  assign n50233 = n50232 ^ n35039 ^ 1'b0 ;
  assign n50234 = n11080 & ~n50233 ;
  assign n50235 = n4762 | n46087 ;
  assign n50236 = n1246 & ~n50235 ;
  assign n50237 = n10344 & ~n50236 ;
  assign n50238 = n44549 ^ n11131 ^ n5292 ;
  assign n50239 = n279 | n29634 ;
  assign n50240 = n15017 ^ n10738 ^ 1'b0 ;
  assign n50241 = ~n2314 & n9016 ;
  assign n50242 = n50240 & n50241 ;
  assign n50243 = n50242 ^ n15463 ^ n9473 ;
  assign n50244 = n50243 ^ n46680 ^ n27116 ;
  assign n50245 = n30183 | n38018 ;
  assign n50246 = n50245 ^ n15321 ^ 1'b0 ;
  assign n50247 = ( ~n50239 & n50244 ) | ( ~n50239 & n50246 ) | ( n50244 & n50246 ) ;
  assign n50248 = n35096 ^ n738 ^ 1'b0 ;
  assign n50249 = n1105 & n50248 ;
  assign n50250 = ( n17441 & ~n33717 ) | ( n17441 & n50249 ) | ( ~n33717 & n50249 ) ;
  assign n50251 = ( n2151 & ~n39622 ) | ( n2151 & n50250 ) | ( ~n39622 & n50250 ) ;
  assign n50252 = ( n15432 & n26128 ) | ( n15432 & ~n28005 ) | ( n26128 & ~n28005 ) ;
  assign n50253 = ( n3805 & ~n8542 ) | ( n3805 & n50252 ) | ( ~n8542 & n50252 ) ;
  assign n50254 = n26305 ^ n5115 ^ 1'b0 ;
  assign n50255 = n12137 & ~n50254 ;
  assign n50256 = n2925 & ~n45602 ;
  assign n50257 = n24937 & n50256 ;
  assign n50258 = n6083 ^ n520 ^ 1'b0 ;
  assign n50259 = n21220 & n28138 ;
  assign n50260 = ~n16507 & n50259 ;
  assign n50261 = ~n50258 & n50260 ;
  assign n50262 = n6803 | n38645 ;
  assign n50263 = n10844 & ~n50262 ;
  assign n50264 = n23129 ^ n20244 ^ 1'b0 ;
  assign n50267 = ( n2341 & n5733 ) | ( n2341 & ~n6556 ) | ( n5733 & ~n6556 ) ;
  assign n50266 = n16096 & ~n18327 ;
  assign n50268 = n50267 ^ n50266 ^ 1'b0 ;
  assign n50265 = ( n3366 & n37817 ) | ( n3366 & n38263 ) | ( n37817 & n38263 ) ;
  assign n50269 = n50268 ^ n50265 ^ n39688 ;
  assign n50273 = n9969 | n15530 ;
  assign n50274 = n38905 ^ n2494 ^ 1'b0 ;
  assign n50275 = n50273 & n50274 ;
  assign n50276 = ~n2345 & n16600 ;
  assign n50277 = ~n50275 & n50276 ;
  assign n50270 = n39750 ^ n13590 ^ 1'b0 ;
  assign n50271 = n11221 & n50270 ;
  assign n50272 = ~n3141 & n50271 ;
  assign n50278 = n50277 ^ n50272 ^ 1'b0 ;
  assign n50284 = ~n9999 & n15777 ;
  assign n50285 = n19689 & n50284 ;
  assign n50281 = n35643 ^ n15296 ^ n10489 ;
  assign n50282 = n50281 ^ n43460 ^ n9855 ;
  assign n50280 = ~n15153 & n38508 ;
  assign n50279 = ( ~n11389 & n38274 ) | ( ~n11389 & n41936 ) | ( n38274 & n41936 ) ;
  assign n50283 = n50282 ^ n50280 ^ n50279 ;
  assign n50286 = n50285 ^ n50283 ^ 1'b0 ;
  assign n50287 = n50147 ^ n18253 ^ n8893 ;
  assign n50288 = n10406 & n14237 ;
  assign n50289 = n10209 ^ n8370 ^ n2160 ;
  assign n50290 = n41164 & ~n50289 ;
  assign n50291 = n50290 ^ n808 ^ 1'b0 ;
  assign n50292 = n11571 | n50291 ;
  assign n50293 = n40385 & ~n50292 ;
  assign n50294 = n22013 ^ n14780 ^ 1'b0 ;
  assign n50295 = n12484 ^ n5158 ^ 1'b0 ;
  assign n50296 = n50294 & n50295 ;
  assign n50297 = n16114 | n50296 ;
  assign n50299 = n37953 & n40039 ;
  assign n50300 = ~n14255 & n50299 ;
  assign n50298 = ~n5647 & n28488 ;
  assign n50301 = n50300 ^ n50298 ^ 1'b0 ;
  assign n50302 = n28107 ^ n13129 ^ 1'b0 ;
  assign n50303 = n23092 ^ n2440 ^ 1'b0 ;
  assign n50304 = n43206 & ~n50303 ;
  assign n50305 = n29305 ^ n6160 ^ 1'b0 ;
  assign n50306 = n50305 ^ n17754 ^ n2507 ;
  assign n50307 = n18320 ^ n18112 ^ 1'b0 ;
  assign n50308 = n44472 | n50307 ;
  assign n50309 = n50306 | n50308 ;
  assign n50310 = n44669 | n50309 ;
  assign n50311 = ~n12063 & n18146 ;
  assign n50312 = n50311 ^ n41213 ^ 1'b0 ;
  assign n50313 = n15513 | n50312 ;
  assign n50314 = n26551 ^ n21370 ^ 1'b0 ;
  assign n50315 = ~n37452 & n38956 ;
  assign n50316 = n9666 ^ n1372 ^ x92 ;
  assign n50317 = n9619 | n50316 ;
  assign n50318 = ~n50315 & n50317 ;
  assign n50319 = ~n19365 & n42616 ;
  assign n50320 = n32657 ^ x78 ^ 1'b0 ;
  assign n50321 = n8477 & n50320 ;
  assign n50322 = n40216 ^ n29117 ^ n2502 ;
  assign n50323 = n21014 ^ n17977 ^ 1'b0 ;
  assign n50324 = n50322 & n50323 ;
  assign n50325 = ( ~n8626 & n49576 ) | ( ~n8626 & n50324 ) | ( n49576 & n50324 ) ;
  assign n50326 = n14548 ^ x78 ^ 1'b0 ;
  assign n50327 = ( n35049 & n43577 ) | ( n35049 & ~n50326 ) | ( n43577 & ~n50326 ) ;
  assign n50328 = ( ~n1616 & n14481 ) | ( ~n1616 & n18497 ) | ( n14481 & n18497 ) ;
  assign n50329 = n50328 ^ n49843 ^ n27428 ;
  assign n50330 = ( n10289 & n33461 ) | ( n10289 & n39537 ) | ( n33461 & n39537 ) ;
  assign n50331 = n14931 | n17286 ;
  assign n50332 = n41780 ^ n40751 ^ 1'b0 ;
  assign n50333 = n18463 ^ n11181 ^ n8083 ;
  assign n50334 = ~n50332 & n50333 ;
  assign n50335 = n3209 & n18268 ;
  assign n50336 = n50335 ^ n21233 ^ 1'b0 ;
  assign n50337 = n735 & n3680 ;
  assign n50338 = ~n13236 & n50337 ;
  assign n50339 = ( ~x162 & n1494 ) | ( ~x162 & n20991 ) | ( n1494 & n20991 ) ;
  assign n50340 = n12777 & n13214 ;
  assign n50341 = n50339 & n50340 ;
  assign n50342 = ( n5741 & ~n14381 ) | ( n5741 & n50341 ) | ( ~n14381 & n50341 ) ;
  assign n50343 = ~n16971 & n27899 ;
  assign n50344 = ( n18666 & n29820 ) | ( n18666 & ~n50343 ) | ( n29820 & ~n50343 ) ;
  assign n50345 = n8669 & n17409 ;
  assign n50346 = n22605 ^ n15660 ^ 1'b0 ;
  assign n50347 = ( n48468 & n50345 ) | ( n48468 & ~n50346 ) | ( n50345 & ~n50346 ) ;
  assign n50348 = ( n3268 & n25293 ) | ( n3268 & ~n27995 ) | ( n25293 & ~n27995 ) ;
  assign n50349 = n17592 ^ n11656 ^ n2082 ;
  assign n50350 = n50349 ^ n2525 ^ 1'b0 ;
  assign n50352 = ( n12672 & n19236 ) | ( n12672 & ~n34808 ) | ( n19236 & ~n34808 ) ;
  assign n50351 = ~n4514 & n11513 ;
  assign n50353 = n50352 ^ n50351 ^ 1'b0 ;
  assign n50354 = n37248 ^ n22125 ^ 1'b0 ;
  assign n50355 = ~n50353 & n50354 ;
  assign n50358 = n17884 ^ n14284 ^ 1'b0 ;
  assign n50356 = n18891 ^ n11070 ^ 1'b0 ;
  assign n50357 = n17334 | n50356 ;
  assign n50359 = n50358 ^ n50357 ^ 1'b0 ;
  assign n50360 = n39575 ^ x14 ^ 1'b0 ;
  assign n50361 = n2444 | n40334 ;
  assign n50362 = ~n25482 & n35994 ;
  assign n50363 = n28387 & n50362 ;
  assign n50364 = n50363 ^ x47 ^ 1'b0 ;
  assign n50365 = n23402 ^ n15309 ^ 1'b0 ;
  assign n50366 = ~n4027 & n14544 ;
  assign n50367 = ~n50365 & n50366 ;
  assign n50368 = n15600 & n50367 ;
  assign n50369 = n13703 & n26693 ;
  assign n50370 = n1652 & n50369 ;
  assign n50371 = ~n21599 & n28818 ;
  assign n50372 = n50371 ^ n15875 ^ 1'b0 ;
  assign n50373 = n11619 & n18968 ;
  assign n50374 = n50373 ^ n5043 ^ 1'b0 ;
  assign n50375 = n24791 ^ n16746 ^ 1'b0 ;
  assign n50376 = x107 & ~n50375 ;
  assign n50377 = n15377 & ~n15969 ;
  assign n50378 = n46027 & n50377 ;
  assign n50379 = n28823 ^ n19424 ^ 1'b0 ;
  assign n50380 = ( n736 & n932 ) | ( n736 & ~n22035 ) | ( n932 & ~n22035 ) ;
  assign n50381 = ( ~x227 & n11869 ) | ( ~x227 & n49223 ) | ( n11869 & n49223 ) ;
  assign n50382 = n50381 ^ n41887 ^ 1'b0 ;
  assign n50383 = x89 & ~n50382 ;
  assign n50384 = n548 | n24985 ;
  assign n50385 = n15722 ^ n9870 ^ 1'b0 ;
  assign n50386 = n2127 & ~n26089 ;
  assign n50387 = ( n7250 & n15290 ) | ( n7250 & n37161 ) | ( n15290 & n37161 ) ;
  assign n50388 = n13373 & n50387 ;
  assign n50389 = ( ~n5633 & n13354 ) | ( ~n5633 & n19931 ) | ( n13354 & n19931 ) ;
  assign n50390 = n2586 & ~n48053 ;
  assign n50391 = ~n50389 & n50390 ;
  assign n50392 = n10353 & ~n44477 ;
  assign n50393 = n1975 & ~n23677 ;
  assign n50394 = ~n303 & n50393 ;
  assign n50395 = n939 & ~n14722 ;
  assign n50396 = n11823 | n50395 ;
  assign n50397 = n50394 & ~n50396 ;
  assign n50398 = ~n8383 & n17352 ;
  assign n50399 = ( n11808 & ~n41238 ) | ( n11808 & n50398 ) | ( ~n41238 & n50398 ) ;
  assign n50404 = ( n12223 & n15701 ) | ( n12223 & n28702 ) | ( n15701 & n28702 ) ;
  assign n50400 = n9759 ^ n9130 ^ 1'b0 ;
  assign n50401 = n5327 & n50400 ;
  assign n50402 = ~n1578 & n50401 ;
  assign n50403 = n50402 ^ n48514 ^ 1'b0 ;
  assign n50405 = n50404 ^ n50403 ^ n48610 ;
  assign n50406 = ( n2218 & n12992 ) | ( n2218 & ~n20208 ) | ( n12992 & ~n20208 ) ;
  assign n50407 = n43227 ^ n35445 ^ 1'b0 ;
  assign n50408 = ( ~n26663 & n30502 ) | ( ~n26663 & n43128 ) | ( n30502 & n43128 ) ;
  assign n50409 = n12516 & n23185 ;
  assign n50410 = n50409 ^ n44130 ^ 1'b0 ;
  assign n50411 = n20377 ^ n14769 ^ n3636 ;
  assign n50412 = x118 & ~n45655 ;
  assign n50413 = ~n35265 & n50412 ;
  assign n50417 = ( n5470 & n21451 ) | ( n5470 & n27023 ) | ( n21451 & n27023 ) ;
  assign n50414 = ( n2340 & n17242 ) | ( n2340 & ~n19485 ) | ( n17242 & ~n19485 ) ;
  assign n50415 = n50414 ^ n17150 ^ 1'b0 ;
  assign n50416 = ( n35594 & n42359 ) | ( n35594 & n50415 ) | ( n42359 & n50415 ) ;
  assign n50418 = n50417 ^ n50416 ^ n38543 ;
  assign n50419 = n6943 ^ n3716 ^ 1'b0 ;
  assign n50420 = n3611 & ~n50419 ;
  assign n50421 = ( n8703 & n26907 ) | ( n8703 & ~n50420 ) | ( n26907 & ~n50420 ) ;
  assign n50422 = n28099 ^ n26743 ^ n24371 ;
  assign n50423 = n32834 & ~n39589 ;
  assign n50424 = n50423 ^ n869 ^ 1'b0 ;
  assign n50425 = n50424 ^ n11627 ^ 1'b0 ;
  assign n50426 = ( n14053 & n14640 ) | ( n14053 & n35009 ) | ( n14640 & n35009 ) ;
  assign n50427 = n29355 ^ n10987 ^ n1600 ;
  assign n50431 = n17038 & n43350 ;
  assign n50432 = n50431 ^ n3133 ^ 1'b0 ;
  assign n50428 = ( n6138 & n17733 ) | ( n6138 & ~n28065 ) | ( n17733 & ~n28065 ) ;
  assign n50429 = n15968 | n50428 ;
  assign n50430 = n41741 & ~n50429 ;
  assign n50433 = n50432 ^ n50430 ^ 1'b0 ;
  assign n50434 = n48682 ^ n4005 ^ 1'b0 ;
  assign n50435 = n43298 ^ n11124 ^ 1'b0 ;
  assign n50436 = n37967 & n50435 ;
  assign n50437 = ~n23414 & n50436 ;
  assign n50438 = ~n23042 & n50437 ;
  assign n50439 = n28265 ^ n21107 ^ n20874 ;
  assign n50440 = ( n13693 & ~n17533 ) | ( n13693 & n18125 ) | ( ~n17533 & n18125 ) ;
  assign n50441 = n50440 ^ n2173 ^ n999 ;
  assign n50442 = n41667 ^ n15333 ^ n14047 ;
  assign n50443 = n39587 ^ n18438 ^ 1'b0 ;
  assign n50444 = ~n6797 & n50443 ;
  assign n50445 = n4910 ^ n2361 ^ 1'b0 ;
  assign n50446 = n726 | n33276 ;
  assign n50447 = n50445 | n50446 ;
  assign n50448 = ( n6225 & n7370 ) | ( n6225 & n23036 ) | ( n7370 & n23036 ) ;
  assign n50449 = n21561 & ~n50448 ;
  assign n50453 = n18245 & n25736 ;
  assign n50450 = n20781 ^ n11332 ^ n6124 ;
  assign n50451 = n50450 ^ n47775 ^ 1'b0 ;
  assign n50452 = ~n3281 & n50451 ;
  assign n50454 = n50453 ^ n50452 ^ n23738 ;
  assign n50455 = n50454 ^ n26093 ^ 1'b0 ;
  assign n50456 = n26802 & ~n50455 ;
  assign n50457 = n27289 ^ n3360 ^ 1'b0 ;
  assign n50458 = n33638 ^ n21838 ^ 1'b0 ;
  assign n50459 = ( n33495 & n38437 ) | ( n33495 & ~n45057 ) | ( n38437 & ~n45057 ) ;
  assign n50460 = n13916 | n18512 ;
  assign n50461 = x156 & n50460 ;
  assign n50462 = n50461 ^ n40839 ^ n26008 ;
  assign n50463 = ( n8942 & n11337 ) | ( n8942 & ~n49380 ) | ( n11337 & ~n49380 ) ;
  assign n50464 = n9387 & ~n26991 ;
  assign n50465 = n9393 & ~n22798 ;
  assign n50466 = ~n31404 & n50465 ;
  assign n50467 = ( x238 & ~n6553 ) | ( x238 & n17201 ) | ( ~n6553 & n17201 ) ;
  assign n50468 = n50467 ^ n13724 ^ 1'b0 ;
  assign n50469 = n50468 ^ n32826 ^ 1'b0 ;
  assign n50470 = n1524 | n9376 ;
  assign n50471 = n11147 & ~n50470 ;
  assign n50472 = n50471 ^ n31005 ^ 1'b0 ;
  assign n50473 = n37738 & n50472 ;
  assign n50474 = n4526 & ~n14249 ;
  assign n50475 = n45492 ^ n18896 ^ n13089 ;
  assign n50476 = ( n11107 & ~n15925 ) | ( n11107 & n50475 ) | ( ~n15925 & n50475 ) ;
  assign n50477 = n50476 ^ n2153 ^ 1'b0 ;
  assign n50478 = n17984 & ~n38254 ;
  assign n50479 = n21229 & n34029 ;
  assign n50480 = n1746 & n5169 ;
  assign n50485 = n41521 ^ n36301 ^ 1'b0 ;
  assign n50483 = n35135 ^ n18603 ^ 1'b0 ;
  assign n50484 = n48744 | n50483 ;
  assign n50481 = n9943 & n34868 ;
  assign n50482 = n50481 ^ n2143 ^ 1'b0 ;
  assign n50486 = n50485 ^ n50484 ^ n50482 ;
  assign n50487 = n50486 ^ n7870 ^ 1'b0 ;
  assign n50488 = n24084 | n50487 ;
  assign n50489 = n21646 & ~n50488 ;
  assign n50490 = ~n20479 & n49566 ;
  assign n50491 = ~n15190 & n50490 ;
  assign n50492 = n9394 ^ n4707 ^ 1'b0 ;
  assign n50493 = n12020 & ~n50492 ;
  assign n50494 = ( n3013 & n4844 ) | ( n3013 & n5936 ) | ( n4844 & n5936 ) ;
  assign n50495 = n11828 | n50494 ;
  assign n50496 = n50495 ^ n7332 ^ 1'b0 ;
  assign n50497 = n50496 ^ n46171 ^ n4918 ;
  assign n50498 = n9623 & ~n10308 ;
  assign n50499 = ~n17937 & n50498 ;
  assign n50500 = n50499 ^ n23240 ^ n19902 ;
  assign n50501 = n44545 ^ n13096 ^ n1945 ;
  assign n50502 = ( n5338 & n6931 ) | ( n5338 & ~n14963 ) | ( n6931 & ~n14963 ) ;
  assign n50503 = ( n9552 & ~n26229 ) | ( n9552 & n50502 ) | ( ~n26229 & n50502 ) ;
  assign n50504 = n17071 ^ n14255 ^ 1'b0 ;
  assign n50505 = n8980 & ~n10949 ;
  assign n50506 = ~n34309 & n50505 ;
  assign n50507 = n41768 ^ n10045 ^ n6982 ;
  assign n50508 = n22567 ^ n3584 ^ 1'b0 ;
  assign n50509 = n50507 | n50508 ;
  assign n50510 = ~n5724 & n7622 ;
  assign n50511 = n50510 ^ n12640 ^ 1'b0 ;
  assign n50512 = ~n20289 & n50511 ;
  assign n50513 = n50512 ^ n18746 ^ 1'b0 ;
  assign n50514 = n19561 & ~n19854 ;
  assign n50515 = n50514 ^ n39495 ^ 1'b0 ;
  assign n50516 = ~n6685 & n8825 ;
  assign n50517 = ~n42302 & n50516 ;
  assign n50518 = n11291 & ~n50517 ;
  assign n50519 = n20626 ^ n8385 ^ 1'b0 ;
  assign n50520 = n4337 | n23477 ;
  assign n50521 = n50520 ^ n13910 ^ 1'b0 ;
  assign n50522 = n50521 ^ n35366 ^ n19606 ;
  assign n50523 = n50522 ^ n44768 ^ n26134 ;
  assign n50524 = n33075 & ~n35693 ;
  assign n50526 = ~n5431 & n27532 ;
  assign n50525 = ~n1742 & n36277 ;
  assign n50527 = n50526 ^ n50525 ^ 1'b0 ;
  assign n50528 = ( n25275 & n32074 ) | ( n25275 & ~n50527 ) | ( n32074 & ~n50527 ) ;
  assign n50529 = n10865 & n34382 ;
  assign n50530 = n44766 ^ n27433 ^ n21061 ;
  assign n50531 = n24976 | n50530 ;
  assign n50532 = n38685 & ~n50531 ;
  assign n50533 = n49413 ^ n41754 ^ n25530 ;
  assign n50534 = n12020 & n50533 ;
  assign n50535 = n48648 ^ n12159 ^ 1'b0 ;
  assign n50536 = n20316 & n50535 ;
  assign n50537 = n50536 ^ n17502 ^ 1'b0 ;
  assign n50539 = ~n13418 & n16072 ;
  assign n50540 = n50539 ^ n12411 ^ 1'b0 ;
  assign n50538 = n7031 | n16446 ;
  assign n50541 = n50540 ^ n50538 ^ 1'b0 ;
  assign n50542 = n30271 & ~n50541 ;
  assign n50543 = n46721 ^ n41159 ^ n1091 ;
  assign n50544 = n45294 ^ n28792 ^ 1'b0 ;
  assign n50545 = n9949 ^ n7102 ^ n1969 ;
  assign n50546 = n19649 & n40115 ;
  assign n50547 = n4522 & ~n16415 ;
  assign n50548 = n50546 & n50547 ;
  assign n50549 = ~n1239 & n1924 ;
  assign n50550 = n50549 ^ n2538 ^ 1'b0 ;
  assign n50551 = n50550 ^ n14913 ^ n10161 ;
  assign n50552 = n13909 ^ n2500 ^ 1'b0 ;
  assign n50553 = n50551 & n50552 ;
  assign n50554 = n33775 ^ n18691 ^ n13444 ;
  assign n50555 = n6575 & n50554 ;
  assign n50556 = n50555 ^ n40334 ^ n8713 ;
  assign n50557 = ~n10881 & n50556 ;
  assign n50558 = n50557 ^ n41404 ^ 1'b0 ;
  assign n50561 = ( n12801 & n13423 ) | ( n12801 & ~n30144 ) | ( n13423 & ~n30144 ) ;
  assign n50559 = n12151 | n23811 ;
  assign n50560 = n7321 & ~n50559 ;
  assign n50562 = n50561 ^ n50560 ^ n2251 ;
  assign n50565 = x185 & ~n13499 ;
  assign n50563 = n13609 ^ n6377 ^ 1'b0 ;
  assign n50564 = n16754 & ~n50563 ;
  assign n50566 = n50565 ^ n50564 ^ n22559 ;
  assign n50567 = n17971 | n19857 ;
  assign n50568 = n47276 & ~n50567 ;
  assign n50569 = n17015 ^ n14342 ^ n9134 ;
  assign n50570 = ( n35916 & n38239 ) | ( n35916 & ~n50569 ) | ( n38239 & ~n50569 ) ;
  assign n50571 = n40167 ^ n4306 ^ 1'b0 ;
  assign n50572 = n50571 ^ n47887 ^ n12182 ;
  assign n50573 = n43075 & n48125 ;
  assign n50574 = n20531 | n21584 ;
  assign n50575 = n50574 ^ n4499 ^ 1'b0 ;
  assign n50576 = n12571 & ~n40179 ;
  assign n50577 = ( n4327 & n10269 ) | ( n4327 & n22202 ) | ( n10269 & n22202 ) ;
  assign n50578 = n50577 ^ n8538 ^ 1'b0 ;
  assign n50579 = n42050 ^ n26680 ^ 1'b0 ;
  assign n50580 = n47630 ^ n8702 ^ 1'b0 ;
  assign n50581 = n38800 & n43918 ;
  assign n50582 = n17554 ^ n10603 ^ 1'b0 ;
  assign n50583 = n8385 & ~n50582 ;
  assign n50584 = n50583 ^ n36886 ^ 1'b0 ;
  assign n50585 = ( n933 & n26116 ) | ( n933 & n34940 ) | ( n26116 & n34940 ) ;
  assign n50586 = n16426 & n19753 ;
  assign n50587 = ~x203 & n50586 ;
  assign n50588 = n9072 | n9334 ;
  assign n50589 = n37955 & n50588 ;
  assign n50590 = ~n272 & n5044 ;
  assign n50591 = n50590 ^ n8275 ^ 1'b0 ;
  assign n50592 = n5173 & n19095 ;
  assign n50593 = ~n17877 & n31249 ;
  assign n50594 = n14244 ^ n9420 ^ n5669 ;
  assign n50595 = n50594 ^ n9808 ^ n687 ;
  assign n50596 = n50595 ^ n44515 ^ n1672 ;
  assign n50597 = ( ~n44641 & n50593 ) | ( ~n44641 & n50596 ) | ( n50593 & n50596 ) ;
  assign n50598 = ( n29211 & ~n50592 ) | ( n29211 & n50597 ) | ( ~n50592 & n50597 ) ;
  assign n50599 = n28325 ^ n27365 ^ n3347 ;
  assign n50600 = n48129 ^ n17518 ^ n10763 ;
  assign n50601 = n27426 | n31831 ;
  assign n50602 = n35612 ^ n4858 ^ 1'b0 ;
  assign n50603 = ~n13421 & n50602 ;
  assign n50604 = n14564 & n17008 ;
  assign n50605 = n50604 ^ n33012 ^ 1'b0 ;
  assign n50606 = n50603 & ~n50605 ;
  assign n50607 = n21319 ^ n14081 ^ 1'b0 ;
  assign n50612 = ( n3246 & ~n6523 ) | ( n3246 & n20296 ) | ( ~n6523 & n20296 ) ;
  assign n50613 = n50612 ^ n16025 ^ n3761 ;
  assign n50608 = n12365 | n24152 ;
  assign n50609 = n6683 & ~n50608 ;
  assign n50610 = n50609 ^ n25359 ^ n20446 ;
  assign n50611 = ( ~n21606 & n23724 ) | ( ~n21606 & n50610 ) | ( n23724 & n50610 ) ;
  assign n50614 = n50613 ^ n50611 ^ 1'b0 ;
  assign n50615 = n26310 & n39233 ;
  assign n50616 = n50615 ^ n19995 ^ 1'b0 ;
  assign n50617 = ~n47399 & n50616 ;
  assign n50618 = n33635 ^ n29353 ^ 1'b0 ;
  assign n50619 = n12886 | n48293 ;
  assign n50620 = n50618 | n50619 ;
  assign n50621 = n13942 ^ n9165 ^ 1'b0 ;
  assign n50622 = n21468 ^ n19659 ^ 1'b0 ;
  assign n50623 = ( n7161 & ~n50621 ) | ( n7161 & n50622 ) | ( ~n50621 & n50622 ) ;
  assign n50624 = n29193 & n39733 ;
  assign n50625 = n50624 ^ n25369 ^ 1'b0 ;
  assign n50626 = n50625 ^ n3136 ^ 1'b0 ;
  assign n50627 = n3742 ^ n2725 ^ 1'b0 ;
  assign n50628 = ~n3510 & n50627 ;
  assign n50629 = n50628 ^ n9161 ^ 1'b0 ;
  assign n50630 = n50629 ^ n39375 ^ n4124 ;
  assign n50631 = n7209 & n18216 ;
  assign n50632 = n50631 ^ n17259 ^ 1'b0 ;
  assign n50633 = n15722 | n50632 ;
  assign n50634 = n43119 ^ n25204 ^ 1'b0 ;
  assign n50635 = ( n20858 & n50633 ) | ( n20858 & ~n50634 ) | ( n50633 & ~n50634 ) ;
  assign n50636 = n3437 | n5208 ;
  assign n50637 = n5307 ^ n5125 ^ 1'b0 ;
  assign n50638 = n15486 & ~n50637 ;
  assign n50639 = n50638 ^ n34712 ^ 1'b0 ;
  assign n50642 = n18769 | n28391 ;
  assign n50640 = n29680 ^ n23728 ^ n7576 ;
  assign n50641 = n33277 & ~n50640 ;
  assign n50643 = n50642 ^ n50641 ^ 1'b0 ;
  assign n50644 = n14113 & n21152 ;
  assign n50645 = n50644 ^ n17943 ^ 1'b0 ;
  assign n50646 = n48743 ^ n39639 ^ 1'b0 ;
  assign n50647 = ~n5440 & n50646 ;
  assign n50648 = n18159 & ~n37395 ;
  assign n50649 = ~n13903 & n50648 ;
  assign n50650 = ~n3960 & n11367 ;
  assign n50651 = ~n5188 & n50650 ;
  assign n50652 = n3901 & n50651 ;
  assign n50653 = n37183 ^ n14776 ^ n14407 ;
  assign n50654 = n27602 & ~n50653 ;
  assign n50655 = ( n18819 & ~n44591 ) | ( n18819 & n50654 ) | ( ~n44591 & n50654 ) ;
  assign n50656 = n50655 ^ n21090 ^ n16441 ;
  assign n50658 = ~n4849 & n34940 ;
  assign n50657 = n19047 | n23114 ;
  assign n50659 = n50658 ^ n50657 ^ n32121 ;
  assign n50660 = n683 & n22092 ;
  assign n50662 = ( n12129 & n19230 ) | ( n12129 & n19951 ) | ( n19230 & n19951 ) ;
  assign n50661 = n49268 ^ n44284 ^ n1178 ;
  assign n50663 = n50662 ^ n50661 ^ n2770 ;
  assign n50664 = n29040 ^ n9174 ^ 1'b0 ;
  assign n50665 = n40759 & n50664 ;
  assign n50666 = n3732 | n50665 ;
  assign n50667 = n9489 & n50666 ;
  assign n50668 = n50667 ^ n1464 ^ 1'b0 ;
  assign n50669 = ~n48417 & n50668 ;
  assign n50670 = n50669 ^ n12726 ^ 1'b0 ;
  assign n50671 = n18115 & ~n24067 ;
  assign n50672 = ~n2944 & n50671 ;
  assign n50673 = ( ~n18595 & n50554 ) | ( ~n18595 & n50672 ) | ( n50554 & n50672 ) ;
  assign n50674 = ~n3012 & n6518 ;
  assign n50675 = n26637 & n50674 ;
  assign n50676 = n50675 ^ n26994 ^ 1'b0 ;
  assign n50677 = ~n50673 & n50676 ;
  assign n50678 = n13456 ^ n8560 ^ 1'b0 ;
  assign n50679 = n50678 ^ n35572 ^ n18070 ;
  assign n50680 = n50679 ^ n34703 ^ 1'b0 ;
  assign n50681 = n31111 & ~n50680 ;
  assign n50682 = ~n22798 & n28936 ;
  assign n50683 = n12353 ^ n8200 ^ n6336 ;
  assign n50684 = n48206 ^ n37441 ^ 1'b0 ;
  assign n50685 = n5874 & n13024 ;
  assign n50686 = n50685 ^ n317 ^ 1'b0 ;
  assign n50687 = n50686 ^ n49415 ^ n2339 ;
  assign n50688 = n50687 ^ n21844 ^ n18222 ;
  assign n50689 = n50688 ^ n28252 ^ n12617 ;
  assign n50690 = n13856 ^ n13352 ^ 1'b0 ;
  assign n50692 = ~n10325 & n26184 ;
  assign n50693 = ~n10922 & n50692 ;
  assign n50691 = ~n17533 & n32106 ;
  assign n50694 = n50693 ^ n50691 ^ 1'b0 ;
  assign n50695 = ( ~n11132 & n50690 ) | ( ~n11132 & n50694 ) | ( n50690 & n50694 ) ;
  assign n50696 = n46371 ^ n10550 ^ n9018 ;
  assign n50697 = n44115 | n50696 ;
  assign n50698 = n9881 & ~n50697 ;
  assign n50699 = n50698 ^ n35352 ^ n4423 ;
  assign n50700 = ( n21470 & ~n21706 ) | ( n21470 & n42093 ) | ( ~n21706 & n42093 ) ;
  assign n50701 = n8220 ^ n912 ^ 1'b0 ;
  assign n50702 = ~n50700 & n50701 ;
  assign n50703 = ~n6083 & n50358 ;
  assign n50704 = ~n11568 & n17679 ;
  assign n50705 = n50703 & n50704 ;
  assign n50706 = ~n9956 & n26708 ;
  assign n50707 = ( n1903 & n37076 ) | ( n1903 & n38712 ) | ( n37076 & n38712 ) ;
  assign n50708 = n19395 & ~n50707 ;
  assign n50709 = n50708 ^ n3716 ^ 1'b0 ;
  assign n50710 = n17703 ^ n12113 ^ 1'b0 ;
  assign n50711 = n5074 & n50710 ;
  assign n50712 = ~n4192 & n12163 ;
  assign n50713 = n50711 & n50712 ;
  assign n50714 = n46921 ^ n19319 ^ n12899 ;
  assign n50715 = ~n10661 & n11419 ;
  assign n50716 = n9956 & n50715 ;
  assign n50717 = ( n5044 & n5082 ) | ( n5044 & n50716 ) | ( n5082 & n50716 ) ;
  assign n50718 = n47844 ^ n39316 ^ n20889 ;
  assign n50719 = n12254 & ~n14467 ;
  assign n50720 = n22415 | n50719 ;
  assign n50721 = ( n31871 & n50718 ) | ( n31871 & ~n50720 ) | ( n50718 & ~n50720 ) ;
  assign n50722 = n35625 ^ n3565 ^ n1822 ;
  assign n50723 = n8096 & ~n29983 ;
  assign n50724 = n24750 & n50723 ;
  assign n50725 = n19531 ^ n9665 ^ 1'b0 ;
  assign n50726 = n22421 & ~n50725 ;
  assign n50727 = n50724 & n50726 ;
  assign n50728 = ( n1645 & ~n15170 ) | ( n1645 & n16458 ) | ( ~n15170 & n16458 ) ;
  assign n50729 = ( n25715 & n29914 ) | ( n25715 & ~n50728 ) | ( n29914 & ~n50728 ) ;
  assign n50730 = n50729 ^ n3605 ^ 1'b0 ;
  assign n50731 = n36527 | n50730 ;
  assign n50732 = n27855 ^ n14678 ^ 1'b0 ;
  assign n50733 = n42754 | n50732 ;
  assign n50734 = n50733 ^ n8159 ^ 1'b0 ;
  assign n50735 = n43433 ^ n39152 ^ n5650 ;
  assign n50736 = ( n15558 & n32953 ) | ( n15558 & ~n41003 ) | ( n32953 & ~n41003 ) ;
  assign n50737 = n8726 ^ n757 ^ 1'b0 ;
  assign n50738 = n5331 & n45708 ;
  assign n50739 = n41741 | n50289 ;
  assign n50740 = n50739 ^ n8271 ^ 1'b0 ;
  assign n50741 = n20660 | n28893 ;
  assign n50742 = n50741 ^ n487 ^ 1'b0 ;
  assign n50743 = n37760 ^ n11512 ^ 1'b0 ;
  assign n50744 = ~x14 & n8339 ;
  assign n50745 = n38188 ^ n21816 ^ 1'b0 ;
  assign n50746 = n32548 | n50745 ;
  assign n50747 = ( ~n13969 & n50744 ) | ( ~n13969 & n50746 ) | ( n50744 & n50746 ) ;
  assign n50748 = n34600 ^ n15433 ^ 1'b0 ;
  assign n50749 = n44774 ^ n41041 ^ 1'b0 ;
  assign n50750 = n50147 & n50749 ;
  assign n50751 = n9851 ^ n6101 ^ 1'b0 ;
  assign n50752 = n17169 | n50751 ;
  assign n50753 = n50752 ^ n48602 ^ 1'b0 ;
  assign n50754 = ( ~n13667 & n34078 ) | ( ~n13667 & n37332 ) | ( n34078 & n37332 ) ;
  assign n50755 = n5639 & n39273 ;
  assign n50756 = n50179 ^ n2965 ^ 1'b0 ;
  assign n50757 = n5811 | n46917 ;
  assign n50758 = n50757 ^ n9590 ^ 1'b0 ;
  assign n50759 = ~n38020 & n38466 ;
  assign n50760 = n39276 ^ n12018 ^ 1'b0 ;
  assign n50761 = n50759 | n50760 ;
  assign n50762 = n50761 ^ n11536 ^ n4421 ;
  assign n50763 = n16836 ^ n16488 ^ 1'b0 ;
  assign n50764 = n50762 & ~n50763 ;
  assign n50765 = n15072 ^ n14244 ^ 1'b0 ;
  assign n50766 = n5231 & n50765 ;
  assign n50767 = n43173 ^ n27854 ^ n26799 ;
  assign n50768 = n43532 ^ n24353 ^ n16526 ;
  assign n50769 = n901 | n3982 ;
  assign n50770 = ~n13299 & n50769 ;
  assign n50771 = n11147 | n16707 ;
  assign n50772 = ( ~n1266 & n4544 ) | ( ~n1266 & n50771 ) | ( n4544 & n50771 ) ;
  assign n50773 = n50772 ^ n30679 ^ n9340 ;
  assign n50774 = n2623 & ~n9911 ;
  assign n50775 = n14944 & n40963 ;
  assign n50776 = n31164 & n50775 ;
  assign n50777 = n31854 ^ n19184 ^ 1'b0 ;
  assign n50778 = n20229 | n50777 ;
  assign n50779 = n43499 ^ n30882 ^ n10806 ;
  assign n50780 = ( ~n17049 & n18063 ) | ( ~n17049 & n47055 ) | ( n18063 & n47055 ) ;
  assign n50781 = n43484 ^ n33687 ^ n11146 ;
  assign n50782 = n17237 ^ x144 ^ 1'b0 ;
  assign n50783 = n24235 ^ n22977 ^ 1'b0 ;
  assign n50784 = n16001 & ~n50783 ;
  assign n50785 = ~n7846 & n50784 ;
  assign n50786 = n50785 ^ n21046 ^ 1'b0 ;
  assign n50787 = n44109 ^ n7383 ^ 1'b0 ;
  assign n50788 = ( n13291 & ~n14062 ) | ( n13291 & n27058 ) | ( ~n14062 & n27058 ) ;
  assign n50789 = n50788 ^ n34925 ^ n1639 ;
  assign n50790 = n50789 ^ n7890 ^ 1'b0 ;
  assign n50791 = ( x72 & n2490 ) | ( x72 & ~n18652 ) | ( n2490 & ~n18652 ) ;
  assign n50792 = n50791 ^ n41537 ^ n24080 ;
  assign n50793 = n37464 ^ n17614 ^ n311 ;
  assign n50794 = ( n4435 & ~n11490 ) | ( n4435 & n17614 ) | ( ~n11490 & n17614 ) ;
  assign n50795 = x82 & ~n29324 ;
  assign n50796 = n50795 ^ n20826 ^ n11208 ;
  assign n50797 = n40321 ^ n30116 ^ 1'b0 ;
  assign n50798 = n4248 & n43507 ;
  assign n50799 = n15766 | n21590 ;
  assign n50800 = n50799 ^ n13843 ^ 1'b0 ;
  assign n50801 = n50800 ^ n12572 ^ 1'b0 ;
  assign n50802 = ~n40922 & n50801 ;
  assign n50803 = n23640 ^ n23059 ^ 1'b0 ;
  assign n50804 = n21229 ^ n3431 ^ 1'b0 ;
  assign n50805 = ~n50803 & n50804 ;
  assign n50806 = n50019 ^ n31836 ^ 1'b0 ;
  assign n50807 = n5189 & n50806 ;
  assign n50808 = n5244 ^ n2354 ^ 1'b0 ;
  assign n50809 = n6064 | n50808 ;
  assign n50810 = ( n18085 & n36176 ) | ( n18085 & ~n39721 ) | ( n36176 & ~n39721 ) ;
  assign n50811 = n23882 | n36479 ;
  assign n50812 = n50811 ^ n35529 ^ n28853 ;
  assign n50817 = n5320 & n12685 ;
  assign n50818 = n50817 ^ n3732 ^ 1'b0 ;
  assign n50815 = n31916 ^ n1356 ^ 1'b0 ;
  assign n50813 = n7966 & ~n18916 ;
  assign n50814 = ~n20817 & n50813 ;
  assign n50816 = n50815 ^ n50814 ^ 1'b0 ;
  assign n50819 = n50818 ^ n50816 ^ n7998 ;
  assign n50820 = n39170 ^ n23644 ^ n5264 ;
  assign n50821 = x56 & ~n14826 ;
  assign n50822 = ~n50820 & n50821 ;
  assign n50823 = ( n2782 & n22083 ) | ( n2782 & ~n50822 ) | ( n22083 & ~n50822 ) ;
  assign n50824 = ~n3257 & n19976 ;
  assign n50825 = n16804 | n50824 ;
  assign n50826 = n50825 ^ n37904 ^ 1'b0 ;
  assign n50827 = x69 & ~n15864 ;
  assign n50828 = ~n13208 & n50827 ;
  assign n50829 = n37681 | n50828 ;
  assign n50830 = n50829 ^ n36473 ^ 1'b0 ;
  assign n50832 = ~n10599 & n20146 ;
  assign n50831 = ~n37384 & n49155 ;
  assign n50833 = n50832 ^ n50831 ^ 1'b0 ;
  assign n50835 = n43122 ^ n13951 ^ n1229 ;
  assign n50836 = n50835 ^ n14611 ^ n4256 ;
  assign n50837 = n20683 ^ n15904 ^ 1'b0 ;
  assign n50838 = ( n16276 & ~n50836 ) | ( n16276 & n50837 ) | ( ~n50836 & n50837 ) ;
  assign n50834 = n10571 | n17696 ;
  assign n50839 = n50838 ^ n50834 ^ 1'b0 ;
  assign n50840 = n7555 & ~n10792 ;
  assign n50845 = n7786 ^ n5604 ^ 1'b0 ;
  assign n50841 = x214 & ~n7127 ;
  assign n50842 = n5500 & n50841 ;
  assign n50843 = ( n38285 & n39784 ) | ( n38285 & n40834 ) | ( n39784 & n40834 ) ;
  assign n50844 = ( n33994 & n50842 ) | ( n33994 & ~n50843 ) | ( n50842 & ~n50843 ) ;
  assign n50846 = n50845 ^ n50844 ^ n28972 ;
  assign n50847 = n27764 & ~n28680 ;
  assign n50848 = n50847 ^ n9866 ^ 1'b0 ;
  assign n50849 = ~n289 & n50848 ;
  assign n50850 = n50849 ^ n7246 ^ 1'b0 ;
  assign n50851 = n50850 ^ n34422 ^ 1'b0 ;
  assign n50852 = n11599 | n19643 ;
  assign n50853 = n50852 ^ x64 ^ 1'b0 ;
  assign n50854 = n50853 ^ n25167 ^ n4975 ;
  assign n50855 = n50854 ^ n3268 ^ 1'b0 ;
  assign n50856 = n50855 ^ n20220 ^ n6864 ;
  assign n50857 = ~n28649 & n46920 ;
  assign n50858 = n30093 & n50857 ;
  assign n50859 = n2542 & ~n16244 ;
  assign n50860 = n18667 | n42616 ;
  assign n50861 = ~n19507 & n24565 ;
  assign n50862 = n50861 ^ n469 ^ 1'b0 ;
  assign n50863 = n27549 & ~n50862 ;
  assign n50864 = n2807 ^ n468 ^ 1'b0 ;
  assign n50865 = ~n7534 & n50864 ;
  assign n50866 = n6401 & n50865 ;
  assign n50867 = ~n12233 & n50866 ;
  assign n50868 = n18354 & ~n31069 ;
  assign n50869 = ~n31259 & n50868 ;
  assign n50870 = n11169 ^ n1785 ^ 1'b0 ;
  assign n50871 = ~n23868 & n50870 ;
  assign n50872 = n50871 ^ n38758 ^ 1'b0 ;
  assign n50873 = n49788 ^ n20192 ^ n9262 ;
  assign n50874 = n50873 ^ n22297 ^ n18000 ;
  assign n50875 = n35180 ^ n32068 ^ n4046 ;
  assign n50876 = n23279 ^ n2761 ^ 1'b0 ;
  assign n50877 = ( n13613 & ~n21245 ) | ( n13613 & n23247 ) | ( ~n21245 & n23247 ) ;
  assign n50878 = n46994 ^ n9501 ^ 1'b0 ;
  assign n50879 = n50877 & ~n50878 ;
  assign n50880 = ( n1806 & n11723 ) | ( n1806 & ~n21818 ) | ( n11723 & ~n21818 ) ;
  assign n50881 = n50880 ^ n853 ^ 1'b0 ;
  assign n50882 = n10772 ^ n6962 ^ 1'b0 ;
  assign n50883 = n597 & n50882 ;
  assign n50884 = n9275 | n24318 ;
  assign n50885 = n1656 & ~n50884 ;
  assign n50886 = ( n2284 & ~n21869 ) | ( n2284 & n50885 ) | ( ~n21869 & n50885 ) ;
  assign n50887 = n50886 ^ n25008 ^ 1'b0 ;
  assign n50888 = n50883 & ~n50887 ;
  assign n50889 = x3 & ~n10829 ;
  assign n50890 = n13798 | n45801 ;
  assign n50891 = n21382 & ~n46329 ;
  assign n50892 = n18638 & n50891 ;
  assign n50893 = ( n32362 & n36843 ) | ( n32362 & ~n50892 ) | ( n36843 & ~n50892 ) ;
  assign n50894 = ( ~n11609 & n35648 ) | ( ~n11609 & n41751 ) | ( n35648 & n41751 ) ;
  assign n50895 = n9475 & n17315 ;
  assign n50896 = n50895 ^ n48477 ^ n29652 ;
  assign n50897 = n20332 ^ n6995 ^ 1'b0 ;
  assign n50898 = n36350 & ~n50897 ;
  assign n50899 = n50898 ^ n10483 ^ 1'b0 ;
  assign n50900 = n50899 ^ n19773 ^ n7264 ;
  assign n50901 = ( n3923 & ~n14501 ) | ( n3923 & n23146 ) | ( ~n14501 & n23146 ) ;
  assign n50902 = ( ~n9293 & n22633 ) | ( ~n9293 & n23114 ) | ( n22633 & n23114 ) ;
  assign n50903 = n50901 | n50902 ;
  assign n50904 = ( ~n13161 & n16716 ) | ( ~n13161 & n34355 ) | ( n16716 & n34355 ) ;
  assign n50905 = n50904 ^ n40494 ^ 1'b0 ;
  assign n50906 = n30222 ^ n3571 ^ 1'b0 ;
  assign n50907 = n50905 & n50906 ;
  assign n50908 = n973 & ~n12556 ;
  assign n50909 = n9951 | n50908 ;
  assign n50910 = n46129 ^ n6252 ^ 1'b0 ;
  assign n50911 = n9861 ^ n9287 ^ 1'b0 ;
  assign n50912 = n50910 | n50911 ;
  assign n50913 = n16336 | n22082 ;
  assign n50914 = ( n1345 & n17442 ) | ( n1345 & ~n50913 ) | ( n17442 & ~n50913 ) ;
  assign n50915 = n50914 ^ n13297 ^ 1'b0 ;
  assign n50916 = n50915 ^ n25318 ^ n23701 ;
  assign n50917 = n50088 ^ n34260 ^ n1166 ;
  assign n50918 = ( ~n17806 & n27012 ) | ( ~n17806 & n50917 ) | ( n27012 & n50917 ) ;
  assign n50919 = ( n48408 & n49104 ) | ( n48408 & ~n50918 ) | ( n49104 & ~n50918 ) ;
  assign n50920 = ~n2771 & n19587 ;
  assign n50921 = n50920 ^ n20417 ^ 1'b0 ;
  assign n50922 = ( n28659 & ~n38772 ) | ( n28659 & n50921 ) | ( ~n38772 & n50921 ) ;
  assign n50923 = n11605 & ~n24619 ;
  assign n50924 = n41954 ^ n39058 ^ 1'b0 ;
  assign n50925 = n50923 & n50924 ;
  assign n50926 = n50925 ^ n36381 ^ n30630 ;
  assign n50927 = n20742 ^ n14725 ^ 1'b0 ;
  assign n50928 = n6949 ^ n6005 ^ 1'b0 ;
  assign n50929 = n19462 & n50928 ;
  assign n50930 = ( n8080 & ~n21488 ) | ( n8080 & n50929 ) | ( ~n21488 & n50929 ) ;
  assign n50931 = n50927 & n50930 ;
  assign n50932 = n44507 ^ n43344 ^ 1'b0 ;
  assign n50933 = ~n2135 & n18896 ;
  assign n50934 = n50933 ^ n12007 ^ 1'b0 ;
  assign n50935 = n20096 & ~n40902 ;
  assign n50936 = ~n23472 & n50935 ;
  assign n50937 = n37034 & ~n44937 ;
  assign n50938 = n50937 ^ n49126 ^ 1'b0 ;
  assign n50939 = n21565 ^ n10386 ^ 1'b0 ;
  assign n50940 = ~n6307 & n8122 ;
  assign n50941 = ~n50939 & n50940 ;
  assign n50942 = n48210 ^ n36391 ^ n25669 ;
  assign n50943 = n10835 ^ n7801 ^ n6376 ;
  assign n50944 = n4984 | n26578 ;
  assign n50945 = n50944 ^ n29177 ^ n12060 ;
  assign n50946 = n49759 ^ n12780 ^ n9330 ;
  assign n50947 = n26348 ^ n7929 ^ 1'b0 ;
  assign n50948 = n13659 | n29851 ;
  assign n50949 = n50948 ^ n5302 ^ 1'b0 ;
  assign n50950 = n8212 & ~n21724 ;
  assign n50951 = n37518 ^ n11901 ^ 1'b0 ;
  assign n50952 = n12607 & n50951 ;
  assign n50953 = n17947 & n50952 ;
  assign n50954 = ~n521 & n50953 ;
  assign n50955 = ~n13840 & n18497 ;
  assign n50959 = n11086 & n19233 ;
  assign n50960 = n50959 ^ n19724 ^ 1'b0 ;
  assign n50956 = n8030 | n21456 ;
  assign n50957 = n50956 ^ n16381 ^ 1'b0 ;
  assign n50958 = ~n7322 & n50957 ;
  assign n50961 = n50960 ^ n50958 ^ n14892 ;
  assign n50962 = n3322 & n10142 ;
  assign n50963 = n23477 ^ n19621 ^ 1'b0 ;
  assign n50964 = ( n45673 & n50962 ) | ( n45673 & n50963 ) | ( n50962 & n50963 ) ;
  assign n50965 = ( n1359 & n3569 ) | ( n1359 & ~n3717 ) | ( n3569 & ~n3717 ) ;
  assign n50966 = n13065 ^ n8894 ^ n3345 ;
  assign n50967 = ( n40761 & ~n50965 ) | ( n40761 & n50966 ) | ( ~n50965 & n50966 ) ;
  assign n50968 = ( ~n5516 & n21340 ) | ( ~n5516 & n35008 ) | ( n21340 & n35008 ) ;
  assign n50969 = n50968 ^ n25091 ^ n13059 ;
  assign n50970 = ( n5054 & ~n26552 ) | ( n5054 & n32316 ) | ( ~n26552 & n32316 ) ;
  assign n50972 = n24760 & n35452 ;
  assign n50973 = n35938 | n50972 ;
  assign n50971 = ~n12936 & n23467 ;
  assign n50974 = n50973 ^ n50971 ^ 1'b0 ;
  assign n50975 = n46224 | n49375 ;
  assign n50976 = n4304 & n45634 ;
  assign n50977 = ~n13849 & n29304 ;
  assign n50978 = ~n6442 & n50977 ;
  assign n50979 = n5104 & ~n25697 ;
  assign n50980 = n50978 & n50979 ;
  assign n50981 = n8560 & ~n30215 ;
  assign n50982 = n1854 & n45044 ;
  assign n50983 = n50982 ^ n41360 ^ 1'b0 ;
  assign n50984 = n50983 ^ n27487 ^ n6468 ;
  assign n50985 = n39731 ^ n14758 ^ n5003 ;
  assign n50986 = ~n11057 & n50985 ;
  assign n50987 = ( n1166 & n30166 ) | ( n1166 & n35819 ) | ( n30166 & n35819 ) ;
  assign n50988 = n37574 ^ n2548 ^ 1'b0 ;
  assign n50989 = n12179 & ~n14019 ;
  assign n50990 = n32269 ^ n5125 ^ n4037 ;
  assign n50991 = n32369 | n33463 ;
  assign n50992 = n50990 | n50991 ;
  assign n50993 = n38922 ^ n20867 ^ 1'b0 ;
  assign n50994 = n6849 & n50993 ;
  assign n50995 = n15406 ^ n3377 ^ 1'b0 ;
  assign n50996 = n43442 ^ n23383 ^ 1'b0 ;
  assign n51001 = ~n2197 & n7860 ;
  assign n51002 = ~n7518 & n51001 ;
  assign n51003 = ( n2585 & ~n40960 ) | ( n2585 & n51002 ) | ( ~n40960 & n51002 ) ;
  assign n50999 = ~n3402 & n13689 ;
  assign n50997 = n39522 ^ n19347 ^ n15969 ;
  assign n50998 = n27538 & ~n50997 ;
  assign n51000 = n50999 ^ n50998 ^ 1'b0 ;
  assign n51004 = n51003 ^ n51000 ^ n24997 ;
  assign n51006 = ~n429 & n7957 ;
  assign n51007 = ~n7957 & n51006 ;
  assign n51008 = n51007 ^ x156 ^ 1'b0 ;
  assign n51009 = n51008 ^ n19870 ^ n512 ;
  assign n51010 = ( n330 & n6800 ) | ( n330 & n51009 ) | ( n6800 & n51009 ) ;
  assign n51005 = n50965 ^ n5697 ^ n3220 ;
  assign n51011 = n51010 ^ n51005 ^ n4524 ;
  assign n51012 = n32377 & n51011 ;
  assign n51013 = n39238 ^ n18384 ^ n11803 ;
  assign n51014 = ( x171 & ~n6913 ) | ( x171 & n51013 ) | ( ~n6913 & n51013 ) ;
  assign n51015 = n18725 ^ n5685 ^ 1'b0 ;
  assign n51016 = ~n15596 & n51015 ;
  assign n51017 = ( n3205 & n15921 ) | ( n3205 & ~n51016 ) | ( n15921 & ~n51016 ) ;
  assign n51018 = n40761 ^ n24670 ^ 1'b0 ;
  assign n51019 = n18338 & ~n51018 ;
  assign n51020 = n37586 ^ n2403 ^ n832 ;
  assign n51021 = n51020 ^ n1840 ^ 1'b0 ;
  assign n51022 = ( n25433 & n33183 ) | ( n25433 & n49099 ) | ( n33183 & n49099 ) ;
  assign n51023 = n10735 | n51022 ;
  assign n51024 = n51023 ^ n21187 ^ 1'b0 ;
  assign n51025 = n42462 ^ n29965 ^ 1'b0 ;
  assign n51026 = ~n3502 & n7395 ;
  assign n51027 = n11741 & n51026 ;
  assign n51028 = ( n17240 & ~n20896 ) | ( n17240 & n51027 ) | ( ~n20896 & n51027 ) ;
  assign n51029 = n51028 ^ n24263 ^ 1'b0 ;
  assign n51030 = ~n51025 & n51029 ;
  assign n51031 = x123 & n18079 ;
  assign n51032 = n9366 & n51031 ;
  assign n51033 = n49866 ^ n45684 ^ n25957 ;
  assign n51034 = n42952 | n43075 ;
  assign n51035 = ( n4363 & n6739 ) | ( n4363 & ~n36797 ) | ( n6739 & ~n36797 ) ;
  assign n51036 = n836 | n16298 ;
  assign n51037 = n51035 | n51036 ;
  assign n51038 = n9420 & n51037 ;
  assign n51039 = n32453 ^ n13391 ^ 1'b0 ;
  assign n51040 = ~n45497 & n51039 ;
  assign n51041 = ~n49235 & n51040 ;
  assign n51042 = n3381 & ~n29963 ;
  assign n51043 = ~n4639 & n51042 ;
  assign n51044 = n5675 | n45348 ;
  assign n51045 = n51044 ^ n45211 ^ 1'b0 ;
  assign n51046 = ( ~n22348 & n23434 ) | ( ~n22348 & n51045 ) | ( n23434 & n51045 ) ;
  assign n51047 = n15220 | n22694 ;
  assign n51048 = n1804 | n51047 ;
  assign n51049 = ( n51043 & n51046 ) | ( n51043 & n51048 ) | ( n51046 & n51048 ) ;
  assign n51050 = n12845 | n42392 ;
  assign n51051 = n51050 ^ n7921 ^ 1'b0 ;
  assign n51052 = n51051 ^ n13527 ^ 1'b0 ;
  assign n51053 = n1124 | n16523 ;
  assign n51054 = n47155 & n48327 ;
  assign n51055 = n51054 ^ n21094 ^ 1'b0 ;
  assign n51056 = n2573 & ~n14130 ;
  assign n51057 = n51056 ^ n47763 ^ 1'b0 ;
  assign n51058 = n11681 & ~n51057 ;
  assign n51059 = n51058 ^ n10242 ^ n5941 ;
  assign n51060 = ~n44344 & n51059 ;
  assign n51061 = n30001 & n51060 ;
  assign n51062 = n33901 & n43998 ;
  assign n51063 = ( n24094 & n28358 ) | ( n24094 & ~n31929 ) | ( n28358 & ~n31929 ) ;
  assign n51064 = n13964 ^ n10481 ^ n8408 ;
  assign n51065 = n37250 & ~n50791 ;
  assign n51066 = n24518 & n46505 ;
  assign n51067 = ( n6001 & n28611 ) | ( n6001 & n51066 ) | ( n28611 & n51066 ) ;
  assign n51068 = n16152 ^ n4003 ^ 1'b0 ;
  assign n51069 = n49606 & ~n51068 ;
  assign n51070 = n18191 ^ n6076 ^ 1'b0 ;
  assign n51071 = n16966 ^ n6390 ^ 1'b0 ;
  assign n51072 = ~n30684 & n36553 ;
  assign n51073 = ( n33844 & n51071 ) | ( n33844 & ~n51072 ) | ( n51071 & ~n51072 ) ;
  assign n51074 = n28574 ^ n2877 ^ 1'b0 ;
  assign n51075 = n16037 ^ n15166 ^ 1'b0 ;
  assign n51076 = n34574 & ~n51075 ;
  assign n51077 = n36012 | n51076 ;
  assign n51078 = n51071 ^ n41892 ^ 1'b0 ;
  assign n51079 = n32284 ^ n8405 ^ 1'b0 ;
  assign n51080 = n5932 | n28477 ;
  assign n51081 = n7802 | n51080 ;
  assign n51082 = n29301 ^ n20191 ^ n10542 ;
  assign n51084 = n13642 & n21431 ;
  assign n51083 = ~n28199 & n44048 ;
  assign n51085 = n51084 ^ n51083 ^ n31974 ;
  assign n51086 = n9359 ^ n4930 ^ 1'b0 ;
  assign n51087 = n10483 & ~n11437 ;
  assign n51088 = n51087 ^ n13711 ^ 1'b0 ;
  assign n51089 = n30915 & ~n51088 ;
  assign n51090 = ( n9799 & n51086 ) | ( n9799 & ~n51089 ) | ( n51086 & ~n51089 ) ;
  assign n51091 = ( n10303 & ~n23841 ) | ( n10303 & n51090 ) | ( ~n23841 & n51090 ) ;
  assign n51092 = n21118 ^ n14803 ^ n11454 ;
  assign n51093 = ( n2958 & n10976 ) | ( n2958 & ~n51092 ) | ( n10976 & ~n51092 ) ;
  assign n51094 = n3444 & ~n34077 ;
  assign n51095 = n23968 ^ n5262 ^ n1943 ;
  assign n51096 = n7837 & ~n51095 ;
  assign n51097 = n51096 ^ n24421 ^ 1'b0 ;
  assign n51098 = ( n26593 & n51094 ) | ( n26593 & ~n51097 ) | ( n51094 & ~n51097 ) ;
  assign n51099 = n14404 & n51098 ;
  assign n51100 = n36811 ^ n22796 ^ n21299 ;
  assign n51101 = ~n39016 & n51100 ;
  assign n51102 = n51101 ^ n42806 ^ 1'b0 ;
  assign n51103 = n9197 | n26949 ;
  assign n51104 = n51103 ^ n19304 ^ 1'b0 ;
  assign n51105 = n20088 ^ n15941 ^ 1'b0 ;
  assign n51106 = n46689 ^ n7201 ^ 1'b0 ;
  assign n51107 = n51105 & n51106 ;
  assign n51108 = n13208 ^ n3474 ^ n2489 ;
  assign n51109 = n51108 ^ n40005 ^ n14273 ;
  assign n51110 = ~n15590 & n16896 ;
  assign n51111 = ~n14137 & n51110 ;
  assign n51112 = n29035 ^ n26187 ^ n1877 ;
  assign n51113 = n51112 ^ n44107 ^ n11216 ;
  assign n51114 = n33779 & n51113 ;
  assign n51115 = ~n18008 & n51114 ;
  assign n51116 = ~n51111 & n51115 ;
  assign n51117 = n11639 ^ n2522 ^ 1'b0 ;
  assign n51118 = n17234 & n29684 ;
  assign n51119 = n51118 ^ n3754 ^ 1'b0 ;
  assign n51120 = ( x239 & n13241 ) | ( x239 & n22992 ) | ( n13241 & n22992 ) ;
  assign n51121 = ( n10542 & n51119 ) | ( n10542 & n51120 ) | ( n51119 & n51120 ) ;
  assign n51122 = n31380 ^ n1840 ^ 1'b0 ;
  assign n51123 = n15056 | n51122 ;
  assign n51124 = n51123 ^ n36885 ^ 1'b0 ;
  assign n51125 = n51124 ^ n5059 ^ 1'b0 ;
  assign n51126 = n47744 | n51125 ;
  assign n51127 = n51126 ^ n47405 ^ n9037 ;
  assign n51128 = n28024 ^ n14758 ^ n13920 ;
  assign n51129 = n18770 & ~n27510 ;
  assign n51130 = n51129 ^ n10102 ^ 1'b0 ;
  assign n51131 = ~n1372 & n51130 ;
  assign n51132 = ~n51128 & n51131 ;
  assign n51133 = n27446 ^ x248 ^ 1'b0 ;
  assign n51134 = ~n4825 & n29961 ;
  assign n51135 = n51133 & n51134 ;
  assign n51136 = n51135 ^ n46770 ^ 1'b0 ;
  assign n51137 = n3718 | n51136 ;
  assign n51138 = n13071 | n43713 ;
  assign n51139 = n29652 & ~n51138 ;
  assign n51140 = n15790 ^ n3175 ^ n1524 ;
  assign n51141 = n51140 ^ n15414 ^ n11237 ;
  assign n51142 = n6267 & ~n11157 ;
  assign n51143 = n7902 ^ n3970 ^ 1'b0 ;
  assign n51144 = n51143 ^ n37734 ^ n34395 ;
  assign n51145 = n20974 ^ n8233 ^ 1'b0 ;
  assign n51147 = ( n2760 & n3430 ) | ( n2760 & ~n19822 ) | ( n3430 & ~n19822 ) ;
  assign n51146 = ~n20882 & n26107 ;
  assign n51148 = n51147 ^ n51146 ^ n33873 ;
  assign n51149 = n26630 ^ n24884 ^ 1'b0 ;
  assign n51150 = n5662 & n51149 ;
  assign n51151 = n2397 & ~n35888 ;
  assign n51152 = n31427 & n51151 ;
  assign n51153 = n13011 & n17057 ;
  assign n51154 = n21423 ^ n6176 ^ 1'b0 ;
  assign n51155 = n51153 | n51154 ;
  assign n51156 = n21030 & ~n51155 ;
  assign n51157 = n43303 ^ n23950 ^ 1'b0 ;
  assign n51158 = n51156 & ~n51157 ;
  assign n51159 = ~n18671 & n51158 ;
  assign n51160 = n51159 ^ n49102 ^ 1'b0 ;
  assign n51161 = n14517 & n25996 ;
  assign n51162 = n18720 & n51161 ;
  assign n51163 = ( n13107 & ~n42006 ) | ( n13107 & n45972 ) | ( ~n42006 & n45972 ) ;
  assign n51164 = n35005 ^ n1956 ^ 1'b0 ;
  assign n51165 = n51163 & ~n51164 ;
  assign n51166 = n51165 ^ n4434 ^ 1'b0 ;
  assign n51167 = ~n51162 & n51166 ;
  assign n51168 = n26212 ^ n14470 ^ 1'b0 ;
  assign n51169 = n3474 & ~n15424 ;
  assign n51170 = n6959 & n51169 ;
  assign n51171 = n36434 ^ n31228 ^ n14304 ;
  assign n51172 = ( n10141 & n22973 ) | ( n10141 & n51171 ) | ( n22973 & n51171 ) ;
  assign n51173 = n51172 ^ n33912 ^ n28315 ;
  assign n51174 = n51173 ^ n6805 ^ 1'b0 ;
  assign n51175 = n26895 ^ n9124 ^ n3062 ;
  assign n51176 = n25164 ^ n9703 ^ 1'b0 ;
  assign n51177 = n51175 | n51176 ;
  assign n51178 = n51177 ^ n28109 ^ 1'b0 ;
  assign n51179 = ( n7282 & n17060 ) | ( n7282 & ~n36442 ) | ( n17060 & ~n36442 ) ;
  assign n51181 = n11092 | n13316 ;
  assign n51182 = n23045 | n51181 ;
  assign n51183 = n51182 ^ n24080 ^ n17685 ;
  assign n51180 = n7142 | n44974 ;
  assign n51184 = n51183 ^ n51180 ^ 1'b0 ;
  assign n51185 = n5390 & ~n48407 ;
  assign n51186 = n51185 ^ n7621 ^ 1'b0 ;
  assign n51187 = n8619 ^ n5251 ^ 1'b0 ;
  assign n51188 = n43474 ^ n38057 ^ 1'b0 ;
  assign n51189 = ~n5292 & n15715 ;
  assign n51190 = n51189 ^ n15727 ^ 1'b0 ;
  assign n51191 = ( ~n8122 & n10349 ) | ( ~n8122 & n17042 ) | ( n10349 & n17042 ) ;
  assign n51192 = ~n3592 & n12280 ;
  assign n51193 = n7546 & n51192 ;
  assign n51194 = n16111 | n51193 ;
  assign n51195 = ( n13516 & n16510 ) | ( n13516 & ~n51194 ) | ( n16510 & ~n51194 ) ;
  assign n51196 = n18541 ^ n15068 ^ n14539 ;
  assign n51197 = n28247 & ~n51196 ;
  assign n51198 = n9339 | n31746 ;
  assign n51199 = n51198 ^ n25453 ^ 1'b0 ;
  assign n51200 = n11382 & ~n51199 ;
  assign n51201 = n51200 ^ n43703 ^ 1'b0 ;
  assign n51203 = n1353 ^ n441 ^ 1'b0 ;
  assign n51204 = ~n19832 & n51203 ;
  assign n51205 = n10496 & n51204 ;
  assign n51202 = n15392 & ~n25205 ;
  assign n51206 = n51205 ^ n51202 ^ 1'b0 ;
  assign n51207 = ~n13186 & n18320 ;
  assign n51208 = n51207 ^ n27623 ^ 1'b0 ;
  assign n51209 = n33756 ^ n25056 ^ 1'b0 ;
  assign n51210 = n6553 & ~n51209 ;
  assign n51211 = n47486 ^ n5271 ^ 1'b0 ;
  assign n51212 = ( n13460 & ~n21757 ) | ( n13460 & n39658 ) | ( ~n21757 & n39658 ) ;
  assign n51213 = ( n12045 & ~n13065 ) | ( n12045 & n49653 ) | ( ~n13065 & n49653 ) ;
  assign n51214 = n51213 ^ n44304 ^ n31972 ;
  assign n51215 = n16942 ^ n5158 ^ 1'b0 ;
  assign n51216 = n14483 | n51215 ;
  assign n51217 = n51216 ^ n1766 ^ 1'b0 ;
  assign n51218 = n51217 ^ n14099 ^ 1'b0 ;
  assign n51219 = ~n5912 & n39922 ;
  assign n51220 = n48410 ^ n47671 ^ 1'b0 ;
  assign n51221 = n19772 ^ n19421 ^ 1'b0 ;
  assign n51222 = n7966 & ~n51221 ;
  assign n51223 = n33683 & ~n39836 ;
  assign n51224 = n709 & n16665 ;
  assign n51225 = ~n16811 & n51224 ;
  assign n51226 = n51225 ^ n9727 ^ 1'b0 ;
  assign n51227 = n51223 | n51226 ;
  assign n51228 = ~n13848 & n25501 ;
  assign n51229 = n51228 ^ n5418 ^ 1'b0 ;
  assign n51230 = n23017 ^ n10857 ^ n7649 ;
  assign n51231 = n1607 & n3206 ;
  assign n51232 = n51230 & n51231 ;
  assign n51233 = n31089 & ~n51232 ;
  assign n51234 = n51233 ^ n4163 ^ 1'b0 ;
  assign n51235 = n36243 ^ n30494 ^ n30339 ;
  assign n51236 = n5030 | n45355 ;
  assign n51237 = n27903 & ~n51236 ;
  assign n51238 = n51237 ^ n22075 ^ 1'b0 ;
  assign n51239 = ( n14981 & ~n41050 ) | ( n14981 & n51238 ) | ( ~n41050 & n51238 ) ;
  assign n51240 = n24431 ^ n23561 ^ n3365 ;
  assign n51241 = n39317 ^ n4838 ^ n2077 ;
  assign n51242 = n9454 | n33883 ;
  assign n51243 = n9364 | n51242 ;
  assign n51244 = ( n16004 & n41672 ) | ( n16004 & ~n51243 ) | ( n41672 & ~n51243 ) ;
  assign n51245 = n20432 & n40061 ;
  assign n51246 = n30948 & n51245 ;
  assign n51247 = n49525 ^ x201 ^ 1'b0 ;
  assign n51248 = n50454 & n51247 ;
  assign n51249 = n9941 | n38107 ;
  assign n51250 = n48160 & ~n51249 ;
  assign n51251 = n27426 ^ n13062 ^ 1'b0 ;
  assign n51252 = n7520 | n21810 ;
  assign n51253 = ( n4848 & n19649 ) | ( n4848 & ~n51252 ) | ( n19649 & ~n51252 ) ;
  assign n51254 = ( ~n14618 & n28108 ) | ( ~n14618 & n46249 ) | ( n28108 & n46249 ) ;
  assign n51255 = n33656 ^ n7488 ^ 1'b0 ;
  assign n51256 = ~n33446 & n51255 ;
  assign n51257 = n51256 ^ n6782 ^ n6339 ;
  assign n51258 = n26927 & ~n43543 ;
  assign n51259 = n12343 & n51258 ;
  assign n51260 = n51259 ^ n25183 ^ n6574 ;
  assign n51261 = ( ~n6939 & n12996 ) | ( ~n6939 & n51260 ) | ( n12996 & n51260 ) ;
  assign n51262 = ~n1148 & n20343 ;
  assign n51263 = ~n29020 & n51262 ;
  assign n51264 = n51263 ^ n46511 ^ n26157 ;
  assign n51265 = n1709 | n46283 ;
  assign n51266 = n51265 ^ n10179 ^ 1'b0 ;
  assign n51267 = n7474 & ~n13522 ;
  assign n51268 = x142 & ~n9770 ;
  assign n51269 = ~n25695 & n51268 ;
  assign n51270 = ( n10176 & n51267 ) | ( n10176 & n51269 ) | ( n51267 & n51269 ) ;
  assign n51271 = n16401 | n51270 ;
  assign n51272 = n51271 ^ n33652 ^ 1'b0 ;
  assign n51273 = ~n34161 & n44398 ;
  assign n51274 = n23210 & n35715 ;
  assign n51275 = n13723 & n42977 ;
  assign n51276 = ( n16503 & n18770 ) | ( n16503 & n50675 ) | ( n18770 & n50675 ) ;
  assign n51277 = n35094 | n48049 ;
  assign n51278 = n51277 ^ n46165 ^ n6486 ;
  assign n51279 = n34544 ^ n14899 ^ 1'b0 ;
  assign n51280 = n5068 & n51279 ;
  assign n51281 = n17511 ^ n11961 ^ 1'b0 ;
  assign n51282 = ( ~n45224 & n51280 ) | ( ~n45224 & n51281 ) | ( n51280 & n51281 ) ;
  assign n51283 = n16935 ^ n6405 ^ 1'b0 ;
  assign n51284 = n51283 ^ n44117 ^ 1'b0 ;
  assign n51285 = n17350 ^ n6736 ^ 1'b0 ;
  assign n51286 = ( n10249 & n15340 ) | ( n10249 & n19195 ) | ( n15340 & n19195 ) ;
  assign n51287 = n51286 ^ n34715 ^ n9101 ;
  assign n51288 = n51285 & ~n51287 ;
  assign n51289 = n39593 ^ n23810 ^ 1'b0 ;
  assign n51290 = n50588 & ~n51289 ;
  assign n51291 = n436 & n7513 ;
  assign n51292 = ( n14259 & n16565 ) | ( n14259 & n26593 ) | ( n16565 & n26593 ) ;
  assign n51293 = n36525 & ~n39131 ;
  assign n51294 = n51292 & n51293 ;
  assign n51295 = n3659 & ~n9890 ;
  assign n51296 = n10030 & ~n25314 ;
  assign n51297 = n27647 & ~n42083 ;
  assign n51298 = n51297 ^ n14351 ^ 1'b0 ;
  assign n51299 = n51296 & n51298 ;
  assign n51300 = n44645 ^ n41164 ^ x204 ;
  assign n51301 = n50259 ^ n8335 ^ 1'b0 ;
  assign n51302 = n49286 & ~n50031 ;
  assign n51303 = n17737 & n51302 ;
  assign n51304 = n3042 | n34156 ;
  assign n51305 = n25592 ^ n14924 ^ n14786 ;
  assign n51306 = n4250 & n51305 ;
  assign n51307 = n3907 ^ n1280 ^ 1'b0 ;
  assign n51308 = n51306 & ~n51307 ;
  assign n51309 = n7838 & n45083 ;
  assign n51310 = n36184 ^ n2955 ^ 1'b0 ;
  assign n51311 = n34079 ^ n7615 ^ 1'b0 ;
  assign n51312 = n40935 ^ n18533 ^ 1'b0 ;
  assign n51313 = n12012 ^ n5301 ^ n4254 ;
  assign n51314 = n49924 ^ n39923 ^ 1'b0 ;
  assign n51315 = ~n9562 & n51314 ;
  assign n51316 = ( n51312 & n51313 ) | ( n51312 & n51315 ) | ( n51313 & n51315 ) ;
  assign n51317 = n31360 ^ n20595 ^ 1'b0 ;
  assign n51318 = n51316 & n51317 ;
  assign n51320 = ( ~n21179 & n32785 ) | ( ~n21179 & n50665 ) | ( n32785 & n50665 ) ;
  assign n51321 = n19290 | n51320 ;
  assign n51319 = ~n21327 & n38075 ;
  assign n51322 = n51321 ^ n51319 ^ 1'b0 ;
  assign n51324 = ~n8465 & n10714 ;
  assign n51325 = n4844 & n51324 ;
  assign n51326 = ( n9555 & n17647 ) | ( n9555 & ~n51325 ) | ( n17647 & ~n51325 ) ;
  assign n51323 = n7777 & n40052 ;
  assign n51327 = n51326 ^ n51323 ^ 1'b0 ;
  assign n51328 = n51327 ^ n13714 ^ 1'b0 ;
  assign n51329 = n51322 & ~n51328 ;
  assign n51330 = ( n1658 & n13871 ) | ( n1658 & n34154 ) | ( n13871 & n34154 ) ;
  assign n51331 = n40360 | n51330 ;
  assign n51332 = n51331 ^ n25652 ^ 1'b0 ;
  assign n51333 = ~n1943 & n51332 ;
  assign n51334 = n17880 & n51333 ;
  assign n51335 = n10740 & ~n46778 ;
  assign n51336 = n50429 & n51335 ;
  assign n51340 = n21586 & n36643 ;
  assign n51341 = n51340 ^ n12894 ^ 1'b0 ;
  assign n51337 = n27996 ^ n24303 ^ 1'b0 ;
  assign n51338 = ~n20055 & n51337 ;
  assign n51339 = ( ~n10152 & n43757 ) | ( ~n10152 & n51338 ) | ( n43757 & n51338 ) ;
  assign n51342 = n51341 ^ n51339 ^ n7597 ;
  assign n51343 = n29357 ^ n21560 ^ 1'b0 ;
  assign n51344 = n51343 ^ n5574 ^ n4298 ;
  assign n51345 = n46909 ^ n9302 ^ 1'b0 ;
  assign n51346 = n30818 ^ n2221 ^ 1'b0 ;
  assign n51347 = ~n31369 & n50590 ;
  assign n51348 = n51347 ^ n37390 ^ 1'b0 ;
  assign n51349 = ~n19781 & n44821 ;
  assign n51350 = n26405 & n51349 ;
  assign n51351 = n23691 ^ n17203 ^ 1'b0 ;
  assign n51352 = ~n51350 & n51351 ;
  assign n51353 = n15641 & ~n27811 ;
  assign n51354 = n51353 ^ n35255 ^ 1'b0 ;
  assign n51355 = n11193 & ~n11571 ;
  assign n51356 = n20486 & n51355 ;
  assign n51357 = n12270 ^ n7921 ^ 1'b0 ;
  assign n51358 = n9249 & ~n11992 ;
  assign n51359 = ~n20567 & n51358 ;
  assign n51360 = ( n23965 & ~n36151 ) | ( n23965 & n51359 ) | ( ~n36151 & n51359 ) ;
  assign n51361 = ( n22079 & n23963 ) | ( n22079 & ~n51360 ) | ( n23963 & ~n51360 ) ;
  assign n51362 = ( n25125 & n51357 ) | ( n25125 & ~n51361 ) | ( n51357 & ~n51361 ) ;
  assign n51363 = ( n5492 & n11193 ) | ( n5492 & ~n14482 ) | ( n11193 & ~n14482 ) ;
  assign n51364 = n50471 ^ n39979 ^ n14683 ;
  assign n51365 = n1421 | n21335 ;
  assign n51366 = n713 | n5954 ;
  assign n51367 = n6035 & ~n51366 ;
  assign n51368 = n834 & n51367 ;
  assign n51369 = n9151 | n18505 ;
  assign n51370 = n50023 & ~n51369 ;
  assign n51371 = n8785 & ~n10430 ;
  assign n51372 = n51371 ^ n5709 ^ 1'b0 ;
  assign n51373 = n51372 ^ n16112 ^ 1'b0 ;
  assign n51374 = n2001 | n39485 ;
  assign n51375 = ( n6996 & n32107 ) | ( n6996 & n33505 ) | ( n32107 & n33505 ) ;
  assign n51376 = n51375 ^ n24139 ^ n9765 ;
  assign n51377 = n4480 | n19435 ;
  assign n51378 = n1771 & ~n51377 ;
  assign n51379 = n23887 | n51378 ;
  assign n51380 = n51379 ^ n26708 ^ n2860 ;
  assign n51381 = n15621 & ~n25056 ;
  assign n51382 = ~n45322 & n51381 ;
  assign n51383 = n4109 ^ n3231 ^ 1'b0 ;
  assign n51384 = n29835 | n51383 ;
  assign n51385 = n51384 ^ n48266 ^ 1'b0 ;
  assign n51386 = ~n12790 & n51385 ;
  assign n51387 = n14922 | n15727 ;
  assign n51388 = n25639 | n51387 ;
  assign n51389 = n45556 ^ n15731 ^ n3465 ;
  assign n51390 = n13984 & n18242 ;
  assign n51391 = ~n51389 & n51390 ;
  assign n51392 = n11387 | n39541 ;
  assign n51393 = n17823 ^ n10998 ^ 1'b0 ;
  assign n51394 = n6721 & n51393 ;
  assign n51395 = ~n3136 & n51394 ;
  assign n51396 = n51392 & n51395 ;
  assign n51397 = n13227 ^ n7869 ^ n2623 ;
  assign n51398 = n14897 & n51397 ;
  assign n51399 = n51398 ^ n18721 ^ n7013 ;
  assign n51400 = n18165 ^ n5494 ^ n3920 ;
  assign n51401 = n51400 ^ n44247 ^ 1'b0 ;
  assign n51402 = ( ~n13927 & n51399 ) | ( ~n13927 & n51401 ) | ( n51399 & n51401 ) ;
  assign n51403 = n48439 ^ n31188 ^ 1'b0 ;
  assign n51404 = ~n14924 & n35778 ;
  assign n51405 = n51203 ^ n3235 ^ 1'b0 ;
  assign n51406 = n6173 | n51405 ;
  assign n51407 = n2899 | n17424 ;
  assign n51408 = n51407 ^ n11197 ^ 1'b0 ;
  assign n51409 = ( n4150 & ~n5388 ) | ( n4150 & n51408 ) | ( ~n5388 & n51408 ) ;
  assign n51410 = n2108 & ~n2412 ;
  assign n51411 = n23434 & n26466 ;
  assign n51412 = n27104 & n51411 ;
  assign n51413 = n51412 ^ n21222 ^ 1'b0 ;
  assign n51414 = n48312 ^ n24080 ^ 1'b0 ;
  assign n51415 = ( n3830 & ~n17994 ) | ( n3830 & n46341 ) | ( ~n17994 & n46341 ) ;
  assign n51416 = n51415 ^ n24968 ^ 1'b0 ;
  assign n51417 = n25541 | n42731 ;
  assign n51418 = ( n22634 & n48129 ) | ( n22634 & n51417 ) | ( n48129 & n51417 ) ;
  assign n51419 = n45621 & n48497 ;
  assign n51420 = n12805 ^ n9673 ^ 1'b0 ;
  assign n51421 = ( n35361 & n51419 ) | ( n35361 & n51420 ) | ( n51419 & n51420 ) ;
  assign n51422 = n31383 ^ n13273 ^ 1'b0 ;
  assign n51423 = ~n5193 & n51422 ;
  assign n51424 = n18104 & n51423 ;
  assign n51425 = n51424 ^ n26661 ^ 1'b0 ;
  assign n51426 = x155 & n25598 ;
  assign n51427 = ~n51425 & n51426 ;
  assign n51428 = n40163 | n45449 ;
  assign n51429 = n20731 | n51428 ;
  assign n51430 = n35630 ^ n5678 ^ 1'b0 ;
  assign n51431 = n39097 ^ n35475 ^ n17929 ;
  assign n51432 = n30346 ^ n26344 ^ n5371 ;
  assign n51433 = n51432 ^ n25060 ^ 1'b0 ;
  assign n51434 = ( n12800 & ~n13804 ) | ( n12800 & n15816 ) | ( ~n13804 & n15816 ) ;
  assign n51435 = n51434 ^ n47351 ^ n19815 ;
  assign n51436 = ( n4307 & n8429 ) | ( n4307 & n26888 ) | ( n8429 & n26888 ) ;
  assign n51437 = n51436 ^ n46761 ^ n23318 ;
  assign n51438 = n51437 ^ n15189 ^ n13686 ;
  assign n51439 = n35063 ^ n23167 ^ 1'b0 ;
  assign n51440 = n19098 & n51439 ;
  assign n51441 = ~n30704 & n38572 ;
  assign n51442 = n51441 ^ n18243 ^ 1'b0 ;
  assign n51447 = ~n28255 & n50281 ;
  assign n51443 = x219 | n4820 ;
  assign n51444 = n534 & ~n51443 ;
  assign n51445 = n17188 & n51444 ;
  assign n51446 = n51445 ^ n10265 ^ n5126 ;
  assign n51448 = n51447 ^ n51446 ^ n5813 ;
  assign n51449 = n24778 ^ n2545 ^ 1'b0 ;
  assign n51450 = n51449 ^ n33088 ^ 1'b0 ;
  assign n51451 = ( n362 & n4823 ) | ( n362 & ~n8710 ) | ( n4823 & ~n8710 ) ;
  assign n51452 = ( n4970 & n40951 ) | ( n4970 & n51451 ) | ( n40951 & n51451 ) ;
  assign n51453 = ~n4015 & n9927 ;
  assign n51454 = n2229 & ~n7141 ;
  assign n51455 = ( n12573 & n51453 ) | ( n12573 & n51454 ) | ( n51453 & n51454 ) ;
  assign n51456 = ( n5898 & n36517 ) | ( n5898 & ~n51455 ) | ( n36517 & ~n51455 ) ;
  assign n51457 = n8051 ^ n4283 ^ 1'b0 ;
  assign n51458 = n16915 & ~n51457 ;
  assign n51459 = n51458 ^ n8187 ^ 1'b0 ;
  assign n51468 = n30900 ^ n26219 ^ n18226 ;
  assign n51460 = n37361 ^ n4801 ^ 1'b0 ;
  assign n51461 = ~n15413 & n51460 ;
  assign n51462 = n51461 ^ n27295 ^ 1'b0 ;
  assign n51463 = n30235 & n51462 ;
  assign n51464 = ( n14258 & n42661 ) | ( n14258 & ~n51463 ) | ( n42661 & ~n51463 ) ;
  assign n51465 = n51464 ^ n10928 ^ n3591 ;
  assign n51466 = n19627 ^ n1311 ^ 1'b0 ;
  assign n51467 = n51465 & n51466 ;
  assign n51469 = n51468 ^ n51467 ^ 1'b0 ;
  assign n51470 = n46583 ^ n2179 ^ 1'b0 ;
  assign n51471 = ( n51459 & n51469 ) | ( n51459 & ~n51470 ) | ( n51469 & ~n51470 ) ;
  assign n51472 = ~n18242 & n37786 ;
  assign n51473 = n26390 ^ n22968 ^ 1'b0 ;
  assign n51474 = n9878 & ~n21570 ;
  assign n51475 = ( n14660 & n26952 ) | ( n14660 & ~n39117 ) | ( n26952 & ~n39117 ) ;
  assign n51476 = n8514 | n51475 ;
  assign n51477 = n4714 & ~n11850 ;
  assign n51478 = n51477 ^ n2847 ^ 1'b0 ;
  assign n51479 = ( n14804 & ~n45501 ) | ( n14804 & n51478 ) | ( ~n45501 & n51478 ) ;
  assign n51480 = ( n13924 & n24089 ) | ( n13924 & ~n41232 ) | ( n24089 & ~n41232 ) ;
  assign n51481 = n49564 ^ n34829 ^ 1'b0 ;
  assign n51487 = n12612 ^ n2867 ^ 1'b0 ;
  assign n51488 = ~n25262 & n51487 ;
  assign n51482 = n4049 & n25189 ;
  assign n51483 = n51482 ^ n11239 ^ 1'b0 ;
  assign n51484 = n32453 ^ n1843 ^ 1'b0 ;
  assign n51485 = ~n51483 & n51484 ;
  assign n51486 = n8680 & n51485 ;
  assign n51489 = n51488 ^ n51486 ^ 1'b0 ;
  assign n51490 = n7042 | n10776 ;
  assign n51491 = n26877 & ~n51490 ;
  assign n51492 = n17414 ^ n7644 ^ 1'b0 ;
  assign n51493 = n38216 ^ n29241 ^ 1'b0 ;
  assign n51494 = ~n8523 & n19630 ;
  assign n51495 = n51494 ^ n49145 ^ 1'b0 ;
  assign n51496 = n32873 ^ n17466 ^ n13190 ;
  assign n51497 = n16707 & n51496 ;
  assign n51498 = n41537 & n51497 ;
  assign n51499 = n14849 ^ n9881 ^ 1'b0 ;
  assign n51500 = ( n15588 & n48779 ) | ( n15588 & ~n51499 ) | ( n48779 & ~n51499 ) ;
  assign n51501 = n51500 ^ n47386 ^ 1'b0 ;
  assign n51502 = ( n5916 & ~n25010 ) | ( n5916 & n51501 ) | ( ~n25010 & n51501 ) ;
  assign n51503 = n25169 ^ n14273 ^ 1'b0 ;
  assign n51504 = n32051 ^ n27373 ^ 1'b0 ;
  assign n51505 = n48092 ^ n28558 ^ 1'b0 ;
  assign n51506 = n39043 ^ n35946 ^ n19233 ;
  assign n51507 = n22332 ^ n17962 ^ n17257 ;
  assign n51508 = ( n16114 & ~n51506 ) | ( n16114 & n51507 ) | ( ~n51506 & n51507 ) ;
  assign n51510 = n17225 ^ n500 ^ 1'b0 ;
  assign n51509 = n31114 ^ n29190 ^ n15415 ;
  assign n51511 = n51510 ^ n51509 ^ n6164 ;
  assign n51512 = ( n8995 & n18543 ) | ( n8995 & n23115 ) | ( n18543 & n23115 ) ;
  assign n51513 = n2143 & ~n51512 ;
  assign n51514 = n22205 ^ n12531 ^ 1'b0 ;
  assign n51515 = n51514 ^ n41637 ^ n5768 ;
  assign n51516 = n43853 ^ n24880 ^ n23276 ;
  assign n51517 = ( ~n1250 & n13859 ) | ( ~n1250 & n48348 ) | ( n13859 & n48348 ) ;
  assign n51518 = n42051 ^ n41398 ^ n15175 ;
  assign n51519 = n400 & ~n15094 ;
  assign n51520 = n50622 ^ n19577 ^ n14614 ;
  assign n51521 = ( n18157 & n51519 ) | ( n18157 & n51520 ) | ( n51519 & n51520 ) ;
  assign n51522 = ( ~n4669 & n20465 ) | ( ~n4669 & n34702 ) | ( n20465 & n34702 ) ;
  assign n51523 = n51522 ^ n2967 ^ 1'b0 ;
  assign n51524 = n6856 | n51523 ;
  assign n51525 = n22144 & n24336 ;
  assign n51526 = ~n3002 & n51525 ;
  assign n51527 = x80 & ~n30960 ;
  assign n51528 = n51526 & n51527 ;
  assign n51529 = n45442 ^ n24857 ^ 1'b0 ;
  assign n51530 = ~n1346 & n3945 ;
  assign n51531 = ~n4516 & n51530 ;
  assign n51532 = ~n10806 & n43785 ;
  assign n51533 = n51532 ^ n33645 ^ 1'b0 ;
  assign n51534 = ( n6433 & n25184 ) | ( n6433 & ~n27118 ) | ( n25184 & ~n27118 ) ;
  assign n51535 = n19349 & n51534 ;
  assign n51536 = n51535 ^ n20940 ^ 1'b0 ;
  assign n51537 = n27948 & ~n51536 ;
  assign n51538 = ( n9299 & n9961 ) | ( n9299 & ~n10169 ) | ( n9961 & ~n10169 ) ;
  assign n51539 = ( n6014 & ~n24473 ) | ( n6014 & n51538 ) | ( ~n24473 & n51538 ) ;
  assign n51540 = n4190 ^ n3095 ^ n1607 ;
  assign n51541 = n3632 | n51540 ;
  assign n51542 = n9662 | n32763 ;
  assign n51543 = n19012 & ~n51542 ;
  assign n51544 = n51543 ^ n18772 ^ 1'b0 ;
  assign n51545 = n3563 | n11283 ;
  assign n51546 = n51545 ^ n14654 ^ 1'b0 ;
  assign n51547 = ( ~n18162 & n41626 ) | ( ~n18162 & n51546 ) | ( n41626 & n51546 ) ;
  assign n51548 = n13257 ^ n7217 ^ n989 ;
  assign n51549 = ~n2063 & n51548 ;
  assign n51550 = ~n38135 & n51549 ;
  assign n51551 = n7007 | n8630 ;
  assign n51552 = n24923 & ~n51551 ;
  assign n51553 = n25776 | n51552 ;
  assign n51554 = n36577 | n51553 ;
  assign n51555 = ~n7254 & n43298 ;
  assign n51556 = n51555 ^ n34839 ^ 1'b0 ;
  assign n51557 = n1325 & ~n51556 ;
  assign n51558 = n34945 | n38301 ;
  assign n51559 = n51558 ^ n9642 ^ 1'b0 ;
  assign n51564 = n22989 & ~n45673 ;
  assign n51562 = n24399 ^ n5461 ^ 1'b0 ;
  assign n51560 = n693 | n36623 ;
  assign n51561 = n6027 & ~n51560 ;
  assign n51563 = n51562 ^ n51561 ^ n39773 ;
  assign n51565 = n51564 ^ n51563 ^ n6854 ;
  assign n51566 = n3136 | n5193 ;
  assign n51567 = n5193 & ~n51566 ;
  assign n51568 = n25858 & n51567 ;
  assign n51569 = n25452 & n29956 ;
  assign n51570 = ~n25452 & n51569 ;
  assign n51571 = n51568 | n51570 ;
  assign n51572 = n51571 ^ n1030 ^ x72 ;
  assign n51573 = ( n12572 & n34339 ) | ( n12572 & n51572 ) | ( n34339 & n51572 ) ;
  assign n51574 = n51573 ^ n13804 ^ n4470 ;
  assign n51575 = n15153 ^ n13870 ^ 1'b0 ;
  assign n51576 = n9841 & ~n51575 ;
  assign n51577 = ( ~n8751 & n31539 ) | ( ~n8751 & n45490 ) | ( n31539 & n45490 ) ;
  assign n51578 = n51577 ^ n45100 ^ n17606 ;
  assign n51579 = n26645 ^ n22926 ^ 1'b0 ;
  assign n51580 = n9394 & n33199 ;
  assign n51581 = n40617 ^ n37081 ^ 1'b0 ;
  assign n51582 = n4034 & ~n51581 ;
  assign n51583 = n35754 | n42769 ;
  assign n51584 = n15337 | n51583 ;
  assign n51588 = n277 & ~n1989 ;
  assign n51586 = n14657 & ~n15071 ;
  assign n51587 = ~n15214 & n51586 ;
  assign n51589 = n51588 ^ n51587 ^ n40132 ;
  assign n51585 = n10388 & n13738 ;
  assign n51590 = n51589 ^ n51585 ^ 1'b0 ;
  assign n51591 = n27679 ^ n19560 ^ n10315 ;
  assign n51593 = n17154 ^ n16568 ^ n1524 ;
  assign n51592 = n5253 & ~n10403 ;
  assign n51594 = n51593 ^ n51592 ^ 1'b0 ;
  assign n51595 = n51594 ^ n37464 ^ n30150 ;
  assign n51596 = n46677 ^ n9917 ^ 1'b0 ;
  assign n51597 = ~n20794 & n37763 ;
  assign n51598 = n43770 ^ n35294 ^ 1'b0 ;
  assign n51599 = n28314 | n45014 ;
  assign n51600 = n1390 & ~n51599 ;
  assign n51601 = n25476 | n38197 ;
  assign n51602 = n32816 & ~n51601 ;
  assign n51603 = n40690 & ~n51602 ;
  assign n51604 = ( n4705 & n11319 ) | ( n4705 & n17544 ) | ( n11319 & n17544 ) ;
  assign n51605 = n51604 ^ n40689 ^ 1'b0 ;
  assign n51606 = n29165 ^ n11487 ^ n3569 ;
  assign n51607 = n20351 & n51606 ;
  assign n51608 = ( n11650 & n26012 ) | ( n11650 & ~n37137 ) | ( n26012 & ~n37137 ) ;
  assign n51609 = ~n8541 & n28813 ;
  assign n51610 = ~n23105 & n51609 ;
  assign n51611 = ( n584 & n10660 ) | ( n584 & n51610 ) | ( n10660 & n51610 ) ;
  assign n51612 = ( n39660 & n51608 ) | ( n39660 & n51611 ) | ( n51608 & n51611 ) ;
  assign n51613 = n7104 & ~n11029 ;
  assign n51614 = n50141 | n51613 ;
  assign n51616 = n33541 ^ n9041 ^ n4272 ;
  assign n51617 = ( n13264 & n39169 ) | ( n13264 & n51616 ) | ( n39169 & n51616 ) ;
  assign n51615 = n9191 & ~n10074 ;
  assign n51618 = n51617 ^ n51615 ^ n25156 ;
  assign n51619 = ( n7215 & ~n9093 ) | ( n7215 & n38368 ) | ( ~n9093 & n38368 ) ;
  assign n51620 = x71 & ~n11817 ;
  assign n51621 = n51620 ^ n45187 ^ 1'b0 ;
  assign n51622 = n12795 | n23589 ;
  assign n51623 = n36141 & n51622 ;
  assign n51624 = n51623 ^ n46781 ^ 1'b0 ;
  assign n51626 = n20423 ^ n16488 ^ 1'b0 ;
  assign n51627 = n51626 ^ n28695 ^ n23475 ;
  assign n51625 = n3328 | n30651 ;
  assign n51628 = n51627 ^ n51625 ^ 1'b0 ;
  assign n51629 = n13327 ^ n12071 ^ n1934 ;
  assign n51630 = ~n5517 & n51629 ;
  assign n51631 = n51630 ^ x36 ^ 1'b0 ;
  assign n51632 = n6329 & ~n14956 ;
  assign n51633 = n9605 & ~n40672 ;
  assign n51634 = n29669 & ~n50640 ;
  assign n51635 = n33924 ^ n7516 ^ 1'b0 ;
  assign n51636 = n36430 ^ n32987 ^ n15262 ;
  assign n51637 = ( n36728 & n38644 ) | ( n36728 & n50814 ) | ( n38644 & n50814 ) ;
  assign n51638 = n21770 ^ n12449 ^ n6306 ;
  assign n51639 = n3358 ^ n1036 ^ n773 ;
  assign n51640 = n51639 ^ n12595 ^ n2944 ;
  assign n51641 = n26016 & ~n51640 ;
  assign n51642 = n23301 & n51641 ;
  assign n51645 = n18078 ^ n13969 ^ n355 ;
  assign n51646 = n2194 & n51645 ;
  assign n51643 = ( ~n13697 & n40202 ) | ( ~n13697 & n45676 ) | ( n40202 & n45676 ) ;
  assign n51644 = n51643 ^ n16995 ^ n6090 ;
  assign n51647 = n51646 ^ n51644 ^ n14470 ;
  assign n51648 = n36205 ^ n6621 ^ n5116 ;
  assign n51649 = ( n16031 & ~n17404 ) | ( n16031 & n37571 ) | ( ~n17404 & n37571 ) ;
  assign n51650 = n45297 & ~n51649 ;
  assign n51651 = n30883 & n38556 ;
  assign n51652 = n7094 | n43315 ;
  assign n51653 = ~n33730 & n35107 ;
  assign n51654 = n51653 ^ n49253 ^ 1'b0 ;
  assign n51655 = ~n7234 & n28464 ;
  assign n51656 = n51655 ^ n7711 ^ 1'b0 ;
  assign n51657 = n269 & n12046 ;
  assign n51658 = n24819 & n51657 ;
  assign n51659 = n36285 ^ n13665 ^ 1'b0 ;
  assign n51660 = n3420 | n51659 ;
  assign n51661 = n29252 ^ n9782 ^ 1'b0 ;
  assign n51662 = n16945 ^ n2490 ^ n1232 ;
  assign n51663 = n8117 ^ n3315 ^ 1'b0 ;
  assign n51664 = n18462 & n51663 ;
  assign n51665 = ( ~n15713 & n51662 ) | ( ~n15713 & n51664 ) | ( n51662 & n51664 ) ;
  assign n51666 = ( n3647 & n51661 ) | ( n3647 & ~n51665 ) | ( n51661 & ~n51665 ) ;
  assign n51669 = n19580 ^ n10245 ^ 1'b0 ;
  assign n51667 = x142 & ~n11838 ;
  assign n51668 = ~n37937 & n51667 ;
  assign n51670 = n51669 ^ n51668 ^ 1'b0 ;
  assign n51671 = n22695 ^ n16273 ^ 1'b0 ;
  assign n51672 = n35441 ^ n27023 ^ n26308 ;
  assign n51674 = n11894 & n23329 ;
  assign n51675 = ~n34777 & n51674 ;
  assign n51673 = n18067 | n34467 ;
  assign n51676 = n51675 ^ n51673 ^ 1'b0 ;
  assign n51677 = n33518 ^ n4382 ^ 1'b0 ;
  assign n51678 = ~n51676 & n51677 ;
  assign n51679 = n37567 | n46588 ;
  assign n51683 = ( ~n9843 & n15820 ) | ( ~n9843 & n23857 ) | ( n15820 & n23857 ) ;
  assign n51680 = n27832 ^ n17062 ^ n14403 ;
  assign n51681 = n27185 | n51680 ;
  assign n51682 = n21598 & ~n51681 ;
  assign n51684 = n51683 ^ n51682 ^ 1'b0 ;
  assign n51685 = n13129 & n24138 ;
  assign n51686 = n9624 & ~n13339 ;
  assign n51687 = n756 & ~n3520 ;
  assign n51688 = n51687 ^ n14281 ^ n2134 ;
  assign n51689 = n44272 ^ n21759 ^ n4461 ;
  assign n51690 = ( n26198 & n33490 ) | ( n26198 & ~n39268 ) | ( n33490 & ~n39268 ) ;
  assign n51691 = n12919 | n29130 ;
  assign n51692 = n51691 ^ n34112 ^ n14320 ;
  assign n51693 = n22473 & ~n26032 ;
  assign n51694 = ~n22928 & n51693 ;
  assign n51695 = n24495 & ~n51694 ;
  assign n51696 = n51695 ^ n15781 ^ 1'b0 ;
  assign n51697 = ( n2489 & n31456 ) | ( n2489 & ~n35560 ) | ( n31456 & ~n35560 ) ;
  assign n51698 = n51697 ^ n7119 ^ 1'b0 ;
  assign n51699 = n45632 ^ n24560 ^ n14436 ;
  assign n51700 = ~n9297 & n40555 ;
  assign n51701 = ( n22395 & ~n50564 ) | ( n22395 & n51700 ) | ( ~n50564 & n51700 ) ;
  assign n51702 = n42731 ^ n31881 ^ n5324 ;
  assign n51703 = ( n1538 & n3725 ) | ( n1538 & n40906 ) | ( n3725 & n40906 ) ;
  assign n51704 = n51703 ^ n43483 ^ x107 ;
  assign n51705 = n4765 & ~n18620 ;
  assign n51706 = n11264 | n29042 ;
  assign n51707 = n24507 & ~n51706 ;
  assign n51708 = n34097 ^ n25262 ^ n2036 ;
  assign n51709 = n51708 ^ n21684 ^ 1'b0 ;
  assign n51710 = n35244 & n51709 ;
  assign n51711 = n36122 ^ n26308 ^ 1'b0 ;
  assign n51712 = x47 & ~n51711 ;
  assign n51713 = ( n9930 & n18847 ) | ( n9930 & n51712 ) | ( n18847 & n51712 ) ;
  assign n51714 = n12748 & ~n37039 ;
  assign n51715 = ( ~n704 & n38596 ) | ( ~n704 & n41030 ) | ( n38596 & n41030 ) ;
  assign n51716 = ( n1782 & n6718 ) | ( n1782 & ~n29163 ) | ( n6718 & ~n29163 ) ;
  assign n51717 = n12396 ^ n8786 ^ n7048 ;
  assign n51718 = ( n24748 & ~n32705 ) | ( n24748 & n51717 ) | ( ~n32705 & n51717 ) ;
  assign n51719 = ( n11242 & ~n51716 ) | ( n11242 & n51718 ) | ( ~n51716 & n51718 ) ;
  assign n51720 = n9442 & ~n32575 ;
  assign n51721 = ~n1447 & n51720 ;
  assign n51722 = n8332 | n35906 ;
  assign n51723 = n51722 ^ n8292 ^ 1'b0 ;
  assign n51724 = n25917 ^ n12212 ^ 1'b0 ;
  assign n51725 = n34376 & n51724 ;
  assign n51726 = n17763 ^ n9512 ^ 1'b0 ;
  assign n51727 = n17848 & ~n51726 ;
  assign n51728 = n40404 ^ n9424 ^ 1'b0 ;
  assign n51729 = n51727 & ~n51728 ;
  assign n51730 = n290 & n7571 ;
  assign n51731 = n51730 ^ n1403 ^ 1'b0 ;
  assign n51732 = n12526 ^ n2750 ^ n737 ;
  assign n51733 = n51732 ^ n36105 ^ 1'b0 ;
  assign n51734 = n51731 & n51733 ;
  assign n51735 = n5188 & n8713 ;
  assign n51736 = n51735 ^ n12590 ^ 1'b0 ;
  assign n51737 = ( ~n791 & n3490 ) | ( ~n791 & n9910 ) | ( n3490 & n9910 ) ;
  assign n51738 = n32828 ^ n22912 ^ 1'b0 ;
  assign n51739 = n51737 & n51738 ;
  assign n51740 = n51739 ^ n49689 ^ n15152 ;
  assign n51741 = n42568 ^ n21432 ^ n18933 ;
  assign n51742 = n13985 ^ n12433 ^ n4537 ;
  assign n51743 = n1118 ^ n553 ^ 1'b0 ;
  assign n51744 = n5720 & n51743 ;
  assign n51745 = ~n51742 & n51744 ;
  assign n51746 = n51745 ^ n15003 ^ 1'b0 ;
  assign n51747 = n24803 ^ n13776 ^ 1'b0 ;
  assign n51748 = n29746 & ~n51747 ;
  assign n51749 = n51748 ^ n28816 ^ 1'b0 ;
  assign n51750 = n26120 ^ n10189 ^ n8196 ;
  assign n51751 = ( n4766 & n11781 ) | ( n4766 & n51750 ) | ( n11781 & n51750 ) ;
  assign n51752 = n51751 ^ n6100 ^ 1'b0 ;
  assign n51753 = ( n26227 & n51749 ) | ( n26227 & n51752 ) | ( n51749 & n51752 ) ;
  assign n51754 = n6367 & n25642 ;
  assign n51755 = n51754 ^ n33724 ^ 1'b0 ;
  assign n51756 = n51755 ^ n9033 ^ n5488 ;
  assign n51757 = n14972 ^ n4865 ^ 1'b0 ;
  assign n51758 = n9271 & ~n51757 ;
  assign n51759 = n32529 & ~n51680 ;
  assign n51760 = n5052 & ~n51759 ;
  assign n51761 = n24598 & ~n51760 ;
  assign n51762 = n51761 ^ n15722 ^ 1'b0 ;
  assign n51763 = n50814 ^ n15703 ^ 1'b0 ;
  assign n51764 = n31980 & n51763 ;
  assign n51765 = ( ~n1372 & n2631 ) | ( ~n1372 & n16363 ) | ( n2631 & n16363 ) ;
  assign n51766 = n51765 ^ n30921 ^ 1'b0 ;
  assign n51767 = n51680 | n51766 ;
  assign n51768 = n35097 ^ n24431 ^ 1'b0 ;
  assign n51769 = ( n3268 & n21900 ) | ( n3268 & ~n34502 ) | ( n21900 & ~n34502 ) ;
  assign n51770 = n40707 & ~n40900 ;
  assign n51771 = ~n51769 & n51770 ;
  assign n51772 = ( ~n18533 & n23898 ) | ( ~n18533 & n26603 ) | ( n23898 & n26603 ) ;
  assign n51773 = ( n28358 & n51675 ) | ( n28358 & n51772 ) | ( n51675 & n51772 ) ;
  assign n51774 = n468 & ~n6404 ;
  assign n51775 = ~n9999 & n14459 ;
  assign n51776 = n3709 & n51775 ;
  assign n51777 = n2485 & n22352 ;
  assign n51778 = n51777 ^ n11794 ^ 1'b0 ;
  assign n51779 = n5490 & n51778 ;
  assign n51780 = n51776 & n51779 ;
  assign n51784 = ~x230 & n34307 ;
  assign n51785 = n51784 ^ n4754 ^ 1'b0 ;
  assign n51786 = n5431 & ~n19355 ;
  assign n51787 = n51786 ^ n21028 ^ 1'b0 ;
  assign n51788 = n51785 | n51787 ;
  assign n51781 = n3026 & n9920 ;
  assign n51782 = ~n1739 & n51781 ;
  assign n51783 = n12936 | n51782 ;
  assign n51789 = n51788 ^ n51783 ^ 1'b0 ;
  assign n51790 = n46125 | n46377 ;
  assign n51791 = n19106 | n51790 ;
  assign n51792 = n40380 ^ n6798 ^ n2945 ;
  assign n51793 = ~n44353 & n51792 ;
  assign n51794 = n3205 & ~n6952 ;
  assign n51795 = n23092 & n51794 ;
  assign n51796 = ~n13704 & n39415 ;
  assign n51797 = ~n25784 & n51796 ;
  assign n51798 = ( n30179 & ~n34146 ) | ( n30179 & n51797 ) | ( ~n34146 & n51797 ) ;
  assign n51799 = ( n3970 & n15350 ) | ( n3970 & ~n43347 ) | ( n15350 & ~n43347 ) ;
  assign n51800 = n19665 & n33187 ;
  assign n51801 = ~n40065 & n51800 ;
  assign n51802 = n51801 ^ n40486 ^ n25339 ;
  assign n51803 = n6907 | n41915 ;
  assign n51804 = n35470 & ~n51803 ;
  assign n51805 = n51804 ^ n31178 ^ n30411 ;
  assign n51806 = n50965 ^ n44836 ^ n3258 ;
  assign n51807 = n51806 ^ n36582 ^ n585 ;
  assign n51808 = n21990 & n42860 ;
  assign n51809 = n51808 ^ n23960 ^ 1'b0 ;
  assign n51810 = n3786 & n12281 ;
  assign n51811 = n49930 & n51810 ;
  assign n51812 = n16486 | n17160 ;
  assign n51813 = n18978 & ~n51812 ;
  assign n51814 = n4832 & n25549 ;
  assign n51815 = n51814 ^ n29510 ^ n14898 ;
  assign n51816 = n1483 & n51815 ;
  assign n51817 = n51816 ^ n29320 ^ 1'b0 ;
  assign n51818 = n6640 & ~n19626 ;
  assign n51819 = n51818 ^ n32910 ^ 1'b0 ;
  assign n51820 = n4206 ^ n3056 ^ 1'b0 ;
  assign n51821 = n1568 & n51820 ;
  assign n51822 = n7743 & n51821 ;
  assign n51823 = n51822 ^ n4446 ^ 1'b0 ;
  assign n51824 = n9868 & ~n51823 ;
  assign n51825 = n4237 ^ n2049 ^ 1'b0 ;
  assign n51826 = n25995 & ~n51825 ;
  assign n51827 = ( n11298 & n27803 ) | ( n11298 & n51826 ) | ( n27803 & n51826 ) ;
  assign n51828 = n31923 ^ n10804 ^ n8885 ;
  assign n51829 = ( ~x111 & x128 ) | ( ~x111 & n51828 ) | ( x128 & n51828 ) ;
  assign n51831 = ( n3888 & n8457 ) | ( n3888 & n51434 ) | ( n8457 & n51434 ) ;
  assign n51830 = n1874 | n47798 ;
  assign n51832 = n51831 ^ n51830 ^ n51512 ;
  assign n51833 = n17721 ^ n10680 ^ 1'b0 ;
  assign n51834 = n3951 & ~n13958 ;
  assign n51835 = n50795 ^ n4250 ^ 1'b0 ;
  assign n51836 = n35997 & n51835 ;
  assign n51837 = n2408 & n14706 ;
  assign n51838 = n51837 ^ n3105 ^ 1'b0 ;
  assign n51839 = n47860 ^ n25100 ^ n12470 ;
  assign n51840 = n21116 ^ n20269 ^ n543 ;
  assign n51841 = n51840 ^ n30485 ^ n7621 ;
  assign n51842 = ~n3375 & n12270 ;
  assign n51843 = n51842 ^ n37923 ^ n3525 ;
  assign n51844 = ( n4548 & ~n23510 ) | ( n4548 & n32575 ) | ( ~n23510 & n32575 ) ;
  assign n51845 = ( n21778 & n45164 ) | ( n21778 & ~n51844 ) | ( n45164 & ~n51844 ) ;
  assign n51846 = n19071 & ~n40094 ;
  assign n51847 = n1088 & n8278 ;
  assign n51848 = n18010 & n51847 ;
  assign n51849 = n38564 ^ n17739 ^ 1'b0 ;
  assign n51850 = ~n18484 & n51849 ;
  assign n51851 = n23295 ^ n14079 ^ 1'b0 ;
  assign n51852 = n31928 | n45872 ;
  assign n51853 = n51851 & ~n51852 ;
  assign n51854 = n1340 | n6438 ;
  assign n51855 = n10820 & ~n51854 ;
  assign n51856 = n37300 ^ n7782 ^ 1'b0 ;
  assign n51857 = n14298 | n24802 ;
  assign n51858 = n51857 ^ n14813 ^ 1'b0 ;
  assign n51859 = n5541 & n51858 ;
  assign n51862 = n33218 ^ n17411 ^ 1'b0 ;
  assign n51860 = n769 & ~n39033 ;
  assign n51861 = n51860 ^ n19983 ^ 1'b0 ;
  assign n51863 = n51862 ^ n51861 ^ n18993 ;
  assign n51865 = n33419 ^ n11807 ^ n2036 ;
  assign n51864 = n44750 ^ n16616 ^ n13495 ;
  assign n51866 = n51865 ^ n51864 ^ n4038 ;
  assign n51868 = n14428 & ~n19649 ;
  assign n51867 = n36682 ^ n17516 ^ n5332 ;
  assign n51869 = n51868 ^ n51867 ^ n17164 ;
  assign n51870 = ~n7420 & n25992 ;
  assign n51871 = n51870 ^ n44577 ^ n21268 ;
  assign n51872 = ( n18349 & ~n51869 ) | ( n18349 & n51871 ) | ( ~n51869 & n51871 ) ;
  assign n51873 = n4714 | n38517 ;
  assign n51874 = x237 & ~n1891 ;
  assign n51875 = ~n51873 & n51874 ;
  assign n51876 = n34750 ^ n30963 ^ n2258 ;
  assign n51877 = n4532 & ~n27906 ;
  assign n51878 = ~n51876 & n51877 ;
  assign n51879 = n5780 ^ x59 ^ 1'b0 ;
  assign n51880 = n28323 | n51879 ;
  assign n51881 = n16721 & ~n51880 ;
  assign n51882 = n23868 & n51881 ;
  assign n51884 = n6066 & n24529 ;
  assign n51885 = n51884 ^ n19153 ^ 1'b0 ;
  assign n51883 = n13145 & ~n23477 ;
  assign n51886 = n51885 ^ n51883 ^ 1'b0 ;
  assign n51887 = n6019 & n9266 ;
  assign n51888 = n51887 ^ n21286 ^ 1'b0 ;
  assign n51889 = n11138 | n51888 ;
  assign n51890 = n756 & ~n51889 ;
  assign n51891 = n14852 & ~n43852 ;
  assign n51892 = ~n28918 & n51891 ;
  assign n51893 = n3261 | n18028 ;
  assign n51894 = n29143 | n51893 ;
  assign n51895 = ~n16179 & n51894 ;
  assign n51896 = n38016 ^ n8680 ^ n5430 ;
  assign n51897 = n48585 & ~n51896 ;
  assign n51898 = n5829 ^ n3264 ^ n2876 ;
  assign n51899 = n51898 ^ n2290 ^ 1'b0 ;
  assign n51900 = ( n482 & n961 ) | ( n482 & n22416 ) | ( n961 & n22416 ) ;
  assign n51901 = n51786 ^ n48340 ^ 1'b0 ;
  assign n51903 = ~n1986 & n2291 ;
  assign n51904 = n51903 ^ n8263 ^ 1'b0 ;
  assign n51902 = ~n27956 & n32839 ;
  assign n51905 = n51904 ^ n51902 ^ 1'b0 ;
  assign n51906 = n35632 ^ n25222 ^ n17807 ;
  assign n51907 = n39433 | n51906 ;
  assign n51908 = n51907 ^ n26567 ^ 1'b0 ;
  assign n51909 = n11244 ^ n4272 ^ n1961 ;
  assign n51910 = n32636 | n51909 ;
  assign n51911 = ~x170 & n23488 ;
  assign n51912 = n42324 ^ n34096 ^ 1'b0 ;
  assign n51913 = ( ~n26069 & n51911 ) | ( ~n26069 & n51912 ) | ( n51911 & n51912 ) ;
  assign n51914 = n46741 ^ n12365 ^ n1806 ;
  assign n51915 = n15507 & ~n36135 ;
  assign n51916 = ( ~n6139 & n50571 ) | ( ~n6139 & n51915 ) | ( n50571 & n51915 ) ;
  assign n51917 = n30719 & n51299 ;
  assign n51918 = ~n47451 & n51917 ;
  assign n51919 = ( n8913 & ~n31175 ) | ( n8913 & n35003 ) | ( ~n31175 & n35003 ) ;
  assign n51920 = n51919 ^ n25495 ^ 1'b0 ;
  assign n51921 = ~n23465 & n51920 ;
  assign n51922 = ~n4750 & n41610 ;
  assign n51923 = n22643 | n51922 ;
  assign n51924 = n51923 ^ n47295 ^ 1'b0 ;
  assign n51925 = n6723 & ~n35006 ;
  assign n51926 = n51556 & n51925 ;
  assign n51927 = n47538 ^ n13071 ^ n13021 ;
  assign n51928 = n41049 ^ n10384 ^ 1'b0 ;
  assign n51929 = ~n51927 & n51928 ;
  assign n51930 = n26120 ^ n25628 ^ n18977 ;
  assign n51931 = ( ~n19634 & n44951 ) | ( ~n19634 & n51930 ) | ( n44951 & n51930 ) ;
  assign n51932 = ~n12583 & n19595 ;
  assign n51933 = n12483 & ~n22042 ;
  assign n51934 = n21405 ^ n1030 ^ 1'b0 ;
  assign n51935 = n15783 & ~n27391 ;
  assign n51936 = n43191 ^ n42740 ^ 1'b0 ;
  assign n51937 = n12971 & n51936 ;
  assign n51938 = n20491 ^ n12798 ^ n2970 ;
  assign n51939 = n41673 ^ n11921 ^ n1409 ;
  assign n51940 = n16317 & ~n51939 ;
  assign n51941 = n51938 & n51940 ;
  assign n51942 = n18419 ^ n12788 ^ n8306 ;
  assign n51943 = n47424 ^ n12933 ^ 1'b0 ;
  assign n51944 = n51942 & n51943 ;
  assign n51945 = n1163 & n51944 ;
  assign n51946 = ~n11849 & n46643 ;
  assign n51947 = ~n39923 & n51946 ;
  assign n51948 = n39281 ^ n26786 ^ n16213 ;
  assign n51949 = n2386 & n3677 ;
  assign n51950 = ~n51948 & n51949 ;
  assign n51951 = n30826 & ~n36746 ;
  assign n51952 = n38521 ^ n23194 ^ n3074 ;
  assign n51953 = n26069 ^ n17628 ^ n1345 ;
  assign n51954 = ~n423 & n51953 ;
  assign n51955 = n51954 ^ n19929 ^ 1'b0 ;
  assign n51956 = ( n13019 & n21538 ) | ( n13019 & ~n51955 ) | ( n21538 & ~n51955 ) ;
  assign n51957 = ( n12861 & ~n51952 ) | ( n12861 & n51956 ) | ( ~n51952 & n51956 ) ;
  assign n51958 = n16369 ^ n10289 ^ 1'b0 ;
  assign n51959 = ~n7548 & n31924 ;
  assign n51960 = n15745 ^ n9357 ^ x76 ;
  assign n51961 = n11995 & ~n12245 ;
  assign n51962 = n9032 & ~n46027 ;
  assign n51963 = ~n7710 & n51962 ;
  assign n51964 = n5741 & ~n51963 ;
  assign n51965 = ~x218 & n24710 ;
  assign n51966 = ~n4396 & n51965 ;
  assign n51967 = n18098 ^ n12479 ^ 1'b0 ;
  assign n51968 = n9282 & n51967 ;
  assign n51969 = n32960 ^ n9740 ^ 1'b0 ;
  assign n51970 = n38407 | n51969 ;
  assign n51971 = n51970 ^ n45348 ^ n35029 ;
  assign n51972 = ( ~n23873 & n27764 ) | ( ~n23873 & n51971 ) | ( n27764 & n51971 ) ;
  assign n51973 = n39969 ^ n25992 ^ n13859 ;
  assign n51974 = n10802 ^ n830 ^ 1'b0 ;
  assign n51975 = n5452 & ~n43006 ;
  assign n51976 = n1806 & ~n51975 ;
  assign n51977 = n30336 ^ n10370 ^ 1'b0 ;
  assign n51978 = n19443 ^ n4253 ^ 1'b0 ;
  assign n51979 = ~n8411 & n51978 ;
  assign n51980 = n51977 & n51979 ;
  assign n51981 = ~n16250 & n33094 ;
  assign n51982 = ~n47131 & n51981 ;
  assign n51983 = n4307 & n10083 ;
  assign n51984 = n18672 & n51983 ;
  assign n51985 = ~n3227 & n31929 ;
  assign n51986 = n51985 ^ n10562 ^ 1'b0 ;
  assign n51987 = ~n23543 & n51986 ;
  assign n51988 = n44099 ^ n25249 ^ n3697 ;
  assign n51989 = n6013 & n8917 ;
  assign n51990 = ( ~n12862 & n25143 ) | ( ~n12862 & n51989 ) | ( n25143 & n51989 ) ;
  assign n51991 = ( n25808 & n47765 ) | ( n25808 & n51990 ) | ( n47765 & n51990 ) ;
  assign n51992 = n13856 | n23092 ;
  assign n51993 = n51992 ^ n41370 ^ n39412 ;
  assign n51994 = n32562 ^ n16143 ^ 1'b0 ;
  assign n51995 = n15624 ^ n9616 ^ 1'b0 ;
  assign n51996 = ~n51676 & n51995 ;
  assign n51997 = n51996 ^ n42473 ^ 1'b0 ;
  assign n51999 = n403 & ~n14680 ;
  assign n51998 = n14371 | n20060 ;
  assign n52000 = n51999 ^ n51998 ^ 1'b0 ;
  assign n52001 = n11581 ^ n4883 ^ x10 ;
  assign n52002 = n9699 & ~n52001 ;
  assign n52003 = n23320 ^ n3114 ^ 1'b0 ;
  assign n52004 = ~n14596 & n52003 ;
  assign n52005 = ~n20250 & n24295 ;
  assign n52006 = n15094 & ~n41541 ;
  assign n52007 = ~n52005 & n52006 ;
  assign n52008 = n23226 & ~n32339 ;
  assign n52009 = n15144 & n52008 ;
  assign n52010 = n52009 ^ n6917 ^ 1'b0 ;
  assign n52011 = n1924 & n38196 ;
  assign n52012 = n23270 ^ n20090 ^ 1'b0 ;
  assign n52013 = n52012 ^ n25563 ^ n23578 ;
  assign n52014 = n52013 ^ n10027 ^ n8917 ;
  assign n52015 = x132 | n3288 ;
  assign n52016 = n52015 ^ n20821 ^ 1'b0 ;
  assign n52017 = n52016 ^ n29930 ^ n6269 ;
  assign n52018 = ( x123 & n20424 ) | ( x123 & ~n20904 ) | ( n20424 & ~n20904 ) ;
  assign n52019 = n41035 ^ n28733 ^ 1'b0 ;
  assign n52020 = n20940 & ~n52019 ;
  assign n52021 = n14492 & ~n17152 ;
  assign n52022 = n33614 & n52021 ;
  assign n52023 = n30853 & n32496 ;
  assign n52024 = n42063 & n52023 ;
  assign n52025 = n47618 ^ n3404 ^ 1'b0 ;
  assign n52026 = n6204 ^ n2682 ^ 1'b0 ;
  assign n52027 = n52026 ^ n42567 ^ 1'b0 ;
  assign n52028 = n5470 | n52027 ;
  assign n52029 = n3810 ^ n3058 ^ 1'b0 ;
  assign n52032 = n12013 | n32264 ;
  assign n52033 = n10792 & ~n52032 ;
  assign n52030 = n3532 ^ n3521 ^ 1'b0 ;
  assign n52031 = n29927 & ~n52030 ;
  assign n52034 = n52033 ^ n52031 ^ n3754 ;
  assign n52035 = n315 & ~n11909 ;
  assign n52036 = n9997 | n17999 ;
  assign n52037 = n52036 ^ n20664 ^ 1'b0 ;
  assign n52038 = ( n20276 & n37880 ) | ( n20276 & ~n46206 ) | ( n37880 & ~n46206 ) ;
  assign n52039 = ( n2610 & n30715 ) | ( n2610 & n52038 ) | ( n30715 & n52038 ) ;
  assign n52040 = ( n879 & n52037 ) | ( n879 & n52039 ) | ( n52037 & n52039 ) ;
  assign n52041 = n38896 & ~n52040 ;
  assign n52042 = n2561 & ~n5037 ;
  assign n52043 = ( ~n4163 & n5251 ) | ( ~n4163 & n12472 ) | ( n5251 & n12472 ) ;
  assign n52044 = n52043 ^ n47870 ^ 1'b0 ;
  assign n52045 = n52042 & n52044 ;
  assign n52046 = n22826 ^ n20368 ^ 1'b0 ;
  assign n52047 = n40216 ^ n26781 ^ 1'b0 ;
  assign n52048 = n4435 | n52047 ;
  assign n52049 = n52048 ^ n25879 ^ 1'b0 ;
  assign n52050 = n10346 & ~n19522 ;
  assign n52051 = n15908 & ~n26907 ;
  assign n52052 = n27077 ^ n2241 ^ 1'b0 ;
  assign n52053 = ~n9975 & n28967 ;
  assign n52054 = n30339 & n52053 ;
  assign n52055 = ( ~n14080 & n22256 ) | ( ~n14080 & n52054 ) | ( n22256 & n52054 ) ;
  assign n52056 = n9391 ^ n8754 ^ 1'b0 ;
  assign n52057 = n37379 ^ n28127 ^ n8937 ;
  assign n52058 = ( n9127 & n44630 ) | ( n9127 & n52057 ) | ( n44630 & n52057 ) ;
  assign n52059 = ~n3129 & n10601 ;
  assign n52060 = n46681 ^ n41391 ^ 1'b0 ;
  assign n52061 = n11907 & n26644 ;
  assign n52062 = ~n41434 & n52061 ;
  assign n52063 = n19060 ^ n10702 ^ 1'b0 ;
  assign n52064 = n7750 | n52063 ;
  assign n52065 = ~n1745 & n16122 ;
  assign n52066 = n18327 & n52065 ;
  assign n52067 = n14111 & n27998 ;
  assign n52068 = n3775 & n52067 ;
  assign n52069 = ~n8988 & n32245 ;
  assign n52070 = n52069 ^ n35290 ^ 1'b0 ;
  assign n52071 = n40617 ^ n29563 ^ n15002 ;
  assign n52072 = ( n52068 & n52070 ) | ( n52068 & n52071 ) | ( n52070 & n52071 ) ;
  assign n52073 = n47553 ^ n20515 ^ n16188 ;
  assign n52074 = n15673 ^ n14863 ^ n10733 ;
  assign n52075 = n28127 ^ n12869 ^ n10265 ;
  assign n52076 = ( n2528 & ~n9504 ) | ( n2528 & n27679 ) | ( ~n9504 & n27679 ) ;
  assign n52077 = n27999 & n52076 ;
  assign n52078 = n4863 & n33074 ;
  assign n52079 = n996 | n46082 ;
  assign n52085 = n17279 ^ n4267 ^ 1'b0 ;
  assign n52086 = n4124 & n52085 ;
  assign n52084 = ~n2092 & n30195 ;
  assign n52087 = n52086 ^ n52084 ^ 1'b0 ;
  assign n52080 = n13416 ^ n12323 ^ n6831 ;
  assign n52081 = n52080 ^ n47538 ^ n2965 ;
  assign n52082 = n7257 & n52081 ;
  assign n52083 = n12730 & n52082 ;
  assign n52088 = n52087 ^ n52083 ^ 1'b0 ;
  assign n52089 = ( n20384 & n33205 ) | ( n20384 & n52088 ) | ( n33205 & n52088 ) ;
  assign n52090 = ~n15664 & n25590 ;
  assign n52091 = n4412 & ~n52090 ;
  assign n52092 = n7935 | n14196 ;
  assign n52093 = n38859 ^ n34911 ^ 1'b0 ;
  assign n52094 = n52093 ^ n39076 ^ n36029 ;
  assign n52095 = n52094 ^ n40887 ^ n15426 ;
  assign n52100 = ( n9076 & n16707 ) | ( n9076 & n35353 ) | ( n16707 & n35353 ) ;
  assign n52101 = n22910 ^ n9603 ^ n4895 ;
  assign n52102 = ( n12640 & ~n52100 ) | ( n12640 & n52101 ) | ( ~n52100 & n52101 ) ;
  assign n52096 = n22576 & ~n41701 ;
  assign n52097 = n52096 ^ n8242 ^ 1'b0 ;
  assign n52098 = ~n47265 & n52097 ;
  assign n52099 = n52098 ^ n30741 ^ 1'b0 ;
  assign n52103 = n52102 ^ n52099 ^ n41232 ;
  assign n52104 = n3683 | n13950 ;
  assign n52105 = n3683 & ~n52104 ;
  assign n52106 = ( n1903 & n3543 ) | ( n1903 & n52105 ) | ( n3543 & n52105 ) ;
  assign n52107 = n27097 & ~n52106 ;
  assign n52108 = n19592 & n52107 ;
  assign n52109 = ( n8536 & n20507 ) | ( n8536 & ~n52108 ) | ( n20507 & ~n52108 ) ;
  assign n52110 = ~n3722 & n52109 ;
  assign n52111 = ~n11542 & n24326 ;
  assign n52112 = n52111 ^ n31304 ^ 1'b0 ;
  assign n52113 = n47355 | n50645 ;
  assign n52114 = n52113 ^ n33137 ^ 1'b0 ;
  assign n52115 = n25926 & ~n36508 ;
  assign n52116 = n52115 ^ n6463 ^ 1'b0 ;
  assign n52118 = n9496 | n22174 ;
  assign n52119 = n52118 ^ n8569 ^ 1'b0 ;
  assign n52120 = ( x77 & n33799 ) | ( x77 & n52119 ) | ( n33799 & n52119 ) ;
  assign n52117 = n4533 & ~n18389 ;
  assign n52121 = n52120 ^ n52117 ^ 1'b0 ;
  assign n52122 = n32798 ^ n28770 ^ 1'b0 ;
  assign n52123 = n7383 & ~n52122 ;
  assign n52124 = n12037 | n27850 ;
  assign n52125 = n14396 | n52124 ;
  assign n52126 = n17710 & n52125 ;
  assign n52127 = n24448 ^ n15019 ^ n2638 ;
  assign n52128 = ( x92 & n4134 ) | ( x92 & n18229 ) | ( n4134 & n18229 ) ;
  assign n52129 = n26570 ^ n15586 ^ 1'b0 ;
  assign n52130 = n52128 & n52129 ;
  assign n52131 = n7166 & n52130 ;
  assign n52132 = n37557 ^ n23740 ^ n2408 ;
  assign n52133 = ( n14504 & ~n19275 ) | ( n14504 & n52132 ) | ( ~n19275 & n52132 ) ;
  assign n52134 = n45826 ^ n2215 ^ 1'b0 ;
  assign n52135 = n25244 & n32374 ;
  assign n52136 = n52135 ^ n12296 ^ 1'b0 ;
  assign n52137 = n31375 ^ n18026 ^ n3790 ;
  assign n52138 = n5308 & ~n52137 ;
  assign n52139 = ~n40080 & n52138 ;
  assign n52140 = n10007 & ~n33497 ;
  assign n52141 = n52140 ^ n15081 ^ 1'b0 ;
  assign n52142 = n7105 & n52141 ;
  assign n52143 = n40292 ^ n20185 ^ 1'b0 ;
  assign n52144 = n52142 | n52143 ;
  assign n52145 = ( ~n13255 & n28728 ) | ( ~n13255 & n28866 ) | ( n28728 & n28866 ) ;
  assign n52146 = n16572 ^ n8315 ^ x123 ;
  assign n52147 = ( ~n5624 & n6785 ) | ( ~n5624 & n52146 ) | ( n6785 & n52146 ) ;
  assign n52149 = n16473 ^ n6395 ^ n739 ;
  assign n52148 = ~n782 & n48667 ;
  assign n52150 = n52149 ^ n52148 ^ n10445 ;
  assign n52152 = n5208 & n10545 ;
  assign n52151 = x92 & ~x159 ;
  assign n52153 = n52152 ^ n52151 ^ 1'b0 ;
  assign n52154 = ( ~n24099 & n52150 ) | ( ~n24099 & n52153 ) | ( n52150 & n52153 ) ;
  assign n52155 = n22817 ^ n7523 ^ n7198 ;
  assign n52156 = n27947 & n36517 ;
  assign n52157 = ~n32374 & n52156 ;
  assign n52158 = n52157 ^ n32542 ^ 1'b0 ;
  assign n52159 = ~n4527 & n52158 ;
  assign n52160 = n18243 & n52159 ;
  assign n52161 = n33445 ^ n10434 ^ 1'b0 ;
  assign n52162 = n4986 & ~n28142 ;
  assign n52163 = n35558 & n52162 ;
  assign n52164 = ~n14086 & n52163 ;
  assign n52165 = ( n3878 & n24751 ) | ( n3878 & ~n42067 ) | ( n24751 & ~n42067 ) ;
  assign n52166 = n16219 & n52165 ;
  assign n52167 = n30253 ^ n21161 ^ 1'b0 ;
  assign n52168 = n52167 ^ n21759 ^ n8271 ;
  assign n52174 = ( n1043 & n22992 ) | ( n1043 & n49151 ) | ( n22992 & n49151 ) ;
  assign n52175 = ( n6463 & n30190 ) | ( n6463 & ~n52174 ) | ( n30190 & ~n52174 ) ;
  assign n52172 = n20629 & n26035 ;
  assign n52173 = ~n1398 & n52172 ;
  assign n52169 = ( ~n4790 & n26976 ) | ( ~n4790 & n41720 ) | ( n26976 & n41720 ) ;
  assign n52170 = n15868 ^ n15370 ^ 1'b0 ;
  assign n52171 = n52169 & ~n52170 ;
  assign n52176 = n52175 ^ n52173 ^ n52171 ;
  assign n52177 = n52176 ^ n37108 ^ 1'b0 ;
  assign n52180 = n5796 ^ n2100 ^ n1216 ;
  assign n52178 = n1384 & ~n7526 ;
  assign n52179 = n52178 ^ n19171 ^ n11550 ;
  assign n52181 = n52180 ^ n52179 ^ n4350 ;
  assign n52182 = n52181 ^ n44649 ^ n26530 ;
  assign n52183 = ( n3228 & n6171 ) | ( n3228 & n23995 ) | ( n6171 & n23995 ) ;
  assign n52184 = n31668 ^ n3109 ^ 1'b0 ;
  assign n52185 = ~n13441 & n32247 ;
  assign n52186 = n34245 & n52185 ;
  assign n52187 = ~n12041 & n50823 ;
  assign n52188 = n52187 ^ n30671 ^ 1'b0 ;
  assign n52189 = n3940 & n4281 ;
  assign n52190 = ~n4281 & n52189 ;
  assign n52191 = n12041 | n52190 ;
  assign n52192 = ~n4632 & n44705 ;
  assign n52193 = n52191 & n52192 ;
  assign n52194 = n25571 ^ n5138 ^ 1'b0 ;
  assign n52195 = ~n52193 & n52194 ;
  assign n52196 = n11233 ^ n579 ^ 1'b0 ;
  assign n52197 = n52196 ^ n34168 ^ 1'b0 ;
  assign n52202 = n4794 ^ n2325 ^ 1'b0 ;
  assign n52203 = n24235 & n52202 ;
  assign n52204 = n5949 & ~n52203 ;
  assign n52205 = n28640 & ~n52204 ;
  assign n52206 = n7544 & n52205 ;
  assign n52198 = n13255 ^ n10958 ^ n9742 ;
  assign n52199 = n52198 ^ n19716 ^ n8619 ;
  assign n52200 = n21382 ^ n14779 ^ 1'b0 ;
  assign n52201 = n52199 & n52200 ;
  assign n52207 = n52206 ^ n52201 ^ n39442 ;
  assign n52208 = n52207 ^ n49500 ^ n7482 ;
  assign n52209 = n13774 | n26653 ;
  assign n52210 = n11727 & ~n52209 ;
  assign n52211 = n52210 ^ n6382 ^ n4673 ;
  assign n52212 = ( n2321 & n28188 ) | ( n2321 & ~n52211 ) | ( n28188 & ~n52211 ) ;
  assign n52213 = n537 | n1780 ;
  assign n52214 = n537 & ~n52213 ;
  assign n52215 = n2825 & ~n52214 ;
  assign n52216 = n52215 ^ n13490 ^ n831 ;
  assign n52217 = n52216 ^ n19397 ^ n5059 ;
  assign n52218 = n28861 ^ n21052 ^ n15743 ;
  assign n52219 = ~n8522 & n25852 ;
  assign n52220 = ~n50162 & n52219 ;
  assign n52221 = ~n1909 & n21157 ;
  assign n52222 = n52220 & n52221 ;
  assign n52223 = n51357 ^ n23588 ^ 1'b0 ;
  assign n52224 = ~n45642 & n52223 ;
  assign n52225 = n45600 ^ n36755 ^ 1'b0 ;
  assign n52226 = n34842 ^ n28198 ^ n12988 ;
  assign n52227 = n7190 | n52226 ;
  assign n52228 = n52225 & ~n52227 ;
  assign n52229 = n42341 ^ n3371 ^ 1'b0 ;
  assign n52230 = n22814 & ~n52229 ;
  assign n52231 = n16729 ^ n10573 ^ 1'b0 ;
  assign n52232 = n1467 | n45475 ;
  assign n52233 = n52232 ^ n24666 ^ 1'b0 ;
  assign n52234 = n52233 ^ n20319 ^ 1'b0 ;
  assign n52235 = n26112 | n26708 ;
  assign n52236 = ( ~n20191 & n38520 ) | ( ~n20191 & n52235 ) | ( n38520 & n52235 ) ;
  assign n52237 = ( n31285 & n46820 ) | ( n31285 & ~n52236 ) | ( n46820 & ~n52236 ) ;
  assign n52238 = n40210 ^ n20575 ^ n11245 ;
  assign n52239 = ~n15898 & n18415 ;
  assign n52240 = n52239 ^ n7007 ^ 1'b0 ;
  assign n52241 = ( n2101 & ~n52238 ) | ( n2101 & n52240 ) | ( ~n52238 & n52240 ) ;
  assign n52242 = n52241 ^ n19239 ^ n6705 ;
  assign n52243 = ( n8039 & n8045 ) | ( n8039 & n15405 ) | ( n8045 & n15405 ) ;
  assign n52244 = ~n9379 & n49099 ;
  assign n52245 = n2039 ^ n812 ^ 1'b0 ;
  assign n52246 = x31 & n52245 ;
  assign n52247 = n52246 ^ n36081 ^ n17507 ;
  assign n52248 = n11588 & n52247 ;
  assign n52249 = n52248 ^ n43519 ^ 1'b0 ;
  assign n52250 = n28870 | n49069 ;
  assign n52251 = n7159 & n24274 ;
  assign n52252 = n52250 & n52251 ;
  assign n52253 = n12389 & n23073 ;
  assign n52254 = n1921 & ~n52253 ;
  assign n52255 = ( n22362 & n38616 ) | ( n22362 & n52254 ) | ( n38616 & n52254 ) ;
  assign n52257 = n33850 ^ n9784 ^ 1'b0 ;
  assign n52258 = n29060 | n52257 ;
  assign n52256 = n16981 & n52042 ;
  assign n52259 = n52258 ^ n52256 ^ 1'b0 ;
  assign n52260 = n52259 ^ n11438 ^ n6739 ;
  assign n52261 = ~n5975 & n18862 ;
  assign n52262 = n33877 & ~n39914 ;
  assign n52263 = ( n22904 & n36556 ) | ( n22904 & ~n52262 ) | ( n36556 & ~n52262 ) ;
  assign n52264 = ( n8908 & ~n16276 ) | ( n8908 & n27415 ) | ( ~n16276 & n27415 ) ;
  assign n52265 = n52264 ^ n31424 ^ n3532 ;
  assign n52266 = n2613 & n25067 ;
  assign n52267 = n11766 & ~n19948 ;
  assign n52268 = n52267 ^ n25167 ^ 1'b0 ;
  assign n52269 = ~n2397 & n15694 ;
  assign n52270 = n52269 ^ n34838 ^ 1'b0 ;
  assign n52271 = ~n20598 & n28307 ;
  assign n52272 = n32198 ^ n21036 ^ n14194 ;
  assign n52273 = n52271 & ~n52272 ;
  assign n52274 = ( n14995 & n33075 ) | ( n14995 & n52273 ) | ( n33075 & n52273 ) ;
  assign n52275 = n52274 ^ n44456 ^ n37048 ;
  assign n52276 = ( ~n8814 & n11654 ) | ( ~n8814 & n18195 ) | ( n11654 & n18195 ) ;
  assign n52277 = ( n26946 & ~n28087 ) | ( n26946 & n52276 ) | ( ~n28087 & n52276 ) ;
  assign n52278 = n27753 ^ n13145 ^ 1'b0 ;
  assign n52279 = ( ~n14617 & n15283 ) | ( ~n14617 & n47372 ) | ( n15283 & n47372 ) ;
  assign n52280 = n615 | n47669 ;
  assign n52283 = n8555 | n16021 ;
  assign n52284 = n15829 | n52283 ;
  assign n52282 = n10492 | n20196 ;
  assign n52285 = n52284 ^ n52282 ^ 1'b0 ;
  assign n52286 = ( n2832 & ~n30575 ) | ( n2832 & n52285 ) | ( ~n30575 & n52285 ) ;
  assign n52281 = n7653 & n10767 ;
  assign n52287 = n52286 ^ n52281 ^ 1'b0 ;
  assign n52288 = ~n41612 & n49951 ;
  assign n52289 = n7694 ^ n7493 ^ 1'b0 ;
  assign n52290 = n27107 & ~n52289 ;
  assign n52291 = ~n28062 & n52290 ;
  assign n52292 = n7289 ^ n4417 ^ 1'b0 ;
  assign n52293 = n44066 | n52292 ;
  assign n52294 = n17719 ^ n16062 ^ 1'b0 ;
  assign n52295 = ( n23249 & n28800 ) | ( n23249 & n52294 ) | ( n28800 & n52294 ) ;
  assign n52296 = ~n33855 & n52295 ;
  assign n52297 = n52296 ^ n8861 ^ 1'b0 ;
  assign n52298 = n45940 & n52297 ;
  assign n52299 = n16260 | n18010 ;
  assign n52300 = n52298 & ~n52299 ;
  assign n52301 = n52293 & n52300 ;
  assign n52302 = n45782 ^ n28179 ^ n10114 ;
  assign n52303 = n11762 ^ n6763 ^ n2767 ;
  assign n52304 = n20461 & ~n40524 ;
  assign n52305 = n52304 ^ n34131 ^ n32828 ;
  assign n52306 = n3208 | n22418 ;
  assign n52307 = n52306 ^ n22934 ^ 1'b0 ;
  assign n52308 = n52307 ^ n36392 ^ n10562 ;
  assign n52309 = n15414 ^ n1231 ^ 1'b0 ;
  assign n52310 = ~n3101 & n52309 ;
  assign n52311 = n1393 | n39514 ;
  assign n52312 = n46620 & ~n52311 ;
  assign n52313 = n52312 ^ n3980 ^ 1'b0 ;
  assign n52314 = n37450 ^ n7482 ^ 1'b0 ;
  assign n52315 = n26626 & n52314 ;
  assign n52316 = n19465 & ~n39385 ;
  assign n52317 = n17681 & n51770 ;
  assign n52318 = ~n52316 & n52317 ;
  assign n52319 = ~n25736 & n32661 ;
  assign n52320 = n34519 & n52319 ;
  assign n52321 = n6865 | n21295 ;
  assign n52322 = n52321 ^ n30442 ^ 1'b0 ;
  assign n52323 = n14364 & n14991 ;
  assign n52324 = n18636 & n52323 ;
  assign n52325 = n52324 ^ n12193 ^ 1'b0 ;
  assign n52326 = n3258 | n23184 ;
  assign n52327 = n24057 & ~n52326 ;
  assign n52328 = ( n27965 & ~n36589 ) | ( n27965 & n52327 ) | ( ~n36589 & n52327 ) ;
  assign n52329 = n25520 ^ n13666 ^ 1'b0 ;
  assign n52330 = n2651 | n39901 ;
  assign n52331 = n52330 ^ n31139 ^ n10500 ;
  assign n52332 = n16860 | n31861 ;
  assign n52333 = n31279 ^ n1024 ^ 1'b0 ;
  assign n52334 = n14810 | n52333 ;
  assign n52335 = n3716 & n38664 ;
  assign n52336 = n52335 ^ n37682 ^ 1'b0 ;
  assign n52337 = n266 & n30382 ;
  assign n52338 = n9078 | n16826 ;
  assign n52339 = n36991 | n52338 ;
  assign n52340 = ~n5000 & n52339 ;
  assign n52341 = ~n52337 & n52340 ;
  assign n52342 = n3665 & n10464 ;
  assign n52343 = n6274 & n52342 ;
  assign n52344 = n4819 & n28967 ;
  assign n52345 = n52344 ^ n23995 ^ 1'b0 ;
  assign n52346 = ( n3639 & n12607 ) | ( n3639 & ~n22096 ) | ( n12607 & ~n22096 ) ;
  assign n52347 = n41559 ^ n9907 ^ 1'b0 ;
  assign n52353 = n30776 ^ n23922 ^ 1'b0 ;
  assign n52354 = n13623 & ~n52353 ;
  assign n52351 = n29621 ^ n12596 ^ n5604 ;
  assign n52348 = n41698 ^ n26153 ^ n18676 ;
  assign n52349 = n23258 & ~n52348 ;
  assign n52350 = ~n13040 & n52349 ;
  assign n52352 = n52351 ^ n52350 ^ 1'b0 ;
  assign n52355 = n52354 ^ n52352 ^ 1'b0 ;
  assign n52356 = ( n52346 & ~n52347 ) | ( n52346 & n52355 ) | ( ~n52347 & n52355 ) ;
  assign n52357 = n52356 ^ n50454 ^ n45983 ;
  assign n52358 = n1501 | n28397 ;
  assign n52359 = ( n13239 & n21375 ) | ( n13239 & ~n52358 ) | ( n21375 & ~n52358 ) ;
  assign n52360 = n11188 & n33006 ;
  assign n52361 = n52360 ^ n29571 ^ 1'b0 ;
  assign n52363 = n26886 ^ n6242 ^ 1'b0 ;
  assign n52364 = n13066 & ~n52363 ;
  assign n52362 = ( n818 & ~n22206 ) | ( n818 & n24284 ) | ( ~n22206 & n24284 ) ;
  assign n52365 = n52364 ^ n52362 ^ 1'b0 ;
  assign n52366 = ~n6795 & n20844 ;
  assign n52367 = n52366 ^ n23623 ^ 1'b0 ;
  assign n52368 = n18203 & n52367 ;
  assign n52369 = ( ~n20804 & n21914 ) | ( ~n20804 & n29241 ) | ( n21914 & n29241 ) ;
  assign n52370 = n19124 & n47612 ;
  assign n52371 = ( n32420 & ~n52369 ) | ( n32420 & n52370 ) | ( ~n52369 & n52370 ) ;
  assign n52372 = n23200 ^ n2252 ^ 1'b0 ;
  assign n52373 = n28792 ^ n19639 ^ 1'b0 ;
  assign n52374 = n38016 & ~n44844 ;
  assign n52375 = n52374 ^ n9700 ^ 1'b0 ;
  assign n52376 = n52375 ^ n10555 ^ 1'b0 ;
  assign n52377 = ( n15714 & n17842 ) | ( n15714 & n28541 ) | ( n17842 & n28541 ) ;
  assign n52378 = n5357 & n29419 ;
  assign n52380 = n41030 ^ n34559 ^ n15734 ;
  assign n52379 = n3169 & ~n5701 ;
  assign n52381 = n52380 ^ n52379 ^ 1'b0 ;
  assign n52383 = n6595 & ~n30805 ;
  assign n52382 = ~n4242 & n26182 ;
  assign n52384 = n52383 ^ n52382 ^ 1'b0 ;
  assign n52385 = n8211 ^ n4187 ^ 1'b0 ;
  assign n52386 = x97 & n916 ;
  assign n52387 = n2865 & n12160 ;
  assign n52388 = n52386 & n52387 ;
  assign n52389 = n327 & ~n22191 ;
  assign n52390 = n52389 ^ n25105 ^ 1'b0 ;
  assign n52391 = n36473 & n52390 ;
  assign n52392 = n29745 ^ n2444 ^ 1'b0 ;
  assign n52393 = n5608 & ~n52392 ;
  assign n52394 = ( n15104 & ~n16631 ) | ( n15104 & n52393 ) | ( ~n16631 & n52393 ) ;
  assign n52395 = n32208 ^ n29063 ^ 1'b0 ;
  assign n52396 = n35883 ^ n12796 ^ n7499 ;
  assign n52397 = ( n19797 & n26381 ) | ( n19797 & n52396 ) | ( n26381 & n52396 ) ;
  assign n52398 = n28950 ^ n21417 ^ 1'b0 ;
  assign n52399 = ~n36730 & n52398 ;
  assign n52400 = ( n18781 & ~n52397 ) | ( n18781 & n52399 ) | ( ~n52397 & n52399 ) ;
  assign n52401 = n24575 ^ n14147 ^ n7970 ;
  assign n52402 = n2923 & n18523 ;
  assign n52403 = n20551 & n52402 ;
  assign n52404 = n2750 & n18352 ;
  assign n52405 = n9787 | n52404 ;
  assign n52406 = n47701 ^ n20842 ^ 1'b0 ;
  assign n52407 = n14139 & n52406 ;
  assign n52408 = n52407 ^ n2662 ^ 1'b0 ;
  assign n52409 = n52405 & n52408 ;
  assign n52410 = ( n516 & n52403 ) | ( n516 & n52409 ) | ( n52403 & n52409 ) ;
  assign n52411 = ~n27504 & n29217 ;
  assign n52412 = ~n52410 & n52411 ;
  assign n52414 = n11437 ^ n9940 ^ n5528 ;
  assign n52415 = ~n11864 & n52414 ;
  assign n52413 = n22670 & ~n52258 ;
  assign n52416 = n52415 ^ n52413 ^ 1'b0 ;
  assign n52417 = n4294 & ~n20630 ;
  assign n52418 = n52417 ^ n2499 ^ 1'b0 ;
  assign n52419 = n52418 ^ n34460 ^ 1'b0 ;
  assign n52420 = n34746 ^ n1554 ^ 1'b0 ;
  assign n52421 = n32516 | n52420 ;
  assign n52422 = ~n11340 & n44529 ;
  assign n52423 = n2907 ^ n1149 ^ 1'b0 ;
  assign n52424 = n34766 | n52423 ;
  assign n52425 = n29824 ^ n3468 ^ 1'b0 ;
  assign n52426 = n25268 & ~n25923 ;
  assign n52427 = n52426 ^ n36447 ^ n22873 ;
  assign n52428 = n28168 & ~n34729 ;
  assign n52429 = ~n9280 & n52428 ;
  assign n52430 = n52429 ^ n41786 ^ x137 ;
  assign n52431 = n10774 ^ n10755 ^ n8823 ;
  assign n52432 = n52431 ^ n18855 ^ n9178 ;
  assign n52433 = ( x49 & n2031 ) | ( x49 & n52432 ) | ( n2031 & n52432 ) ;
  assign n52434 = n17964 ^ n2788 ^ 1'b0 ;
  assign n52435 = n52433 & n52434 ;
  assign n52436 = n4217 | n31570 ;
  assign n52437 = n26080 ^ n22398 ^ n10665 ;
  assign n52438 = n5439 & ~n13054 ;
  assign n52439 = ( n9289 & n19206 ) | ( n9289 & n52438 ) | ( n19206 & n52438 ) ;
  assign n52440 = n52439 ^ n48197 ^ 1'b0 ;
  assign n52441 = n5196 | n52440 ;
  assign n52442 = n52437 & ~n52441 ;
  assign n52443 = ( ~n4274 & n38808 ) | ( ~n4274 & n50762 ) | ( n38808 & n50762 ) ;
  assign n52444 = ( ~n9015 & n42277 ) | ( ~n9015 & n44909 ) | ( n42277 & n44909 ) ;
  assign n52445 = n22310 ^ n17035 ^ n12492 ;
  assign n52446 = n47090 ^ n16659 ^ n4996 ;
  assign n52447 = n33153 & ~n37571 ;
  assign n52448 = n52447 ^ n36204 ^ 1'b0 ;
  assign n52449 = n7120 & n33438 ;
  assign n52450 = ~n19650 & n52449 ;
  assign n52453 = ( n4003 & n7957 ) | ( n4003 & ~n19604 ) | ( n7957 & ~n19604 ) ;
  assign n52451 = n24414 ^ n21624 ^ n15698 ;
  assign n52452 = ~n27435 & n52451 ;
  assign n52454 = n52453 ^ n52452 ^ 1'b0 ;
  assign n52455 = n15172 & n18534 ;
  assign n52456 = n52455 ^ n12491 ^ 1'b0 ;
  assign n52457 = n48512 ^ n27978 ^ n18410 ;
  assign n52458 = ~n692 & n36197 ;
  assign n52459 = ( n3123 & n14796 ) | ( n3123 & ~n41157 ) | ( n14796 & ~n41157 ) ;
  assign n52460 = n27108 ^ n9623 ^ n6393 ;
  assign n52461 = n50970 & ~n52460 ;
  assign n52462 = n52461 ^ n27314 ^ 1'b0 ;
  assign n52463 = n28896 | n43430 ;
  assign n52464 = n52463 ^ n21389 ^ 1'b0 ;
  assign n52465 = n44821 ^ n44774 ^ n14758 ;
  assign n52466 = ~n6480 & n52465 ;
  assign n52467 = ~n25974 & n35533 ;
  assign n52468 = n52467 ^ n514 ^ 1'b0 ;
  assign n52469 = n50595 ^ n12174 ^ 1'b0 ;
  assign n52470 = n52469 ^ n51088 ^ n10258 ;
  assign n52471 = n15552 ^ n10534 ^ 1'b0 ;
  assign n52472 = ( n9745 & ~n15862 ) | ( n9745 & n52471 ) | ( ~n15862 & n52471 ) ;
  assign n52473 = n12466 & ~n31283 ;
  assign n52474 = ~n52472 & n52473 ;
  assign n52475 = n16250 ^ n15016 ^ 1'b0 ;
  assign n52476 = ( ~n11373 & n23337 ) | ( ~n11373 & n50030 ) | ( n23337 & n50030 ) ;
  assign n52477 = ( n16468 & ~n22256 ) | ( n16468 & n52476 ) | ( ~n22256 & n52476 ) ;
  assign n52478 = n6425 & n29902 ;
  assign n52479 = n29364 ^ n19619 ^ 1'b0 ;
  assign n52480 = n1524 & n27703 ;
  assign n52481 = n52480 ^ n27231 ^ 1'b0 ;
  assign n52482 = n12905 ^ n4232 ^ 1'b0 ;
  assign n52483 = n13310 ^ n3510 ^ 1'b0 ;
  assign n52484 = ( n9855 & n14817 ) | ( n9855 & ~n18026 ) | ( n14817 & ~n18026 ) ;
  assign n52485 = n52484 ^ n26984 ^ n16542 ;
  assign n52486 = ~n2689 & n52485 ;
  assign n52487 = ( n1468 & n15747 ) | ( n1468 & n40343 ) | ( n15747 & n40343 ) ;
  assign n52489 = n9498 | n31360 ;
  assign n52490 = n8659 & ~n52489 ;
  assign n52491 = n52490 ^ n35092 ^ 1'b0 ;
  assign n52488 = n23156 ^ n21572 ^ n13452 ;
  assign n52492 = n52491 ^ n52488 ^ n14421 ;
  assign n52493 = ( ~n8835 & n11710 ) | ( ~n8835 & n28738 ) | ( n11710 & n28738 ) ;
  assign n52494 = ( n7166 & n17273 ) | ( n7166 & ~n23833 ) | ( n17273 & ~n23833 ) ;
  assign n52495 = ( n52380 & ~n52493 ) | ( n52380 & n52494 ) | ( ~n52493 & n52494 ) ;
  assign n52496 = n688 | n12541 ;
  assign n52497 = n21500 | n52496 ;
  assign n52498 = n36933 ^ n27457 ^ 1'b0 ;
  assign n52499 = n46179 ^ n21904 ^ n15337 ;
  assign n52500 = n52499 ^ n28506 ^ 1'b0 ;
  assign n52501 = n52498 | n52500 ;
  assign n52502 = n39275 ^ n21026 ^ 1'b0 ;
  assign n52503 = n13989 & n52502 ;
  assign n52504 = n52503 ^ n13299 ^ 1'b0 ;
  assign n52505 = n25334 ^ n11692 ^ 1'b0 ;
  assign n52506 = x159 & n52505 ;
  assign n52507 = n38140 ^ n3404 ^ 1'b0 ;
  assign n52508 = n4958 ^ n2326 ^ 1'b0 ;
  assign n52509 = n9098 | n52508 ;
  assign n52510 = ( ~n25284 & n28905 ) | ( ~n25284 & n52509 ) | ( n28905 & n52509 ) ;
  assign n52511 = ( n32637 & n39098 ) | ( n32637 & ~n42246 ) | ( n39098 & ~n42246 ) ;
  assign n52512 = ( n2610 & n9966 ) | ( n2610 & ~n49546 ) | ( n9966 & ~n49546 ) ;
  assign n52513 = n52512 ^ n3449 ^ 1'b0 ;
  assign n52514 = ~n22878 & n30109 ;
  assign n52515 = n52514 ^ n11976 ^ n4386 ;
  assign n52516 = n5995 & ~n7727 ;
  assign n52517 = n52516 ^ n44810 ^ n39125 ;
  assign n52518 = n9095 & ~n52517 ;
  assign n52519 = ~n24868 & n32554 ;
  assign n52520 = n9501 | n30705 ;
  assign n52521 = n22053 & ~n52520 ;
  assign n52522 = n12739 | n49402 ;
  assign n52523 = n35094 | n52522 ;
  assign n52524 = n12897 | n26644 ;
  assign n52525 = n52472 ^ n21012 ^ n8031 ;
  assign n52526 = ( n41026 & ~n52524 ) | ( n41026 & n52525 ) | ( ~n52524 & n52525 ) ;
  assign n52527 = n21108 ^ n14432 ^ 1'b0 ;
  assign n52528 = ( n20546 & n22884 ) | ( n20546 & ~n24080 ) | ( n22884 & ~n24080 ) ;
  assign n52529 = ( n11050 & ~n11587 ) | ( n11050 & n23474 ) | ( ~n11587 & n23474 ) ;
  assign n52530 = n4005 & ~n52529 ;
  assign n52531 = n52530 ^ n27395 ^ 1'b0 ;
  assign n52532 = n1385 & n52531 ;
  assign n52533 = ~n17162 & n48050 ;
  assign n52534 = n33443 ^ n7675 ^ 1'b0 ;
  assign n52535 = n33896 | n52534 ;
  assign n52536 = ~n6838 & n8483 ;
  assign n52537 = n52535 & n52536 ;
  assign n52538 = n21851 & ~n49235 ;
  assign n52539 = n52538 ^ n24749 ^ 1'b0 ;
  assign n52540 = n19446 | n52539 ;
  assign n52541 = n52540 ^ n34703 ^ 1'b0 ;
  assign n52543 = n12254 ^ n8209 ^ 1'b0 ;
  assign n52542 = n14797 & ~n25941 ;
  assign n52544 = n52543 ^ n52542 ^ 1'b0 ;
  assign n52545 = n8783 & n19900 ;
  assign n52546 = ~n17314 & n52545 ;
  assign n52547 = n50901 ^ n27978 ^ n13205 ;
  assign n52548 = n7250 & ~n52547 ;
  assign n52549 = n52548 ^ n22662 ^ 1'b0 ;
  assign n52550 = n52549 ^ n16062 ^ 1'b0 ;
  assign n52551 = ~n1411 & n52550 ;
  assign n52552 = ( n20023 & n52546 ) | ( n20023 & n52551 ) | ( n52546 & n52551 ) ;
  assign n52554 = ~n28928 & n38708 ;
  assign n52553 = ( ~n11157 & n14436 ) | ( ~n11157 & n19822 ) | ( n14436 & n19822 ) ;
  assign n52555 = n52554 ^ n52553 ^ n52351 ;
  assign n52556 = n8841 & n30176 ;
  assign n52557 = n52556 ^ n9541 ^ 1'b0 ;
  assign n52558 = n52557 ^ n10799 ^ 1'b0 ;
  assign n52559 = n48797 ^ n48154 ^ n14021 ;
  assign n52560 = ( n15651 & n34483 ) | ( n15651 & n46217 ) | ( n34483 & n46217 ) ;
  assign n52561 = ~n25941 & n31572 ;
  assign n52562 = ~n52560 & n52561 ;
  assign n52564 = n6075 & n28473 ;
  assign n52563 = n337 & n3429 ;
  assign n52565 = n52564 ^ n52563 ^ 1'b0 ;
  assign n52566 = n14899 & n44915 ;
  assign n52567 = n52565 & n52566 ;
  assign n52568 = n26860 & n52567 ;
  assign n52569 = x210 & ~n28771 ;
  assign n52570 = ~n16258 & n52569 ;
  assign n52571 = ~n13664 & n38969 ;
  assign n52572 = n52570 & n52571 ;
  assign n52573 = n50792 ^ n40211 ^ 1'b0 ;
  assign n52574 = n46179 & ~n52573 ;
  assign n52575 = n16074 | n46262 ;
  assign n52576 = n21460 | n52575 ;
  assign n52577 = ( ~n3318 & n9959 ) | ( ~n3318 & n21161 ) | ( n9959 & n21161 ) ;
  assign n52578 = n52577 ^ n34432 ^ 1'b0 ;
  assign n52579 = n25033 & n44631 ;
  assign n52580 = n52579 ^ n51894 ^ 1'b0 ;
  assign n52581 = n52580 ^ n31295 ^ n7324 ;
  assign n52582 = ( n1885 & ~n36330 ) | ( n1885 & n52120 ) | ( ~n36330 & n52120 ) ;
  assign n52583 = ( n2243 & n7166 ) | ( n2243 & ~n15422 ) | ( n7166 & ~n15422 ) ;
  assign n52586 = n28535 ^ n27066 ^ n21783 ;
  assign n52584 = n34940 ^ n22141 ^ 1'b0 ;
  assign n52585 = n8280 & n52584 ;
  assign n52587 = n52586 ^ n52585 ^ 1'b0 ;
  assign n52588 = n30856 ^ n5686 ^ 1'b0 ;
  assign n52589 = n34876 & ~n52588 ;
  assign n52590 = n48172 ^ n28592 ^ n11704 ;
  assign n52591 = ~n43587 & n52590 ;
  assign n52592 = ~n360 & n8004 ;
  assign n52593 = n52592 ^ n6620 ^ 1'b0 ;
  assign n52594 = ( n4045 & n10071 ) | ( n4045 & n24730 ) | ( n10071 & n24730 ) ;
  assign n52595 = ( n17048 & n52593 ) | ( n17048 & n52594 ) | ( n52593 & n52594 ) ;
  assign n52596 = n46749 ^ n10185 ^ n6274 ;
  assign n52597 = n50317 & n52596 ;
  assign n52598 = ( n13116 & n52595 ) | ( n13116 & n52597 ) | ( n52595 & n52597 ) ;
  assign n52599 = n17189 ^ n1450 ^ 1'b0 ;
  assign n52600 = n50836 | n52599 ;
  assign n52601 = n52600 ^ n36198 ^ 1'b0 ;
  assign n52602 = n42927 ^ n9760 ^ n8493 ;
  assign n52603 = ( n9809 & n35069 ) | ( n9809 & n37171 ) | ( n35069 & n37171 ) ;
  assign n52604 = ( ~n7986 & n28313 ) | ( ~n7986 & n52603 ) | ( n28313 & n52603 ) ;
  assign n52605 = ( n49883 & n52602 ) | ( n49883 & ~n52604 ) | ( n52602 & ~n52604 ) ;
  assign n52606 = ( ~n3551 & n32319 ) | ( ~n3551 & n45554 ) | ( n32319 & n45554 ) ;
  assign n52607 = n5303 ^ n487 ^ 1'b0 ;
  assign n52608 = n23913 & n52607 ;
  assign n52609 = ~n3933 & n40254 ;
  assign n52610 = n34351 & n52609 ;
  assign n52611 = n21053 & ~n23909 ;
  assign n52612 = n52610 & ~n52611 ;
  assign n52613 = ~n1154 & n1512 ;
  assign n52614 = ( n33840 & n34556 ) | ( n33840 & ~n47141 ) | ( n34556 & ~n47141 ) ;
  assign n52615 = n1948 & ~n26578 ;
  assign n52616 = ~n52614 & n52615 ;
  assign n52617 = n27330 ^ n5221 ^ 1'b0 ;
  assign n52618 = ~n16865 & n52617 ;
  assign n52619 = n2180 & n36809 ;
  assign n52620 = ~n52618 & n52619 ;
  assign n52621 = ( n7357 & ~n13713 ) | ( n7357 & n18295 ) | ( ~n13713 & n18295 ) ;
  assign n52622 = ( ~n2818 & n9703 ) | ( ~n2818 & n16797 ) | ( n9703 & n16797 ) ;
  assign n52623 = n52622 ^ n25064 ^ n5363 ;
  assign n52624 = n18281 & ~n45490 ;
  assign n52625 = n35149 ^ n4961 ^ 1'b0 ;
  assign n52626 = ~n6431 & n43915 ;
  assign n52627 = n52626 ^ n26708 ^ 1'b0 ;
  assign n52628 = ~n34994 & n51187 ;
  assign n52629 = ~n5183 & n52628 ;
  assign n52630 = ~n4868 & n47352 ;
  assign n52631 = n13929 & n52630 ;
  assign n52632 = n16908 ^ n14347 ^ 1'b0 ;
  assign n52633 = ( ~n1984 & n10005 ) | ( ~n1984 & n52632 ) | ( n10005 & n52632 ) ;
  assign n52634 = n52633 ^ n39422 ^ n11100 ;
  assign n52635 = n12780 ^ n5882 ^ n4478 ;
  assign n52636 = ( n8337 & n9312 ) | ( n8337 & n52635 ) | ( n9312 & n52635 ) ;
  assign n52637 = n42111 ^ n35552 ^ 1'b0 ;
  assign n52638 = ~n52636 & n52637 ;
  assign n52639 = ( ~n18960 & n52634 ) | ( ~n18960 & n52638 ) | ( n52634 & n52638 ) ;
  assign n52640 = n27961 & n30366 ;
  assign n52641 = n23001 ^ n3235 ^ 1'b0 ;
  assign n52642 = n20871 & n52641 ;
  assign n52643 = n52642 ^ n13810 ^ 1'b0 ;
  assign n52644 = n52643 ^ n33668 ^ n9118 ;
  assign n52645 = n7237 ^ n7073 ^ 1'b0 ;
  assign n52646 = n26600 & n52645 ;
  assign n52647 = ( n5466 & ~n7136 ) | ( n5466 & n52646 ) | ( ~n7136 & n52646 ) ;
  assign n52648 = n13527 & ~n37307 ;
  assign n52649 = n13079 ^ n2995 ^ 1'b0 ;
  assign n52650 = n21347 ^ n8386 ^ 1'b0 ;
  assign n52651 = n41687 ^ n21341 ^ n19545 ;
  assign n52652 = n38788 & ~n52651 ;
  assign n52653 = n9250 & n52652 ;
  assign n52654 = ( n52649 & n52650 ) | ( n52649 & ~n52653 ) | ( n52650 & ~n52653 ) ;
  assign n52655 = n7294 & n8981 ;
  assign n52656 = ~n52654 & n52655 ;
  assign n52657 = n9162 & ~n49943 ;
  assign n52658 = n52657 ^ n40227 ^ 1'b0 ;
  assign n52659 = ( n1981 & ~n5315 ) | ( n1981 & n49906 ) | ( ~n5315 & n49906 ) ;
  assign n52660 = n7752 & ~n52659 ;
  assign n52661 = n16381 ^ n13752 ^ 1'b0 ;
  assign n52662 = n25486 & n52661 ;
  assign n52663 = n50699 & n52662 ;
  assign n52664 = n52663 ^ n25882 ^ 1'b0 ;
  assign n52665 = n5029 | n8133 ;
  assign n52666 = n33658 & ~n39055 ;
  assign n52667 = n36239 & n52666 ;
  assign n52668 = ( ~n27643 & n52665 ) | ( ~n27643 & n52667 ) | ( n52665 & n52667 ) ;
  assign n52669 = n51739 ^ n44453 ^ n26952 ;
  assign n52670 = n13813 ^ n11560 ^ 1'b0 ;
  assign n52671 = ( n40404 & n41353 ) | ( n40404 & ~n52670 ) | ( n41353 & ~n52670 ) ;
  assign n52672 = ( n4939 & ~n12262 ) | ( n4939 & n16760 ) | ( ~n12262 & n16760 ) ;
  assign n52673 = n52672 ^ n39548 ^ n6483 ;
  assign n52674 = ( n8919 & n52671 ) | ( n8919 & n52673 ) | ( n52671 & n52673 ) ;
  assign n52675 = ( ~n18200 & n27057 ) | ( ~n18200 & n48476 ) | ( n27057 & n48476 ) ;
  assign n52679 = ( n11354 & n13158 ) | ( n11354 & ~n18470 ) | ( n13158 & ~n18470 ) ;
  assign n52676 = n7181 & ~n15771 ;
  assign n52677 = n7827 & n52676 ;
  assign n52678 = n52677 ^ n26294 ^ n13417 ;
  assign n52680 = n52679 ^ n52678 ^ n11367 ;
  assign n52681 = n34192 ^ n17735 ^ 1'b0 ;
  assign n52682 = n39937 ^ n37847 ^ 1'b0 ;
  assign n52683 = n5226 & ~n18793 ;
  assign n52684 = ~n3535 & n5996 ;
  assign n52685 = n52684 ^ n12278 ^ 1'b0 ;
  assign n52686 = n30018 ^ n25801 ^ 1'b0 ;
  assign n52687 = n52685 | n52686 ;
  assign n52688 = n11658 | n19711 ;
  assign n52689 = ( n8282 & n29391 ) | ( n8282 & ~n36193 ) | ( n29391 & ~n36193 ) ;
  assign n52690 = ( ~n31134 & n35229 ) | ( ~n31134 & n52689 ) | ( n35229 & n52689 ) ;
  assign n52691 = n52690 ^ n46244 ^ n22785 ;
  assign n52692 = n48090 ^ n29368 ^ n23632 ;
  assign n52693 = ( n4373 & ~n9910 ) | ( n4373 & n9919 ) | ( ~n9910 & n9919 ) ;
  assign n52694 = n25442 & n52693 ;
  assign n52695 = ( n13621 & n36440 ) | ( n13621 & ~n52429 ) | ( n36440 & ~n52429 ) ;
  assign n52696 = n42361 | n48500 ;
  assign n52697 = ~n10968 & n14979 ;
  assign n52698 = ~n7177 & n52697 ;
  assign n52699 = ~n1098 & n17683 ;
  assign n52700 = n52698 & n52699 ;
  assign n52703 = n48212 & n51446 ;
  assign n52704 = n22569 & n52703 ;
  assign n52701 = n45100 ^ n25173 ^ n23375 ;
  assign n52702 = ~n42793 & n52701 ;
  assign n52705 = n52704 ^ n52702 ^ 1'b0 ;
  assign n52706 = ( n9505 & n15875 ) | ( n9505 & ~n38097 ) | ( n15875 & ~n38097 ) ;
  assign n52707 = ( n5082 & n17106 ) | ( n5082 & ~n52706 ) | ( n17106 & ~n52706 ) ;
  assign n52708 = n14682 ^ n9953 ^ 1'b0 ;
  assign n52709 = ~n52707 & n52708 ;
  assign n52710 = ~n3578 & n8881 ;
  assign n52711 = n52710 ^ n1437 ^ 1'b0 ;
  assign n52712 = ( n8055 & n30523 ) | ( n8055 & ~n52711 ) | ( n30523 & ~n52711 ) ;
  assign n52713 = n29743 ^ n25815 ^ n281 ;
  assign n52714 = ( n14707 & n42361 ) | ( n14707 & n46541 ) | ( n42361 & n46541 ) ;
  assign n52715 = ( n1635 & ~n16485 ) | ( n1635 & n29111 ) | ( ~n16485 & n29111 ) ;
  assign n52716 = ( n4998 & n12161 ) | ( n4998 & n20191 ) | ( n12161 & n20191 ) ;
  assign n52717 = ( ~n24029 & n52715 ) | ( ~n24029 & n52716 ) | ( n52715 & n52716 ) ;
  assign n52722 = n37034 ^ n15736 ^ 1'b0 ;
  assign n52719 = n40194 ^ n34370 ^ 1'b0 ;
  assign n52720 = n52719 ^ n3427 ^ n2247 ;
  assign n52721 = n52720 ^ n45713 ^ n38187 ;
  assign n52718 = n25190 ^ n7762 ^ 1'b0 ;
  assign n52723 = n52722 ^ n52721 ^ n52718 ;
  assign n52724 = n19465 & n26118 ;
  assign n52725 = n20259 & n28029 ;
  assign n52726 = n12475 | n33938 ;
  assign n52727 = n9254 & ~n52726 ;
  assign n52728 = n52727 ^ n28478 ^ 1'b0 ;
  assign n52729 = n52728 ^ n26589 ^ 1'b0 ;
  assign n52730 = ~n52725 & n52729 ;
  assign n52731 = ~n29929 & n34336 ;
  assign n52732 = n1475 | n42961 ;
  assign n52733 = n52732 ^ n44551 ^ 1'b0 ;
  assign n52734 = n17735 ^ n11696 ^ 1'b0 ;
  assign n52735 = x15 & n52734 ;
  assign n52736 = ~n15996 & n52735 ;
  assign n52737 = ( ~n14745 & n42495 ) | ( ~n14745 & n52736 ) | ( n42495 & n52736 ) ;
  assign n52739 = ( n14805 & n35936 ) | ( n14805 & ~n45861 ) | ( n35936 & ~n45861 ) ;
  assign n52738 = n35328 ^ n18733 ^ 1'b0 ;
  assign n52740 = n52739 ^ n52738 ^ 1'b0 ;
  assign n52741 = n46562 ^ n40981 ^ 1'b0 ;
  assign n52742 = n11476 ^ n9531 ^ n1297 ;
  assign n52743 = n24956 ^ n2139 ^ 1'b0 ;
  assign n52744 = n735 | n7563 ;
  assign n52745 = n39756 & ~n52744 ;
  assign n52746 = n7300 ^ n7256 ^ 1'b0 ;
  assign n52747 = n12123 | n52746 ;
  assign n52748 = ~n2812 & n25589 ;
  assign n52749 = n47578 ^ n13450 ^ 1'b0 ;
  assign n52750 = n8127 | n36921 ;
  assign n52751 = n22726 ^ n5895 ^ 1'b0 ;
  assign n52752 = n47539 ^ n22188 ^ 1'b0 ;
  assign n52753 = n262 & n32636 ;
  assign n52754 = n52753 ^ n21141 ^ 1'b0 ;
  assign n52755 = ( n50415 & n52752 ) | ( n50415 & n52754 ) | ( n52752 & n52754 ) ;
  assign n52756 = n1598 & n8888 ;
  assign n52757 = n11321 & n52756 ;
  assign n52758 = n21235 & ~n50532 ;
  assign n52759 = n52758 ^ n44597 ^ 1'b0 ;
  assign n52760 = n9623 & n12024 ;
  assign n52761 = n33080 & n52760 ;
  assign n52762 = n6326 ^ n5171 ^ n2007 ;
  assign n52763 = ~n20150 & n52762 ;
  assign n52764 = n28152 & n52763 ;
  assign n52767 = ~n7187 & n14072 ;
  assign n52768 = n12702 & n52767 ;
  assign n52769 = n6823 & ~n52768 ;
  assign n52770 = ( n13518 & n20130 ) | ( n13518 & n33637 ) | ( n20130 & n33637 ) ;
  assign n52771 = n52770 ^ n23287 ^ 1'b0 ;
  assign n52772 = n52769 | n52771 ;
  assign n52765 = n14568 ^ n6368 ^ 1'b0 ;
  assign n52766 = n52765 ^ n34129 ^ n1893 ;
  assign n52773 = n52772 ^ n52766 ^ n16062 ;
  assign n52774 = n15859 & n52773 ;
  assign n52775 = ( n8813 & n30786 ) | ( n8813 & ~n51784 ) | ( n30786 & ~n51784 ) ;
  assign n52776 = n25971 ^ n20550 ^ 1'b0 ;
  assign n52777 = n6312 & n52776 ;
  assign n52778 = n52777 ^ n37987 ^ 1'b0 ;
  assign n52779 = ( ~n10835 & n25848 ) | ( ~n10835 & n52778 ) | ( n25848 & n52778 ) ;
  assign n52780 = n24408 ^ n11977 ^ 1'b0 ;
  assign n52781 = n30178 ^ n4826 ^ 1'b0 ;
  assign n52782 = ( n7364 & n50615 ) | ( n7364 & ~n52781 ) | ( n50615 & ~n52781 ) ;
  assign n52783 = n15818 ^ n7173 ^ n358 ;
  assign n52784 = ( n9238 & n15021 ) | ( n9238 & n33944 ) | ( n15021 & n33944 ) ;
  assign n52785 = ~n34148 & n52784 ;
  assign n52786 = ~n52783 & n52785 ;
  assign n52787 = n7698 & ~n51801 ;
  assign n52788 = n5597 ^ n5440 ^ 1'b0 ;
  assign n52789 = n19428 & n52788 ;
  assign n52790 = n52789 ^ n6788 ^ 1'b0 ;
  assign n52791 = n34936 ^ n10045 ^ 1'b0 ;
  assign n52792 = n22226 & ~n52791 ;
  assign n52793 = n12421 ^ x1 ^ 1'b0 ;
  assign n52794 = n29432 | n41752 ;
  assign n52795 = ( ~n4720 & n28773 ) | ( ~n4720 & n34443 ) | ( n28773 & n34443 ) ;
  assign n52796 = n28792 & n41393 ;
  assign n52797 = n42841 ^ n13256 ^ 1'b0 ;
  assign n52798 = n40777 ^ n22310 ^ n4977 ;
  assign n52799 = ( n13034 & n20999 ) | ( n13034 & ~n52179 ) | ( n20999 & ~n52179 ) ;
  assign n52800 = n18218 ^ n6331 ^ 1'b0 ;
  assign n52801 = n29002 | n52800 ;
  assign n52802 = n16999 | n43468 ;
  assign n52803 = n52802 ^ n41091 ^ 1'b0 ;
  assign n52804 = n11901 ^ n11043 ^ 1'b0 ;
  assign n52805 = n39893 ^ n25576 ^ n21878 ;
  assign n52806 = n52805 ^ n45531 ^ n19313 ;
  assign n52807 = ~n9593 & n52806 ;
  assign n52808 = n34181 ^ n20384 ^ n9274 ;
  assign n52809 = n30931 ^ n11687 ^ 1'b0 ;
  assign n52810 = n52809 ^ n15394 ^ n551 ;
  assign n52811 = n52810 ^ n6101 ^ 1'b0 ;
  assign n52812 = n52811 ^ n51468 ^ 1'b0 ;
  assign n52813 = n8410 & n16940 ;
  assign n52814 = n52813 ^ n22675 ^ n13748 ;
  assign n52815 = n10166 | n23974 ;
  assign n52816 = n52815 ^ n4383 ^ 1'b0 ;
  assign n52817 = n52816 ^ n41631 ^ n8964 ;
  assign n52818 = n13667 | n39337 ;
  assign n52819 = n52818 ^ n42788 ^ 1'b0 ;
  assign n52820 = n52819 ^ n23618 ^ n22643 ;
  assign n52821 = n39575 & n52820 ;
  assign n52822 = n52817 & n52821 ;
  assign n52823 = n27491 ^ n5408 ^ 1'b0 ;
  assign n52824 = n25259 ^ n17216 ^ 1'b0 ;
  assign n52825 = ~n27009 & n52824 ;
  assign n52826 = n3306 & n52825 ;
  assign n52827 = n52823 & n52826 ;
  assign n52828 = n41233 ^ n31304 ^ n2974 ;
  assign n52829 = n5289 | n52828 ;
  assign n52830 = n4085 & ~n52829 ;
  assign n52831 = ~n22871 & n43393 ;
  assign n52832 = n21707 & ~n26106 ;
  assign n52833 = n52832 ^ n6562 ^ 1'b0 ;
  assign n52834 = ( n22674 & n34395 ) | ( n22674 & ~n52833 ) | ( n34395 & ~n52833 ) ;
  assign n52835 = n11860 ^ n3082 ^ 1'b0 ;
  assign n52836 = n52835 ^ n47151 ^ 1'b0 ;
  assign n52837 = n16302 & n29071 ;
  assign n52838 = ~n13731 & n52837 ;
  assign n52839 = n52838 ^ n29431 ^ n20794 ;
  assign n52840 = ~n15415 & n49238 ;
  assign n52841 = n52840 ^ x116 ^ 1'b0 ;
  assign n52842 = ( ~n25108 & n50268 ) | ( ~n25108 & n52841 ) | ( n50268 & n52841 ) ;
  assign n52843 = n31980 ^ n27643 ^ n11868 ;
  assign n52844 = n1199 | n14530 ;
  assign n52845 = n27457 | n52844 ;
  assign y0 = x9 ;
  assign y1 = x10 ;
  assign y2 = x11 ;
  assign y3 = x13 ;
  assign y4 = x18 ;
  assign y5 = x20 ;
  assign y6 = x29 ;
  assign y7 = x38 ;
  assign y8 = x43 ;
  assign y9 = x60 ;
  assign y10 = x62 ;
  assign y11 = x67 ;
  assign y12 = x69 ;
  assign y13 = x70 ;
  assign y14 = x71 ;
  assign y15 = x80 ;
  assign y16 = x88 ;
  assign y17 = x91 ;
  assign y18 = x92 ;
  assign y19 = x96 ;
  assign y20 = x101 ;
  assign y21 = x102 ;
  assign y22 = x124 ;
  assign y23 = x125 ;
  assign y24 = x135 ;
  assign y25 = x136 ;
  assign y26 = x146 ;
  assign y27 = x150 ;
  assign y28 = x154 ;
  assign y29 = x160 ;
  assign y30 = x167 ;
  assign y31 = x172 ;
  assign y32 = x175 ;
  assign y33 = x176 ;
  assign y34 = x188 ;
  assign y35 = x200 ;
  assign y36 = x210 ;
  assign y37 = x218 ;
  assign y38 = x219 ;
  assign y39 = x224 ;
  assign y40 = x226 ;
  assign y41 = x231 ;
  assign y42 = x233 ;
  assign y43 = x242 ;
  assign y44 = x244 ;
  assign y45 = x245 ;
  assign y46 = x246 ;
  assign y47 = x247 ;
  assign y48 = n256 ;
  assign y49 = n257 ;
  assign y50 = ~n258 ;
  assign y51 = ~n259 ;
  assign y52 = ~1'b0 ;
  assign y53 = ~1'b0 ;
  assign y54 = ~n261 ;
  assign y55 = ~n262 ;
  assign y56 = n264 ;
  assign y57 = n266 ;
  assign y58 = ~n268 ;
  assign y59 = n269 ;
  assign y60 = ~n271 ;
  assign y61 = ~1'b0 ;
  assign y62 = ~n272 ;
  assign y63 = ~n276 ;
  assign y64 = ~n279 ;
  assign y65 = ~n280 ;
  assign y66 = n282 ;
  assign y67 = n285 ;
  assign y68 = ~n287 ;
  assign y69 = ~n289 ;
  assign y70 = n290 ;
  assign y71 = ~1'b0 ;
  assign y72 = n291 ;
  assign y73 = n293 ;
  assign y74 = n294 ;
  assign y75 = ~n299 ;
  assign y76 = ~n301 ;
  assign y77 = ~n305 ;
  assign y78 = n306 ;
  assign y79 = ~1'b0 ;
  assign y80 = n307 ;
  assign y81 = n310 ;
  assign y82 = n313 ;
  assign y83 = ~n318 ;
  assign y84 = ~1'b0 ;
  assign y85 = n321 ;
  assign y86 = ~n322 ;
  assign y87 = ~n325 ;
  assign y88 = n327 ;
  assign y89 = n332 ;
  assign y90 = n333 ;
  assign y91 = ~1'b0 ;
  assign y92 = n335 ;
  assign y93 = n336 ;
  assign y94 = n337 ;
  assign y95 = ~n340 ;
  assign y96 = n341 ;
  assign y97 = n345 ;
  assign y98 = ~n346 ;
  assign y99 = n348 ;
  assign y100 = n353 ;
  assign y101 = ~1'b0 ;
  assign y102 = ~n354 ;
  assign y103 = n355 ;
  assign y104 = ~1'b0 ;
  assign y105 = ~n361 ;
  assign y106 = n365 ;
  assign y107 = ~n370 ;
  assign y108 = ~n372 ;
  assign y109 = n373 ;
  assign y110 = ~1'b0 ;
  assign y111 = ~1'b0 ;
  assign y112 = ~1'b0 ;
  assign y113 = ~n379 ;
  assign y114 = n382 ;
  assign y115 = ~n384 ;
  assign y116 = ~n386 ;
  assign y117 = n389 ;
  assign y118 = n391 ;
  assign y119 = n392 ;
  assign y120 = n393 ;
  assign y121 = ~n396 ;
  assign y122 = ~n398 ;
  assign y123 = ~n402 ;
  assign y124 = ~1'b0 ;
  assign y125 = n404 ;
  assign y126 = n405 ;
  assign y127 = ~n409 ;
  assign y128 = ~n421 ;
  assign y129 = ~n423 ;
  assign y130 = n426 ;
  assign y131 = ~1'b0 ;
  assign y132 = ~n429 ;
  assign y133 = n434 ;
  assign y134 = n435 ;
  assign y135 = n436 ;
  assign y136 = ~1'b0 ;
  assign y137 = n438 ;
  assign y138 = ~n445 ;
  assign y139 = ~n447 ;
  assign y140 = n450 ;
  assign y141 = ~n457 ;
  assign y142 = ~1'b0 ;
  assign y143 = n459 ;
  assign y144 = ~n469 ;
  assign y145 = ~n470 ;
  assign y146 = ~n473 ;
  assign y147 = n479 ;
  assign y148 = ~1'b0 ;
  assign y149 = n480 ;
  assign y150 = ~1'b0 ;
  assign y151 = ~n483 ;
  assign y152 = ~n487 ;
  assign y153 = n488 ;
  assign y154 = n500 ;
  assign y155 = ~1'b0 ;
  assign y156 = n511 ;
  assign y157 = ~n512 ;
  assign y158 = ~1'b0 ;
  assign y159 = ~1'b0 ;
  assign y160 = n515 ;
  assign y161 = ~n518 ;
  assign y162 = ~1'b0 ;
  assign y163 = n520 ;
  assign y164 = n524 ;
  assign y165 = ~n530 ;
  assign y166 = n534 ;
  assign y167 = x207 ;
  assign y168 = ~n536 ;
  assign y169 = ~1'b0 ;
  assign y170 = ~n543 ;
  assign y171 = ~x5 ;
  assign y172 = n544 ;
  assign y173 = ~n553 ;
  assign y174 = ~n554 ;
  assign y175 = ~n555 ;
  assign y176 = n558 ;
  assign y177 = n561 ;
  assign y178 = ~n564 ;
  assign y179 = n568 ;
  assign y180 = n574 ;
  assign y181 = ~n577 ;
  assign y182 = ~n581 ;
  assign y183 = ~n583 ;
  assign y184 = ~n586 ;
  assign y185 = ~n602 ;
  assign y186 = ~n607 ;
  assign y187 = ~1'b0 ;
  assign y188 = n614 ;
  assign y189 = n616 ;
  assign y190 = n618 ;
  assign y191 = ~n632 ;
  assign y192 = ~n642 ;
  assign y193 = ~n645 ;
  assign y194 = n656 ;
  assign y195 = ~n657 ;
  assign y196 = ~1'b0 ;
  assign y197 = ~n660 ;
  assign y198 = n666 ;
  assign y199 = ~1'b0 ;
  assign y200 = n668 ;
  assign y201 = ~n669 ;
  assign y202 = ~n673 ;
  assign y203 = ~n678 ;
  assign y204 = ~n681 ;
  assign y205 = ~n686 ;
  assign y206 = ~n687 ;
  assign y207 = ~n688 ;
  assign y208 = ~n689 ;
  assign y209 = ~n693 ;
  assign y210 = n709 ;
  assign y211 = ~n713 ;
  assign y212 = ~n720 ;
  assign y213 = n725 ;
  assign y214 = n728 ;
  assign y215 = ~n732 ;
  assign y216 = ~n733 ;
  assign y217 = ~1'b0 ;
  assign y218 = n738 ;
  assign y219 = n749 ;
  assign y220 = ~n751 ;
  assign y221 = ~1'b0 ;
  assign y222 = ~x81 ;
  assign y223 = n755 ;
  assign y224 = n756 ;
  assign y225 = ~n757 ;
  assign y226 = ~n763 ;
  assign y227 = ~1'b0 ;
  assign y228 = n769 ;
  assign y229 = ~n771 ;
  assign y230 = ~n773 ;
  assign y231 = ~n785 ;
  assign y232 = ~n284 ;
  assign y233 = ~n793 ;
  assign y234 = ~n799 ;
  assign y235 = n800 ;
  assign y236 = ~n802 ;
  assign y237 = ~n806 ;
  assign y238 = ~n807 ;
  assign y239 = n809 ;
  assign y240 = n816 ;
  assign y241 = n821 ;
  assign y242 = ~1'b0 ;
  assign y243 = ~n827 ;
  assign y244 = n829 ;
  assign y245 = ~1'b0 ;
  assign y246 = ~n834 ;
  assign y247 = ~n840 ;
  assign y248 = ~n843 ;
  assign y249 = ~n845 ;
  assign y250 = n851 ;
  assign y251 = n853 ;
  assign y252 = ~n855 ;
  assign y253 = ~n863 ;
  assign y254 = n864 ;
  assign y255 = ~1'b0 ;
  assign y256 = n865 ;
  assign y257 = ~n869 ;
  assign y258 = ~n871 ;
  assign y259 = n872 ;
  assign y260 = ~n873 ;
  assign y261 = n875 ;
  assign y262 = ~n883 ;
  assign y263 = n889 ;
  assign y264 = ~n891 ;
  assign y265 = n893 ;
  assign y266 = ~n894 ;
  assign y267 = n903 ;
  assign y268 = ~n905 ;
  assign y269 = n912 ;
  assign y270 = ~n921 ;
  assign y271 = ~n925 ;
  assign y272 = ~n930 ;
  assign y273 = ~1'b0 ;
  assign y274 = n936 ;
  assign y275 = n939 ;
  assign y276 = n940 ;
  assign y277 = n941 ;
  assign y278 = ~n943 ;
  assign y279 = ~n950 ;
  assign y280 = ~n951 ;
  assign y281 = n955 ;
  assign y282 = ~n964 ;
  assign y283 = ~1'b0 ;
  assign y284 = n966 ;
  assign y285 = ~n967 ;
  assign y286 = n979 ;
  assign y287 = n983 ;
  assign y288 = n984 ;
  assign y289 = n989 ;
  assign y290 = ~n993 ;
  assign y291 = ~n995 ;
  assign y292 = n998 ;
  assign y293 = ~n1001 ;
  assign y294 = ~1'b0 ;
  assign y295 = 1'b0 ;
  assign y296 = ~n1009 ;
  assign y297 = ~n1014 ;
  assign y298 = ~n905 ;
  assign y299 = n1018 ;
  assign y300 = ~1'b0 ;
  assign y301 = ~1'b0 ;
  assign y302 = ~n1029 ;
  assign y303 = ~1'b0 ;
  assign y304 = n1034 ;
  assign y305 = ~n1036 ;
  assign y306 = ~n1040 ;
  assign y307 = n1042 ;
  assign y308 = n1046 ;
  assign y309 = ~n1047 ;
  assign y310 = ~n1049 ;
  assign y311 = ~n1050 ;
  assign y312 = n1052 ;
  assign y313 = ~n1053 ;
  assign y314 = n1063 ;
  assign y315 = ~n1068 ;
  assign y316 = n1077 ;
  assign y317 = ~n1087 ;
  assign y318 = ~n1092 ;
  assign y319 = ~n1106 ;
  assign y320 = ~1'b0 ;
  assign y321 = ~1'b0 ;
  assign y322 = n1108 ;
  assign y323 = ~1'b0 ;
  assign y324 = ~n1111 ;
  assign y325 = n1112 ;
  assign y326 = n1114 ;
  assign y327 = ~n1118 ;
  assign y328 = ~n1120 ;
  assign y329 = ~n1125 ;
  assign y330 = ~n1130 ;
  assign y331 = n1133 ;
  assign y332 = n1136 ;
  assign y333 = ~n1148 ;
  assign y334 = ~n1149 ;
  assign y335 = ~n1150 ;
  assign y336 = n1153 ;
  assign y337 = n1158 ;
  assign y338 = ~n1159 ;
  assign y339 = ~n1162 ;
  assign y340 = n1169 ;
  assign y341 = ~n1180 ;
  assign y342 = ~n1183 ;
  assign y343 = ~n1184 ;
  assign y344 = ~n1186 ;
  assign y345 = ~n1187 ;
  assign y346 = n1198 ;
  assign y347 = ~n1199 ;
  assign y348 = n1204 ;
  assign y349 = ~1'b0 ;
  assign y350 = n1208 ;
  assign y351 = n1212 ;
  assign y352 = n1218 ;
  assign y353 = n1223 ;
  assign y354 = n1228 ;
  assign y355 = ~n1235 ;
  assign y356 = ~n1236 ;
  assign y357 = ~n1240 ;
  assign y358 = ~n1241 ;
  assign y359 = ~n331 ;
  assign y360 = n1243 ;
  assign y361 = ~n1247 ;
  assign y362 = ~n1249 ;
  assign y363 = ~1'b0 ;
  assign y364 = n1251 ;
  assign y365 = ~1'b0 ;
  assign y366 = n1255 ;
  assign y367 = n1256 ;
  assign y368 = ~n1258 ;
  assign y369 = n1264 ;
  assign y370 = n1266 ;
  assign y371 = n1270 ;
  assign y372 = n1274 ;
  assign y373 = n1279 ;
  assign y374 = n1287 ;
  assign y375 = n1292 ;
  assign y376 = ~n1296 ;
  assign y377 = ~n1297 ;
  assign y378 = ~n1303 ;
  assign y379 = ~1'b0 ;
  assign y380 = n290 ;
  assign y381 = n1308 ;
  assign y382 = ~n1311 ;
  assign y383 = ~n1314 ;
  assign y384 = ~n1317 ;
  assign y385 = n1323 ;
  assign y386 = n1324 ;
  assign y387 = ~n1325 ;
  assign y388 = n1328 ;
  assign y389 = ~1'b0 ;
  assign y390 = ~n1331 ;
  assign y391 = ~n1342 ;
  assign y392 = ~1'b0 ;
  assign y393 = ~n1346 ;
  assign y394 = ~n1348 ;
  assign y395 = n1349 ;
  assign y396 = ~1'b0 ;
  assign y397 = ~n1351 ;
  assign y398 = n1354 ;
  assign y399 = ~n1355 ;
  assign y400 = ~1'b0 ;
  assign y401 = ~1'b0 ;
  assign y402 = ~n1362 ;
  assign y403 = ~1'b0 ;
  assign y404 = n1365 ;
  assign y405 = n1370 ;
  assign y406 = ~1'b0 ;
  assign y407 = ~n1372 ;
  assign y408 = ~n1379 ;
  assign y409 = ~1'b0 ;
  assign y410 = ~n1383 ;
  assign y411 = ~1'b0 ;
  assign y412 = n1384 ;
  assign y413 = n1387 ;
  assign y414 = ~n1388 ;
  assign y415 = n1392 ;
  assign y416 = ~n1396 ;
  assign y417 = ~n1401 ;
  assign y418 = ~n1408 ;
  assign y419 = ~n1410 ;
  assign y420 = ~1'b0 ;
  assign y421 = ~n1412 ;
  assign y422 = ~n1417 ;
  assign y423 = ~n1423 ;
  assign y424 = ~n1429 ;
  assign y425 = n1443 ;
  assign y426 = ~n1444 ;
  assign y427 = n1451 ;
  assign y428 = n1458 ;
  assign y429 = ~1'b0 ;
  assign y430 = ~n1467 ;
  assign y431 = n1468 ;
  assign y432 = ~1'b0 ;
  assign y433 = ~1'b0 ;
  assign y434 = ~n1470 ;
  assign y435 = ~n1475 ;
  assign y436 = ~n1477 ;
  assign y437 = n1483 ;
  assign y438 = n1484 ;
  assign y439 = n1489 ;
  assign y440 = ~n1496 ;
  assign y441 = ~n1499 ;
  assign y442 = ~n1505 ;
  assign y443 = ~n1513 ;
  assign y444 = n1518 ;
  assign y445 = ~1'b0 ;
  assign y446 = ~1'b0 ;
  assign y447 = n1524 ;
  assign y448 = ~1'b0 ;
  assign y449 = n1529 ;
  assign y450 = n1533 ;
  assign y451 = ~n1541 ;
  assign y452 = ~n1551 ;
  assign y453 = n1552 ;
  assign y454 = ~n1555 ;
  assign y455 = ~n1557 ;
  assign y456 = ~1'b0 ;
  assign y457 = n1558 ;
  assign y458 = ~n1567 ;
  assign y459 = n1568 ;
  assign y460 = ~1'b0 ;
  assign y461 = ~1'b0 ;
  assign y462 = n1573 ;
  assign y463 = ~n1578 ;
  assign y464 = n1580 ;
  assign y465 = n1581 ;
  assign y466 = n1583 ;
  assign y467 = n1598 ;
  assign y468 = n1601 ;
  assign y469 = ~1'b0 ;
  assign y470 = ~1'b0 ;
  assign y471 = ~n1608 ;
  assign y472 = ~n1619 ;
  assign y473 = ~1'b0 ;
  assign y474 = n1622 ;
  assign y475 = n1623 ;
  assign y476 = ~n1634 ;
  assign y477 = ~n1637 ;
  assign y478 = n1639 ;
  assign y479 = ~n1641 ;
  assign y480 = ~n1643 ;
  assign y481 = ~1'b0 ;
  assign y482 = ~n1645 ;
  assign y483 = n1654 ;
  assign y484 = ~1'b0 ;
  assign y485 = ~n1659 ;
  assign y486 = ~n1660 ;
  assign y487 = n1662 ;
  assign y488 = ~n1663 ;
  assign y489 = n1667 ;
  assign y490 = ~n1673 ;
  assign y491 = ~n1674 ;
  assign y492 = ~1'b0 ;
  assign y493 = n1675 ;
  assign y494 = n1676 ;
  assign y495 = n1678 ;
  assign y496 = ~n1685 ;
  assign y497 = ~n1687 ;
  assign y498 = ~n1688 ;
  assign y499 = ~n1695 ;
  assign y500 = n1698 ;
  assign y501 = ~n1704 ;
  assign y502 = ~n1709 ;
  assign y503 = n1710 ;
  assign y504 = ~1'b0 ;
  assign y505 = ~n1720 ;
  assign y506 = ~n1721 ;
  assign y507 = ~1'b0 ;
  assign y508 = n1730 ;
  assign y509 = ~1'b0 ;
  assign y510 = n1735 ;
  assign y511 = ~n1738 ;
  assign y512 = n1739 ;
  assign y513 = ~n1742 ;
  assign y514 = ~n1744 ;
  assign y515 = ~1'b0 ;
  assign y516 = ~1'b0 ;
  assign y517 = ~n1752 ;
  assign y518 = ~n1753 ;
  assign y519 = ~1'b0 ;
  assign y520 = n1758 ;
  assign y521 = ~n1771 ;
  assign y522 = ~1'b0 ;
  assign y523 = n1775 ;
  assign y524 = ~n1776 ;
  assign y525 = n1786 ;
  assign y526 = ~1'b0 ;
  assign y527 = ~1'b0 ;
  assign y528 = ~n1789 ;
  assign y529 = ~n1796 ;
  assign y530 = ~n1800 ;
  assign y531 = n1802 ;
  assign y532 = n1807 ;
  assign y533 = n1813 ;
  assign y534 = n1828 ;
  assign y535 = ~1'b0 ;
  assign y536 = n1838 ;
  assign y537 = n1840 ;
  assign y538 = n1843 ;
  assign y539 = ~n1845 ;
  assign y540 = ~n1852 ;
  assign y541 = ~n1857 ;
  assign y542 = ~1'b0 ;
  assign y543 = n1866 ;
  assign y544 = ~1'b0 ;
  assign y545 = n1874 ;
  assign y546 = n1877 ;
  assign y547 = n1881 ;
  assign y548 = ~n1883 ;
  assign y549 = ~n1884 ;
  assign y550 = n1886 ;
  assign y551 = ~1'b0 ;
  assign y552 = ~n1889 ;
  assign y553 = ~1'b0 ;
  assign y554 = ~n1891 ;
  assign y555 = ~1'b0 ;
  assign y556 = ~n1894 ;
  assign y557 = ~n1898 ;
  assign y558 = ~1'b0 ;
  assign y559 = n1901 ;
  assign y560 = ~n1904 ;
  assign y561 = ~1'b0 ;
  assign y562 = ~n1909 ;
  assign y563 = n1917 ;
  assign y564 = n1921 ;
  assign y565 = ~n1933 ;
  assign y566 = ~1'b0 ;
  assign y567 = ~n1935 ;
  assign y568 = ~n1943 ;
  assign y569 = ~n1947 ;
  assign y570 = ~1'b0 ;
  assign y571 = n1950 ;
  assign y572 = ~n1952 ;
  assign y573 = ~1'b0 ;
  assign y574 = ~1'b0 ;
  assign y575 = n1956 ;
  assign y576 = n1958 ;
  assign y577 = n1959 ;
  assign y578 = n1964 ;
  assign y579 = ~1'b0 ;
  assign y580 = n1973 ;
  assign y581 = ~n1974 ;
  assign y582 = ~1'b0 ;
  assign y583 = ~n1981 ;
  assign y584 = ~n1998 ;
  assign y585 = ~n2000 ;
  assign y586 = n2006 ;
  assign y587 = n2007 ;
  assign y588 = ~1'b0 ;
  assign y589 = ~n2009 ;
  assign y590 = ~1'b0 ;
  assign y591 = ~n2016 ;
  assign y592 = ~1'b0 ;
  assign y593 = ~n1916 ;
  assign y594 = n2020 ;
  assign y595 = ~1'b0 ;
  assign y596 = ~n2028 ;
  assign y597 = n2030 ;
  assign y598 = ~n2038 ;
  assign y599 = n2041 ;
  assign y600 = n1524 ;
  assign y601 = ~1'b0 ;
  assign y602 = ~1'b0 ;
  assign y603 = n2047 ;
  assign y604 = n1438 ;
  assign y605 = n2048 ;
  assign y606 = n2049 ;
  assign y607 = ~1'b0 ;
  assign y608 = n2052 ;
  assign y609 = ~1'b0 ;
  assign y610 = n2056 ;
  assign y611 = ~n2062 ;
  assign y612 = ~1'b0 ;
  assign y613 = ~n2063 ;
  assign y614 = n2070 ;
  assign y615 = ~n2082 ;
  assign y616 = n2085 ;
  assign y617 = ~1'b0 ;
  assign y618 = ~n2094 ;
  assign y619 = n2096 ;
  assign y620 = n2104 ;
  assign y621 = ~n2105 ;
  assign y622 = n2106 ;
  assign y623 = n2110 ;
  assign y624 = ~n2124 ;
  assign y625 = ~n2130 ;
  assign y626 = n2131 ;
  assign y627 = n2140 ;
  assign y628 = ~n2142 ;
  assign y629 = n2155 ;
  assign y630 = n2158 ;
  assign y631 = ~n2163 ;
  assign y632 = n2164 ;
  assign y633 = ~n2167 ;
  assign y634 = ~1'b0 ;
  assign y635 = n2170 ;
  assign y636 = n2175 ;
  assign y637 = ~1'b0 ;
  assign y638 = 1'b0 ;
  assign y639 = ~1'b0 ;
  assign y640 = ~n2177 ;
  assign y641 = ~n2192 ;
  assign y642 = n2194 ;
  assign y643 = ~n2197 ;
  assign y644 = n2201 ;
  assign y645 = ~n2205 ;
  assign y646 = ~1'b0 ;
  assign y647 = ~n2208 ;
  assign y648 = n2211 ;
  assign y649 = ~n2226 ;
  assign y650 = ~n2232 ;
  assign y651 = ~n2233 ;
  assign y652 = n2247 ;
  assign y653 = ~1'b0 ;
  assign y654 = ~1'b0 ;
  assign y655 = ~n2249 ;
  assign y656 = ~n2254 ;
  assign y657 = n2261 ;
  assign y658 = n2263 ;
  assign y659 = ~n2267 ;
  assign y660 = n2268 ;
  assign y661 = ~n2273 ;
  assign y662 = n2276 ;
  assign y663 = n2281 ;
  assign y664 = n2282 ;
  assign y665 = n2283 ;
  assign y666 = n2295 ;
  assign y667 = ~n2303 ;
  assign y668 = ~n2308 ;
  assign y669 = n2310 ;
  assign y670 = ~n2322 ;
  assign y671 = n2330 ;
  assign y672 = n2338 ;
  assign y673 = ~n2339 ;
  assign y674 = ~n2349 ;
  assign y675 = ~n2356 ;
  assign y676 = ~n2359 ;
  assign y677 = ~n2364 ;
  assign y678 = n2372 ;
  assign y679 = ~n2379 ;
  assign y680 = ~1'b0 ;
  assign y681 = n2380 ;
  assign y682 = n2384 ;
  assign y683 = n2386 ;
  assign y684 = ~n2388 ;
  assign y685 = ~1'b0 ;
  assign y686 = ~n2389 ;
  assign y687 = n2390 ;
  assign y688 = n2401 ;
  assign y689 = n2409 ;
  assign y690 = ~n2415 ;
  assign y691 = ~n2417 ;
  assign y692 = n2419 ;
  assign y693 = n2421 ;
  assign y694 = 1'b0 ;
  assign y695 = n2427 ;
  assign y696 = ~1'b0 ;
  assign y697 = ~n1873 ;
  assign y698 = n2430 ;
  assign y699 = ~n2445 ;
  assign y700 = ~n2447 ;
  assign y701 = n2448 ;
  assign y702 = n2456 ;
  assign y703 = n2460 ;
  assign y704 = ~n2469 ;
  assign y705 = ~1'b0 ;
  assign y706 = ~n2476 ;
  assign y707 = n2479 ;
  assign y708 = n2481 ;
  assign y709 = ~n2494 ;
  assign y710 = ~n2498 ;
  assign y711 = n2500 ;
  assign y712 = n2502 ;
  assign y713 = n2506 ;
  assign y714 = n2508 ;
  assign y715 = ~n2509 ;
  assign y716 = ~1'b0 ;
  assign y717 = n2512 ;
  assign y718 = ~n2515 ;
  assign y719 = ~n1475 ;
  assign y720 = ~n2517 ;
  assign y721 = ~n2518 ;
  assign y722 = n2520 ;
  assign y723 = n2530 ;
  assign y724 = ~n2536 ;
  assign y725 = ~n2557 ;
  assign y726 = ~1'b0 ;
  assign y727 = ~n2561 ;
  assign y728 = ~1'b0 ;
  assign y729 = n2562 ;
  assign y730 = ~1'b0 ;
  assign y731 = ~n2565 ;
  assign y732 = n2575 ;
  assign y733 = n2576 ;
  assign y734 = ~n2582 ;
  assign y735 = n2585 ;
  assign y736 = n2594 ;
  assign y737 = n2597 ;
  assign y738 = n2601 ;
  assign y739 = ~n2602 ;
  assign y740 = n2611 ;
  assign y741 = ~n2613 ;
  assign y742 = ~1'b0 ;
  assign y743 = ~n2614 ;
  assign y744 = n2615 ;
  assign y745 = n2616 ;
  assign y746 = n2620 ;
  assign y747 = n2624 ;
  assign y748 = ~n2631 ;
  assign y749 = n2634 ;
  assign y750 = ~n2637 ;
  assign y751 = n2639 ;
  assign y752 = n2642 ;
  assign y753 = ~n2646 ;
  assign y754 = n2651 ;
  assign y755 = n2655 ;
  assign y756 = n2662 ;
  assign y757 = ~1'b0 ;
  assign y758 = n2663 ;
  assign y759 = ~n2666 ;
  assign y760 = n2672 ;
  assign y761 = ~n2673 ;
  assign y762 = n2675 ;
  assign y763 = ~1'b0 ;
  assign y764 = ~n2676 ;
  assign y765 = ~1'b0 ;
  assign y766 = n2679 ;
  assign y767 = n2683 ;
  assign y768 = n2688 ;
  assign y769 = ~n2691 ;
  assign y770 = n2693 ;
  assign y771 = n2695 ;
  assign y772 = ~1'b0 ;
  assign y773 = n2699 ;
  assign y774 = ~n2704 ;
  assign y775 = n2712 ;
  assign y776 = ~n2716 ;
  assign y777 = ~1'b0 ;
  assign y778 = ~n2719 ;
  assign y779 = ~n2721 ;
  assign y780 = ~n2722 ;
  assign y781 = n2726 ;
  assign y782 = ~n2730 ;
  assign y783 = ~n2732 ;
  assign y784 = n2733 ;
  assign y785 = ~n2735 ;
  assign y786 = ~n2741 ;
  assign y787 = n2744 ;
  assign y788 = ~n2745 ;
  assign y789 = ~n2748 ;
  assign y790 = ~1'b0 ;
  assign y791 = n2753 ;
  assign y792 = ~n2755 ;
  assign y793 = ~n2760 ;
  assign y794 = n2766 ;
  assign y795 = ~n2768 ;
  assign y796 = ~n2771 ;
  assign y797 = n2775 ;
  assign y798 = ~1'b0 ;
  assign y799 = ~n2782 ;
  assign y800 = ~n2794 ;
  assign y801 = ~n426 ;
  assign y802 = ~n2800 ;
  assign y803 = ~n2805 ;
  assign y804 = n2807 ;
  assign y805 = ~n2808 ;
  assign y806 = ~1'b0 ;
  assign y807 = n2814 ;
  assign y808 = n2815 ;
  assign y809 = ~n2818 ;
  assign y810 = n2822 ;
  assign y811 = n2824 ;
  assign y812 = n2834 ;
  assign y813 = ~1'b0 ;
  assign y814 = ~n2835 ;
  assign y815 = n2836 ;
  assign y816 = ~n2838 ;
  assign y817 = n2849 ;
  assign y818 = n2854 ;
  assign y819 = ~n2862 ;
  assign y820 = ~1'b0 ;
  assign y821 = ~n2867 ;
  assign y822 = n2869 ;
  assign y823 = ~1'b0 ;
  assign y824 = ~n2870 ;
  assign y825 = ~n2871 ;
  assign y826 = ~n2872 ;
  assign y827 = n2887 ;
  assign y828 = ~n2889 ;
  assign y829 = n2892 ;
  assign y830 = ~n2897 ;
  assign y831 = n2901 ;
  assign y832 = 1'b0 ;
  assign y833 = n2908 ;
  assign y834 = n2917 ;
  assign y835 = ~1'b0 ;
  assign y836 = ~n2919 ;
  assign y837 = n2921 ;
  assign y838 = ~n2929 ;
  assign y839 = ~n2935 ;
  assign y840 = ~n2937 ;
  assign y841 = ~n2946 ;
  assign y842 = ~n2947 ;
  assign y843 = ~n2949 ;
  assign y844 = ~n2965 ;
  assign y845 = n2967 ;
  assign y846 = n2971 ;
  assign y847 = n2972 ;
  assign y848 = ~1'b0 ;
  assign y849 = ~n2975 ;
  assign y850 = n2977 ;
  assign y851 = ~1'b0 ;
  assign y852 = n2978 ;
  assign y853 = ~n2983 ;
  assign y854 = n2985 ;
  assign y855 = ~n2986 ;
  assign y856 = ~n2987 ;
  assign y857 = n2993 ;
  assign y858 = n2997 ;
  assign y859 = ~n3001 ;
  assign y860 = ~n3003 ;
  assign y861 = ~1'b0 ;
  assign y862 = n3004 ;
  assign y863 = n3010 ;
  assign y864 = ~1'b0 ;
  assign y865 = ~n3012 ;
  assign y866 = ~n3013 ;
  assign y867 = ~n1953 ;
  assign y868 = ~n3016 ;
  assign y869 = ~n3022 ;
  assign y870 = ~n3023 ;
  assign y871 = ~n3027 ;
  assign y872 = n3031 ;
  assign y873 = n3033 ;
  assign y874 = n3037 ;
  assign y875 = ~1'b0 ;
  assign y876 = n3038 ;
  assign y877 = n3055 ;
  assign y878 = ~n3059 ;
  assign y879 = n3060 ;
  assign y880 = ~1'b0 ;
  assign y881 = n3063 ;
  assign y882 = ~n3069 ;
  assign y883 = n3070 ;
  assign y884 = ~n3075 ;
  assign y885 = n3077 ;
  assign y886 = ~1'b0 ;
  assign y887 = n637 ;
  assign y888 = ~n3083 ;
  assign y889 = n3085 ;
  assign y890 = n855 ;
  assign y891 = ~n1284 ;
  assign y892 = n3089 ;
  assign y893 = n3091 ;
  assign y894 = n3093 ;
  assign y895 = n3094 ;
  assign y896 = n3096 ;
  assign y897 = ~n3100 ;
  assign y898 = ~n3103 ;
  assign y899 = n3106 ;
  assign y900 = ~n3107 ;
  assign y901 = n3110 ;
  assign y902 = ~1'b0 ;
  assign y903 = ~n3113 ;
  assign y904 = n3120 ;
  assign y905 = n3121 ;
  assign y906 = ~n3133 ;
  assign y907 = 1'b0 ;
  assign y908 = n3135 ;
  assign y909 = ~n3136 ;
  assign y910 = n3138 ;
  assign y911 = n3142 ;
  assign y912 = n3146 ;
  assign y913 = n3147 ;
  assign y914 = ~n3159 ;
  assign y915 = ~n3161 ;
  assign y916 = ~n3170 ;
  assign y917 = ~n3171 ;
  assign y918 = n3173 ;
  assign y919 = ~n3177 ;
  assign y920 = ~1'b0 ;
  assign y921 = ~n3197 ;
  assign y922 = n3204 ;
  assign y923 = ~1'b0 ;
  assign y924 = n3209 ;
  assign y925 = ~n3210 ;
  assign y926 = ~n3212 ;
  assign y927 = ~1'b0 ;
  assign y928 = ~n3219 ;
  assign y929 = n3223 ;
  assign y930 = n3225 ;
  assign y931 = ~1'b0 ;
  assign y932 = ~n3227 ;
  assign y933 = n3230 ;
  assign y934 = n3231 ;
  assign y935 = ~n3232 ;
  assign y936 = ~n3235 ;
  assign y937 = ~n3238 ;
  assign y938 = n3243 ;
  assign y939 = ~n3245 ;
  assign y940 = n3246 ;
  assign y941 = ~1'b0 ;
  assign y942 = n3253 ;
  assign y943 = n3257 ;
  assign y944 = n3262 ;
  assign y945 = ~n3274 ;
  assign y946 = n3278 ;
  assign y947 = ~1'b0 ;
  assign y948 = ~n3280 ;
  assign y949 = n3286 ;
  assign y950 = ~1'b0 ;
  assign y951 = n3290 ;
  assign y952 = n3294 ;
  assign y953 = ~n3298 ;
  assign y954 = ~n3299 ;
  assign y955 = n3301 ;
  assign y956 = n3306 ;
  assign y957 = n3313 ;
  assign y958 = ~1'b0 ;
  assign y959 = ~1'b0 ;
  assign y960 = n3314 ;
  assign y961 = ~n3315 ;
  assign y962 = ~1'b0 ;
  assign y963 = n3320 ;
  assign y964 = n3321 ;
  assign y965 = n3324 ;
  assign y966 = n1403 ;
  assign y967 = ~n3328 ;
  assign y968 = ~n3339 ;
  assign y969 = ~n3346 ;
  assign y970 = ~1'b0 ;
  assign y971 = n3361 ;
  assign y972 = n3364 ;
  assign y973 = n3368 ;
  assign y974 = ~1'b0 ;
  assign y975 = n3371 ;
  assign y976 = ~1'b0 ;
  assign y977 = n3375 ;
  assign y978 = ~1'b0 ;
  assign y979 = ~n3378 ;
  assign y980 = n3381 ;
  assign y981 = ~n3385 ;
  assign y982 = ~n3391 ;
  assign y983 = ~n3392 ;
  assign y984 = ~n3397 ;
  assign y985 = ~1'b0 ;
  assign y986 = ~n3402 ;
  assign y987 = ~1'b0 ;
  assign y988 = ~n3409 ;
  assign y989 = n3415 ;
  assign y990 = n3419 ;
  assign y991 = ~1'b0 ;
  assign y992 = ~n3422 ;
  assign y993 = ~n3432 ;
  assign y994 = ~n3440 ;
  assign y995 = n3441 ;
  assign y996 = ~n3442 ;
  assign y997 = ~n3457 ;
  assign y998 = n3460 ;
  assign y999 = ~n3465 ;
  assign y1000 = n3466 ;
  assign y1001 = ~n3471 ;
  assign y1002 = n3475 ;
  assign y1003 = n3479 ;
  assign y1004 = ~n3481 ;
  assign y1005 = n3487 ;
  assign y1006 = n3490 ;
  assign y1007 = ~1'b0 ;
  assign y1008 = ~n3496 ;
  assign y1009 = n3504 ;
  assign y1010 = ~n3506 ;
  assign y1011 = ~n3510 ;
  assign y1012 = ~n3512 ;
  assign y1013 = ~1'b0 ;
  assign y1014 = ~n3515 ;
  assign y1015 = ~n3518 ;
  assign y1016 = ~n3521 ;
  assign y1017 = n3523 ;
  assign y1018 = n3528 ;
  assign y1019 = n3534 ;
  assign y1020 = ~1'b0 ;
  assign y1021 = ~n3541 ;
  assign y1022 = n3026 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = n3549 ;
  assign y1025 = n3559 ;
  assign y1026 = n3561 ;
  assign y1027 = ~n3565 ;
  assign y1028 = ~n3571 ;
  assign y1029 = n3573 ;
  assign y1030 = ~n3578 ;
  assign y1031 = n3579 ;
  assign y1032 = ~n3580 ;
  assign y1033 = n3584 ;
  assign y1034 = ~1'b0 ;
  assign y1035 = ~n3585 ;
  assign y1036 = 1'b0 ;
  assign y1037 = ~n3592 ;
  assign y1038 = n2234 ;
  assign y1039 = n3601 ;
  assign y1040 = ~1'b0 ;
  assign y1041 = n3602 ;
  assign y1042 = n3605 ;
  assign y1043 = ~n3609 ;
  assign y1044 = n3616 ;
  assign y1045 = ~n3617 ;
  assign y1046 = n3621 ;
  assign y1047 = ~n3625 ;
  assign y1048 = ~n3633 ;
  assign y1049 = n3639 ;
  assign y1050 = ~n3640 ;
  assign y1051 = n3651 ;
  assign y1052 = n3653 ;
  assign y1053 = ~n3656 ;
  assign y1054 = ~1'b0 ;
  assign y1055 = n3661 ;
  assign y1056 = n3666 ;
  assign y1057 = ~n3668 ;
  assign y1058 = ~1'b0 ;
  assign y1059 = ~n3672 ;
  assign y1060 = ~n3673 ;
  assign y1061 = n3676 ;
  assign y1062 = ~1'b0 ;
  assign y1063 = n3680 ;
  assign y1064 = n3684 ;
  assign y1065 = ~n3685 ;
  assign y1066 = ~n3688 ;
  assign y1067 = n3689 ;
  assign y1068 = n3693 ;
  assign y1069 = ~1'b0 ;
  assign y1070 = ~n3694 ;
  assign y1071 = ~n3701 ;
  assign y1072 = ~n3706 ;
  assign y1073 = n3713 ;
  assign y1074 = n3715 ;
  assign y1075 = n3716 ;
  assign y1076 = n3721 ;
  assign y1077 = ~n3722 ;
  assign y1078 = ~n3725 ;
  assign y1079 = n3737 ;
  assign y1080 = n3738 ;
  assign y1081 = n3739 ;
  assign y1082 = ~n3744 ;
  assign y1083 = n3748 ;
  assign y1084 = ~n3751 ;
  assign y1085 = n3757 ;
  assign y1086 = n3763 ;
  assign y1087 = n3765 ;
  assign y1088 = ~n3767 ;
  assign y1089 = n3769 ;
  assign y1090 = n3771 ;
  assign y1091 = ~n3772 ;
  assign y1092 = n3774 ;
  assign y1093 = ~n3776 ;
  assign y1094 = n3783 ;
  assign y1095 = ~n3784 ;
  assign y1096 = n3786 ;
  assign y1097 = n3792 ;
  assign y1098 = n3797 ;
  assign y1099 = n3798 ;
  assign y1100 = ~1'b0 ;
  assign y1101 = ~n3802 ;
  assign y1102 = n3805 ;
  assign y1103 = ~n3809 ;
  assign y1104 = n3811 ;
  assign y1105 = ~n3824 ;
  assign y1106 = n3829 ;
  assign y1107 = n3832 ;
  assign y1108 = n3834 ;
  assign y1109 = ~n3835 ;
  assign y1110 = n3841 ;
  assign y1111 = ~n3847 ;
  assign y1112 = n3859 ;
  assign y1113 = ~n3863 ;
  assign y1114 = n3868 ;
  assign y1115 = ~n3872 ;
  assign y1116 = ~n3876 ;
  assign y1117 = ~n3880 ;
  assign y1118 = ~1'b0 ;
  assign y1119 = ~n3885 ;
  assign y1120 = ~n3892 ;
  assign y1121 = ~n3903 ;
  assign y1122 = ~n3905 ;
  assign y1123 = n3907 ;
  assign y1124 = ~1'b0 ;
  assign y1125 = ~n3909 ;
  assign y1126 = n3911 ;
  assign y1127 = n3921 ;
  assign y1128 = n3935 ;
  assign y1129 = n3940 ;
  assign y1130 = ~n3943 ;
  assign y1131 = ~n3946 ;
  assign y1132 = ~n3947 ;
  assign y1133 = ~n3958 ;
  assign y1134 = n3962 ;
  assign y1135 = ~1'b0 ;
  assign y1136 = ~1'b0 ;
  assign y1137 = n3964 ;
  assign y1138 = n3965 ;
  assign y1139 = ~n3966 ;
  assign y1140 = n1405 ;
  assign y1141 = ~1'b0 ;
  assign y1142 = ~n3968 ;
  assign y1143 = n3973 ;
  assign y1144 = n3974 ;
  assign y1145 = n3979 ;
  assign y1146 = n3980 ;
  assign y1147 = n3986 ;
  assign y1148 = n3987 ;
  assign y1149 = n3989 ;
  assign y1150 = n3991 ;
  assign y1151 = n3994 ;
  assign y1152 = ~1'b0 ;
  assign y1153 = n3995 ;
  assign y1154 = n3999 ;
  assign y1155 = n4001 ;
  assign y1156 = ~n4002 ;
  assign y1157 = n4004 ;
  assign y1158 = ~n4008 ;
  assign y1159 = ~1'b0 ;
  assign y1160 = n4009 ;
  assign y1161 = ~1'b0 ;
  assign y1162 = ~n4013 ;
  assign y1163 = n4016 ;
  assign y1164 = n4026 ;
  assign y1165 = ~n4027 ;
  assign y1166 = ~n4028 ;
  assign y1167 = ~n4030 ;
  assign y1168 = ~1'b0 ;
  assign y1169 = ~1'b0 ;
  assign y1170 = ~n4032 ;
  assign y1171 = n4042 ;
  assign y1172 = n4043 ;
  assign y1173 = n4046 ;
  assign y1174 = n3858 ;
  assign y1175 = ~n4053 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = n1390 ;
  assign y1178 = n4056 ;
  assign y1179 = ~n4069 ;
  assign y1180 = n4079 ;
  assign y1181 = n4081 ;
  assign y1182 = n4086 ;
  assign y1183 = n4087 ;
  assign y1184 = n4089 ;
  assign y1185 = ~n4095 ;
  assign y1186 = ~1'b0 ;
  assign y1187 = n4100 ;
  assign y1188 = ~n4106 ;
  assign y1189 = ~n4108 ;
  assign y1190 = n4114 ;
  assign y1191 = ~n4116 ;
  assign y1192 = ~n4123 ;
  assign y1193 = ~n4125 ;
  assign y1194 = ~n4129 ;
  assign y1195 = ~n4134 ;
  assign y1196 = ~n4137 ;
  assign y1197 = ~1'b0 ;
  assign y1198 = n4138 ;
  assign y1199 = n4147 ;
  assign y1200 = ~1'b0 ;
  assign y1201 = n4151 ;
  assign y1202 = n4154 ;
  assign y1203 = ~n4157 ;
  assign y1204 = ~1'b0 ;
  assign y1205 = n4158 ;
  assign y1206 = ~n4166 ;
  assign y1207 = n4168 ;
  assign y1208 = n4180 ;
  assign y1209 = ~n4183 ;
  assign y1210 = ~n4189 ;
  assign y1211 = ~n4190 ;
  assign y1212 = ~n4194 ;
  assign y1213 = ~n4201 ;
  assign y1214 = ~n4202 ;
  assign y1215 = ~n4211 ;
  assign y1216 = ~1'b0 ;
  assign y1217 = ~1'b0 ;
  assign y1218 = ~1'b0 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~1'b0 ;
  assign y1221 = ~n4212 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = n4218 ;
  assign y1224 = ~n4227 ;
  assign y1225 = ~1'b0 ;
  assign y1226 = ~n4235 ;
  assign y1227 = ~1'b0 ;
  assign y1228 = ~n4237 ;
  assign y1229 = n4238 ;
  assign y1230 = n1662 ;
  assign y1231 = ~1'b0 ;
  assign y1232 = n4241 ;
  assign y1233 = ~n4242 ;
  assign y1234 = ~n4244 ;
  assign y1235 = ~n4248 ;
  assign y1236 = ~n4253 ;
  assign y1237 = n4257 ;
  assign y1238 = n4260 ;
  assign y1239 = ~n4266 ;
  assign y1240 = ~n4270 ;
  assign y1241 = n3138 ;
  assign y1242 = n4278 ;
  assign y1243 = n4283 ;
  assign y1244 = n4292 ;
  assign y1245 = n4294 ;
  assign y1246 = n4300 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = n4304 ;
  assign y1249 = n4314 ;
  assign y1250 = n4318 ;
  assign y1251 = ~n4325 ;
  assign y1252 = ~1'b0 ;
  assign y1253 = ~n4334 ;
  assign y1254 = ~n4345 ;
  assign y1255 = ~n4346 ;
  assign y1256 = ~1'b0 ;
  assign y1257 = n4349 ;
  assign y1258 = n4350 ;
  assign y1259 = ~n4353 ;
  assign y1260 = n4356 ;
  assign y1261 = n4359 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = n4360 ;
  assign y1264 = n4366 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = n4374 ;
  assign y1267 = n4379 ;
  assign y1268 = ~n4381 ;
  assign y1269 = n4389 ;
  assign y1270 = ~n4391 ;
  assign y1271 = n4394 ;
  assign y1272 = ~n4404 ;
  assign y1273 = ~n4409 ;
  assign y1274 = n4424 ;
  assign y1275 = ~n4425 ;
  assign y1276 = ~n4432 ;
  assign y1277 = ~n4433 ;
  assign y1278 = n4434 ;
  assign y1279 = ~n4435 ;
  assign y1280 = n4436 ;
  assign y1281 = ~n4439 ;
  assign y1282 = ~n4440 ;
  assign y1283 = n4442 ;
  assign y1284 = ~1'b0 ;
  assign y1285 = ~n4443 ;
  assign y1286 = n355 ;
  assign y1287 = ~1'b0 ;
  assign y1288 = ~n4445 ;
  assign y1289 = ~1'b0 ;
  assign y1290 = n4453 ;
  assign y1291 = ~n4454 ;
  assign y1292 = ~n4455 ;
  assign y1293 = ~n4460 ;
  assign y1294 = ~n4467 ;
  assign y1295 = ~1'b0 ;
  assign y1296 = ~n4472 ;
  assign y1297 = n4474 ;
  assign y1298 = ~1'b0 ;
  assign y1299 = ~n4476 ;
  assign y1300 = ~n4482 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = n4484 ;
  assign y1304 = ~n4490 ;
  assign y1305 = n4492 ;
  assign y1306 = ~n4494 ;
  assign y1307 = ~1'b0 ;
  assign y1308 = n4506 ;
  assign y1309 = ~n4509 ;
  assign y1310 = n4510 ;
  assign y1311 = ~n4512 ;
  assign y1312 = ~n4513 ;
  assign y1313 = n4517 ;
  assign y1314 = ~n4521 ;
  assign y1315 = ~1'b0 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = ~1'b0 ;
  assign y1318 = ~n4526 ;
  assign y1319 = ~n4527 ;
  assign y1320 = ~n4528 ;
  assign y1321 = n4532 ;
  assign y1322 = ~n4535 ;
  assign y1323 = ~n4543 ;
  assign y1324 = ~n4546 ;
  assign y1325 = n4551 ;
  assign y1326 = ~1'b0 ;
  assign y1327 = n4558 ;
  assign y1328 = ~1'b0 ;
  assign y1329 = ~1'b0 ;
  assign y1330 = ~n4559 ;
  assign y1331 = ~1'b0 ;
  assign y1332 = ~n4560 ;
  assign y1333 = ~1'b0 ;
  assign y1334 = n4562 ;
  assign y1335 = ~n4568 ;
  assign y1336 = ~n4574 ;
  assign y1337 = n4575 ;
  assign y1338 = n4577 ;
  assign y1339 = ~n4581 ;
  assign y1340 = ~n4582 ;
  assign y1341 = n4587 ;
  assign y1342 = ~1'b0 ;
  assign y1343 = ~n4592 ;
  assign y1344 = n4595 ;
  assign y1345 = n4598 ;
  assign y1346 = n4601 ;
  assign y1347 = ~n4603 ;
  assign y1348 = n330 ;
  assign y1349 = n4605 ;
  assign y1350 = ~n4606 ;
  assign y1351 = n1385 ;
  assign y1352 = n4612 ;
  assign y1353 = n4618 ;
  assign y1354 = ~n4624 ;
  assign y1355 = ~n4626 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = n4627 ;
  assign y1358 = ~n4630 ;
  assign y1359 = ~n4634 ;
  assign y1360 = n4637 ;
  assign y1361 = n4642 ;
  assign y1362 = n4644 ;
  assign y1363 = n4653 ;
  assign y1364 = ~1'b0 ;
  assign y1365 = n4659 ;
  assign y1366 = ~n4660 ;
  assign y1367 = n4662 ;
  assign y1368 = n4675 ;
  assign y1369 = ~1'b0 ;
  assign y1370 = n4678 ;
  assign y1371 = ~n4680 ;
  assign y1372 = ~n4682 ;
  assign y1373 = n4688 ;
  assign y1374 = ~n4689 ;
  assign y1375 = ~1'b0 ;
  assign y1376 = ~n4690 ;
  assign y1377 = ~n4694 ;
  assign y1378 = ~n4695 ;
  assign y1379 = n4698 ;
  assign y1380 = n4701 ;
  assign y1381 = ~n4705 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = n4706 ;
  assign y1384 = ~n4714 ;
  assign y1385 = n4715 ;
  assign y1386 = n4719 ;
  assign y1387 = ~n4725 ;
  assign y1388 = ~1'b0 ;
  assign y1389 = n4726 ;
  assign y1390 = ~n4730 ;
  assign y1391 = n4733 ;
  assign y1392 = ~n4735 ;
  assign y1393 = ~n4740 ;
  assign y1394 = ~n4745 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = n4754 ;
  assign y1397 = n4758 ;
  assign y1398 = ~n4760 ;
  assign y1399 = ~n4762 ;
  assign y1400 = n4765 ;
  assign y1401 = n4769 ;
  assign y1402 = ~1'b0 ;
  assign y1403 = ~n4770 ;
  assign y1404 = ~n4771 ;
  assign y1405 = n4775 ;
  assign y1406 = ~1'b0 ;
  assign y1407 = ~n4779 ;
  assign y1408 = ~n4781 ;
  assign y1409 = ~1'b0 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = n4787 ;
  assign y1412 = ~n4788 ;
  assign y1413 = ~n4789 ;
  assign y1414 = ~n4790 ;
  assign y1415 = n4797 ;
  assign y1416 = ~1'b0 ;
  assign y1417 = ~n4801 ;
  assign y1418 = ~1'b0 ;
  assign y1419 = n4809 ;
  assign y1420 = ~n4811 ;
  assign y1421 = n4819 ;
  assign y1422 = ~n4822 ;
  assign y1423 = ~n4823 ;
  assign y1424 = ~n4825 ;
  assign y1425 = ~n4828 ;
  assign y1426 = ~n4834 ;
  assign y1427 = ~n4837 ;
  assign y1428 = ~1'b0 ;
  assign y1429 = ~n4847 ;
  assign y1430 = ~1'b0 ;
  assign y1431 = ~n4859 ;
  assign y1432 = n4860 ;
  assign y1433 = n4863 ;
  assign y1434 = ~n4865 ;
  assign y1435 = ~n4868 ;
  assign y1436 = n4869 ;
  assign y1437 = n4874 ;
  assign y1438 = n4892 ;
  assign y1439 = ~n4893 ;
  assign y1440 = n4895 ;
  assign y1441 = ~n4900 ;
  assign y1442 = n4905 ;
  assign y1443 = n4907 ;
  assign y1444 = ~n4910 ;
  assign y1445 = n4916 ;
  assign y1446 = n4924 ;
  assign y1447 = ~n4930 ;
  assign y1448 = n4939 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = ~n4942 ;
  assign y1451 = ~1'b0 ;
  assign y1452 = ~n4947 ;
  assign y1453 = n4950 ;
  assign y1454 = ~n4956 ;
  assign y1455 = n4959 ;
  assign y1456 = ~n3765 ;
  assign y1457 = n4962 ;
  assign y1458 = n4963 ;
  assign y1459 = n4965 ;
  assign y1460 = ~1'b0 ;
  assign y1461 = n4975 ;
  assign y1462 = ~n4976 ;
  assign y1463 = ~n4979 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = ~n4983 ;
  assign y1466 = ~n5000 ;
  assign y1467 = ~n5004 ;
  assign y1468 = ~n5009 ;
  assign y1469 = ~n5014 ;
  assign y1470 = ~n5016 ;
  assign y1471 = n5019 ;
  assign y1472 = n5020 ;
  assign y1473 = n5026 ;
  assign y1474 = n5029 ;
  assign y1475 = ~n5030 ;
  assign y1476 = n5035 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = ~n5039 ;
  assign y1479 = n5050 ;
  assign y1480 = ~n2369 ;
  assign y1481 = n5051 ;
  assign y1482 = ~n5053 ;
  assign y1483 = ~1'b0 ;
  assign y1484 = n5064 ;
  assign y1485 = ~n5065 ;
  assign y1486 = ~1'b0 ;
  assign y1487 = n5066 ;
  assign y1488 = n5074 ;
  assign y1489 = ~n5081 ;
  assign y1490 = n5087 ;
  assign y1491 = ~n5088 ;
  assign y1492 = ~n3699 ;
  assign y1493 = ~1'b0 ;
  assign y1494 = n2519 ;
  assign y1495 = n5090 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = ~1'b0 ;
  assign y1498 = ~1'b0 ;
  assign y1499 = ~n5091 ;
  assign y1500 = ~1'b0 ;
  assign y1501 = ~n5094 ;
  assign y1502 = ~n5096 ;
  assign y1503 = ~n5097 ;
  assign y1504 = ~n5098 ;
  assign y1505 = n5107 ;
  assign y1506 = ~n5110 ;
  assign y1507 = ~n5114 ;
  assign y1508 = ~n5115 ;
  assign y1509 = ~1'b0 ;
  assign y1510 = ~1'b0 ;
  assign y1511 = n5121 ;
  assign y1512 = n5123 ;
  assign y1513 = n5127 ;
  assign y1514 = n5136 ;
  assign y1515 = ~n2878 ;
  assign y1516 = ~n5149 ;
  assign y1517 = n5150 ;
  assign y1518 = ~n436 ;
  assign y1519 = ~n5151 ;
  assign y1520 = n5153 ;
  assign y1521 = ~1'b0 ;
  assign y1522 = ~n5157 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~n5166 ;
  assign y1525 = n5167 ;
  assign y1526 = n5168 ;
  assign y1527 = n5172 ;
  assign y1528 = n5173 ;
  assign y1529 = ~1'b0 ;
  assign y1530 = ~n5176 ;
  assign y1531 = ~n5179 ;
  assign y1532 = ~n5195 ;
  assign y1533 = ~1'b0 ;
  assign y1534 = ~n5196 ;
  assign y1535 = ~n5199 ;
  assign y1536 = n5202 ;
  assign y1537 = n5205 ;
  assign y1538 = n5208 ;
  assign y1539 = ~n5212 ;
  assign y1540 = n5214 ;
  assign y1541 = ~n5217 ;
  assign y1542 = n5222 ;
  assign y1543 = ~n5225 ;
  assign y1544 = ~n5231 ;
  assign y1545 = ~n5235 ;
  assign y1546 = n5236 ;
  assign y1547 = ~n5242 ;
  assign y1548 = ~n5244 ;
  assign y1549 = n5246 ;
  assign y1550 = ~n5250 ;
  assign y1551 = n5252 ;
  assign y1552 = n5254 ;
  assign y1553 = ~n5256 ;
  assign y1554 = n5257 ;
  assign y1555 = ~n5261 ;
  assign y1556 = ~n5263 ;
  assign y1557 = n5265 ;
  assign y1558 = ~n5268 ;
  assign y1559 = n5272 ;
  assign y1560 = n5275 ;
  assign y1561 = ~n2945 ;
  assign y1562 = ~n5277 ;
  assign y1563 = ~n5279 ;
  assign y1564 = n1348 ;
  assign y1565 = n5286 ;
  assign y1566 = n5288 ;
  assign y1567 = ~n5289 ;
  assign y1568 = n5291 ;
  assign y1569 = ~1'b0 ;
  assign y1570 = ~n5298 ;
  assign y1571 = n5308 ;
  assign y1572 = ~n5310 ;
  assign y1573 = ~n5313 ;
  assign y1574 = ~n5316 ;
  assign y1575 = n5320 ;
  assign y1576 = n5321 ;
  assign y1577 = n5326 ;
  assign y1578 = n5331 ;
  assign y1579 = ~n5333 ;
  assign y1580 = ~n5334 ;
  assign y1581 = n5341 ;
  assign y1582 = ~x10 ;
  assign y1583 = n5344 ;
  assign y1584 = n5365 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = ~1'b0 ;
  assign y1587 = n5367 ;
  assign y1588 = n5368 ;
  assign y1589 = n5372 ;
  assign y1590 = ~n5376 ;
  assign y1591 = ~n5381 ;
  assign y1592 = ~n5383 ;
  assign y1593 = ~1'b0 ;
  assign y1594 = ~n305 ;
  assign y1595 = n5386 ;
  assign y1596 = n5387 ;
  assign y1597 = n5390 ;
  assign y1598 = ~n3148 ;
  assign y1599 = ~n5393 ;
  assign y1600 = ~n5397 ;
  assign y1601 = ~1'b0 ;
  assign y1602 = n5399 ;
  assign y1603 = ~n5406 ;
  assign y1604 = n5415 ;
  assign y1605 = n5427 ;
  assign y1606 = n5428 ;
  assign y1607 = n5436 ;
  assign y1608 = ~n5438 ;
  assign y1609 = n1743 ;
  assign y1610 = n5442 ;
  assign y1611 = ~n5448 ;
  assign y1612 = ~1'b0 ;
  assign y1613 = ~n5459 ;
  assign y1614 = ~n5484 ;
  assign y1615 = n5486 ;
  assign y1616 = n5490 ;
  assign y1617 = ~1'b0 ;
  assign y1618 = ~1'b0 ;
  assign y1619 = ~n5496 ;
  assign y1620 = ~1'b0 ;
  assign y1621 = ~n5497 ;
  assign y1622 = ~n5498 ;
  assign y1623 = n4429 ;
  assign y1624 = ~n5508 ;
  assign y1625 = ~n5510 ;
  assign y1626 = ~n5513 ;
  assign y1627 = ~n5517 ;
  assign y1628 = ~n5524 ;
  assign y1629 = n5526 ;
  assign y1630 = ~1'b0 ;
  assign y1631 = n5530 ;
  assign y1632 = ~n5533 ;
  assign y1633 = n5536 ;
  assign y1634 = ~n5538 ;
  assign y1635 = ~1'b0 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = n5539 ;
  assign y1638 = n5544 ;
  assign y1639 = ~1'b0 ;
  assign y1640 = ~n5551 ;
  assign y1641 = ~n5556 ;
  assign y1642 = ~n5564 ;
  assign y1643 = ~n5566 ;
  assign y1644 = n5570 ;
  assign y1645 = n5573 ;
  assign y1646 = ~n5579 ;
  assign y1647 = n5581 ;
  assign y1648 = n5582 ;
  assign y1649 = ~n5589 ;
  assign y1650 = n5595 ;
  assign y1651 = ~n5598 ;
  assign y1652 = n5607 ;
  assign y1653 = n5608 ;
  assign y1654 = n5613 ;
  assign y1655 = ~n5620 ;
  assign y1656 = n5627 ;
  assign y1657 = n5631 ;
  assign y1658 = ~n5637 ;
  assign y1659 = ~n5640 ;
  assign y1660 = ~n5647 ;
  assign y1661 = n5652 ;
  assign y1662 = n5653 ;
  assign y1663 = n5663 ;
  assign y1664 = ~n5667 ;
  assign y1665 = ~n5668 ;
  assign y1666 = ~n5671 ;
  assign y1667 = n5672 ;
  assign y1668 = ~n5676 ;
  assign y1669 = ~n5677 ;
  assign y1670 = ~n5681 ;
  assign y1671 = n5686 ;
  assign y1672 = n5689 ;
  assign y1673 = n3499 ;
  assign y1674 = ~n5691 ;
  assign y1675 = n5693 ;
  assign y1676 = ~n5701 ;
  assign y1677 = ~n5703 ;
  assign y1678 = ~n5707 ;
  assign y1679 = n5709 ;
  assign y1680 = n5710 ;
  assign y1681 = n5720 ;
  assign y1682 = ~n5722 ;
  assign y1683 = ~n5723 ;
  assign y1684 = ~n5726 ;
  assign y1685 = ~n5733 ;
  assign y1686 = n5735 ;
  assign y1687 = n5741 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = ~1'b0 ;
  assign y1690 = ~n5744 ;
  assign y1691 = n5746 ;
  assign y1692 = n5748 ;
  assign y1693 = ~n5750 ;
  assign y1694 = ~n5754 ;
  assign y1695 = ~n5757 ;
  assign y1696 = n5758 ;
  assign y1697 = ~n5759 ;
  assign y1698 = n5760 ;
  assign y1699 = n5763 ;
  assign y1700 = ~n5770 ;
  assign y1701 = ~n5773 ;
  assign y1702 = 1'b0 ;
  assign y1703 = ~n5780 ;
  assign y1704 = ~n5783 ;
  assign y1705 = n5785 ;
  assign y1706 = n5789 ;
  assign y1707 = n5795 ;
  assign y1708 = n5803 ;
  assign y1709 = n5804 ;
  assign y1710 = n5805 ;
  assign y1711 = ~n5811 ;
  assign y1712 = ~n5816 ;
  assign y1713 = ~1'b0 ;
  assign y1714 = n5819 ;
  assign y1715 = n5822 ;
  assign y1716 = n5823 ;
  assign y1717 = n5827 ;
  assign y1718 = ~n5834 ;
  assign y1719 = ~1'b0 ;
  assign y1720 = ~n5839 ;
  assign y1721 = ~n5842 ;
  assign y1722 = ~1'b0 ;
  assign y1723 = n5843 ;
  assign y1724 = n5849 ;
  assign y1725 = n5851 ;
  assign y1726 = ~n5857 ;
  assign y1727 = ~n5863 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = n5866 ;
  assign y1730 = n5872 ;
  assign y1731 = ~n5873 ;
  assign y1732 = ~n5876 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = ~n5879 ;
  assign y1735 = n5884 ;
  assign y1736 = ~n5887 ;
  assign y1737 = n5889 ;
  assign y1738 = ~n5894 ;
  assign y1739 = ~1'b0 ;
  assign y1740 = ~1'b0 ;
  assign y1741 = n5896 ;
  assign y1742 = n5900 ;
  assign y1743 = n5901 ;
  assign y1744 = ~n5903 ;
  assign y1745 = n5909 ;
  assign y1746 = n5917 ;
  assign y1747 = n5930 ;
  assign y1748 = n5931 ;
  assign y1749 = ~1'b0 ;
  assign y1750 = ~n5935 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = ~n5938 ;
  assign y1753 = n5942 ;
  assign y1754 = ~1'b0 ;
  assign y1755 = ~n5946 ;
  assign y1756 = n5949 ;
  assign y1757 = ~n5950 ;
  assign y1758 = ~1'b0 ;
  assign y1759 = ~n5958 ;
  assign y1760 = ~1'b0 ;
  assign y1761 = ~n5961 ;
  assign y1762 = n5970 ;
  assign y1763 = n5978 ;
  assign y1764 = ~n5981 ;
  assign y1765 = ~n5982 ;
  assign y1766 = ~1'b0 ;
  assign y1767 = n5983 ;
  assign y1768 = ~1'b0 ;
  assign y1769 = n5988 ;
  assign y1770 = ~n5989 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = n5991 ;
  assign y1773 = n5996 ;
  assign y1774 = n5998 ;
  assign y1775 = ~n6003 ;
  assign y1776 = ~1'b0 ;
  assign y1777 = ~n6008 ;
  assign y1778 = ~n6009 ;
  assign y1779 = n6019 ;
  assign y1780 = n6030 ;
  assign y1781 = ~n6032 ;
  assign y1782 = ~n6038 ;
  assign y1783 = ~1'b0 ;
  assign y1784 = n6044 ;
  assign y1785 = ~1'b0 ;
  assign y1786 = n6051 ;
  assign y1787 = ~n6055 ;
  assign y1788 = n6060 ;
  assign y1789 = ~1'b0 ;
  assign y1790 = n6066 ;
  assign y1791 = ~n6068 ;
  assign y1792 = n6075 ;
  assign y1793 = ~n6077 ;
  assign y1794 = n6081 ;
  assign y1795 = n6083 ;
  assign y1796 = ~n6085 ;
  assign y1797 = ~n6091 ;
  assign y1798 = n6096 ;
  assign y1799 = ~n6105 ;
  assign y1800 = ~n6108 ;
  assign y1801 = ~n6113 ;
  assign y1802 = n6117 ;
  assign y1803 = ~n6121 ;
  assign y1804 = ~n6123 ;
  assign y1805 = ~n6125 ;
  assign y1806 = ~n6146 ;
  assign y1807 = ~n6155 ;
  assign y1808 = ~n6156 ;
  assign y1809 = n6159 ;
  assign y1810 = ~n6170 ;
  assign y1811 = ~n6178 ;
  assign y1812 = n6179 ;
  assign y1813 = ~n6182 ;
  assign y1814 = n6191 ;
  assign y1815 = n6196 ;
  assign y1816 = ~n6199 ;
  assign y1817 = n6201 ;
  assign y1818 = n6203 ;
  assign y1819 = n6207 ;
  assign y1820 = ~n6220 ;
  assign y1821 = ~1'b0 ;
  assign y1822 = ~n6227 ;
  assign y1823 = ~n6228 ;
  assign y1824 = n6233 ;
  assign y1825 = n6237 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~n6241 ;
  assign y1828 = n6242 ;
  assign y1829 = ~n6244 ;
  assign y1830 = ~n6245 ;
  assign y1831 = n6249 ;
  assign y1832 = n1607 ;
  assign y1833 = ~n6250 ;
  assign y1834 = n6253 ;
  assign y1835 = n1475 ;
  assign y1836 = ~n6262 ;
  assign y1837 = ~1'b0 ;
  assign y1838 = ~n6265 ;
  assign y1839 = ~1'b0 ;
  assign y1840 = ~1'b0 ;
  assign y1841 = n6266 ;
  assign y1842 = ~1'b0 ;
  assign y1843 = n6271 ;
  assign y1844 = n6273 ;
  assign y1845 = n6276 ;
  assign y1846 = n6288 ;
  assign y1847 = n6291 ;
  assign y1848 = ~1'b0 ;
  assign y1849 = ~n6294 ;
  assign y1850 = ~n6295 ;
  assign y1851 = n6299 ;
  assign y1852 = n6301 ;
  assign y1853 = ~n6307 ;
  assign y1854 = n6308 ;
  assign y1855 = ~n6310 ;
  assign y1856 = ~n6312 ;
  assign y1857 = ~1'b0 ;
  assign y1858 = n5507 ;
  assign y1859 = ~n6318 ;
  assign y1860 = ~n6319 ;
  assign y1861 = n6325 ;
  assign y1862 = n6329 ;
  assign y1863 = n6330 ;
  assign y1864 = n6331 ;
  assign y1865 = n6332 ;
  assign y1866 = ~n6337 ;
  assign y1867 = ~n6344 ;
  assign y1868 = ~n6345 ;
  assign y1869 = n6351 ;
  assign y1870 = ~n6353 ;
  assign y1871 = n6357 ;
  assign y1872 = n6361 ;
  assign y1873 = n6365 ;
  assign y1874 = n6374 ;
  assign y1875 = n6381 ;
  assign y1876 = ~n6386 ;
  assign y1877 = ~n6388 ;
  assign y1878 = ~1'b0 ;
  assign y1879 = ~n6394 ;
  assign y1880 = ~n6397 ;
  assign y1881 = n6398 ;
  assign y1882 = n6401 ;
  assign y1883 = n6402 ;
  assign y1884 = ~n6405 ;
  assign y1885 = ~n6411 ;
  assign y1886 = ~n6417 ;
  assign y1887 = n6427 ;
  assign y1888 = n6428 ;
  assign y1889 = ~n6432 ;
  assign y1890 = ~1'b0 ;
  assign y1891 = ~n6434 ;
  assign y1892 = ~n6437 ;
  assign y1893 = ~1'b0 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = ~1'b0 ;
  assign y1896 = ~n6438 ;
  assign y1897 = n6440 ;
  assign y1898 = n6444 ;
  assign y1899 = ~n6455 ;
  assign y1900 = ~n6456 ;
  assign y1901 = n6459 ;
  assign y1902 = ~n6465 ;
  assign y1903 = ~1'b0 ;
  assign y1904 = n6484 ;
  assign y1905 = ~n6506 ;
  assign y1906 = ~n6508 ;
  assign y1907 = ~1'b0 ;
  assign y1908 = n6509 ;
  assign y1909 = n6510 ;
  assign y1910 = ~1'b0 ;
  assign y1911 = ~1'b0 ;
  assign y1912 = ~n6515 ;
  assign y1913 = n6521 ;
  assign y1914 = ~n6524 ;
  assign y1915 = ~n6527 ;
  assign y1916 = ~n6528 ;
  assign y1917 = ~1'b0 ;
  assign y1918 = n6530 ;
  assign y1919 = ~1'b0 ;
  assign y1920 = ~n6536 ;
  assign y1921 = n6538 ;
  assign y1922 = ~n6542 ;
  assign y1923 = ~n6543 ;
  assign y1924 = ~n6548 ;
  assign y1925 = n6553 ;
  assign y1926 = ~n6555 ;
  assign y1927 = n6565 ;
  assign y1928 = n6568 ;
  assign y1929 = ~n6574 ;
  assign y1930 = n6577 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = ~1'b0 ;
  assign y1933 = n6579 ;
  assign y1934 = n6594 ;
  assign y1935 = ~n6596 ;
  assign y1936 = ~1'b0 ;
  assign y1937 = n6599 ;
  assign y1938 = ~n6610 ;
  assign y1939 = n6613 ;
  assign y1940 = n6615 ;
  assign y1941 = n6619 ;
  assign y1942 = n6621 ;
  assign y1943 = ~n6627 ;
  assign y1944 = ~n6637 ;
  assign y1945 = ~n6639 ;
  assign y1946 = n6642 ;
  assign y1947 = ~n6643 ;
  assign y1948 = n6645 ;
  assign y1949 = ~1'b0 ;
  assign y1950 = ~1'b0 ;
  assign y1951 = ~n6659 ;
  assign y1952 = n6660 ;
  assign y1953 = ~n6664 ;
  assign y1954 = n4250 ;
  assign y1955 = n6669 ;
  assign y1956 = ~n6670 ;
  assign y1957 = ~1'b0 ;
  assign y1958 = ~n6674 ;
  assign y1959 = n6677 ;
  assign y1960 = ~1'b0 ;
  assign y1961 = ~1'b0 ;
  assign y1962 = ~n6679 ;
  assign y1963 = ~n6681 ;
  assign y1964 = ~n6687 ;
  assign y1965 = ~n6695 ;
  assign y1966 = ~1'b0 ;
  assign y1967 = ~1'b0 ;
  assign y1968 = ~n3771 ;
  assign y1969 = n6696 ;
  assign y1970 = ~n6698 ;
  assign y1971 = n6707 ;
  assign y1972 = n6708 ;
  assign y1973 = ~n6716 ;
  assign y1974 = n6723 ;
  assign y1975 = n6725 ;
  assign y1976 = n6730 ;
  assign y1977 = ~n6735 ;
  assign y1978 = n4152 ;
  assign y1979 = ~n6736 ;
  assign y1980 = n6742 ;
  assign y1981 = n6743 ;
  assign y1982 = n6745 ;
  assign y1983 = ~n6750 ;
  assign y1984 = n6757 ;
  assign y1985 = ~n6758 ;
  assign y1986 = n6759 ;
  assign y1987 = ~n3479 ;
  assign y1988 = ~n6761 ;
  assign y1989 = ~n6767 ;
  assign y1990 = ~1'b0 ;
  assign y1991 = n6781 ;
  assign y1992 = ~n6782 ;
  assign y1993 = n6784 ;
  assign y1994 = n6786 ;
  assign y1995 = ~n6787 ;
  assign y1996 = ~1'b0 ;
  assign y1997 = ~n6792 ;
  assign y1998 = ~n6799 ;
  assign y1999 = ~1'b0 ;
  assign y2000 = n6800 ;
  assign y2001 = ~n6803 ;
  assign y2002 = n6806 ;
  assign y2003 = ~n6808 ;
  assign y2004 = ~n6811 ;
  assign y2005 = n6820 ;
  assign y2006 = n2860 ;
  assign y2007 = ~n6824 ;
  assign y2008 = n6825 ;
  assign y2009 = ~1'b0 ;
  assign y2010 = ~1'b0 ;
  assign y2011 = ~n6829 ;
  assign y2012 = n6831 ;
  assign y2013 = ~n6833 ;
  assign y2014 = ~n6838 ;
  assign y2015 = n6841 ;
  assign y2016 = n6849 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = ~n6850 ;
  assign y2019 = n6858 ;
  assign y2020 = n6871 ;
  assign y2021 = ~n6879 ;
  assign y2022 = ~n6893 ;
  assign y2023 = ~1'b0 ;
  assign y2024 = n6903 ;
  assign y2025 = ~n6905 ;
  assign y2026 = ~n6907 ;
  assign y2027 = ~n6908 ;
  assign y2028 = n6912 ;
  assign y2029 = n6915 ;
  assign y2030 = n6919 ;
  assign y2031 = ~n6925 ;
  assign y2032 = n6930 ;
  assign y2033 = ~n6933 ;
  assign y2034 = n6937 ;
  assign y2035 = ~n6940 ;
  assign y2036 = ~n6943 ;
  assign y2037 = ~n6949 ;
  assign y2038 = ~n6952 ;
  assign y2039 = ~n6954 ;
  assign y2040 = ~n6956 ;
  assign y2041 = n6973 ;
  assign y2042 = ~n6977 ;
  assign y2043 = ~n6978 ;
  assign y2044 = n6981 ;
  assign y2045 = n6983 ;
  assign y2046 = ~1'b0 ;
  assign y2047 = ~n6984 ;
  assign y2048 = ~n6988 ;
  assign y2049 = ~1'b0 ;
  assign y2050 = ~n6989 ;
  assign y2051 = ~n6995 ;
  assign y2052 = ~1'b0 ;
  assign y2053 = ~1'b0 ;
  assign y2054 = ~n7001 ;
  assign y2055 = ~n7003 ;
  assign y2056 = ~n7004 ;
  assign y2057 = n7009 ;
  assign y2058 = ~n7016 ;
  assign y2059 = ~n7017 ;
  assign y2060 = ~1'b0 ;
  assign y2061 = n7021 ;
  assign y2062 = ~n7023 ;
  assign y2063 = ~n7024 ;
  assign y2064 = ~1'b0 ;
  assign y2065 = ~n7025 ;
  assign y2066 = n7026 ;
  assign y2067 = ~n7029 ;
  assign y2068 = ~1'b0 ;
  assign y2069 = ~n7031 ;
  assign y2070 = n7032 ;
  assign y2071 = ~n7040 ;
  assign y2072 = ~n7042 ;
  assign y2073 = n7048 ;
  assign y2074 = n7051 ;
  assign y2075 = n7052 ;
  assign y2076 = n7062 ;
  assign y2077 = n5509 ;
  assign y2078 = n7063 ;
  assign y2079 = n7071 ;
  assign y2080 = ~n7073 ;
  assign y2081 = n7075 ;
  assign y2082 = ~n7080 ;
  assign y2083 = ~n7081 ;
  assign y2084 = ~n7086 ;
  assign y2085 = n7092 ;
  assign y2086 = ~n7096 ;
  assign y2087 = ~n7098 ;
  assign y2088 = ~n7099 ;
  assign y2089 = ~n7101 ;
  assign y2090 = ~1'b0 ;
  assign y2091 = ~n7103 ;
  assign y2092 = ~n7107 ;
  assign y2093 = ~1'b0 ;
  assign y2094 = ~n7112 ;
  assign y2095 = ~n7117 ;
  assign y2096 = ~n7118 ;
  assign y2097 = n7119 ;
  assign y2098 = ~n7122 ;
  assign y2099 = n7123 ;
  assign y2100 = 1'b0 ;
  assign y2101 = n7129 ;
  assign y2102 = ~n7130 ;
  assign y2103 = n7131 ;
  assign y2104 = n7133 ;
  assign y2105 = n7134 ;
  assign y2106 = n7136 ;
  assign y2107 = ~n7142 ;
  assign y2108 = 1'b0 ;
  assign y2109 = n7148 ;
  assign y2110 = n7149 ;
  assign y2111 = n7156 ;
  assign y2112 = 1'b0 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = ~1'b0 ;
  assign y2115 = n7159 ;
  assign y2116 = 1'b0 ;
  assign y2117 = ~1'b0 ;
  assign y2118 = ~n7168 ;
  assign y2119 = n7174 ;
  assign y2120 = ~n7176 ;
  assign y2121 = n7180 ;
  assign y2122 = n7181 ;
  assign y2123 = ~n7190 ;
  assign y2124 = ~n7204 ;
  assign y2125 = n7209 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = n7214 ;
  assign y2128 = n7218 ;
  assign y2129 = ~1'b0 ;
  assign y2130 = n7220 ;
  assign y2131 = n7222 ;
  assign y2132 = ~n7223 ;
  assign y2133 = n7225 ;
  assign y2134 = ~n7234 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = n7235 ;
  assign y2137 = ~n7248 ;
  assign y2138 = n7250 ;
  assign y2139 = n7256 ;
  assign y2140 = n7257 ;
  assign y2141 = n7260 ;
  assign y2142 = n5025 ;
  assign y2143 = n7263 ;
  assign y2144 = n7265 ;
  assign y2145 = n7266 ;
  assign y2146 = n5500 ;
  assign y2147 = ~n7272 ;
  assign y2148 = n7278 ;
  assign y2149 = ~n7280 ;
  assign y2150 = n7281 ;
  assign y2151 = ~n7283 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = n7291 ;
  assign y2154 = ~n7296 ;
  assign y2155 = ~1'b0 ;
  assign y2156 = n7298 ;
  assign y2157 = ~n7302 ;
  assign y2158 = n7304 ;
  assign y2159 = ~1'b0 ;
  assign y2160 = ~n7311 ;
  assign y2161 = ~n7313 ;
  assign y2162 = n7322 ;
  assign y2163 = n7323 ;
  assign y2164 = n7331 ;
  assign y2165 = ~1'b0 ;
  assign y2166 = n7336 ;
  assign y2167 = ~n7341 ;
  assign y2168 = n7345 ;
  assign y2169 = ~1'b0 ;
  assign y2170 = n7349 ;
  assign y2171 = ~n7354 ;
  assign y2172 = ~n7355 ;
  assign y2173 = n7359 ;
  assign y2174 = n7361 ;
  assign y2175 = ~1'b0 ;
  assign y2176 = n7371 ;
  assign y2177 = ~n7374 ;
  assign y2178 = n7382 ;
  assign y2179 = ~n7390 ;
  assign y2180 = ~n7392 ;
  assign y2181 = ~n7395 ;
  assign y2182 = n7396 ;
  assign y2183 = n7402 ;
  assign y2184 = n7408 ;
  assign y2185 = n7409 ;
  assign y2186 = ~n7412 ;
  assign y2187 = n7417 ;
  assign y2188 = n7419 ;
  assign y2189 = n7421 ;
  assign y2190 = n7427 ;
  assign y2191 = n7428 ;
  assign y2192 = n7434 ;
  assign y2193 = n7436 ;
  assign y2194 = ~n7444 ;
  assign y2195 = ~n7445 ;
  assign y2196 = n7446 ;
  assign y2197 = ~n7448 ;
  assign y2198 = ~n7449 ;
  assign y2199 = ~1'b0 ;
  assign y2200 = n7466 ;
  assign y2201 = ~n7473 ;
  assign y2202 = ~n7475 ;
  assign y2203 = n7477 ;
  assign y2204 = n7478 ;
  assign y2205 = n7481 ;
  assign y2206 = n7488 ;
  assign y2207 = ~n7490 ;
  assign y2208 = ~n7496 ;
  assign y2209 = n7498 ;
  assign y2210 = ~1'b0 ;
  assign y2211 = ~1'b0 ;
  assign y2212 = n7499 ;
  assign y2213 = ~n7500 ;
  assign y2214 = ~n7501 ;
  assign y2215 = n7503 ;
  assign y2216 = n7505 ;
  assign y2217 = ~n7508 ;
  assign y2218 = ~n7510 ;
  assign y2219 = ~1'b0 ;
  assign y2220 = ~n7520 ;
  assign y2221 = ~n7524 ;
  assign y2222 = ~n7528 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = n7541 ;
  assign y2225 = ~1'b0 ;
  assign y2226 = n7544 ;
  assign y2227 = ~n7547 ;
  assign y2228 = ~n393 ;
  assign y2229 = n7549 ;
  assign y2230 = ~n7551 ;
  assign y2231 = n7553 ;
  assign y2232 = ~n7557 ;
  assign y2233 = ~n7561 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = ~1'b0 ;
  assign y2236 = n7572 ;
  assign y2237 = ~n7574 ;
  assign y2238 = ~n5928 ;
  assign y2239 = ~1'b0 ;
  assign y2240 = ~n7583 ;
  assign y2241 = n7584 ;
  assign y2242 = ~1'b0 ;
  assign y2243 = ~n7590 ;
  assign y2244 = n7592 ;
  assign y2245 = n7593 ;
  assign y2246 = ~1'b0 ;
  assign y2247 = ~n7605 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = n7610 ;
  assign y2250 = ~n7616 ;
  assign y2251 = n7622 ;
  assign y2252 = n7628 ;
  assign y2253 = n7639 ;
  assign y2254 = ~n7646 ;
  assign y2255 = ~n7656 ;
  assign y2256 = n7663 ;
  assign y2257 = ~n7668 ;
  assign y2258 = n7672 ;
  assign y2259 = n7674 ;
  assign y2260 = n7676 ;
  assign y2261 = n1795 ;
  assign y2262 = n7679 ;
  assign y2263 = ~1'b0 ;
  assign y2264 = ~n7681 ;
  assign y2265 = ~n7685 ;
  assign y2266 = ~n7691 ;
  assign y2267 = ~n7694 ;
  assign y2268 = ~n7705 ;
  assign y2269 = n7706 ;
  assign y2270 = ~1'b0 ;
  assign y2271 = ~n7712 ;
  assign y2272 = n7718 ;
  assign y2273 = ~n7727 ;
  assign y2274 = n7729 ;
  assign y2275 = n7743 ;
  assign y2276 = ~n7745 ;
  assign y2277 = n7746 ;
  assign y2278 = ~n7754 ;
  assign y2279 = ~1'b0 ;
  assign y2280 = ~n7757 ;
  assign y2281 = n7763 ;
  assign y2282 = ~n7767 ;
  assign y2283 = ~n7773 ;
  assign y2284 = n7775 ;
  assign y2285 = n7777 ;
  assign y2286 = ~n7779 ;
  assign y2287 = ~n7785 ;
  assign y2288 = n7788 ;
  assign y2289 = n7795 ;
  assign y2290 = ~n7796 ;
  assign y2291 = ~1'b0 ;
  assign y2292 = n7798 ;
  assign y2293 = ~n7815 ;
  assign y2294 = ~n7826 ;
  assign y2295 = n7831 ;
  assign y2296 = n7837 ;
  assign y2297 = n7840 ;
  assign y2298 = ~n7846 ;
  assign y2299 = n7848 ;
  assign y2300 = ~1'b0 ;
  assign y2301 = n7850 ;
  assign y2302 = n7854 ;
  assign y2303 = n7857 ;
  assign y2304 = n7864 ;
  assign y2305 = n7869 ;
  assign y2306 = ~n7871 ;
  assign y2307 = ~1'b0 ;
  assign y2308 = ~n7873 ;
  assign y2309 = n7884 ;
  assign y2310 = ~n7887 ;
  assign y2311 = ~n7889 ;
  assign y2312 = ~1'b0 ;
  assign y2313 = ~n7890 ;
  assign y2314 = n7894 ;
  assign y2315 = n7908 ;
  assign y2316 = n7909 ;
  assign y2317 = ~n7912 ;
  assign y2318 = n7919 ;
  assign y2319 = ~n7920 ;
  assign y2320 = ~n7930 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = ~n7932 ;
  assign y2323 = ~n7934 ;
  assign y2324 = ~n7939 ;
  assign y2325 = ~n7944 ;
  assign y2326 = ~n7952 ;
  assign y2327 = n7961 ;
  assign y2328 = n7969 ;
  assign y2329 = ~1'b0 ;
  assign y2330 = ~n7971 ;
  assign y2331 = ~n7974 ;
  assign y2332 = n7987 ;
  assign y2333 = ~n7988 ;
  assign y2334 = n7989 ;
  assign y2335 = ~n7992 ;
  assign y2336 = n7999 ;
  assign y2337 = ~n8000 ;
  assign y2338 = n8001 ;
  assign y2339 = ~n8007 ;
  assign y2340 = ~1'b0 ;
  assign y2341 = n8010 ;
  assign y2342 = ~n8012 ;
  assign y2343 = n8013 ;
  assign y2344 = n8015 ;
  assign y2345 = n8018 ;
  assign y2346 = ~1'b0 ;
  assign y2347 = ~n8020 ;
  assign y2348 = ~n8023 ;
  assign y2349 = n8024 ;
  assign y2350 = n8025 ;
  assign y2351 = n8036 ;
  assign y2352 = n8042 ;
  assign y2353 = ~n8044 ;
  assign y2354 = n8050 ;
  assign y2355 = ~n8051 ;
  assign y2356 = n8057 ;
  assign y2357 = ~n8060 ;
  assign y2358 = n8064 ;
  assign y2359 = n8069 ;
  assign y2360 = ~n8073 ;
  assign y2361 = n8078 ;
  assign y2362 = ~n8082 ;
  assign y2363 = n8084 ;
  assign y2364 = n8085 ;
  assign y2365 = n8088 ;
  assign y2366 = ~n8090 ;
  assign y2367 = ~1'b0 ;
  assign y2368 = n8096 ;
  assign y2369 = n8100 ;
  assign y2370 = n8101 ;
  assign y2371 = ~n8104 ;
  assign y2372 = ~1'b0 ;
  assign y2373 = n8105 ;
  assign y2374 = ~1'b0 ;
  assign y2375 = ~n8111 ;
  assign y2376 = ~n8112 ;
  assign y2377 = ~n8117 ;
  assign y2378 = ~n8131 ;
  assign y2379 = ~n8136 ;
  assign y2380 = ~n8146 ;
  assign y2381 = ~n8148 ;
  assign y2382 = ~n8152 ;
  assign y2383 = n8154 ;
  assign y2384 = n8158 ;
  assign y2385 = n8159 ;
  assign y2386 = n8163 ;
  assign y2387 = ~n8167 ;
  assign y2388 = ~1'b0 ;
  assign y2389 = ~1'b0 ;
  assign y2390 = ~1'b0 ;
  assign y2391 = ~n8170 ;
  assign y2392 = ~n8171 ;
  assign y2393 = n8174 ;
  assign y2394 = n8177 ;
  assign y2395 = ~n8178 ;
  assign y2396 = ~1'b0 ;
  assign y2397 = n8182 ;
  assign y2398 = n8186 ;
  assign y2399 = ~n8187 ;
  assign y2400 = n8194 ;
  assign y2401 = n8195 ;
  assign y2402 = n8201 ;
  assign y2403 = n8208 ;
  assign y2404 = n8209 ;
  assign y2405 = ~n8211 ;
  assign y2406 = ~1'b0 ;
  assign y2407 = ~n8215 ;
  assign y2408 = ~n8217 ;
  assign y2409 = ~1'b0 ;
  assign y2410 = ~n8230 ;
  assign y2411 = ~n8234 ;
  assign y2412 = ~n8237 ;
  assign y2413 = ~1'b0 ;
  assign y2414 = 1'b0 ;
  assign y2415 = ~n8239 ;
  assign y2416 = n8240 ;
  assign y2417 = n8253 ;
  assign y2418 = ~n8257 ;
  assign y2419 = ~n8258 ;
  assign y2420 = n8267 ;
  assign y2421 = n8270 ;
  assign y2422 = n8272 ;
  assign y2423 = ~1'b0 ;
  assign y2424 = n8278 ;
  assign y2425 = n8280 ;
  assign y2426 = ~n8281 ;
  assign y2427 = n8288 ;
  assign y2428 = ~n8293 ;
  assign y2429 = n8294 ;
  assign y2430 = n8296 ;
  assign y2431 = ~n8301 ;
  assign y2432 = ~n8304 ;
  assign y2433 = n3924 ;
  assign y2434 = n8309 ;
  assign y2435 = ~n8314 ;
  assign y2436 = n8316 ;
  assign y2437 = n8319 ;
  assign y2438 = n8320 ;
  assign y2439 = ~1'b0 ;
  assign y2440 = n8325 ;
  assign y2441 = n8328 ;
  assign y2442 = ~n8332 ;
  assign y2443 = n8336 ;
  assign y2444 = ~n8341 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = ~n8343 ;
  assign y2447 = ~1'b0 ;
  assign y2448 = n8344 ;
  assign y2449 = n8345 ;
  assign y2450 = ~n8348 ;
  assign y2451 = ~n8350 ;
  assign y2452 = ~n8352 ;
  assign y2453 = ~n8355 ;
  assign y2454 = ~n8358 ;
  assign y2455 = n8359 ;
  assign y2456 = n6246 ;
  assign y2457 = ~n8363 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = n8365 ;
  assign y2460 = ~1'b0 ;
  assign y2461 = n8375 ;
  assign y2462 = n8376 ;
  assign y2463 = ~n8381 ;
  assign y2464 = ~n8384 ;
  assign y2465 = n8387 ;
  assign y2466 = n8394 ;
  assign y2467 = ~n8401 ;
  assign y2468 = ~n8402 ;
  assign y2469 = ~n8411 ;
  assign y2470 = n8412 ;
  assign y2471 = ~n8421 ;
  assign y2472 = ~1'b0 ;
  assign y2473 = n8422 ;
  assign y2474 = ~n8425 ;
  assign y2475 = ~n8426 ;
  assign y2476 = n8436 ;
  assign y2477 = n8441 ;
  assign y2478 = ~n8444 ;
  assign y2479 = ~1'b0 ;
  assign y2480 = n8448 ;
  assign y2481 = n8449 ;
  assign y2482 = ~1'b0 ;
  assign y2483 = ~n8458 ;
  assign y2484 = ~n8461 ;
  assign y2485 = n1472 ;
  assign y2486 = ~n8462 ;
  assign y2487 = n8464 ;
  assign y2488 = ~n8469 ;
  assign y2489 = ~n1547 ;
  assign y2490 = ~n8475 ;
  assign y2491 = ~n8484 ;
  assign y2492 = n8486 ;
  assign y2493 = ~n8490 ;
  assign y2494 = n8492 ;
  assign y2495 = n8493 ;
  assign y2496 = ~n8496 ;
  assign y2497 = n8500 ;
  assign y2498 = ~n8504 ;
  assign y2499 = n8512 ;
  assign y2500 = n8517 ;
  assign y2501 = n5299 ;
  assign y2502 = n8519 ;
  assign y2503 = ~1'b0 ;
  assign y2504 = ~n8522 ;
  assign y2505 = ~1'b0 ;
  assign y2506 = ~n8523 ;
  assign y2507 = n8531 ;
  assign y2508 = ~n8535 ;
  assign y2509 = ~n8540 ;
  assign y2510 = ~1'b0 ;
  assign y2511 = ~n8541 ;
  assign y2512 = ~n8546 ;
  assign y2513 = ~1'b0 ;
  assign y2514 = n8550 ;
  assign y2515 = n8554 ;
  assign y2516 = ~n8561 ;
  assign y2517 = n8565 ;
  assign y2518 = ~n810 ;
  assign y2519 = n8567 ;
  assign y2520 = ~1'b0 ;
  assign y2521 = n8568 ;
  assign y2522 = ~n8573 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = n8574 ;
  assign y2525 = n8580 ;
  assign y2526 = ~n8581 ;
  assign y2527 = n8582 ;
  assign y2528 = n8589 ;
  assign y2529 = n8595 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~1'b0 ;
  assign y2532 = ~1'b0 ;
  assign y2533 = ~1'b0 ;
  assign y2534 = ~n8598 ;
  assign y2535 = ~n8601 ;
  assign y2536 = n8603 ;
  assign y2537 = ~n8610 ;
  assign y2538 = ~n8617 ;
  assign y2539 = ~n8631 ;
  assign y2540 = ~n8632 ;
  assign y2541 = ~1'b0 ;
  assign y2542 = n8641 ;
  assign y2543 = ~n8647 ;
  assign y2544 = ~n8648 ;
  assign y2545 = n8649 ;
  assign y2546 = n8678 ;
  assign y2547 = ~1'b0 ;
  assign y2548 = n8680 ;
  assign y2549 = ~1'b0 ;
  assign y2550 = n8686 ;
  assign y2551 = n8695 ;
  assign y2552 = ~1'b0 ;
  assign y2553 = ~n8699 ;
  assign y2554 = ~1'b0 ;
  assign y2555 = ~n8704 ;
  assign y2556 = n8713 ;
  assign y2557 = n8718 ;
  assign y2558 = ~n8719 ;
  assign y2559 = ~n8721 ;
  assign y2560 = n8724 ;
  assign y2561 = n8725 ;
  assign y2562 = ~n8732 ;
  assign y2563 = n8733 ;
  assign y2564 = n8744 ;
  assign y2565 = ~n8749 ;
  assign y2566 = n8758 ;
  assign y2567 = ~1'b0 ;
  assign y2568 = ~n8767 ;
  assign y2569 = ~n8769 ;
  assign y2570 = ~n8776 ;
  assign y2571 = ~1'b0 ;
  assign y2572 = ~n8777 ;
  assign y2573 = ~1'b0 ;
  assign y2574 = n8778 ;
  assign y2575 = n8780 ;
  assign y2576 = ~1'b0 ;
  assign y2577 = n8785 ;
  assign y2578 = ~1'b0 ;
  assign y2579 = n8787 ;
  assign y2580 = n8791 ;
  assign y2581 = n8793 ;
  assign y2582 = n8797 ;
  assign y2583 = n8801 ;
  assign y2584 = n7395 ;
  assign y2585 = ~1'b0 ;
  assign y2586 = ~n8809 ;
  assign y2587 = n8816 ;
  assign y2588 = n8823 ;
  assign y2589 = n8825 ;
  assign y2590 = ~n8826 ;
  assign y2591 = n8832 ;
  assign y2592 = n8833 ;
  assign y2593 = n7252 ;
  assign y2594 = n8838 ;
  assign y2595 = n8841 ;
  assign y2596 = ~n8842 ;
  assign y2597 = ~n8844 ;
  assign y2598 = n8847 ;
  assign y2599 = n8849 ;
  assign y2600 = ~n8850 ;
  assign y2601 = ~1'b0 ;
  assign y2602 = ~n8853 ;
  assign y2603 = ~n8856 ;
  assign y2604 = ~n8858 ;
  assign y2605 = n8862 ;
  assign y2606 = ~n8865 ;
  assign y2607 = ~n8866 ;
  assign y2608 = ~n8869 ;
  assign y2609 = ~n8870 ;
  assign y2610 = ~n8875 ;
  assign y2611 = n8877 ;
  assign y2612 = ~n8881 ;
  assign y2613 = ~1'b0 ;
  assign y2614 = ~n8884 ;
  assign y2615 = ~n8886 ;
  assign y2616 = ~n8887 ;
  assign y2617 = n8892 ;
  assign y2618 = ~n8895 ;
  assign y2619 = n8898 ;
  assign y2620 = ~n8899 ;
  assign y2621 = n8906 ;
  assign y2622 = ~n8916 ;
  assign y2623 = n8922 ;
  assign y2624 = n8923 ;
  assign y2625 = ~1'b0 ;
  assign y2626 = n8924 ;
  assign y2627 = ~n8936 ;
  assign y2628 = ~n8943 ;
  assign y2629 = n8951 ;
  assign y2630 = n8956 ;
  assign y2631 = ~n8970 ;
  assign y2632 = n8971 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = ~n8976 ;
  assign y2635 = ~1'b0 ;
  assign y2636 = n8981 ;
  assign y2637 = ~n8983 ;
  assign y2638 = n8984 ;
  assign y2639 = ~n8988 ;
  assign y2640 = ~n9001 ;
  assign y2641 = n9002 ;
  assign y2642 = ~1'b0 ;
  assign y2643 = ~n9004 ;
  assign y2644 = n9008 ;
  assign y2645 = n9012 ;
  assign y2646 = ~n9014 ;
  assign y2647 = n9020 ;
  assign y2648 = ~n9028 ;
  assign y2649 = n9032 ;
  assign y2650 = ~n9034 ;
  assign y2651 = ~n9035 ;
  assign y2652 = ~n9039 ;
  assign y2653 = ~n9048 ;
  assign y2654 = ~n9053 ;
  assign y2655 = ~1'b0 ;
  assign y2656 = ~n9054 ;
  assign y2657 = n9057 ;
  assign y2658 = ~n9059 ;
  assign y2659 = ~1'b0 ;
  assign y2660 = ~1'b0 ;
  assign y2661 = ~1'b0 ;
  assign y2662 = n9061 ;
  assign y2663 = n9063 ;
  assign y2664 = ~n9065 ;
  assign y2665 = ~n9070 ;
  assign y2666 = ~1'b0 ;
  assign y2667 = n9071 ;
  assign y2668 = ~n9076 ;
  assign y2669 = ~n9077 ;
  assign y2670 = ~1'b0 ;
  assign y2671 = n9079 ;
  assign y2672 = ~n9081 ;
  assign y2673 = ~n9088 ;
  assign y2674 = n9091 ;
  assign y2675 = n9095 ;
  assign y2676 = ~n9096 ;
  assign y2677 = ~n9097 ;
  assign y2678 = ~1'b0 ;
  assign y2679 = ~n9105 ;
  assign y2680 = ~n9106 ;
  assign y2681 = ~n9110 ;
  assign y2682 = ~n9114 ;
  assign y2683 = ~1'b0 ;
  assign y2684 = n9122 ;
  assign y2685 = ~n9142 ;
  assign y2686 = n9143 ;
  assign y2687 = ~n9146 ;
  assign y2688 = n9147 ;
  assign y2689 = ~1'b0 ;
  assign y2690 = n9154 ;
  assign y2691 = n9155 ;
  assign y2692 = ~n9158 ;
  assign y2693 = n9162 ;
  assign y2694 = n9163 ;
  assign y2695 = ~1'b0 ;
  assign y2696 = ~n9164 ;
  assign y2697 = ~n9169 ;
  assign y2698 = n9178 ;
  assign y2699 = ~1'b0 ;
  assign y2700 = ~n9184 ;
  assign y2701 = ~n9188 ;
  assign y2702 = 1'b0 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = ~n9196 ;
  assign y2705 = ~1'b0 ;
  assign y2706 = ~n2528 ;
  assign y2707 = n3870 ;
  assign y2708 = n4060 ;
  assign y2709 = n9201 ;
  assign y2710 = n9210 ;
  assign y2711 = ~n9222 ;
  assign y2712 = ~n9230 ;
  assign y2713 = ~1'b0 ;
  assign y2714 = ~n9239 ;
  assign y2715 = ~1'b0 ;
  assign y2716 = ~n9248 ;
  assign y2717 = n9249 ;
  assign y2718 = ~n9251 ;
  assign y2719 = n9254 ;
  assign y2720 = n9257 ;
  assign y2721 = ~n9260 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = ~n9262 ;
  assign y2724 = n9270 ;
  assign y2725 = n9278 ;
  assign y2726 = ~1'b0 ;
  assign y2727 = n9290 ;
  assign y2728 = n9291 ;
  assign y2729 = ~n9292 ;
  assign y2730 = n9301 ;
  assign y2731 = ~1'b0 ;
  assign y2732 = n9314 ;
  assign y2733 = n9316 ;
  assign y2734 = ~n9317 ;
  assign y2735 = ~1'b0 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = ~n9322 ;
  assign y2738 = ~n9323 ;
  assign y2739 = n9325 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = ~n4461 ;
  assign y2742 = ~n9327 ;
  assign y2743 = ~1'b0 ;
  assign y2744 = ~1'b0 ;
  assign y2745 = ~n9332 ;
  assign y2746 = n9334 ;
  assign y2747 = ~n9339 ;
  assign y2748 = n9341 ;
  assign y2749 = ~n9342 ;
  assign y2750 = n9350 ;
  assign y2751 = ~n9356 ;
  assign y2752 = ~n9362 ;
  assign y2753 = n9368 ;
  assign y2754 = ~n9370 ;
  assign y2755 = ~n9376 ;
  assign y2756 = n9380 ;
  assign y2757 = ~1'b0 ;
  assign y2758 = ~n9383 ;
  assign y2759 = ~1'b0 ;
  assign y2760 = ~n9385 ;
  assign y2761 = ~n9386 ;
  assign y2762 = n9393 ;
  assign y2763 = ~n9397 ;
  assign y2764 = n9398 ;
  assign y2765 = n9402 ;
  assign y2766 = n9412 ;
  assign y2767 = ~n9419 ;
  assign y2768 = ~n9422 ;
  assign y2769 = ~n9424 ;
  assign y2770 = n8896 ;
  assign y2771 = n9427 ;
  assign y2772 = ~n9432 ;
  assign y2773 = ~n9434 ;
  assign y2774 = ~n9436 ;
  assign y2775 = ~n9444 ;
  assign y2776 = ~n9448 ;
  assign y2777 = ~n7742 ;
  assign y2778 = ~n9449 ;
  assign y2779 = ~n9450 ;
  assign y2780 = ~n9457 ;
  assign y2781 = ~1'b0 ;
  assign y2782 = ~n9458 ;
  assign y2783 = ~n9460 ;
  assign y2784 = n9461 ;
  assign y2785 = ~n9467 ;
  assign y2786 = ~n9468 ;
  assign y2787 = ~n9472 ;
  assign y2788 = ~n9473 ;
  assign y2789 = ~1'b0 ;
  assign y2790 = ~n9476 ;
  assign y2791 = 1'b0 ;
  assign y2792 = n5470 ;
  assign y2793 = n9480 ;
  assign y2794 = ~n9481 ;
  assign y2795 = n9494 ;
  assign y2796 = ~n9496 ;
  assign y2797 = n9497 ;
  assign y2798 = ~1'b0 ;
  assign y2799 = ~n9498 ;
  assign y2800 = n9500 ;
  assign y2801 = ~n9501 ;
  assign y2802 = n9512 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = ~1'b0 ;
  assign y2805 = n9516 ;
  assign y2806 = ~1'b0 ;
  assign y2807 = ~n9520 ;
  assign y2808 = ~n9522 ;
  assign y2809 = ~n9526 ;
  assign y2810 = ~n9529 ;
  assign y2811 = n9534 ;
  assign y2812 = ~n9536 ;
  assign y2813 = n9544 ;
  assign y2814 = n9545 ;
  assign y2815 = ~n9549 ;
  assign y2816 = n9557 ;
  assign y2817 = ~n9575 ;
  assign y2818 = ~n9578 ;
  assign y2819 = ~n9592 ;
  assign y2820 = n9595 ;
  assign y2821 = ~n9596 ;
  assign y2822 = ~n9597 ;
  assign y2823 = ~n9598 ;
  assign y2824 = ~n9600 ;
  assign y2825 = ~n9607 ;
  assign y2826 = n9611 ;
  assign y2827 = ~n9612 ;
  assign y2828 = ~n9615 ;
  assign y2829 = ~n9616 ;
  assign y2830 = ~n9620 ;
  assign y2831 = ~n9621 ;
  assign y2832 = ~1'b0 ;
  assign y2833 = n9622 ;
  assign y2834 = n9624 ;
  assign y2835 = ~1'b0 ;
  assign y2836 = ~n9631 ;
  assign y2837 = ~n9633 ;
  assign y2838 = n9634 ;
  assign y2839 = n9637 ;
  assign y2840 = ~n9643 ;
  assign y2841 = ~n9151 ;
  assign y2842 = ~n9646 ;
  assign y2843 = ~1'b0 ;
  assign y2844 = ~n9647 ;
  assign y2845 = n9650 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = n9652 ;
  assign y2848 = n9663 ;
  assign y2849 = n9664 ;
  assign y2850 = ~n8422 ;
  assign y2851 = n9665 ;
  assign y2852 = ~n9674 ;
  assign y2853 = ~n9677 ;
  assign y2854 = ~1'b0 ;
  assign y2855 = ~n9678 ;
  assign y2856 = ~n9680 ;
  assign y2857 = n9681 ;
  assign y2858 = ~n9683 ;
  assign y2859 = ~1'b0 ;
  assign y2860 = ~n9688 ;
  assign y2861 = n9691 ;
  assign y2862 = ~n9697 ;
  assign y2863 = n9699 ;
  assign y2864 = ~n5242 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = ~n9703 ;
  assign y2867 = n9711 ;
  assign y2868 = ~n9712 ;
  assign y2869 = ~n9714 ;
  assign y2870 = n9724 ;
  assign y2871 = ~1'b0 ;
  assign y2872 = n9727 ;
  assign y2873 = n9733 ;
  assign y2874 = n9740 ;
  assign y2875 = ~n9751 ;
  assign y2876 = ~n9756 ;
  assign y2877 = ~n9759 ;
  assign y2878 = ~n9761 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~n9770 ;
  assign y2881 = ~n9777 ;
  assign y2882 = n9784 ;
  assign y2883 = ~1'b0 ;
  assign y2884 = ~n9786 ;
  assign y2885 = n9790 ;
  assign y2886 = ~n9793 ;
  assign y2887 = ~n9797 ;
  assign y2888 = ~1'b0 ;
  assign y2889 = n9804 ;
  assign y2890 = ~n9805 ;
  assign y2891 = ~1'b0 ;
  assign y2892 = n9810 ;
  assign y2893 = ~n9814 ;
  assign y2894 = ~n9816 ;
  assign y2895 = ~n9817 ;
  assign y2896 = n9821 ;
  assign y2897 = n9823 ;
  assign y2898 = n9833 ;
  assign y2899 = ~n9840 ;
  assign y2900 = ~n9849 ;
  assign y2901 = ~n9858 ;
  assign y2902 = n9859 ;
  assign y2903 = ~1'b0 ;
  assign y2904 = ~n9861 ;
  assign y2905 = ~n9867 ;
  assign y2906 = n9871 ;
  assign y2907 = n9874 ;
  assign y2908 = ~n9879 ;
  assign y2909 = ~n9882 ;
  assign y2910 = ~1'b0 ;
  assign y2911 = n9888 ;
  assign y2912 = n9889 ;
  assign y2913 = ~n9894 ;
  assign y2914 = ~n9895 ;
  assign y2915 = ~n9896 ;
  assign y2916 = ~n9897 ;
  assign y2917 = ~n9899 ;
  assign y2918 = n9905 ;
  assign y2919 = ~n9909 ;
  assign y2920 = n9914 ;
  assign y2921 = ~n9915 ;
  assign y2922 = n9916 ;
  assign y2923 = n9920 ;
  assign y2924 = n9921 ;
  assign y2925 = ~n9922 ;
  assign y2926 = n9924 ;
  assign y2927 = n9929 ;
  assign y2928 = ~n9931 ;
  assign y2929 = ~n9940 ;
  assign y2930 = ~n9941 ;
  assign y2931 = n9943 ;
  assign y2932 = ~n9944 ;
  assign y2933 = ~1'b0 ;
  assign y2934 = ~n9951 ;
  assign y2935 = ~n9956 ;
  assign y2936 = ~1'b0 ;
  assign y2937 = n9960 ;
  assign y2938 = n9961 ;
  assign y2939 = n9966 ;
  assign y2940 = ~n4860 ;
  assign y2941 = n9971 ;
  assign y2942 = ~n9975 ;
  assign y2943 = ~1'b0 ;
  assign y2944 = ~1'b0 ;
  assign y2945 = ~n9978 ;
  assign y2946 = ~n9981 ;
  assign y2947 = n9986 ;
  assign y2948 = n9995 ;
  assign y2949 = n9996 ;
  assign y2950 = ~n9997 ;
  assign y2951 = ~n10009 ;
  assign y2952 = ~n10012 ;
  assign y2953 = ~n10014 ;
  assign y2954 = ~n10019 ;
  assign y2955 = n10020 ;
  assign y2956 = ~1'b0 ;
  assign y2957 = n10022 ;
  assign y2958 = ~x169 ;
  assign y2959 = ~n10023 ;
  assign y2960 = ~n10024 ;
  assign y2961 = ~n4005 ;
  assign y2962 = ~1'b0 ;
  assign y2963 = n10033 ;
  assign y2964 = n10034 ;
  assign y2965 = n10036 ;
  assign y2966 = n10039 ;
  assign y2967 = ~1'b0 ;
  assign y2968 = ~n10041 ;
  assign y2969 = ~n10044 ;
  assign y2970 = n10045 ;
  assign y2971 = ~n10047 ;
  assign y2972 = n10053 ;
  assign y2973 = ~1'b0 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = ~n1363 ;
  assign y2976 = ~n10057 ;
  assign y2977 = n10058 ;
  assign y2978 = n10060 ;
  assign y2979 = n10066 ;
  assign y2980 = ~n10067 ;
  assign y2981 = n10069 ;
  assign y2982 = ~n10076 ;
  assign y2983 = n10079 ;
  assign y2984 = ~n10080 ;
  assign y2985 = n10083 ;
  assign y2986 = ~n7138 ;
  assign y2987 = ~n10087 ;
  assign y2988 = x3 ;
  assign y2989 = n10088 ;
  assign y2990 = n10089 ;
  assign y2991 = n6708 ;
  assign y2992 = n10090 ;
  assign y2993 = ~n10091 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = ~1'b0 ;
  assign y2996 = ~n10095 ;
  assign y2997 = ~n10096 ;
  assign y2998 = n10109 ;
  assign y2999 = n10113 ;
  assign y3000 = n10126 ;
  assign y3001 = ~n10136 ;
  assign y3002 = n10137 ;
  assign y3003 = ~n10138 ;
  assign y3004 = n10139 ;
  assign y3005 = n10148 ;
  assign y3006 = n10154 ;
  assign y3007 = ~n10155 ;
  assign y3008 = ~1'b0 ;
  assign y3009 = ~n10161 ;
  assign y3010 = ~n9003 ;
  assign y3011 = n10167 ;
  assign y3012 = ~n10171 ;
  assign y3013 = ~n10172 ;
  assign y3014 = ~n10174 ;
  assign y3015 = ~1'b0 ;
  assign y3016 = n10177 ;
  assign y3017 = n10179 ;
  assign y3018 = n10187 ;
  assign y3019 = n10188 ;
  assign y3020 = ~n10193 ;
  assign y3021 = ~n10200 ;
  assign y3022 = n10201 ;
  assign y3023 = ~1'b0 ;
  assign y3024 = n10206 ;
  assign y3025 = ~1'b0 ;
  assign y3026 = ~n10218 ;
  assign y3027 = ~n10220 ;
  assign y3028 = ~1'b0 ;
  assign y3029 = ~n10225 ;
  assign y3030 = ~n10226 ;
  assign y3031 = n10231 ;
  assign y3032 = n10235 ;
  assign y3033 = ~1'b0 ;
  assign y3034 = ~n10236 ;
  assign y3035 = n10240 ;
  assign y3036 = ~n10245 ;
  assign y3037 = ~n10252 ;
  assign y3038 = ~n10255 ;
  assign y3039 = n10261 ;
  assign y3040 = ~1'b0 ;
  assign y3041 = n10270 ;
  assign y3042 = ~1'b0 ;
  assign y3043 = n10273 ;
  assign y3044 = ~n10281 ;
  assign y3045 = ~n10283 ;
  assign y3046 = ~n10286 ;
  assign y3047 = ~n10292 ;
  assign y3048 = ~n10295 ;
  assign y3049 = n10298 ;
  assign y3050 = n3697 ;
  assign y3051 = n10305 ;
  assign y3052 = ~1'b0 ;
  assign y3053 = ~n10307 ;
  assign y3054 = ~n10308 ;
  assign y3055 = ~n10310 ;
  assign y3056 = n10314 ;
  assign y3057 = ~n10316 ;
  assign y3058 = ~n10324 ;
  assign y3059 = ~n10328 ;
  assign y3060 = n10330 ;
  assign y3061 = n10333 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = ~n10347 ;
  assign y3064 = n10348 ;
  assign y3065 = ~n10354 ;
  assign y3066 = ~n10359 ;
  assign y3067 = ~n10360 ;
  assign y3068 = n10361 ;
  assign y3069 = n10364 ;
  assign y3070 = n10365 ;
  assign y3071 = n10373 ;
  assign y3072 = n10378 ;
  assign y3073 = ~n10380 ;
  assign y3074 = n10386 ;
  assign y3075 = n10388 ;
  assign y3076 = n10394 ;
  assign y3077 = ~1'b0 ;
  assign y3078 = ~n10398 ;
  assign y3079 = ~n10401 ;
  assign y3080 = ~1'b0 ;
  assign y3081 = 1'b0 ;
  assign y3082 = n10413 ;
  assign y3083 = n10418 ;
  assign y3084 = ~n10419 ;
  assign y3085 = ~1'b0 ;
  assign y3086 = ~n10425 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~n10434 ;
  assign y3090 = ~n10445 ;
  assign y3091 = ~n10446 ;
  assign y3092 = n10451 ;
  assign y3093 = n10452 ;
  assign y3094 = ~n10460 ;
  assign y3095 = n10464 ;
  assign y3096 = ~n10471 ;
  assign y3097 = ~1'b0 ;
  assign y3098 = n10472 ;
  assign y3099 = n10474 ;
  assign y3100 = ~n10481 ;
  assign y3101 = n10482 ;
  assign y3102 = ~n10487 ;
  assign y3103 = n10488 ;
  assign y3104 = n10489 ;
  assign y3105 = ~1'b0 ;
  assign y3106 = ~n10498 ;
  assign y3107 = n10501 ;
  assign y3108 = ~n10505 ;
  assign y3109 = ~n10506 ;
  assign y3110 = ~n10507 ;
  assign y3111 = n10514 ;
  assign y3112 = ~1'b0 ;
  assign y3113 = n10516 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = n10524 ;
  assign y3116 = 1'b0 ;
  assign y3117 = n8324 ;
  assign y3118 = n10526 ;
  assign y3119 = ~n10528 ;
  assign y3120 = ~n10530 ;
  assign y3121 = ~n10532 ;
  assign y3122 = ~n10545 ;
  assign y3123 = ~n10550 ;
  assign y3124 = ~1'b0 ;
  assign y3125 = n10565 ;
  assign y3126 = ~n10569 ;
  assign y3127 = ~n10575 ;
  assign y3128 = ~n10591 ;
  assign y3129 = n10597 ;
  assign y3130 = n10603 ;
  assign y3131 = n10613 ;
  assign y3132 = ~n10617 ;
  assign y3133 = n10622 ;
  assign y3134 = ~n10624 ;
  assign y3135 = ~n10627 ;
  assign y3136 = n10630 ;
  assign y3137 = n10631 ;
  assign y3138 = n10636 ;
  assign y3139 = ~n10637 ;
  assign y3140 = n10641 ;
  assign y3141 = ~n10646 ;
  assign y3142 = ~1'b0 ;
  assign y3143 = ~1'b0 ;
  assign y3144 = ~n10661 ;
  assign y3145 = ~n10663 ;
  assign y3146 = n10673 ;
  assign y3147 = n10678 ;
  assign y3148 = ~1'b0 ;
  assign y3149 = n10680 ;
  assign y3150 = ~1'b0 ;
  assign y3151 = n10689 ;
  assign y3152 = n10690 ;
  assign y3153 = ~n10699 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = ~n10702 ;
  assign y3156 = ~n10703 ;
  assign y3157 = ~n10710 ;
  assign y3158 = ~n10712 ;
  assign y3159 = n10713 ;
  assign y3160 = ~1'b0 ;
  assign y3161 = ~n10715 ;
  assign y3162 = ~n10723 ;
  assign y3163 = n10724 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = n2573 ;
  assign y3166 = ~n10730 ;
  assign y3167 = ~n10731 ;
  assign y3168 = ~n10735 ;
  assign y3169 = ~n10737 ;
  assign y3170 = ~1'b0 ;
  assign y3171 = n10740 ;
  assign y3172 = ~n10741 ;
  assign y3173 = ~n10742 ;
  assign y3174 = ~n10748 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = n10750 ;
  assign y3177 = n10751 ;
  assign y3178 = n10752 ;
  assign y3179 = n10753 ;
  assign y3180 = ~n10755 ;
  assign y3181 = ~1'b0 ;
  assign y3182 = n10757 ;
  assign y3183 = ~n10759 ;
  assign y3184 = ~1'b0 ;
  assign y3185 = n10767 ;
  assign y3186 = n10770 ;
  assign y3187 = n10775 ;
  assign y3188 = 1'b0 ;
  assign y3189 = n10779 ;
  assign y3190 = n10791 ;
  assign y3191 = ~n10794 ;
  assign y3192 = n10801 ;
  assign y3193 = n10804 ;
  assign y3194 = ~1'b0 ;
  assign y3195 = ~n10806 ;
  assign y3196 = ~1'b0 ;
  assign y3197 = ~1'b0 ;
  assign y3198 = ~n10810 ;
  assign y3199 = ~n10811 ;
  assign y3200 = n10813 ;
  assign y3201 = n10822 ;
  assign y3202 = n10823 ;
  assign y3203 = n10824 ;
  assign y3204 = ~n10826 ;
  assign y3205 = ~1'b0 ;
  assign y3206 = ~n10831 ;
  assign y3207 = ~n10836 ;
  assign y3208 = ~n10838 ;
  assign y3209 = ~n10839 ;
  assign y3210 = ~1'b0 ;
  assign y3211 = ~1'b0 ;
  assign y3212 = ~n10843 ;
  assign y3213 = ~n10852 ;
  assign y3214 = ~1'b0 ;
  assign y3215 = ~n10854 ;
  assign y3216 = ~1'b0 ;
  assign y3217 = 1'b0 ;
  assign y3218 = ~n10857 ;
  assign y3219 = ~n10858 ;
  assign y3220 = ~n10860 ;
  assign y3221 = n10872 ;
  assign y3222 = ~1'b0 ;
  assign y3223 = n10873 ;
  assign y3224 = n10878 ;
  assign y3225 = ~n10880 ;
  assign y3226 = ~n10881 ;
  assign y3227 = n1108 ;
  assign y3228 = ~n10882 ;
  assign y3229 = ~n10883 ;
  assign y3230 = ~n10884 ;
  assign y3231 = n10885 ;
  assign y3232 = n10891 ;
  assign y3233 = ~n10893 ;
  assign y3234 = ~n10902 ;
  assign y3235 = n10908 ;
  assign y3236 = ~n10909 ;
  assign y3237 = ~n10910 ;
  assign y3238 = ~n10913 ;
  assign y3239 = n10920 ;
  assign y3240 = n10922 ;
  assign y3241 = n10925 ;
  assign y3242 = ~n10929 ;
  assign y3243 = n10941 ;
  assign y3244 = ~n10942 ;
  assign y3245 = ~n10949 ;
  assign y3246 = ~n10952 ;
  assign y3247 = n10958 ;
  assign y3248 = n10960 ;
  assign y3249 = ~1'b0 ;
  assign y3250 = n10967 ;
  assign y3251 = n10971 ;
  assign y3252 = ~n10972 ;
  assign y3253 = ~n10973 ;
  assign y3254 = n10974 ;
  assign y3255 = n10994 ;
  assign y3256 = ~n11000 ;
  assign y3257 = ~n11001 ;
  assign y3258 = n11003 ;
  assign y3259 = ~1'b0 ;
  assign y3260 = n11005 ;
  assign y3261 = n11009 ;
  assign y3262 = ~n11026 ;
  assign y3263 = ~1'b0 ;
  assign y3264 = ~n11031 ;
  assign y3265 = n11032 ;
  assign y3266 = ~n11035 ;
  assign y3267 = ~n11047 ;
  assign y3268 = ~n11050 ;
  assign y3269 = n11051 ;
  assign y3270 = n11059 ;
  assign y3271 = n11061 ;
  assign y3272 = ~n11062 ;
  assign y3273 = n11064 ;
  assign y3274 = n11068 ;
  assign y3275 = n11069 ;
  assign y3276 = ~n11070 ;
  assign y3277 = ~n11072 ;
  assign y3278 = ~1'b0 ;
  assign y3279 = n11081 ;
  assign y3280 = n11083 ;
  assign y3281 = ~n11092 ;
  assign y3282 = n11096 ;
  assign y3283 = ~n11100 ;
  assign y3284 = ~n11102 ;
  assign y3285 = n11108 ;
  assign y3286 = ~1'b0 ;
  assign y3287 = n11116 ;
  assign y3288 = ~n11126 ;
  assign y3289 = ~n11135 ;
  assign y3290 = ~n11138 ;
  assign y3291 = n11139 ;
  assign y3292 = ~n11144 ;
  assign y3293 = n11149 ;
  assign y3294 = ~1'b0 ;
  assign y3295 = ~n11151 ;
  assign y3296 = n11158 ;
  assign y3297 = ~n11159 ;
  assign y3298 = n11162 ;
  assign y3299 = n11169 ;
  assign y3300 = n11174 ;
  assign y3301 = ~n11181 ;
  assign y3302 = n11183 ;
  assign y3303 = ~n11187 ;
  assign y3304 = n11190 ;
  assign y3305 = ~n11204 ;
  assign y3306 = n11206 ;
  assign y3307 = ~n11207 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = ~n11211 ;
  assign y3310 = n11216 ;
  assign y3311 = ~n11217 ;
  assign y3312 = n11219 ;
  assign y3313 = n11221 ;
  assign y3314 = n11223 ;
  assign y3315 = ~n11226 ;
  assign y3316 = ~n11230 ;
  assign y3317 = n11233 ;
  assign y3318 = n11245 ;
  assign y3319 = ~n11249 ;
  assign y3320 = ~n11250 ;
  assign y3321 = n11258 ;
  assign y3322 = ~n11260 ;
  assign y3323 = ~1'b0 ;
  assign y3324 = n11261 ;
  assign y3325 = n11263 ;
  assign y3326 = ~1'b0 ;
  assign y3327 = ~n11267 ;
  assign y3328 = ~n11269 ;
  assign y3329 = ~n11271 ;
  assign y3330 = ~1'b0 ;
  assign y3331 = ~1'b0 ;
  assign y3332 = n11272 ;
  assign y3333 = ~n11277 ;
  assign y3334 = ~n11280 ;
  assign y3335 = ~n11283 ;
  assign y3336 = ~n11284 ;
  assign y3337 = ~n11287 ;
  assign y3338 = ~1'b0 ;
  assign y3339 = ~n11288 ;
  assign y3340 = n11290 ;
  assign y3341 = n11292 ;
  assign y3342 = ~n11293 ;
  assign y3343 = ~n11299 ;
  assign y3344 = ~n11310 ;
  assign y3345 = ~n11312 ;
  assign y3346 = ~n11313 ;
  assign y3347 = n11315 ;
  assign y3348 = n11323 ;
  assign y3349 = n11326 ;
  assign y3350 = n11339 ;
  assign y3351 = ~n11341 ;
  assign y3352 = ~n11343 ;
  assign y3353 = ~1'b0 ;
  assign y3354 = n11347 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = n11348 ;
  assign y3357 = n11360 ;
  assign y3358 = n11366 ;
  assign y3359 = ~n11371 ;
  assign y3360 = ~1'b0 ;
  assign y3361 = ~n11379 ;
  assign y3362 = ~1'b0 ;
  assign y3363 = n11382 ;
  assign y3364 = n11383 ;
  assign y3365 = n11385 ;
  assign y3366 = n11386 ;
  assign y3367 = n11392 ;
  assign y3368 = n11394 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = n11398 ;
  assign y3371 = n11401 ;
  assign y3372 = ~n11407 ;
  assign y3373 = ~n11417 ;
  assign y3374 = n11418 ;
  assign y3375 = n11424 ;
  assign y3376 = ~n11426 ;
  assign y3377 = n11433 ;
  assign y3378 = n6721 ;
  assign y3379 = n11435 ;
  assign y3380 = ~1'b0 ;
  assign y3381 = ~n11437 ;
  assign y3382 = ~n11440 ;
  assign y3383 = n11441 ;
  assign y3384 = n11448 ;
  assign y3385 = ~n11449 ;
  assign y3386 = n11458 ;
  assign y3387 = ~1'b0 ;
  assign y3388 = n11461 ;
  assign y3389 = ~n11462 ;
  assign y3390 = ~n11466 ;
  assign y3391 = n11468 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = ~n11475 ;
  assign y3394 = n11479 ;
  assign y3395 = ~n11484 ;
  assign y3396 = ~n11486 ;
  assign y3397 = ~1'b0 ;
  assign y3398 = n11489 ;
  assign y3399 = ~n11496 ;
  assign y3400 = ~n11498 ;
  assign y3401 = ~n11500 ;
  assign y3402 = ~n11502 ;
  assign y3403 = n11505 ;
  assign y3404 = ~n11506 ;
  assign y3405 = n11510 ;
  assign y3406 = ~n11515 ;
  assign y3407 = ~n11518 ;
  assign y3408 = n11525 ;
  assign y3409 = ~n11528 ;
  assign y3410 = ~1'b0 ;
  assign y3411 = ~n11533 ;
  assign y3412 = ~n11537 ;
  assign y3413 = ~n11541 ;
  assign y3414 = n11544 ;
  assign y3415 = n11548 ;
  assign y3416 = 1'b0 ;
  assign y3417 = ~n11553 ;
  assign y3418 = ~1'b0 ;
  assign y3419 = n11554 ;
  assign y3420 = ~n11557 ;
  assign y3421 = ~n11561 ;
  assign y3422 = ~n11565 ;
  assign y3423 = ~n11568 ;
  assign y3424 = ~n11571 ;
  assign y3425 = n11572 ;
  assign y3426 = ~n11578 ;
  assign y3427 = n11583 ;
  assign y3428 = ~1'b0 ;
  assign y3429 = ~n11585 ;
  assign y3430 = n11588 ;
  assign y3431 = ~n11598 ;
  assign y3432 = n11600 ;
  assign y3433 = ~n11605 ;
  assign y3434 = ~n11607 ;
  assign y3435 = n11619 ;
  assign y3436 = ~1'b0 ;
  assign y3437 = n11621 ;
  assign y3438 = ~n11623 ;
  assign y3439 = n11625 ;
  assign y3440 = n11628 ;
  assign y3441 = ~n11629 ;
  assign y3442 = ~1'b0 ;
  assign y3443 = ~n11643 ;
  assign y3444 = ~n11651 ;
  assign y3445 = n11653 ;
  assign y3446 = ~n11662 ;
  assign y3447 = n11664 ;
  assign y3448 = n11669 ;
  assign y3449 = n11670 ;
  assign y3450 = n11672 ;
  assign y3451 = n11673 ;
  assign y3452 = ~n11674 ;
  assign y3453 = ~n11679 ;
  assign y3454 = ~n11680 ;
  assign y3455 = n11681 ;
  assign y3456 = ~n11684 ;
  assign y3457 = n11690 ;
  assign y3458 = ~n11693 ;
  assign y3459 = ~n11694 ;
  assign y3460 = n11698 ;
  assign y3461 = ~n11713 ;
  assign y3462 = n11720 ;
  assign y3463 = ~n11724 ;
  assign y3464 = n11732 ;
  assign y3465 = ~n11734 ;
  assign y3466 = n11738 ;
  assign y3467 = n11744 ;
  assign y3468 = ~n11745 ;
  assign y3469 = n11750 ;
  assign y3470 = ~n11756 ;
  assign y3471 = ~n11764 ;
  assign y3472 = n11773 ;
  assign y3473 = ~n11776 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = ~n11780 ;
  assign y3476 = 1'b0 ;
  assign y3477 = n11781 ;
  assign y3478 = ~n11785 ;
  assign y3479 = ~n11786 ;
  assign y3480 = ~n11787 ;
  assign y3481 = ~n11791 ;
  assign y3482 = ~n11803 ;
  assign y3483 = n11809 ;
  assign y3484 = n11810 ;
  assign y3485 = n11814 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = ~n11817 ;
  assign y3488 = ~1'b0 ;
  assign y3489 = ~n11823 ;
  assign y3490 = ~n11827 ;
  assign y3491 = ~n11828 ;
  assign y3492 = n11840 ;
  assign y3493 = ~n11842 ;
  assign y3494 = n11845 ;
  assign y3495 = ~n11851 ;
  assign y3496 = ~n11857 ;
  assign y3497 = ~n11865 ;
  assign y3498 = ~n11871 ;
  assign y3499 = ~n11873 ;
  assign y3500 = n11878 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = n11880 ;
  assign y3503 = ~n11881 ;
  assign y3504 = ~n11883 ;
  assign y3505 = ~n11885 ;
  assign y3506 = ~n11888 ;
  assign y3507 = n11889 ;
  assign y3508 = ~n11896 ;
  assign y3509 = n11897 ;
  assign y3510 = n11902 ;
  assign y3511 = n11905 ;
  assign y3512 = n11912 ;
  assign y3513 = n11917 ;
  assign y3514 = n11932 ;
  assign y3515 = ~n11934 ;
  assign y3516 = ~1'b0 ;
  assign y3517 = ~n11936 ;
  assign y3518 = ~n11943 ;
  assign y3519 = n11949 ;
  assign y3520 = ~1'b0 ;
  assign y3521 = ~n11951 ;
  assign y3522 = ~n11957 ;
  assign y3523 = ~n11963 ;
  assign y3524 = ~n11964 ;
  assign y3525 = ~n11965 ;
  assign y3526 = ~n11968 ;
  assign y3527 = ~n11969 ;
  assign y3528 = ~n11978 ;
  assign y3529 = ~n11980 ;
  assign y3530 = ~n11984 ;
  assign y3531 = ~1'b0 ;
  assign y3532 = n11986 ;
  assign y3533 = n11988 ;
  assign y3534 = n11989 ;
  assign y3535 = ~n11992 ;
  assign y3536 = n11993 ;
  assign y3537 = ~n11996 ;
  assign y3538 = n12001 ;
  assign y3539 = ~n12008 ;
  assign y3540 = ~1'b0 ;
  assign y3541 = n12009 ;
  assign y3542 = ~n12010 ;
  assign y3543 = n12016 ;
  assign y3544 = ~1'b0 ;
  assign y3545 = n12018 ;
  assign y3546 = ~1'b0 ;
  assign y3547 = ~n12019 ;
  assign y3548 = ~n12021 ;
  assign y3549 = n12024 ;
  assign y3550 = ~n12030 ;
  assign y3551 = ~1'b0 ;
  assign y3552 = n12032 ;
  assign y3553 = ~n12035 ;
  assign y3554 = ~n12037 ;
  assign y3555 = ~n12040 ;
  assign y3556 = ~n12042 ;
  assign y3557 = ~n12043 ;
  assign y3558 = n12047 ;
  assign y3559 = n12052 ;
  assign y3560 = n12058 ;
  assign y3561 = ~1'b0 ;
  assign y3562 = n12061 ;
  assign y3563 = ~1'b0 ;
  assign y3564 = ~n12067 ;
  assign y3565 = ~n12072 ;
  assign y3566 = n12073 ;
  assign y3567 = ~n12076 ;
  assign y3568 = n12077 ;
  assign y3569 = ~1'b0 ;
  assign y3570 = n12078 ;
  assign y3571 = n409 ;
  assign y3572 = n12083 ;
  assign y3573 = ~n12085 ;
  assign y3574 = n12090 ;
  assign y3575 = ~n12103 ;
  assign y3576 = ~n12104 ;
  assign y3577 = n12105 ;
  assign y3578 = n12118 ;
  assign y3579 = n12120 ;
  assign y3580 = n7047 ;
  assign y3581 = n12122 ;
  assign y3582 = n12124 ;
  assign y3583 = n12126 ;
  assign y3584 = n12127 ;
  assign y3585 = ~n12131 ;
  assign y3586 = ~n12140 ;
  assign y3587 = ~n12148 ;
  assign y3588 = ~1'b0 ;
  assign y3589 = ~1'b0 ;
  assign y3590 = n12154 ;
  assign y3591 = ~n12155 ;
  assign y3592 = n12160 ;
  assign y3593 = n12162 ;
  assign y3594 = ~1'b0 ;
  assign y3595 = ~n12167 ;
  assign y3596 = ~n12171 ;
  assign y3597 = ~n12173 ;
  assign y3598 = n12176 ;
  assign y3599 = n12181 ;
  assign y3600 = n12183 ;
  assign y3601 = ~n12188 ;
  assign y3602 = ~n12197 ;
  assign y3603 = ~n12201 ;
  assign y3604 = ~1'b0 ;
  assign y3605 = ~n12204 ;
  assign y3606 = n12212 ;
  assign y3607 = n12213 ;
  assign y3608 = n12216 ;
  assign y3609 = n12221 ;
  assign y3610 = n12223 ;
  assign y3611 = ~n12225 ;
  assign y3612 = n12229 ;
  assign y3613 = ~n12239 ;
  assign y3614 = n12246 ;
  assign y3615 = ~n12256 ;
  assign y3616 = ~n12258 ;
  assign y3617 = ~n12261 ;
  assign y3618 = ~n12265 ;
  assign y3619 = ~1'b0 ;
  assign y3620 = n12267 ;
  assign y3621 = ~n12274 ;
  assign y3622 = ~n12283 ;
  assign y3623 = n12285 ;
  assign y3624 = ~1'b0 ;
  assign y3625 = ~n12288 ;
  assign y3626 = ~1'b0 ;
  assign y3627 = ~n12300 ;
  assign y3628 = ~n12302 ;
  assign y3629 = n12309 ;
  assign y3630 = n12315 ;
  assign y3631 = n12322 ;
  assign y3632 = ~n12325 ;
  assign y3633 = ~n12326 ;
  assign y3634 = ~n12336 ;
  assign y3635 = ~1'b0 ;
  assign y3636 = n12338 ;
  assign y3637 = ~n12339 ;
  assign y3638 = ~n12345 ;
  assign y3639 = ~n12350 ;
  assign y3640 = n12355 ;
  assign y3641 = n12364 ;
  assign y3642 = ~1'b0 ;
  assign y3643 = ~1'b0 ;
  assign y3644 = n12368 ;
  assign y3645 = n12371 ;
  assign y3646 = ~n12374 ;
  assign y3647 = n12389 ;
  assign y3648 = n12391 ;
  assign y3649 = n12393 ;
  assign y3650 = n12397 ;
  assign y3651 = ~n12403 ;
  assign y3652 = n12404 ;
  assign y3653 = n12409 ;
  assign y3654 = ~n12413 ;
  assign y3655 = n12421 ;
  assign y3656 = n12422 ;
  assign y3657 = ~n12432 ;
  assign y3658 = n12436 ;
  assign y3659 = n12438 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = ~n12439 ;
  assign y3662 = n6433 ;
  assign y3663 = ~1'b0 ;
  assign y3664 = n12441 ;
  assign y3665 = n12443 ;
  assign y3666 = ~n12444 ;
  assign y3667 = ~n12446 ;
  assign y3668 = n12447 ;
  assign y3669 = ~n12449 ;
  assign y3670 = ~1'b0 ;
  assign y3671 = ~n12452 ;
  assign y3672 = ~1'b0 ;
  assign y3673 = ~n12455 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = ~n12459 ;
  assign y3676 = ~n12466 ;
  assign y3677 = n12474 ;
  assign y3678 = ~n12476 ;
  assign y3679 = ~n12484 ;
  assign y3680 = n12489 ;
  assign y3681 = n12506 ;
  assign y3682 = ~1'b0 ;
  assign y3683 = ~n12507 ;
  assign y3684 = n12508 ;
  assign y3685 = n12512 ;
  assign y3686 = n12516 ;
  assign y3687 = ~1'b0 ;
  assign y3688 = n12519 ;
  assign y3689 = n12521 ;
  assign y3690 = ~n12524 ;
  assign y3691 = ~1'b0 ;
  assign y3692 = ~n12537 ;
  assign y3693 = ~n12540 ;
  assign y3694 = n12560 ;
  assign y3695 = ~n12561 ;
  assign y3696 = ~n12565 ;
  assign y3697 = n12571 ;
  assign y3698 = n12572 ;
  assign y3699 = n12575 ;
  assign y3700 = ~n12582 ;
  assign y3701 = ~n12585 ;
  assign y3702 = ~n12586 ;
  assign y3703 = ~1'b0 ;
  assign y3704 = n12597 ;
  assign y3705 = ~1'b0 ;
  assign y3706 = ~n12599 ;
  assign y3707 = n12604 ;
  assign y3708 = n12609 ;
  assign y3709 = ~n12611 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = ~1'b0 ;
  assign y3712 = ~n12613 ;
  assign y3713 = ~1'b0 ;
  assign y3714 = ~n12616 ;
  assign y3715 = ~n12618 ;
  assign y3716 = ~n12619 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = ~1'b0 ;
  assign y3719 = ~1'b0 ;
  assign y3720 = n12622 ;
  assign y3721 = ~n12626 ;
  assign y3722 = ~n12628 ;
  assign y3723 = n12630 ;
  assign y3724 = ~n12636 ;
  assign y3725 = n12639 ;
  assign y3726 = n12644 ;
  assign y3727 = ~1'b0 ;
  assign y3728 = ~n12645 ;
  assign y3729 = n12647 ;
  assign y3730 = n12656 ;
  assign y3731 = ~n12657 ;
  assign y3732 = ~n12658 ;
  assign y3733 = n12661 ;
  assign y3734 = ~n12663 ;
  assign y3735 = n12665 ;
  assign y3736 = ~n12674 ;
  assign y3737 = ~1'b0 ;
  assign y3738 = n12679 ;
  assign y3739 = n12686 ;
  assign y3740 = ~n12692 ;
  assign y3741 = ~n12699 ;
  assign y3742 = n12706 ;
  assign y3743 = ~n12707 ;
  assign y3744 = ~n12711 ;
  assign y3745 = n12714 ;
  assign y3746 = n12717 ;
  assign y3747 = n12719 ;
  assign y3748 = ~n12721 ;
  assign y3749 = ~n12725 ;
  assign y3750 = n12730 ;
  assign y3751 = n12735 ;
  assign y3752 = n12737 ;
  assign y3753 = n12739 ;
  assign y3754 = ~1'b0 ;
  assign y3755 = ~n12744 ;
  assign y3756 = n12746 ;
  assign y3757 = ~n12747 ;
  assign y3758 = n12753 ;
  assign y3759 = ~n12754 ;
  assign y3760 = n12755 ;
  assign y3761 = ~n12762 ;
  assign y3762 = n12763 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = ~1'b0 ;
  assign y3765 = n12767 ;
  assign y3766 = ~1'b0 ;
  assign y3767 = ~n12769 ;
  assign y3768 = n12771 ;
  assign y3769 = ~n12781 ;
  assign y3770 = ~1'b0 ;
  assign y3771 = ~n12783 ;
  assign y3772 = ~n12784 ;
  assign y3773 = n12785 ;
  assign y3774 = n12793 ;
  assign y3775 = n12797 ;
  assign y3776 = ~n12801 ;
  assign y3777 = ~n12807 ;
  assign y3778 = n12812 ;
  assign y3779 = n12822 ;
  assign y3780 = ~n12830 ;
  assign y3781 = n12832 ;
  assign y3782 = n12834 ;
  assign y3783 = ~n12845 ;
  assign y3784 = n12850 ;
  assign y3785 = ~1'b0 ;
  assign y3786 = ~n12851 ;
  assign y3787 = n12853 ;
  assign y3788 = ~n12855 ;
  assign y3789 = ~1'b0 ;
  assign y3790 = ~1'b0 ;
  assign y3791 = n12857 ;
  assign y3792 = ~n12860 ;
  assign y3793 = ~n10007 ;
  assign y3794 = n12866 ;
  assign y3795 = n12867 ;
  assign y3796 = n12868 ;
  assign y3797 = ~n12871 ;
  assign y3798 = ~n12874 ;
  assign y3799 = n12875 ;
  assign y3800 = n12880 ;
  assign y3801 = ~1'b0 ;
  assign y3802 = ~1'b0 ;
  assign y3803 = ~n12884 ;
  assign y3804 = ~1'b0 ;
  assign y3805 = ~n12886 ;
  assign y3806 = n12888 ;
  assign y3807 = ~n12903 ;
  assign y3808 = n12905 ;
  assign y3809 = ~n12909 ;
  assign y3810 = ~n12912 ;
  assign y3811 = ~n12913 ;
  assign y3812 = ~n12917 ;
  assign y3813 = ~n12924 ;
  assign y3814 = ~n12928 ;
  assign y3815 = ~n12934 ;
  assign y3816 = ~n12936 ;
  assign y3817 = ~n4307 ;
  assign y3818 = ~n12938 ;
  assign y3819 = ~n12939 ;
  assign y3820 = ~n12943 ;
  assign y3821 = ~n12947 ;
  assign y3822 = n12948 ;
  assign y3823 = ~n12953 ;
  assign y3824 = n12954 ;
  assign y3825 = n12959 ;
  assign y3826 = ~n12962 ;
  assign y3827 = ~n12965 ;
  assign y3828 = n12969 ;
  assign y3829 = ~n12970 ;
  assign y3830 = n12972 ;
  assign y3831 = n12981 ;
  assign y3832 = n12985 ;
  assign y3833 = ~n12988 ;
  assign y3834 = ~n12998 ;
  assign y3835 = n12999 ;
  assign y3836 = n13003 ;
  assign y3837 = n13007 ;
  assign y3838 = ~n13010 ;
  assign y3839 = n13011 ;
  assign y3840 = ~n13015 ;
  assign y3841 = n13016 ;
  assign y3842 = ~n13018 ;
  assign y3843 = ~n13033 ;
  assign y3844 = ~n13038 ;
  assign y3845 = ~n13041 ;
  assign y3846 = ~n13045 ;
  assign y3847 = n13062 ;
  assign y3848 = ~1'b0 ;
  assign y3849 = ~n13064 ;
  assign y3850 = ~n13071 ;
  assign y3851 = ~1'b0 ;
  assign y3852 = ~n13079 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = ~n13084 ;
  assign y3855 = ~n13085 ;
  assign y3856 = n13088 ;
  assign y3857 = ~n13089 ;
  assign y3858 = ~1'b0 ;
  assign y3859 = ~1'b0 ;
  assign y3860 = ~n13091 ;
  assign y3861 = n13103 ;
  assign y3862 = ~1'b0 ;
  assign y3863 = ~1'b0 ;
  assign y3864 = n13104 ;
  assign y3865 = n13109 ;
  assign y3866 = n261 ;
  assign y3867 = n13110 ;
  assign y3868 = ~n13111 ;
  assign y3869 = ~n13113 ;
  assign y3870 = ~n13114 ;
  assign y3871 = ~n13118 ;
  assign y3872 = n13123 ;
  assign y3873 = ~n13125 ;
  assign y3874 = ~n13129 ;
  assign y3875 = ~n13130 ;
  assign y3876 = n13131 ;
  assign y3877 = ~n13137 ;
  assign y3878 = n13138 ;
  assign y3879 = ~n13139 ;
  assign y3880 = n13143 ;
  assign y3881 = n13146 ;
  assign y3882 = n13150 ;
  assign y3883 = n13152 ;
  assign y3884 = n13156 ;
  assign y3885 = n13157 ;
  assign y3886 = ~n13161 ;
  assign y3887 = ~n13162 ;
  assign y3888 = n13163 ;
  assign y3889 = ~n13164 ;
  assign y3890 = ~1'b0 ;
  assign y3891 = n13165 ;
  assign y3892 = ~n13170 ;
  assign y3893 = 1'b0 ;
  assign y3894 = n13176 ;
  assign y3895 = ~n13180 ;
  assign y3896 = ~n13186 ;
  assign y3897 = ~n13188 ;
  assign y3898 = ~n13192 ;
  assign y3899 = ~1'b0 ;
  assign y3900 = n13195 ;
  assign y3901 = n13196 ;
  assign y3902 = ~1'b0 ;
  assign y3903 = ~1'b0 ;
  assign y3904 = ~1'b0 ;
  assign y3905 = n13199 ;
  assign y3906 = ~n13201 ;
  assign y3907 = n13203 ;
  assign y3908 = n13206 ;
  assign y3909 = ~n13207 ;
  assign y3910 = n13209 ;
  assign y3911 = ~n13212 ;
  assign y3912 = n13214 ;
  assign y3913 = ~n13218 ;
  assign y3914 = n13219 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = n13222 ;
  assign y3917 = ~1'b0 ;
  assign y3918 = ~n13225 ;
  assign y3919 = ~n13231 ;
  assign y3920 = ~1'b0 ;
  assign y3921 = n13234 ;
  assign y3922 = n13240 ;
  assign y3923 = ~n13246 ;
  assign y3924 = ~n13258 ;
  assign y3925 = n13259 ;
  assign y3926 = n13266 ;
  assign y3927 = n13268 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = n13273 ;
  assign y3931 = n13277 ;
  assign y3932 = n13287 ;
  assign y3933 = ~1'b0 ;
  assign y3934 = n13290 ;
  assign y3935 = n13294 ;
  assign y3936 = n13297 ;
  assign y3937 = n13299 ;
  assign y3938 = ~n13313 ;
  assign y3939 = ~n13322 ;
  assign y3940 = n13323 ;
  assign y3941 = n13324 ;
  assign y3942 = ~1'b0 ;
  assign y3943 = n13327 ;
  assign y3944 = ~1'b0 ;
  assign y3945 = ~n13328 ;
  assign y3946 = n13332 ;
  assign y3947 = n13338 ;
  assign y3948 = n13340 ;
  assign y3949 = ~n4095 ;
  assign y3950 = ~n13344 ;
  assign y3951 = n11533 ;
  assign y3952 = ~n13349 ;
  assign y3953 = ~n13352 ;
  assign y3954 = ~n13359 ;
  assign y3955 = ~n13364 ;
  assign y3956 = ~1'b0 ;
  assign y3957 = ~1'b0 ;
  assign y3958 = n13365 ;
  assign y3959 = n13369 ;
  assign y3960 = ~n13371 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = ~1'b0 ;
  assign y3963 = ~1'b0 ;
  assign y3964 = ~n13373 ;
  assign y3965 = ~n13377 ;
  assign y3966 = ~n13382 ;
  assign y3967 = n13387 ;
  assign y3968 = n13391 ;
  assign y3969 = n13393 ;
  assign y3970 = n13401 ;
  assign y3971 = ~n13402 ;
  assign y3972 = n13404 ;
  assign y3973 = n13414 ;
  assign y3974 = ~n13417 ;
  assign y3975 = ~n13422 ;
  assign y3976 = n13425 ;
  assign y3977 = ~1'b0 ;
  assign y3978 = n13427 ;
  assign y3979 = n13432 ;
  assign y3980 = ~n13434 ;
  assign y3981 = n13436 ;
  assign y3982 = ~n13444 ;
  assign y3983 = ~n13445 ;
  assign y3984 = n1912 ;
  assign y3985 = ~n13448 ;
  assign y3986 = n13449 ;
  assign y3987 = ~1'b0 ;
  assign y3988 = ~n13454 ;
  assign y3989 = ~n13463 ;
  assign y3990 = n13464 ;
  assign y3991 = ~n13468 ;
  assign y3992 = ~n13473 ;
  assign y3993 = ~1'b0 ;
  assign y3994 = n13474 ;
  assign y3995 = ~1'b0 ;
  assign y3996 = n13476 ;
  assign y3997 = n13479 ;
  assign y3998 = ~1'b0 ;
  assign y3999 = n13482 ;
  assign y4000 = n13487 ;
  assign y4001 = ~n13488 ;
  assign y4002 = ~n13495 ;
  assign y4003 = n13496 ;
  assign y4004 = n13500 ;
  assign y4005 = n13501 ;
  assign y4006 = n13505 ;
  assign y4007 = ~n13507 ;
  assign y4008 = n13508 ;
  assign y4009 = n13512 ;
  assign y4010 = ~n13513 ;
  assign y4011 = ~1'b0 ;
  assign y4012 = n13520 ;
  assign y4013 = n13525 ;
  assign y4014 = ~n13540 ;
  assign y4015 = n13546 ;
  assign y4016 = n13551 ;
  assign y4017 = n13552 ;
  assign y4018 = ~n13553 ;
  assign y4019 = ~n13559 ;
  assign y4020 = n13564 ;
  assign y4021 = n13567 ;
  assign y4022 = ~n13570 ;
  assign y4023 = ~n13572 ;
  assign y4024 = ~n13577 ;
  assign y4025 = ~n13580 ;
  assign y4026 = n13590 ;
  assign y4027 = ~n13596 ;
  assign y4028 = ~n13597 ;
  assign y4029 = ~n13600 ;
  assign y4030 = ~n13603 ;
  assign y4031 = ~1'b0 ;
  assign y4032 = ~n13604 ;
  assign y4033 = n13609 ;
  assign y4034 = ~n13612 ;
  assign y4035 = n13617 ;
  assign y4036 = ~n13625 ;
  assign y4037 = ~n13629 ;
  assign y4038 = ~n13631 ;
  assign y4039 = ~n13633 ;
  assign y4040 = n13636 ;
  assign y4041 = ~1'b0 ;
  assign y4042 = ~n13641 ;
  assign y4043 = n13643 ;
  assign y4044 = ~1'b0 ;
  assign y4045 = ~n13645 ;
  assign y4046 = ~n13651 ;
  assign y4047 = ~n13653 ;
  assign y4048 = ~1'b0 ;
  assign y4049 = ~n13659 ;
  assign y4050 = n13661 ;
  assign y4051 = ~n13662 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = ~1'b0 ;
  assign y4054 = ~n13669 ;
  assign y4055 = ~n13674 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = n13675 ;
  assign y4058 = ~n13681 ;
  assign y4059 = ~n13689 ;
  assign y4060 = ~n13691 ;
  assign y4061 = n13695 ;
  assign y4062 = n13701 ;
  assign y4063 = n13703 ;
  assign y4064 = ~n13704 ;
  assign y4065 = n13712 ;
  assign y4066 = n13714 ;
  assign y4067 = ~1'b0 ;
  assign y4068 = ~n13723 ;
  assign y4069 = ~n13725 ;
  assign y4070 = ~n13726 ;
  assign y4071 = ~n13728 ;
  assign y4072 = n13729 ;
  assign y4073 = n13745 ;
  assign y4074 = ~1'b0 ;
  assign y4075 = ~1'b0 ;
  assign y4076 = ~1'b0 ;
  assign y4077 = n13751 ;
  assign y4078 = n13759 ;
  assign y4079 = ~n13763 ;
  assign y4080 = ~n13774 ;
  assign y4081 = ~1'b0 ;
  assign y4082 = ~n13781 ;
  assign y4083 = ~1'b0 ;
  assign y4084 = ~1'b0 ;
  assign y4085 = ~1'b0 ;
  assign y4086 = n13783 ;
  assign y4087 = n13786 ;
  assign y4088 = n13791 ;
  assign y4089 = n13798 ;
  assign y4090 = n7190 ;
  assign y4091 = ~1'b0 ;
  assign y4092 = n13801 ;
  assign y4093 = ~1'b0 ;
  assign y4094 = ~n13803 ;
  assign y4095 = ~n13807 ;
  assign y4096 = ~1'b0 ;
  assign y4097 = ~1'b0 ;
  assign y4098 = ~n13811 ;
  assign y4099 = ~1'b0 ;
  assign y4100 = ~1'b0 ;
  assign y4101 = ~n13813 ;
  assign y4102 = ~n13815 ;
  assign y4103 = ~1'b0 ;
  assign y4104 = n13820 ;
  assign y4105 = n13835 ;
  assign y4106 = n13836 ;
  assign y4107 = ~n13838 ;
  assign y4108 = ~n13840 ;
  assign y4109 = n13842 ;
  assign y4110 = ~n13846 ;
  assign y4111 = ~n13848 ;
  assign y4112 = ~n13849 ;
  assign y4113 = ~1'b0 ;
  assign y4114 = n13851 ;
  assign y4115 = ~1'b0 ;
  assign y4116 = ~n13852 ;
  assign y4117 = n13853 ;
  assign y4118 = n13854 ;
  assign y4119 = ~n13855 ;
  assign y4120 = n13870 ;
  assign y4121 = n13874 ;
  assign y4122 = ~n13877 ;
  assign y4123 = ~1'b0 ;
  assign y4124 = ~n13878 ;
  assign y4125 = n13881 ;
  assign y4126 = ~n13884 ;
  assign y4127 = ~n13887 ;
  assign y4128 = n13890 ;
  assign y4129 = n13895 ;
  assign y4130 = n13899 ;
  assign y4131 = ~n13901 ;
  assign y4132 = n13906 ;
  assign y4133 = ~n13913 ;
  assign y4134 = n13914 ;
  assign y4135 = ~n13925 ;
  assign y4136 = ~n13936 ;
  assign y4137 = ~n13939 ;
  assign y4138 = n13941 ;
  assign y4139 = n13947 ;
  assign y4140 = ~1'b0 ;
  assign y4141 = ~1'b0 ;
  assign y4142 = n13948 ;
  assign y4143 = ~n13953 ;
  assign y4144 = ~n13954 ;
  assign y4145 = ~1'b0 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = ~n13956 ;
  assign y4148 = n13958 ;
  assign y4149 = ~1'b0 ;
  assign y4150 = ~n13960 ;
  assign y4151 = ~n13961 ;
  assign y4152 = ~n13962 ;
  assign y4153 = n13963 ;
  assign y4154 = n13966 ;
  assign y4155 = ~1'b0 ;
  assign y4156 = ~n13968 ;
  assign y4157 = ~n13972 ;
  assign y4158 = n13977 ;
  assign y4159 = n13978 ;
  assign y4160 = n13983 ;
  assign y4161 = n13984 ;
  assign y4162 = n13989 ;
  assign y4163 = ~n13997 ;
  assign y4164 = ~n13999 ;
  assign y4165 = ~n14004 ;
  assign y4166 = n14006 ;
  assign y4167 = ~n14013 ;
  assign y4168 = n14014 ;
  assign y4169 = ~n14019 ;
  assign y4170 = n14020 ;
  assign y4171 = n14028 ;
  assign y4172 = n14032 ;
  assign y4173 = ~n14036 ;
  assign y4174 = ~n14038 ;
  assign y4175 = ~n14045 ;
  assign y4176 = n14054 ;
  assign y4177 = n14056 ;
  assign y4178 = n14059 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = ~n14060 ;
  assign y4182 = ~n14065 ;
  assign y4183 = n14067 ;
  assign y4184 = ~n14070 ;
  assign y4185 = ~n14075 ;
  assign y4186 = ~1'b0 ;
  assign y4187 = ~n14081 ;
  assign y4188 = n14082 ;
  assign y4189 = ~n14085 ;
  assign y4190 = n14093 ;
  assign y4191 = ~1'b0 ;
  assign y4192 = ~1'b0 ;
  assign y4193 = n14104 ;
  assign y4194 = n14106 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = ~1'b0 ;
  assign y4197 = ~n14108 ;
  assign y4198 = ~n14109 ;
  assign y4199 = n14111 ;
  assign y4200 = ~1'b0 ;
  assign y4201 = n14113 ;
  assign y4202 = n14114 ;
  assign y4203 = ~1'b0 ;
  assign y4204 = n14115 ;
  assign y4205 = ~n14117 ;
  assign y4206 = n14120 ;
  assign y4207 = ~n14121 ;
  assign y4208 = ~n14122 ;
  assign y4209 = n14125 ;
  assign y4210 = n14126 ;
  assign y4211 = ~n14127 ;
  assign y4212 = n11747 ;
  assign y4213 = n14128 ;
  assign y4214 = ~n14129 ;
  assign y4215 = ~n14131 ;
  assign y4216 = ~n14135 ;
  assign y4217 = ~1'b0 ;
  assign y4218 = n14138 ;
  assign y4219 = n14142 ;
  assign y4220 = n14146 ;
  assign y4221 = n14150 ;
  assign y4222 = ~n14157 ;
  assign y4223 = ~n14161 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~n14167 ;
  assign y4226 = n14178 ;
  assign y4227 = ~n14180 ;
  assign y4228 = ~1'b0 ;
  assign y4229 = n5840 ;
  assign y4230 = n14182 ;
  assign y4231 = ~1'b0 ;
  assign y4232 = ~n14184 ;
  assign y4233 = ~n14194 ;
  assign y4234 = ~n14196 ;
  assign y4235 = n14200 ;
  assign y4236 = ~n14201 ;
  assign y4237 = ~1'b0 ;
  assign y4238 = ~1'b0 ;
  assign y4239 = ~n14204 ;
  assign y4240 = n14207 ;
  assign y4241 = ~n14215 ;
  assign y4242 = n14217 ;
  assign y4243 = ~n14218 ;
  assign y4244 = n14223 ;
  assign y4245 = ~n14230 ;
  assign y4246 = ~n14233 ;
  assign y4247 = ~n14241 ;
  assign y4248 = ~n14243 ;
  assign y4249 = n14255 ;
  assign y4250 = ~n14261 ;
  assign y4251 = ~n14268 ;
  assign y4252 = ~n14276 ;
  assign y4253 = n14278 ;
  assign y4254 = ~n14283 ;
  assign y4255 = n14285 ;
  assign y4256 = n14287 ;
  assign y4257 = ~n14297 ;
  assign y4258 = ~n14300 ;
  assign y4259 = ~1'b0 ;
  assign y4260 = ~n14309 ;
  assign y4261 = n14313 ;
  assign y4262 = ~n14323 ;
  assign y4263 = n14324 ;
  assign y4264 = ~n14328 ;
  assign y4265 = ~n14332 ;
  assign y4266 = ~n14333 ;
  assign y4267 = n14334 ;
  assign y4268 = n10000 ;
  assign y4269 = ~n14339 ;
  assign y4270 = n14340 ;
  assign y4271 = n14342 ;
  assign y4272 = n14346 ;
  assign y4273 = n14347 ;
  assign y4274 = n14352 ;
  assign y4275 = ~n14356 ;
  assign y4276 = ~n14362 ;
  assign y4277 = ~n14371 ;
  assign y4278 = n14375 ;
  assign y4279 = n14380 ;
  assign y4280 = ~1'b0 ;
  assign y4281 = n14383 ;
  assign y4282 = n14385 ;
  assign y4283 = ~1'b0 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = ~n14391 ;
  assign y4286 = ~n14399 ;
  assign y4287 = ~n14404 ;
  assign y4288 = ~n14413 ;
  assign y4289 = ~n14415 ;
  assign y4290 = n14417 ;
  assign y4291 = ~1'b0 ;
  assign y4292 = n14419 ;
  assign y4293 = n14422 ;
  assign y4294 = ~n14424 ;
  assign y4295 = ~n14426 ;
  assign y4296 = n14428 ;
  assign y4297 = ~1'b0 ;
  assign y4298 = ~n14438 ;
  assign y4299 = ~n14443 ;
  assign y4300 = n14444 ;
  assign y4301 = ~1'b0 ;
  assign y4302 = ~n14454 ;
  assign y4303 = n14455 ;
  assign y4304 = n14459 ;
  assign y4305 = ~n14460 ;
  assign y4306 = ~x84 ;
  assign y4307 = ~1'b0 ;
  assign y4308 = ~n14461 ;
  assign y4309 = ~n14465 ;
  assign y4310 = n14469 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = ~n2876 ;
  assign y4313 = n14471 ;
  assign y4314 = ~n14472 ;
  assign y4315 = ~n14477 ;
  assign y4316 = n14479 ;
  assign y4317 = n14481 ;
  assign y4318 = ~n14483 ;
  assign y4319 = ~n14486 ;
  assign y4320 = n14501 ;
  assign y4321 = ~n13020 ;
  assign y4322 = ~n14508 ;
  assign y4323 = n14511 ;
  assign y4324 = n14517 ;
  assign y4325 = n14523 ;
  assign y4326 = ~1'b0 ;
  assign y4327 = n14525 ;
  assign y4328 = n14528 ;
  assign y4329 = ~n14529 ;
  assign y4330 = ~1'b0 ;
  assign y4331 = n14530 ;
  assign y4332 = ~n14535 ;
  assign y4333 = ~n14541 ;
  assign y4334 = n14547 ;
  assign y4335 = ~1'b0 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = n14551 ;
  assign y4338 = ~n14552 ;
  assign y4339 = n14555 ;
  assign y4340 = n14558 ;
  assign y4341 = n14561 ;
  assign y4342 = ~n14565 ;
  assign y4343 = n14566 ;
  assign y4344 = ~n14569 ;
  assign y4345 = ~n14571 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = n14582 ;
  assign y4348 = ~n14583 ;
  assign y4349 = ~1'b0 ;
  assign y4350 = ~n14585 ;
  assign y4351 = ~n14588 ;
  assign y4352 = ~n14594 ;
  assign y4353 = n14598 ;
  assign y4354 = ~n14604 ;
  assign y4355 = n14606 ;
  assign y4356 = ~n14609 ;
  assign y4357 = ~n14614 ;
  assign y4358 = n14615 ;
  assign y4359 = ~n14623 ;
  assign y4360 = ~n14630 ;
  assign y4361 = ~n14632 ;
  assign y4362 = ~1'b0 ;
  assign y4363 = n14634 ;
  assign y4364 = n14636 ;
  assign y4365 = ~n14638 ;
  assign y4366 = n14639 ;
  assign y4367 = ~n14642 ;
  assign y4368 = ~1'b0 ;
  assign y4369 = ~n14651 ;
  assign y4370 = ~n14653 ;
  assign y4371 = n14655 ;
  assign y4372 = ~n14656 ;
  assign y4373 = ~n14661 ;
  assign y4374 = ~n14663 ;
  assign y4375 = n14665 ;
  assign y4376 = ~n14666 ;
  assign y4377 = ~1'b0 ;
  assign y4378 = ~n14669 ;
  assign y4379 = ~n14676 ;
  assign y4380 = ~n14677 ;
  assign y4381 = ~n14678 ;
  assign y4382 = n14682 ;
  assign y4383 = n14684 ;
  assign y4384 = n14687 ;
  assign y4385 = ~n14692 ;
  assign y4386 = ~1'b0 ;
  assign y4387 = ~1'b0 ;
  assign y4388 = ~n14696 ;
  assign y4389 = n14702 ;
  assign y4390 = ~1'b0 ;
  assign y4391 = ~1'b0 ;
  assign y4392 = n14706 ;
  assign y4393 = n14712 ;
  assign y4394 = n14718 ;
  assign y4395 = ~n14720 ;
  assign y4396 = ~n14723 ;
  assign y4397 = ~n14728 ;
  assign y4398 = n13188 ;
  assign y4399 = ~n14729 ;
  assign y4400 = ~n14744 ;
  assign y4401 = ~n14755 ;
  assign y4402 = n14765 ;
  assign y4403 = ~1'b0 ;
  assign y4404 = n14769 ;
  assign y4405 = n14779 ;
  assign y4406 = ~n14783 ;
  assign y4407 = n14785 ;
  assign y4408 = n14797 ;
  assign y4409 = n14798 ;
  assign y4410 = ~n14800 ;
  assign y4411 = ~1'b0 ;
  assign y4412 = ~n14805 ;
  assign y4413 = n14813 ;
  assign y4414 = n14822 ;
  assign y4415 = ~n14826 ;
  assign y4416 = n14827 ;
  assign y4417 = n14828 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = ~1'b0 ;
  assign y4420 = ~n14835 ;
  assign y4421 = n14842 ;
  assign y4422 = ~n14846 ;
  assign y4423 = n14847 ;
  assign y4424 = n14851 ;
  assign y4425 = ~n14856 ;
  assign y4426 = n14859 ;
  assign y4427 = ~1'b0 ;
  assign y4428 = n14861 ;
  assign y4429 = ~n14862 ;
  assign y4430 = n14865 ;
  assign y4431 = n14867 ;
  assign y4432 = ~n14869 ;
  assign y4433 = ~n14875 ;
  assign y4434 = n14876 ;
  assign y4435 = ~n1545 ;
  assign y4436 = n14877 ;
  assign y4437 = n14878 ;
  assign y4438 = ~n14880 ;
  assign y4439 = n14885 ;
  assign y4440 = n14887 ;
  assign y4441 = ~n14908 ;
  assign y4442 = ~1'b0 ;
  assign y4443 = ~1'b0 ;
  assign y4444 = n14912 ;
  assign y4445 = ~n14920 ;
  assign y4446 = ~n14922 ;
  assign y4447 = ~n14927 ;
  assign y4448 = ~1'b0 ;
  assign y4449 = ~1'b0 ;
  assign y4450 = n14930 ;
  assign y4451 = n14931 ;
  assign y4452 = ~1'b0 ;
  assign y4453 = ~n14937 ;
  assign y4454 = ~1'b0 ;
  assign y4455 = ~n14940 ;
  assign y4456 = n14942 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = ~n14946 ;
  assign y4459 = n14947 ;
  assign y4460 = n14954 ;
  assign y4461 = n14955 ;
  assign y4462 = ~n14957 ;
  assign y4463 = n14960 ;
  assign y4464 = n14965 ;
  assign y4465 = ~1'b0 ;
  assign y4466 = ~1'b0 ;
  assign y4467 = ~n14966 ;
  assign y4468 = ~n14968 ;
  assign y4469 = n14969 ;
  assign y4470 = ~n14970 ;
  assign y4471 = ~n14973 ;
  assign y4472 = ~n14974 ;
  assign y4473 = ~n14977 ;
  assign y4474 = n14978 ;
  assign y4475 = ~n14982 ;
  assign y4476 = ~n14989 ;
  assign y4477 = ~1'b0 ;
  assign y4478 = n14990 ;
  assign y4479 = ~n14996 ;
  assign y4480 = n14998 ;
  assign y4481 = ~n15004 ;
  assign y4482 = ~n15014 ;
  assign y4483 = n15015 ;
  assign y4484 = n15017 ;
  assign y4485 = ~n15022 ;
  assign y4486 = ~n15023 ;
  assign y4487 = ~n15024 ;
  assign y4488 = ~n15026 ;
  assign y4489 = n15031 ;
  assign y4490 = n15040 ;
  assign y4491 = ~n15049 ;
  assign y4492 = ~1'b0 ;
  assign y4493 = ~1'b0 ;
  assign y4494 = ~1'b0 ;
  assign y4495 = ~n461 ;
  assign y4496 = n15051 ;
  assign y4497 = ~1'b0 ;
  assign y4498 = ~n15058 ;
  assign y4499 = ~n15059 ;
  assign y4500 = n15061 ;
  assign y4501 = ~1'b0 ;
  assign y4502 = n15065 ;
  assign y4503 = ~n15071 ;
  assign y4504 = ~n15072 ;
  assign y4505 = n15075 ;
  assign y4506 = n15080 ;
  assign y4507 = n15085 ;
  assign y4508 = n15086 ;
  assign y4509 = ~n15088 ;
  assign y4510 = ~n15089 ;
  assign y4511 = n15094 ;
  assign y4512 = n15096 ;
  assign y4513 = n15101 ;
  assign y4514 = n15103 ;
  assign y4515 = ~n15106 ;
  assign y4516 = n15107 ;
  assign y4517 = n15109 ;
  assign y4518 = n15111 ;
  assign y4519 = ~n15119 ;
  assign y4520 = n15121 ;
  assign y4521 = n15126 ;
  assign y4522 = ~n15127 ;
  assign y4523 = ~n15128 ;
  assign y4524 = n15129 ;
  assign y4525 = ~n15138 ;
  assign y4526 = ~n15141 ;
  assign y4527 = ~n15146 ;
  assign y4528 = ~n15150 ;
  assign y4529 = ~n15154 ;
  assign y4530 = ~1'b0 ;
  assign y4531 = n15159 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = ~n783 ;
  assign y4534 = n15160 ;
  assign y4535 = ~n15163 ;
  assign y4536 = n15168 ;
  assign y4537 = n15172 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = ~n15178 ;
  assign y4540 = ~n15181 ;
  assign y4541 = ~n15187 ;
  assign y4542 = n15194 ;
  assign y4543 = ~n15197 ;
  assign y4544 = n15198 ;
  assign y4545 = ~1'b0 ;
  assign y4546 = ~n15199 ;
  assign y4547 = n15205 ;
  assign y4548 = n15208 ;
  assign y4549 = ~n15209 ;
  assign y4550 = n15218 ;
  assign y4551 = ~n15225 ;
  assign y4552 = n15233 ;
  assign y4553 = ~n15236 ;
  assign y4554 = n15237 ;
  assign y4555 = n15242 ;
  assign y4556 = ~n15245 ;
  assign y4557 = n15250 ;
  assign y4558 = n15256 ;
  assign y4559 = ~1'b0 ;
  assign y4560 = ~n15264 ;
  assign y4561 = ~n15267 ;
  assign y4562 = ~1'b0 ;
  assign y4563 = ~n15277 ;
  assign y4564 = n15278 ;
  assign y4565 = n15282 ;
  assign y4566 = ~n15284 ;
  assign y4567 = ~n15286 ;
  assign y4568 = ~1'b0 ;
  assign y4569 = ~n15288 ;
  assign y4570 = ~n9805 ;
  assign y4571 = ~n15293 ;
  assign y4572 = ~n15297 ;
  assign y4573 = n15307 ;
  assign y4574 = ~n15310 ;
  assign y4575 = ~n15313 ;
  assign y4576 = ~n15318 ;
  assign y4577 = ~1'b0 ;
  assign y4578 = 1'b0 ;
  assign y4579 = n15326 ;
  assign y4580 = n15328 ;
  assign y4581 = ~n15329 ;
  assign y4582 = ~n15331 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = ~n15332 ;
  assign y4585 = n15333 ;
  assign y4586 = ~n15336 ;
  assign y4587 = ~n15341 ;
  assign y4588 = ~n15342 ;
  assign y4589 = ~n15353 ;
  assign y4590 = ~n15355 ;
  assign y4591 = ~n15356 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = ~n15361 ;
  assign y4594 = ~n15364 ;
  assign y4595 = ~1'b0 ;
  assign y4596 = ~n15368 ;
  assign y4597 = n15370 ;
  assign y4598 = n15373 ;
  assign y4599 = ~1'b0 ;
  assign y4600 = ~1'b0 ;
  assign y4601 = n15379 ;
  assign y4602 = ~n15380 ;
  assign y4603 = ~1'b0 ;
  assign y4604 = n15389 ;
  assign y4605 = ~n15390 ;
  assign y4606 = n15392 ;
  assign y4607 = ~n15395 ;
  assign y4608 = n15398 ;
  assign y4609 = ~n15401 ;
  assign y4610 = ~n15403 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = n15406 ;
  assign y4613 = n15407 ;
  assign y4614 = ~1'b0 ;
  assign y4615 = n15411 ;
  assign y4616 = ~n15415 ;
  assign y4617 = ~1'b0 ;
  assign y4618 = ~n10922 ;
  assign y4619 = n15421 ;
  assign y4620 = ~n15439 ;
  assign y4621 = n15441 ;
  assign y4622 = ~n15444 ;
  assign y4623 = ~1'b0 ;
  assign y4624 = n2127 ;
  assign y4625 = n15451 ;
  assign y4626 = ~n15453 ;
  assign y4627 = ~n15454 ;
  assign y4628 = n15457 ;
  assign y4629 = ~n15459 ;
  assign y4630 = ~n15464 ;
  assign y4631 = ~1'b0 ;
  assign y4632 = n15465 ;
  assign y4633 = ~n15467 ;
  assign y4634 = ~n15468 ;
  assign y4635 = ~n15471 ;
  assign y4636 = ~n15475 ;
  assign y4637 = n15481 ;
  assign y4638 = n15486 ;
  assign y4639 = ~n15487 ;
  assign y4640 = ~1'b0 ;
  assign y4641 = n15489 ;
  assign y4642 = ~n15492 ;
  assign y4643 = n15494 ;
  assign y4644 = ~1'b0 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = n15496 ;
  assign y4647 = ~n15499 ;
  assign y4648 = ~n15500 ;
  assign y4649 = ~n15504 ;
  assign y4650 = ~1'b0 ;
  assign y4651 = n15512 ;
  assign y4652 = n15514 ;
  assign y4653 = n15522 ;
  assign y4654 = ~1'b0 ;
  assign y4655 = n15525 ;
  assign y4656 = n15528 ;
  assign y4657 = n15535 ;
  assign y4658 = n15537 ;
  assign y4659 = ~n15539 ;
  assign y4660 = n15541 ;
  assign y4661 = ~n15545 ;
  assign y4662 = ~n15548 ;
  assign y4663 = ~n15553 ;
  assign y4664 = n15561 ;
  assign y4665 = n15562 ;
  assign y4666 = ~1'b0 ;
  assign y4667 = n15567 ;
  assign y4668 = ~n15576 ;
  assign y4669 = ~1'b0 ;
  assign y4670 = ~n15581 ;
  assign y4671 = n15582 ;
  assign y4672 = ~n15589 ;
  assign y4673 = n15591 ;
  assign y4674 = ~n15597 ;
  assign y4675 = ~1'b0 ;
  assign y4676 = ~n15599 ;
  assign y4677 = ~n15604 ;
  assign y4678 = ~1'b0 ;
  assign y4679 = ~1'b0 ;
  assign y4680 = ~n15605 ;
  assign y4681 = n15610 ;
  assign y4682 = ~n15611 ;
  assign y4683 = n15613 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = n15614 ;
  assign y4686 = ~n15617 ;
  assign y4687 = ~n15618 ;
  assign y4688 = ~1'b0 ;
  assign y4689 = ~1'b0 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = ~1'b0 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = ~n15624 ;
  assign y4695 = ~n15626 ;
  assign y4696 = ~n15628 ;
  assign y4697 = n15634 ;
  assign y4698 = n15639 ;
  assign y4699 = n15647 ;
  assign y4700 = ~n15653 ;
  assign y4701 = ~n15654 ;
  assign y4702 = n15660 ;
  assign y4703 = ~1'b0 ;
  assign y4704 = ~n15663 ;
  assign y4705 = ~n15664 ;
  assign y4706 = ~n15665 ;
  assign y4707 = n15668 ;
  assign y4708 = ~1'b0 ;
  assign y4709 = n15671 ;
  assign y4710 = ~n15672 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = ~n15679 ;
  assign y4714 = ~n15690 ;
  assign y4715 = ~n15691 ;
  assign y4716 = ~1'b0 ;
  assign y4717 = n15694 ;
  assign y4718 = ~n15696 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = ~n15703 ;
  assign y4721 = ~n15711 ;
  assign y4722 = n15715 ;
  assign y4723 = n15718 ;
  assign y4724 = ~n13382 ;
  assign y4725 = n15723 ;
  assign y4726 = ~n15724 ;
  assign y4727 = n15725 ;
  assign y4728 = ~n15736 ;
  assign y4729 = n15738 ;
  assign y4730 = ~n15751 ;
  assign y4731 = n15757 ;
  assign y4732 = n15760 ;
  assign y4733 = ~n15761 ;
  assign y4734 = ~n15763 ;
  assign y4735 = ~1'b0 ;
  assign y4736 = ~n15764 ;
  assign y4737 = n15765 ;
  assign y4738 = ~n15768 ;
  assign y4739 = ~n15769 ;
  assign y4740 = n15775 ;
  assign y4741 = n15777 ;
  assign y4742 = ~1'b0 ;
  assign y4743 = n15779 ;
  assign y4744 = n15786 ;
  assign y4745 = n15788 ;
  assign y4746 = n15792 ;
  assign y4747 = ~n15802 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = n15806 ;
  assign y4750 = n15815 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = n15819 ;
  assign y4754 = ~n15821 ;
  assign y4755 = n15822 ;
  assign y4756 = ~n15828 ;
  assign y4757 = ~n15830 ;
  assign y4758 = ~n15831 ;
  assign y4759 = n15833 ;
  assign y4760 = ~n15834 ;
  assign y4761 = ~n15837 ;
  assign y4762 = n15839 ;
  assign y4763 = ~n15841 ;
  assign y4764 = n15848 ;
  assign y4765 = n15851 ;
  assign y4766 = ~n15853 ;
  assign y4767 = ~1'b0 ;
  assign y4768 = ~n15861 ;
  assign y4769 = n15862 ;
  assign y4770 = n15872 ;
  assign y4771 = ~n15873 ;
  assign y4772 = ~n15876 ;
  assign y4773 = ~n15880 ;
  assign y4774 = ~n15882 ;
  assign y4775 = ~n15885 ;
  assign y4776 = ~n15887 ;
  assign y4777 = ~1'b0 ;
  assign y4778 = n15888 ;
  assign y4779 = ~1'b0 ;
  assign y4780 = n15893 ;
  assign y4781 = ~1'b0 ;
  assign y4782 = ~n15896 ;
  assign y4783 = n15897 ;
  assign y4784 = ~n15898 ;
  assign y4785 = n15900 ;
  assign y4786 = n8399 ;
  assign y4787 = ~n15901 ;
  assign y4788 = n15902 ;
  assign y4789 = ~n15909 ;
  assign y4790 = ~1'b0 ;
  assign y4791 = ~n15910 ;
  assign y4792 = n15920 ;
  assign y4793 = n15921 ;
  assign y4794 = n15929 ;
  assign y4795 = n13895 ;
  assign y4796 = ~n15931 ;
  assign y4797 = ~n15933 ;
  assign y4798 = ~1'b0 ;
  assign y4799 = ~n15937 ;
  assign y4800 = ~n15939 ;
  assign y4801 = ~n15946 ;
  assign y4802 = ~n15950 ;
  assign y4803 = ~1'b0 ;
  assign y4804 = 1'b0 ;
  assign y4805 = ~n15952 ;
  assign y4806 = ~n15954 ;
  assign y4807 = n15959 ;
  assign y4808 = n15960 ;
  assign y4809 = n15962 ;
  assign y4810 = ~n15963 ;
  assign y4811 = ~1'b0 ;
  assign y4812 = ~1'b0 ;
  assign y4813 = ~n15968 ;
  assign y4814 = ~n15969 ;
  assign y4815 = ~n15970 ;
  assign y4816 = ~1'b0 ;
  assign y4817 = ~n15971 ;
  assign y4818 = n15974 ;
  assign y4819 = n15978 ;
  assign y4820 = ~1'b0 ;
  assign y4821 = n15980 ;
  assign y4822 = n15981 ;
  assign y4823 = ~1'b0 ;
  assign y4824 = ~n15983 ;
  assign y4825 = n15986 ;
  assign y4826 = n15988 ;
  assign y4827 = ~1'b0 ;
  assign y4828 = ~n15990 ;
  assign y4829 = ~n15993 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = n15999 ;
  assign y4832 = n16002 ;
  assign y4833 = ~n16003 ;
  assign y4834 = ~1'b0 ;
  assign y4835 = n16005 ;
  assign y4836 = ~n16006 ;
  assign y4837 = ~n16010 ;
  assign y4838 = n16012 ;
  assign y4839 = n16016 ;
  assign y4840 = ~n16018 ;
  assign y4841 = n16020 ;
  assign y4842 = ~n16023 ;
  assign y4843 = ~n16031 ;
  assign y4844 = n15486 ;
  assign y4845 = ~n16039 ;
  assign y4846 = ~n16046 ;
  assign y4847 = n16049 ;
  assign y4848 = ~1'b0 ;
  assign y4849 = ~1'b0 ;
  assign y4850 = n16050 ;
  assign y4851 = ~n16052 ;
  assign y4852 = ~n16056 ;
  assign y4853 = n16057 ;
  assign y4854 = ~1'b0 ;
  assign y4855 = ~1'b0 ;
  assign y4856 = n16060 ;
  assign y4857 = ~n16062 ;
  assign y4858 = ~n16065 ;
  assign y4859 = ~n16066 ;
  assign y4860 = n16068 ;
  assign y4861 = ~n16071 ;
  assign y4862 = ~n16079 ;
  assign y4863 = n16083 ;
  assign y4864 = n16084 ;
  assign y4865 = ~1'b0 ;
  assign y4866 = ~n16086 ;
  assign y4867 = ~n11978 ;
  assign y4868 = ~1'b0 ;
  assign y4869 = n16087 ;
  assign y4870 = n16088 ;
  assign y4871 = ~n16091 ;
  assign y4872 = n16092 ;
  assign y4873 = n16096 ;
  assign y4874 = ~n16099 ;
  assign y4875 = ~1'b0 ;
  assign y4876 = ~n16106 ;
  assign y4877 = ~1'b0 ;
  assign y4878 = ~1'b0 ;
  assign y4879 = ~n16109 ;
  assign y4880 = n16111 ;
  assign y4881 = n16116 ;
  assign y4882 = n16119 ;
  assign y4883 = ~n16121 ;
  assign y4884 = ~n16127 ;
  assign y4885 = ~n16129 ;
  assign y4886 = ~1'b0 ;
  assign y4887 = n16134 ;
  assign y4888 = ~n16139 ;
  assign y4889 = ~n16147 ;
  assign y4890 = n16149 ;
  assign y4891 = n16151 ;
  assign y4892 = ~1'b0 ;
  assign y4893 = n16152 ;
  assign y4894 = ~n16159 ;
  assign y4895 = ~n16160 ;
  assign y4896 = ~n16162 ;
  assign y4897 = ~n16165 ;
  assign y4898 = n16166 ;
  assign y4899 = n16169 ;
  assign y4900 = n16171 ;
  assign y4901 = ~n16173 ;
  assign y4902 = n16175 ;
  assign y4903 = ~n16177 ;
  assign y4904 = n703 ;
  assign y4905 = ~1'b0 ;
  assign y4906 = ~n16186 ;
  assign y4907 = ~n16187 ;
  assign y4908 = ~n16189 ;
  assign y4909 = ~n16192 ;
  assign y4910 = ~1'b0 ;
  assign y4911 = n16193 ;
  assign y4912 = n16194 ;
  assign y4913 = ~n16200 ;
  assign y4914 = ~1'b0 ;
  assign y4915 = n16201 ;
  assign y4916 = ~n16202 ;
  assign y4917 = ~n16203 ;
  assign y4918 = ~n16208 ;
  assign y4919 = ~n12262 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = ~1'b0 ;
  assign y4922 = n16209 ;
  assign y4923 = n3515 ;
  assign y4924 = n16211 ;
  assign y4925 = ~n16214 ;
  assign y4926 = ~n13488 ;
  assign y4927 = n16216 ;
  assign y4928 = n16226 ;
  assign y4929 = ~n16239 ;
  assign y4930 = ~n16241 ;
  assign y4931 = n16242 ;
  assign y4932 = ~n16245 ;
  assign y4933 = ~1'b0 ;
  assign y4934 = n16247 ;
  assign y4935 = n16254 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = ~1'b0 ;
  assign y4938 = ~n16258 ;
  assign y4939 = n16259 ;
  assign y4940 = ~n16260 ;
  assign y4941 = n16262 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = n16267 ;
  assign y4944 = ~n16286 ;
  assign y4945 = n16287 ;
  assign y4946 = ~n16290 ;
  assign y4947 = n16291 ;
  assign y4948 = ~n16292 ;
  assign y4949 = n16293 ;
  assign y4950 = ~n16298 ;
  assign y4951 = n16302 ;
  assign y4952 = ~n16303 ;
  assign y4953 = ~n16308 ;
  assign y4954 = ~n4478 ;
  assign y4955 = n16311 ;
  assign y4956 = ~1'b0 ;
  assign y4957 = n16312 ;
  assign y4958 = n16317 ;
  assign y4959 = n16319 ;
  assign y4960 = n16321 ;
  assign y4961 = ~1'b0 ;
  assign y4962 = ~n16322 ;
  assign y4963 = ~n16323 ;
  assign y4964 = ~n16329 ;
  assign y4965 = n16332 ;
  assign y4966 = n16334 ;
  assign y4967 = ~1'b0 ;
  assign y4968 = ~n16335 ;
  assign y4969 = n16338 ;
  assign y4970 = n16343 ;
  assign y4971 = ~n16346 ;
  assign y4972 = n16349 ;
  assign y4973 = n16353 ;
  assign y4974 = n16357 ;
  assign y4975 = ~1'b0 ;
  assign y4976 = ~n16358 ;
  assign y4977 = ~n16367 ;
  assign y4978 = ~n16368 ;
  assign y4979 = ~n16372 ;
  assign y4980 = ~n16373 ;
  assign y4981 = n16374 ;
  assign y4982 = n16381 ;
  assign y4983 = ~n16385 ;
  assign y4984 = n16387 ;
  assign y4985 = ~n16389 ;
  assign y4986 = ~n16395 ;
  assign y4987 = n16397 ;
  assign y4988 = n16398 ;
  assign y4989 = n16399 ;
  assign y4990 = ~n16400 ;
  assign y4991 = ~n16401 ;
  assign y4992 = ~n16402 ;
  assign y4993 = ~1'b0 ;
  assign y4994 = ~n14758 ;
  assign y4995 = ~n16403 ;
  assign y4996 = ~n16411 ;
  assign y4997 = ~n16415 ;
  assign y4998 = n16419 ;
  assign y4999 = ~1'b0 ;
  assign y5000 = n16421 ;
  assign y5001 = ~n16422 ;
  assign y5002 = ~n16424 ;
  assign y5003 = n16433 ;
  assign y5004 = ~n16437 ;
  assign y5005 = ~n16446 ;
  assign y5006 = n16448 ;
  assign y5007 = n16453 ;
  assign y5008 = ~n16456 ;
  assign y5009 = n16460 ;
  assign y5010 = ~n16462 ;
  assign y5011 = ~n16464 ;
  assign y5012 = n16471 ;
  assign y5013 = ~1'b0 ;
  assign y5014 = ~1'b0 ;
  assign y5015 = ~n16475 ;
  assign y5016 = n16477 ;
  assign y5017 = n16481 ;
  assign y5018 = n16483 ;
  assign y5019 = ~n16486 ;
  assign y5020 = n16491 ;
  assign y5021 = ~1'b0 ;
  assign y5022 = n16492 ;
  assign y5023 = ~n368 ;
  assign y5024 = ~n16493 ;
  assign y5025 = n16496 ;
  assign y5026 = n16497 ;
  assign y5027 = ~n16506 ;
  assign y5028 = ~n16507 ;
  assign y5029 = n16512 ;
  assign y5030 = n16525 ;
  assign y5031 = ~n16535 ;
  assign y5032 = ~n16538 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = ~n16540 ;
  assign y5035 = n16544 ;
  assign y5036 = n16546 ;
  assign y5037 = ~n16551 ;
  assign y5038 = ~n16560 ;
  assign y5039 = n16561 ;
  assign y5040 = ~n16563 ;
  assign y5041 = ~n16566 ;
  assign y5042 = ~n16573 ;
  assign y5043 = n16574 ;
  assign y5044 = ~n16575 ;
  assign y5045 = n16578 ;
  assign y5046 = n16580 ;
  assign y5047 = ~n16581 ;
  assign y5048 = n16582 ;
  assign y5049 = n16586 ;
  assign y5050 = ~n16587 ;
  assign y5051 = ~1'b0 ;
  assign y5052 = ~n16589 ;
  assign y5053 = ~n16593 ;
  assign y5054 = ~n16596 ;
  assign y5055 = n16600 ;
  assign y5056 = n16607 ;
  assign y5057 = n16612 ;
  assign y5058 = ~n16614 ;
  assign y5059 = n16622 ;
  assign y5060 = ~n16624 ;
  assign y5061 = ~n16629 ;
  assign y5062 = ~n16633 ;
  assign y5063 = ~n16635 ;
  assign y5064 = ~n16637 ;
  assign y5065 = ~1'b0 ;
  assign y5066 = ~n16638 ;
  assign y5067 = n16642 ;
  assign y5068 = ~n16644 ;
  assign y5069 = ~n16646 ;
  assign y5070 = ~1'b0 ;
  assign y5071 = 1'b0 ;
  assign y5072 = n16653 ;
  assign y5073 = n16660 ;
  assign y5074 = ~n16668 ;
  assign y5075 = n16671 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = ~n16672 ;
  assign y5078 = n16686 ;
  assign y5079 = ~n16687 ;
  assign y5080 = ~1'b0 ;
  assign y5081 = n5221 ;
  assign y5082 = ~n16688 ;
  assign y5083 = ~n16690 ;
  assign y5084 = n16695 ;
  assign y5085 = n16698 ;
  assign y5086 = n16700 ;
  assign y5087 = n16707 ;
  assign y5088 = ~1'b0 ;
  assign y5089 = ~n16709 ;
  assign y5090 = n16715 ;
  assign y5091 = n16718 ;
  assign y5092 = ~n16719 ;
  assign y5093 = n16721 ;
  assign y5094 = ~n16724 ;
  assign y5095 = n16725 ;
  assign y5096 = n16729 ;
  assign y5097 = n16731 ;
  assign y5098 = 1'b0 ;
  assign y5099 = ~n16732 ;
  assign y5100 = n16736 ;
  assign y5101 = ~n16742 ;
  assign y5102 = ~n16747 ;
  assign y5103 = ~n16750 ;
  assign y5104 = n16755 ;
  assign y5105 = ~n16757 ;
  assign y5106 = n16758 ;
  assign y5107 = ~n16769 ;
  assign y5108 = n16770 ;
  assign y5109 = n16776 ;
  assign y5110 = ~n16779 ;
  assign y5111 = ~n16782 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = n16791 ;
  assign y5114 = ~n16792 ;
  assign y5115 = ~n16794 ;
  assign y5116 = n16798 ;
  assign y5117 = n16801 ;
  assign y5118 = ~n16804 ;
  assign y5119 = n16808 ;
  assign y5120 = ~n16809 ;
  assign y5121 = n16812 ;
  assign y5122 = n16813 ;
  assign y5123 = n16816 ;
  assign y5124 = ~1'b0 ;
  assign y5125 = ~n16824 ;
  assign y5126 = n16829 ;
  assign y5127 = n16832 ;
  assign y5128 = ~n16836 ;
  assign y5129 = ~1'b0 ;
  assign y5130 = n16840 ;
  assign y5131 = ~n16845 ;
  assign y5132 = n16849 ;
  assign y5133 = n16857 ;
  assign y5134 = ~n16860 ;
  assign y5135 = n16861 ;
  assign y5136 = ~1'b0 ;
  assign y5137 = ~n16863 ;
  assign y5138 = n16864 ;
  assign y5139 = ~n16866 ;
  assign y5140 = n16868 ;
  assign y5141 = n16870 ;
  assign y5142 = ~n16871 ;
  assign y5143 = ~n16872 ;
  assign y5144 = ~n16875 ;
  assign y5145 = ~n16877 ;
  assign y5146 = ~n16880 ;
  assign y5147 = n16884 ;
  assign y5148 = ~1'b0 ;
  assign y5149 = n16292 ;
  assign y5150 = n16885 ;
  assign y5151 = ~n16890 ;
  assign y5152 = n16896 ;
  assign y5153 = ~1'b0 ;
  assign y5154 = n16897 ;
  assign y5155 = n16905 ;
  assign y5156 = n16911 ;
  assign y5157 = n16913 ;
  assign y5158 = ~1'b0 ;
  assign y5159 = n16918 ;
  assign y5160 = n16931 ;
  assign y5161 = n16939 ;
  assign y5162 = ~n16944 ;
  assign y5163 = n16946 ;
  assign y5164 = n16948 ;
  assign y5165 = ~1'b0 ;
  assign y5166 = n16950 ;
  assign y5167 = n16953 ;
  assign y5168 = n16956 ;
  assign y5169 = ~1'b0 ;
  assign y5170 = ~n16957 ;
  assign y5171 = n16962 ;
  assign y5172 = ~1'b0 ;
  assign y5173 = ~1'b0 ;
  assign y5174 = ~n16969 ;
  assign y5175 = ~n16977 ;
  assign y5176 = ~n16983 ;
  assign y5177 = ~n16984 ;
  assign y5178 = ~n16986 ;
  assign y5179 = ~1'b0 ;
  assign y5180 = ~n16992 ;
  assign y5181 = ~n16999 ;
  assign y5182 = ~n17007 ;
  assign y5183 = n17008 ;
  assign y5184 = ~1'b0 ;
  assign y5185 = ~n17009 ;
  assign y5186 = ~n17010 ;
  assign y5187 = n17015 ;
  assign y5188 = n17018 ;
  assign y5189 = n15462 ;
  assign y5190 = n17019 ;
  assign y5191 = n17028 ;
  assign y5192 = ~n17030 ;
  assign y5193 = ~1'b0 ;
  assign y5194 = ~n17033 ;
  assign y5195 = ~n17034 ;
  assign y5196 = ~1'b0 ;
  assign y5197 = n17036 ;
  assign y5198 = n17038 ;
  assign y5199 = n17041 ;
  assign y5200 = ~1'b0 ;
  assign y5201 = n17046 ;
  assign y5202 = n17052 ;
  assign y5203 = ~1'b0 ;
  assign y5204 = ~n17056 ;
  assign y5205 = ~1'b0 ;
  assign y5206 = n17067 ;
  assign y5207 = n2325 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = n17075 ;
  assign y5210 = n17081 ;
  assign y5211 = ~1'b0 ;
  assign y5212 = ~1'b0 ;
  assign y5213 = n17082 ;
  assign y5214 = n17087 ;
  assign y5215 = ~n17089 ;
  assign y5216 = n17099 ;
  assign y5217 = ~n17107 ;
  assign y5218 = n17115 ;
  assign y5219 = n17127 ;
  assign y5220 = ~n17128 ;
  assign y5221 = n17130 ;
  assign y5222 = n17139 ;
  assign y5223 = ~1'b0 ;
  assign y5224 = n17142 ;
  assign y5225 = n17144 ;
  assign y5226 = ~n17149 ;
  assign y5227 = n17150 ;
  assign y5228 = ~1'b0 ;
  assign y5229 = ~n17152 ;
  assign y5230 = ~n17156 ;
  assign y5231 = n17157 ;
  assign y5232 = ~n17159 ;
  assign y5233 = 1'b0 ;
  assign y5234 = ~n17172 ;
  assign y5235 = n17174 ;
  assign y5236 = ~n17175 ;
  assign y5237 = n17180 ;
  assign y5238 = ~n17184 ;
  assign y5239 = ~1'b0 ;
  assign y5240 = ~n17189 ;
  assign y5241 = ~1'b0 ;
  assign y5242 = ~n17191 ;
  assign y5243 = ~n17195 ;
  assign y5244 = n17209 ;
  assign y5245 = n17210 ;
  assign y5246 = n17212 ;
  assign y5247 = n17221 ;
  assign y5248 = ~1'b0 ;
  assign y5249 = ~n17230 ;
  assign y5250 = n17234 ;
  assign y5251 = n17238 ;
  assign y5252 = n11178 ;
  assign y5253 = ~n17241 ;
  assign y5254 = n17250 ;
  assign y5255 = ~n17254 ;
  assign y5256 = ~1'b0 ;
  assign y5257 = ~n17258 ;
  assign y5258 = n17260 ;
  assign y5259 = n17261 ;
  assign y5260 = ~n17263 ;
  assign y5261 = ~1'b0 ;
  assign y5262 = ~n17266 ;
  assign y5263 = ~n17267 ;
  assign y5264 = ~n17269 ;
  assign y5265 = n17276 ;
  assign y5266 = ~n17278 ;
  assign y5267 = ~1'b0 ;
  assign y5268 = ~n17279 ;
  assign y5269 = ~n17284 ;
  assign y5270 = n17291 ;
  assign y5271 = ~n17295 ;
  assign y5272 = n17296 ;
  assign y5273 = ~n17298 ;
  assign y5274 = ~n17301 ;
  assign y5275 = n17303 ;
  assign y5276 = ~n17307 ;
  assign y5277 = ~n17318 ;
  assign y5278 = ~n17319 ;
  assign y5279 = ~1'b0 ;
  assign y5280 = ~1'b0 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = ~n17334 ;
  assign y5283 = n17344 ;
  assign y5284 = ~1'b0 ;
  assign y5285 = ~n17349 ;
  assign y5286 = ~n17353 ;
  assign y5287 = ~n17354 ;
  assign y5288 = n17357 ;
  assign y5289 = n17361 ;
  assign y5290 = n17367 ;
  assign y5291 = n17368 ;
  assign y5292 = n17371 ;
  assign y5293 = ~n17372 ;
  assign y5294 = ~n17377 ;
  assign y5295 = n17382 ;
  assign y5296 = ~n17389 ;
  assign y5297 = ~n17400 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = n17401 ;
  assign y5300 = ~n17406 ;
  assign y5301 = ~n17415 ;
  assign y5302 = ~n17417 ;
  assign y5303 = ~1'b0 ;
  assign y5304 = n17422 ;
  assign y5305 = n11669 ;
  assign y5306 = ~n17424 ;
  assign y5307 = ~1'b0 ;
  assign y5308 = ~n17425 ;
  assign y5309 = 1'b0 ;
  assign y5310 = ~n17430 ;
  assign y5311 = ~n17432 ;
  assign y5312 = ~n17436 ;
  assign y5313 = ~n17438 ;
  assign y5314 = ~n17439 ;
  assign y5315 = n17440 ;
  assign y5316 = ~n17444 ;
  assign y5317 = n17447 ;
  assign y5318 = ~n17450 ;
  assign y5319 = ~1'b0 ;
  assign y5320 = ~n17453 ;
  assign y5321 = n17455 ;
  assign y5322 = ~n17456 ;
  assign y5323 = ~n17457 ;
  assign y5324 = n17458 ;
  assign y5325 = ~n17462 ;
  assign y5326 = n17463 ;
  assign y5327 = n17468 ;
  assign y5328 = ~1'b0 ;
  assign y5329 = ~n17474 ;
  assign y5330 = ~n17483 ;
  assign y5331 = n17484 ;
  assign y5332 = ~n17486 ;
  assign y5333 = ~1'b0 ;
  assign y5334 = ~n17488 ;
  assign y5335 = ~n17490 ;
  assign y5336 = n17491 ;
  assign y5337 = ~n17492 ;
  assign y5338 = ~1'b0 ;
  assign y5339 = ~1'b0 ;
  assign y5340 = n17495 ;
  assign y5341 = n17501 ;
  assign y5342 = ~n17508 ;
  assign y5343 = ~1'b0 ;
  assign y5344 = ~n4739 ;
  assign y5345 = ~n17509 ;
  assign y5346 = n17510 ;
  assign y5347 = ~n17513 ;
  assign y5348 = ~1'b0 ;
  assign y5349 = ~n17520 ;
  assign y5350 = ~n17528 ;
  assign y5351 = n17531 ;
  assign y5352 = n17532 ;
  assign y5353 = ~n17533 ;
  assign y5354 = ~1'b0 ;
  assign y5355 = n17536 ;
  assign y5356 = ~n17537 ;
  assign y5357 = ~n17546 ;
  assign y5358 = n17549 ;
  assign y5359 = ~n17550 ;
  assign y5360 = n17551 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = n17555 ;
  assign y5363 = n17557 ;
  assign y5364 = ~n17562 ;
  assign y5365 = ~1'b0 ;
  assign y5366 = n17564 ;
  assign y5367 = n17569 ;
  assign y5368 = ~n17574 ;
  assign y5369 = ~1'b0 ;
  assign y5370 = n17575 ;
  assign y5371 = ~1'b0 ;
  assign y5372 = n16031 ;
  assign y5373 = ~n17578 ;
  assign y5374 = n17579 ;
  assign y5375 = n17580 ;
  assign y5376 = ~n17581 ;
  assign y5377 = ~n17590 ;
  assign y5378 = ~1'b0 ;
  assign y5379 = n17595 ;
  assign y5380 = n17597 ;
  assign y5381 = ~n17599 ;
  assign y5382 = n17600 ;
  assign y5383 = ~n17602 ;
  assign y5384 = n17604 ;
  assign y5385 = ~1'b0 ;
  assign y5386 = n17607 ;
  assign y5387 = ~n17613 ;
  assign y5388 = ~1'b0 ;
  assign y5389 = ~n17627 ;
  assign y5390 = ~n17633 ;
  assign y5391 = ~n17638 ;
  assign y5392 = n17641 ;
  assign y5393 = ~n17645 ;
  assign y5394 = ~n17646 ;
  assign y5395 = n17648 ;
  assign y5396 = ~n17649 ;
  assign y5397 = n17656 ;
  assign y5398 = ~1'b0 ;
  assign y5399 = ~1'b0 ;
  assign y5400 = n17660 ;
  assign y5401 = n17662 ;
  assign y5402 = n17666 ;
  assign y5403 = ~n17668 ;
  assign y5404 = n17677 ;
  assign y5405 = n17681 ;
  assign y5406 = n17683 ;
  assign y5407 = n6683 ;
  assign y5408 = n17689 ;
  assign y5409 = ~n17692 ;
  assign y5410 = n17693 ;
  assign y5411 = ~n17696 ;
  assign y5412 = n17698 ;
  assign y5413 = n17701 ;
  assign y5414 = n17704 ;
  assign y5415 = ~n17706 ;
  assign y5416 = ~n17711 ;
  assign y5417 = ~1'b0 ;
  assign y5418 = n17722 ;
  assign y5419 = n17727 ;
  assign y5420 = n17728 ;
  assign y5421 = ~1'b0 ;
  assign y5422 = ~n17735 ;
  assign y5423 = ~1'b0 ;
  assign y5424 = n17737 ;
  assign y5425 = n17741 ;
  assign y5426 = ~n17742 ;
  assign y5427 = ~n17746 ;
  assign y5428 = ~n17748 ;
  assign y5429 = ~n17755 ;
  assign y5430 = n17757 ;
  assign y5431 = n17759 ;
  assign y5432 = ~n17762 ;
  assign y5433 = ~n17766 ;
  assign y5434 = ~1'b0 ;
  assign y5435 = n17773 ;
  assign y5436 = ~n17778 ;
  assign y5437 = ~n17780 ;
  assign y5438 = n17783 ;
  assign y5439 = n17785 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = ~n17790 ;
  assign y5442 = n17791 ;
  assign y5443 = ~n17794 ;
  assign y5444 = ~n17796 ;
  assign y5445 = n17797 ;
  assign y5446 = ~n17801 ;
  assign y5447 = ~n17802 ;
  assign y5448 = n17809 ;
  assign y5449 = ~n17813 ;
  assign y5450 = ~n17817 ;
  assign y5451 = n17819 ;
  assign y5452 = ~1'b0 ;
  assign y5453 = n17822 ;
  assign y5454 = ~n17825 ;
  assign y5455 = n17826 ;
  assign y5456 = ~1'b0 ;
  assign y5457 = ~n17832 ;
  assign y5458 = n17833 ;
  assign y5459 = ~n17840 ;
  assign y5460 = ~1'b0 ;
  assign y5461 = n17841 ;
  assign y5462 = ~n17847 ;
  assign y5463 = ~n17868 ;
  assign y5464 = ~n17871 ;
  assign y5465 = ~n17873 ;
  assign y5466 = n17874 ;
  assign y5467 = n17876 ;
  assign y5468 = n17878 ;
  assign y5469 = n17884 ;
  assign y5470 = ~n17885 ;
  assign y5471 = ~1'b0 ;
  assign y5472 = ~n17888 ;
  assign y5473 = n17898 ;
  assign y5474 = ~n17899 ;
  assign y5475 = n17902 ;
  assign y5476 = ~n17905 ;
  assign y5477 = ~1'b0 ;
  assign y5478 = ~1'b0 ;
  assign y5479 = ~1'b0 ;
  assign y5480 = n17915 ;
  assign y5481 = ~n17920 ;
  assign y5482 = n17922 ;
  assign y5483 = ~1'b0 ;
  assign y5484 = ~1'b0 ;
  assign y5485 = ~n17925 ;
  assign y5486 = n17938 ;
  assign y5487 = ~n17940 ;
  assign y5488 = ~1'b0 ;
  assign y5489 = ~n17942 ;
  assign y5490 = ~n17944 ;
  assign y5491 = n17947 ;
  assign y5492 = ~n17950 ;
  assign y5493 = ~n17959 ;
  assign y5494 = ~n17964 ;
  assign y5495 = ~1'b0 ;
  assign y5496 = n17967 ;
  assign y5497 = ~1'b0 ;
  assign y5498 = n17968 ;
  assign y5499 = ~1'b0 ;
  assign y5500 = ~n17969 ;
  assign y5501 = n17970 ;
  assign y5502 = ~n17983 ;
  assign y5503 = n17985 ;
  assign y5504 = ~n17989 ;
  assign y5505 = ~n17990 ;
  assign y5506 = ~1'b0 ;
  assign y5507 = n17992 ;
  assign y5508 = n17995 ;
  assign y5509 = ~n18001 ;
  assign y5510 = ~n18003 ;
  assign y5511 = ~n18004 ;
  assign y5512 = ~1'b0 ;
  assign y5513 = ~1'b0 ;
  assign y5514 = ~n18006 ;
  assign y5515 = n18012 ;
  assign y5516 = n18013 ;
  assign y5517 = n18019 ;
  assign y5518 = n18020 ;
  assign y5519 = ~1'b0 ;
  assign y5520 = ~n18024 ;
  assign y5521 = ~1'b0 ;
  assign y5522 = n18027 ;
  assign y5523 = n18031 ;
  assign y5524 = n18034 ;
  assign y5525 = ~1'b0 ;
  assign y5526 = ~n18038 ;
  assign y5527 = ~n18046 ;
  assign y5528 = ~n18050 ;
  assign y5529 = ~n18051 ;
  assign y5530 = ~n18053 ;
  assign y5531 = n18056 ;
  assign y5532 = n18064 ;
  assign y5533 = ~1'b0 ;
  assign y5534 = ~n18067 ;
  assign y5535 = ~1'b0 ;
  assign y5536 = n18069 ;
  assign y5537 = ~n10442 ;
  assign y5538 = n18070 ;
  assign y5539 = ~n18076 ;
  assign y5540 = ~n18077 ;
  assign y5541 = ~1'b0 ;
  assign y5542 = ~1'b0 ;
  assign y5543 = ~n18081 ;
  assign y5544 = ~n18082 ;
  assign y5545 = n18086 ;
  assign y5546 = ~n18087 ;
  assign y5547 = ~1'b0 ;
  assign y5548 = ~n18092 ;
  assign y5549 = ~n1574 ;
  assign y5550 = n18093 ;
  assign y5551 = ~n18094 ;
  assign y5552 = ~1'b0 ;
  assign y5553 = ~1'b0 ;
  assign y5554 = n18096 ;
  assign y5555 = n18100 ;
  assign y5556 = ~n18107 ;
  assign y5557 = ~n18109 ;
  assign y5558 = n18110 ;
  assign y5559 = ~1'b0 ;
  assign y5560 = n18117 ;
  assign y5561 = n18127 ;
  assign y5562 = ~n18129 ;
  assign y5563 = n18133 ;
  assign y5564 = n18137 ;
  assign y5565 = ~n18139 ;
  assign y5566 = ~n18141 ;
  assign y5567 = n18146 ;
  assign y5568 = n18147 ;
  assign y5569 = n18149 ;
  assign y5570 = n18152 ;
  assign y5571 = n18154 ;
  assign y5572 = n18159 ;
  assign y5573 = n18164 ;
  assign y5574 = n18168 ;
  assign y5575 = n18173 ;
  assign y5576 = ~n18175 ;
  assign y5577 = n18177 ;
  assign y5578 = n18180 ;
  assign y5579 = ~n18186 ;
  assign y5580 = ~n18188 ;
  assign y5581 = ~n18196 ;
  assign y5582 = ~1'b0 ;
  assign y5583 = n18197 ;
  assign y5584 = ~n18208 ;
  assign y5585 = ~n18212 ;
  assign y5586 = n18215 ;
  assign y5587 = n18226 ;
  assign y5588 = ~n18228 ;
  assign y5589 = n18235 ;
  assign y5590 = ~n18240 ;
  assign y5591 = ~1'b0 ;
  assign y5592 = 1'b0 ;
  assign y5593 = ~n18252 ;
  assign y5594 = n18257 ;
  assign y5595 = n18258 ;
  assign y5596 = ~n18260 ;
  assign y5597 = ~n18270 ;
  assign y5598 = n18296 ;
  assign y5599 = n18299 ;
  assign y5600 = n18306 ;
  assign y5601 = ~n18312 ;
  assign y5602 = ~1'b0 ;
  assign y5603 = ~n18319 ;
  assign y5604 = n18321 ;
  assign y5605 = n18322 ;
  assign y5606 = ~1'b0 ;
  assign y5607 = ~n18329 ;
  assign y5608 = ~1'b0 ;
  assign y5609 = ~n18332 ;
  assign y5610 = ~1'b0 ;
  assign y5611 = n18336 ;
  assign y5612 = ~1'b0 ;
  assign y5613 = ~n18340 ;
  assign y5614 = 1'b0 ;
  assign y5615 = n18350 ;
  assign y5616 = n18357 ;
  assign y5617 = n18359 ;
  assign y5618 = ~1'b0 ;
  assign y5619 = ~n18360 ;
  assign y5620 = n18364 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = ~n18365 ;
  assign y5623 = n18369 ;
  assign y5624 = ~n18377 ;
  assign y5625 = n18379 ;
  assign y5626 = n18381 ;
  assign y5627 = n18388 ;
  assign y5628 = ~1'b0 ;
  assign y5629 = ~n18389 ;
  assign y5630 = ~n18394 ;
  assign y5631 = ~n18397 ;
  assign y5632 = ~n18398 ;
  assign y5633 = n18406 ;
  assign y5634 = ~n18412 ;
  assign y5635 = ~n18419 ;
  assign y5636 = ~n18425 ;
  assign y5637 = n3059 ;
  assign y5638 = ~1'b0 ;
  assign y5639 = n18427 ;
  assign y5640 = n18429 ;
  assign y5641 = ~n18438 ;
  assign y5642 = n18442 ;
  assign y5643 = n18445 ;
  assign y5644 = ~n18453 ;
  assign y5645 = ~n18454 ;
  assign y5646 = ~n18461 ;
  assign y5647 = ~n18464 ;
  assign y5648 = n18469 ;
  assign y5649 = ~1'b0 ;
  assign y5650 = ~n18472 ;
  assign y5651 = n18473 ;
  assign y5652 = ~n18476 ;
  assign y5653 = ~n18477 ;
  assign y5654 = ~1'b0 ;
  assign y5655 = ~n18478 ;
  assign y5656 = ~1'b0 ;
  assign y5657 = ~1'b0 ;
  assign y5658 = ~1'b0 ;
  assign y5659 = n18485 ;
  assign y5660 = n18486 ;
  assign y5661 = ~1'b0 ;
  assign y5662 = n18487 ;
  assign y5663 = n18491 ;
  assign y5664 = n18496 ;
  assign y5665 = n18499 ;
  assign y5666 = n18502 ;
  assign y5667 = n18504 ;
  assign y5668 = ~n18508 ;
  assign y5669 = ~n18509 ;
  assign y5670 = ~n18513 ;
  assign y5671 = ~n18514 ;
  assign y5672 = ~1'b0 ;
  assign y5673 = ~n18515 ;
  assign y5674 = ~1'b0 ;
  assign y5675 = n18517 ;
  assign y5676 = ~n18520 ;
  assign y5677 = n18522 ;
  assign y5678 = n18523 ;
  assign y5679 = ~n18525 ;
  assign y5680 = ~n18529 ;
  assign y5681 = n18537 ;
  assign y5682 = n18540 ;
  assign y5683 = n11349 ;
  assign y5684 = n18545 ;
  assign y5685 = n18547 ;
  assign y5686 = n18551 ;
  assign y5687 = ~n18557 ;
  assign y5688 = ~n18561 ;
  assign y5689 = n18566 ;
  assign y5690 = ~1'b0 ;
  assign y5691 = n18567 ;
  assign y5692 = n18569 ;
  assign y5693 = ~n18570 ;
  assign y5694 = ~1'b0 ;
  assign y5695 = ~1'b0 ;
  assign y5696 = ~n18571 ;
  assign y5697 = ~1'b0 ;
  assign y5698 = ~n18577 ;
  assign y5699 = ~1'b0 ;
  assign y5700 = n10829 ;
  assign y5701 = ~n18578 ;
  assign y5702 = ~n18579 ;
  assign y5703 = ~1'b0 ;
  assign y5704 = n18583 ;
  assign y5705 = ~n18586 ;
  assign y5706 = ~n18587 ;
  assign y5707 = ~1'b0 ;
  assign y5708 = n18590 ;
  assign y5709 = ~n18592 ;
  assign y5710 = n18593 ;
  assign y5711 = ~1'b0 ;
  assign y5712 = n9988 ;
  assign y5713 = ~n18604 ;
  assign y5714 = n18605 ;
  assign y5715 = ~n18608 ;
  assign y5716 = ~n18609 ;
  assign y5717 = ~n18618 ;
  assign y5718 = ~n18627 ;
  assign y5719 = ~n18634 ;
  assign y5720 = ~1'b0 ;
  assign y5721 = n18644 ;
  assign y5722 = n18645 ;
  assign y5723 = ~n18646 ;
  assign y5724 = n18650 ;
  assign y5725 = ~n18654 ;
  assign y5726 = ~n18655 ;
  assign y5727 = ~1'b0 ;
  assign y5728 = ~n18660 ;
  assign y5729 = ~1'b0 ;
  assign y5730 = n18662 ;
  assign y5731 = ~n18667 ;
  assign y5732 = ~n18671 ;
  assign y5733 = ~n18681 ;
  assign y5734 = n18689 ;
  assign y5735 = n18694 ;
  assign y5736 = n18697 ;
  assign y5737 = ~n18698 ;
  assign y5738 = n18702 ;
  assign y5739 = n18709 ;
  assign y5740 = ~n18712 ;
  assign y5741 = ~n18714 ;
  assign y5742 = ~n18715 ;
  assign y5743 = ~1'b0 ;
  assign y5744 = ~n18718 ;
  assign y5745 = n18719 ;
  assign y5746 = ~n18723 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = ~1'b0 ;
  assign y5749 = ~1'b0 ;
  assign y5750 = n18728 ;
  assign y5751 = n18730 ;
  assign y5752 = ~1'b0 ;
  assign y5753 = n18731 ;
  assign y5754 = ~n18735 ;
  assign y5755 = ~n18737 ;
  assign y5756 = n18741 ;
  assign y5757 = ~n18742 ;
  assign y5758 = ~n18743 ;
  assign y5759 = ~n18745 ;
  assign y5760 = n18747 ;
  assign y5761 = n18749 ;
  assign y5762 = ~n18754 ;
  assign y5763 = n18758 ;
  assign y5764 = n18760 ;
  assign y5765 = ~1'b0 ;
  assign y5766 = ~n18763 ;
  assign y5767 = n18768 ;
  assign y5768 = ~n18772 ;
  assign y5769 = n18783 ;
  assign y5770 = n18787 ;
  assign y5771 = ~1'b0 ;
  assign y5772 = ~n18791 ;
  assign y5773 = n18798 ;
  assign y5774 = ~n18803 ;
  assign y5775 = n18808 ;
  assign y5776 = ~1'b0 ;
  assign y5777 = ~n18811 ;
  assign y5778 = n18812 ;
  assign y5779 = ~1'b0 ;
  assign y5780 = ~n18816 ;
  assign y5781 = ~n18817 ;
  assign y5782 = n18824 ;
  assign y5783 = ~n18826 ;
  assign y5784 = n18827 ;
  assign y5785 = ~1'b0 ;
  assign y5786 = ~n18831 ;
  assign y5787 = ~n10637 ;
  assign y5788 = n18832 ;
  assign y5789 = n18834 ;
  assign y5790 = n18835 ;
  assign y5791 = n18840 ;
  assign y5792 = n18846 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = ~n18858 ;
  assign y5795 = ~1'b0 ;
  assign y5796 = ~n18859 ;
  assign y5797 = ~n18865 ;
  assign y5798 = ~n18868 ;
  assign y5799 = ~1'b0 ;
  assign y5800 = ~n18869 ;
  assign y5801 = ~n18873 ;
  assign y5802 = ~1'b0 ;
  assign y5803 = n9545 ;
  assign y5804 = ~n18876 ;
  assign y5805 = ~n18879 ;
  assign y5806 = ~n18881 ;
  assign y5807 = ~n18882 ;
  assign y5808 = ~n18884 ;
  assign y5809 = n18888 ;
  assign y5810 = n18893 ;
  assign y5811 = n18896 ;
  assign y5812 = ~n18897 ;
  assign y5813 = n18904 ;
  assign y5814 = ~n18907 ;
  assign y5815 = n18913 ;
  assign y5816 = n18915 ;
  assign y5817 = ~n18916 ;
  assign y5818 = ~n18917 ;
  assign y5819 = n18919 ;
  assign y5820 = ~n18933 ;
  assign y5821 = ~n18937 ;
  assign y5822 = ~1'b0 ;
  assign y5823 = n18939 ;
  assign y5824 = ~n18940 ;
  assign y5825 = ~n18945 ;
  assign y5826 = ~n18946 ;
  assign y5827 = n18949 ;
  assign y5828 = n18950 ;
  assign y5829 = ~n18953 ;
  assign y5830 = ~n18956 ;
  assign y5831 = n18957 ;
  assign y5832 = ~1'b0 ;
  assign y5833 = ~1'b0 ;
  assign y5834 = ~n18961 ;
  assign y5835 = n18962 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = n18970 ;
  assign y5838 = n18971 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = ~n18972 ;
  assign y5841 = ~n18977 ;
  assign y5842 = ~n18993 ;
  assign y5843 = ~n19002 ;
  assign y5844 = ~n19008 ;
  assign y5845 = ~1'b0 ;
  assign y5846 = n19013 ;
  assign y5847 = ~1'b0 ;
  assign y5848 = n19014 ;
  assign y5849 = n19015 ;
  assign y5850 = n19017 ;
  assign y5851 = ~n19022 ;
  assign y5852 = ~n19026 ;
  assign y5853 = ~n19031 ;
  assign y5854 = n19032 ;
  assign y5855 = ~1'b0 ;
  assign y5856 = ~1'b0 ;
  assign y5857 = n19033 ;
  assign y5858 = n19034 ;
  assign y5859 = ~n19035 ;
  assign y5860 = ~n19037 ;
  assign y5861 = ~n19039 ;
  assign y5862 = n19040 ;
  assign y5863 = n19041 ;
  assign y5864 = ~n19043 ;
  assign y5865 = n19044 ;
  assign y5866 = ~1'b0 ;
  assign y5867 = ~1'b0 ;
  assign y5868 = x195 ;
  assign y5869 = n19045 ;
  assign y5870 = ~n19047 ;
  assign y5871 = ~n19049 ;
  assign y5872 = n19051 ;
  assign y5873 = ~n19054 ;
  assign y5874 = n19055 ;
  assign y5875 = n19056 ;
  assign y5876 = n19058 ;
  assign y5877 = ~1'b0 ;
  assign y5878 = ~n19063 ;
  assign y5879 = ~n19068 ;
  assign y5880 = ~1'b0 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = n19070 ;
  assign y5883 = ~n19076 ;
  assign y5884 = ~1'b0 ;
  assign y5885 = ~n19081 ;
  assign y5886 = ~n19087 ;
  assign y5887 = ~n19088 ;
  assign y5888 = ~n19089 ;
  assign y5889 = ~1'b0 ;
  assign y5890 = n19094 ;
  assign y5891 = ~n19103 ;
  assign y5892 = ~1'b0 ;
  assign y5893 = n19109 ;
  assign y5894 = n19110 ;
  assign y5895 = n19114 ;
  assign y5896 = ~1'b0 ;
  assign y5897 = n19118 ;
  assign y5898 = ~1'b0 ;
  assign y5899 = ~n19123 ;
  assign y5900 = n19125 ;
  assign y5901 = ~n19126 ;
  assign y5902 = ~n19131 ;
  assign y5903 = n19137 ;
  assign y5904 = n19138 ;
  assign y5905 = ~n19140 ;
  assign y5906 = ~1'b0 ;
  assign y5907 = ~1'b0 ;
  assign y5908 = ~n19142 ;
  assign y5909 = ~n19144 ;
  assign y5910 = ~n19147 ;
  assign y5911 = ~n19150 ;
  assign y5912 = ~n19159 ;
  assign y5913 = ~1'b0 ;
  assign y5914 = n19161 ;
  assign y5915 = n19169 ;
  assign y5916 = ~n19170 ;
  assign y5917 = n19173 ;
  assign y5918 = ~n19174 ;
  assign y5919 = ~n19180 ;
  assign y5920 = n19187 ;
  assign y5921 = ~n19199 ;
  assign y5922 = ~n19203 ;
  assign y5923 = n19204 ;
  assign y5924 = n19212 ;
  assign y5925 = ~1'b0 ;
  assign y5926 = ~n19220 ;
  assign y5927 = n19224 ;
  assign y5928 = n19226 ;
  assign y5929 = n19227 ;
  assign y5930 = n19230 ;
  assign y5931 = n19235 ;
  assign y5932 = ~1'b0 ;
  assign y5933 = ~n19242 ;
  assign y5934 = n19243 ;
  assign y5935 = ~n19245 ;
  assign y5936 = ~n19248 ;
  assign y5937 = n19251 ;
  assign y5938 = n19252 ;
  assign y5939 = n19264 ;
  assign y5940 = n19268 ;
  assign y5941 = ~n19269 ;
  assign y5942 = ~n19272 ;
  assign y5943 = 1'b0 ;
  assign y5944 = ~n19279 ;
  assign y5945 = n19285 ;
  assign y5946 = n19287 ;
  assign y5947 = n19291 ;
  assign y5948 = n19296 ;
  assign y5949 = n19309 ;
  assign y5950 = ~n19312 ;
  assign y5951 = ~n19317 ;
  assign y5952 = n19318 ;
  assign y5953 = ~1'b0 ;
  assign y5954 = ~n19321 ;
  assign y5955 = ~n19322 ;
  assign y5956 = n19327 ;
  assign y5957 = n19351 ;
  assign y5958 = n19354 ;
  assign y5959 = n19358 ;
  assign y5960 = ~n19360 ;
  assign y5961 = ~n19364 ;
  assign y5962 = ~n19365 ;
  assign y5963 = n19370 ;
  assign y5964 = n19381 ;
  assign y5965 = ~n19385 ;
  assign y5966 = n19386 ;
  assign y5967 = n19388 ;
  assign y5968 = ~n19390 ;
  assign y5969 = n9285 ;
  assign y5970 = ~1'b0 ;
  assign y5971 = n19394 ;
  assign y5972 = n19395 ;
  assign y5973 = ~n19398 ;
  assign y5974 = n19400 ;
  assign y5975 = ~n19403 ;
  assign y5976 = ~n19406 ;
  assign y5977 = ~1'b0 ;
  assign y5978 = ~n19408 ;
  assign y5979 = n19412 ;
  assign y5980 = n19416 ;
  assign y5981 = ~1'b0 ;
  assign y5982 = ~n19423 ;
  assign y5983 = n19426 ;
  assign y5984 = ~n19427 ;
  assign y5985 = n19428 ;
  assign y5986 = n19433 ;
  assign y5987 = n19436 ;
  assign y5988 = ~n19444 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = ~n19446 ;
  assign y5991 = n19452 ;
  assign y5992 = ~n19455 ;
  assign y5993 = n19460 ;
  assign y5994 = ~n19468 ;
  assign y5995 = ~1'b0 ;
  assign y5996 = n19472 ;
  assign y5997 = ~n19475 ;
  assign y5998 = ~n19477 ;
  assign y5999 = ~1'b0 ;
  assign y6000 = n19482 ;
  assign y6001 = n19486 ;
  assign y6002 = n19488 ;
  assign y6003 = ~n19489 ;
  assign y6004 = n19491 ;
  assign y6005 = ~n19498 ;
  assign y6006 = n19500 ;
  assign y6007 = ~n19505 ;
  assign y6008 = ~n19510 ;
  assign y6009 = n19515 ;
  assign y6010 = ~n19518 ;
  assign y6011 = ~n19520 ;
  assign y6012 = ~n19522 ;
  assign y6013 = ~n19528 ;
  assign y6014 = ~1'b0 ;
  assign y6015 = n19533 ;
  assign y6016 = ~n19534 ;
  assign y6017 = n19535 ;
  assign y6018 = n19538 ;
  assign y6019 = n19543 ;
  assign y6020 = n19545 ;
  assign y6021 = n19551 ;
  assign y6022 = ~n19554 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = ~1'b0 ;
  assign y6025 = ~n19557 ;
  assign y6026 = ~n19558 ;
  assign y6027 = ~1'b0 ;
  assign y6028 = n19561 ;
  assign y6029 = n19562 ;
  assign y6030 = n19564 ;
  assign y6031 = n19567 ;
  assign y6032 = ~1'b0 ;
  assign y6033 = ~n19574 ;
  assign y6034 = n19577 ;
  assign y6035 = ~1'b0 ;
  assign y6036 = n19578 ;
  assign y6037 = 1'b0 ;
  assign y6038 = ~n9488 ;
  assign y6039 = ~n19581 ;
  assign y6040 = ~n19582 ;
  assign y6041 = n19584 ;
  assign y6042 = ~1'b0 ;
  assign y6043 = ~n19586 ;
  assign y6044 = ~n18934 ;
  assign y6045 = n19589 ;
  assign y6046 = ~n19590 ;
  assign y6047 = ~1'b0 ;
  assign y6048 = ~n19593 ;
  assign y6049 = n19594 ;
  assign y6050 = n19596 ;
  assign y6051 = ~n19599 ;
  assign y6052 = n19608 ;
  assign y6053 = n19620 ;
  assign y6054 = ~n19624 ;
  assign y6055 = ~n19626 ;
  assign y6056 = n19627 ;
  assign y6057 = ~n19636 ;
  assign y6058 = n19646 ;
  assign y6059 = n19662 ;
  assign y6060 = n19663 ;
  assign y6061 = ~1'b0 ;
  assign y6062 = ~n19667 ;
  assign y6063 = n19668 ;
  assign y6064 = ~1'b0 ;
  assign y6065 = ~n19670 ;
  assign y6066 = ~n19676 ;
  assign y6067 = n19681 ;
  assign y6068 = ~n19682 ;
  assign y6069 = ~n19684 ;
  assign y6070 = n19687 ;
  assign y6071 = n19694 ;
  assign y6072 = n19696 ;
  assign y6073 = n19698 ;
  assign y6074 = ~1'b0 ;
  assign y6075 = n19700 ;
  assign y6076 = n19707 ;
  assign y6077 = n19710 ;
  assign y6078 = n19714 ;
  assign y6079 = ~1'b0 ;
  assign y6080 = n19723 ;
  assign y6081 = ~n19728 ;
  assign y6082 = ~1'b0 ;
  assign y6083 = n19734 ;
  assign y6084 = n19741 ;
  assign y6085 = ~n19744 ;
  assign y6086 = ~n19745 ;
  assign y6087 = n19747 ;
  assign y6088 = n19748 ;
  assign y6089 = n19751 ;
  assign y6090 = n19753 ;
  assign y6091 = ~n19754 ;
  assign y6092 = ~n19757 ;
  assign y6093 = ~n19764 ;
  assign y6094 = n19768 ;
  assign y6095 = n19769 ;
  assign y6096 = ~n19772 ;
  assign y6097 = ~n19776 ;
  assign y6098 = ~1'b0 ;
  assign y6099 = n19777 ;
  assign y6100 = ~n19781 ;
  assign y6101 = n19787 ;
  assign y6102 = n19788 ;
  assign y6103 = n19791 ;
  assign y6104 = ~n19792 ;
  assign y6105 = n19796 ;
  assign y6106 = n19798 ;
  assign y6107 = n19802 ;
  assign y6108 = n19803 ;
  assign y6109 = n19808 ;
  assign y6110 = ~n19820 ;
  assign y6111 = n19767 ;
  assign y6112 = ~n19823 ;
  assign y6113 = ~1'b0 ;
  assign y6114 = ~1'b0 ;
  assign y6115 = n19825 ;
  assign y6116 = n19828 ;
  assign y6117 = ~n19830 ;
  assign y6118 = ~n19832 ;
  assign y6119 = ~n19838 ;
  assign y6120 = n19841 ;
  assign y6121 = ~n19843 ;
  assign y6122 = n19852 ;
  assign y6123 = ~n19855 ;
  assign y6124 = ~n19856 ;
  assign y6125 = n19861 ;
  assign y6126 = ~n19864 ;
  assign y6127 = n19873 ;
  assign y6128 = ~n19876 ;
  assign y6129 = ~n19886 ;
  assign y6130 = n19889 ;
  assign y6131 = n19894 ;
  assign y6132 = n19897 ;
  assign y6133 = ~1'b0 ;
  assign y6134 = n19898 ;
  assign y6135 = ~n19901 ;
  assign y6136 = ~1'b0 ;
  assign y6137 = ~1'b0 ;
  assign y6138 = ~n19903 ;
  assign y6139 = n19904 ;
  assign y6140 = ~n19907 ;
  assign y6141 = n19912 ;
  assign y6142 = n16730 ;
  assign y6143 = ~n19914 ;
  assign y6144 = n19915 ;
  assign y6145 = ~n19916 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~n19920 ;
  assign y6148 = ~n19922 ;
  assign y6149 = ~n19923 ;
  assign y6150 = ~n19927 ;
  assign y6151 = ~n19935 ;
  assign y6152 = ~n19938 ;
  assign y6153 = ~n19944 ;
  assign y6154 = n19947 ;
  assign y6155 = ~n19948 ;
  assign y6156 = n19954 ;
  assign y6157 = ~n19958 ;
  assign y6158 = ~n19960 ;
  assign y6159 = n19962 ;
  assign y6160 = ~n19964 ;
  assign y6161 = n19970 ;
  assign y6162 = ~n19975 ;
  assign y6163 = ~n19977 ;
  assign y6164 = ~1'b0 ;
  assign y6165 = ~1'b0 ;
  assign y6166 = ~n19982 ;
  assign y6167 = ~n19987 ;
  assign y6168 = ~1'b0 ;
  assign y6169 = ~n19992 ;
  assign y6170 = ~n19995 ;
  assign y6171 = ~n19996 ;
  assign y6172 = ~1'b0 ;
  assign y6173 = n19998 ;
  assign y6174 = n20003 ;
  assign y6175 = ~n20009 ;
  assign y6176 = n20010 ;
  assign y6177 = ~n20014 ;
  assign y6178 = ~1'b0 ;
  assign y6179 = ~n20016 ;
  assign y6180 = n20020 ;
  assign y6181 = n20024 ;
  assign y6182 = n20025 ;
  assign y6183 = ~1'b0 ;
  assign y6184 = n20029 ;
  assign y6185 = ~n20031 ;
  assign y6186 = n20034 ;
  assign y6187 = n20036 ;
  assign y6188 = ~n20039 ;
  assign y6189 = ~1'b0 ;
  assign y6190 = ~n20043 ;
  assign y6191 = ~n20045 ;
  assign y6192 = ~n20049 ;
  assign y6193 = ~n20051 ;
  assign y6194 = n20052 ;
  assign y6195 = ~n20058 ;
  assign y6196 = n20061 ;
  assign y6197 = n20065 ;
  assign y6198 = ~n20070 ;
  assign y6199 = ~n20072 ;
  assign y6200 = ~n20073 ;
  assign y6201 = n20079 ;
  assign y6202 = n20082 ;
  assign y6203 = n20083 ;
  assign y6204 = ~n20090 ;
  assign y6205 = n20091 ;
  assign y6206 = n20096 ;
  assign y6207 = ~1'b0 ;
  assign y6208 = ~n20101 ;
  assign y6209 = n20103 ;
  assign y6210 = ~n20108 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = ~n20111 ;
  assign y6213 = n20114 ;
  assign y6214 = n20117 ;
  assign y6215 = ~n20122 ;
  assign y6216 = ~1'b0 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = ~n20124 ;
  assign y6219 = ~n20126 ;
  assign y6220 = ~1'b0 ;
  assign y6221 = ~1'b0 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = ~n20129 ;
  assign y6224 = n20135 ;
  assign y6225 = ~n20136 ;
  assign y6226 = ~n20142 ;
  assign y6227 = ~1'b0 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = ~n20150 ;
  assign y6230 = n20151 ;
  assign y6231 = n20153 ;
  assign y6232 = n20156 ;
  assign y6233 = n20161 ;
  assign y6234 = n20162 ;
  assign y6235 = ~n20163 ;
  assign y6236 = ~n20168 ;
  assign y6237 = ~n20169 ;
  assign y6238 = ~n9137 ;
  assign y6239 = ~n20170 ;
  assign y6240 = n20177 ;
  assign y6241 = n20180 ;
  assign y6242 = n20184 ;
  assign y6243 = ~n20185 ;
  assign y6244 = n20189 ;
  assign y6245 = ~n20193 ;
  assign y6246 = n20197 ;
  assign y6247 = ~n20198 ;
  assign y6248 = ~1'b0 ;
  assign y6249 = ~n20200 ;
  assign y6250 = ~n20202 ;
  assign y6251 = n20205 ;
  assign y6252 = ~n20212 ;
  assign y6253 = ~n20213 ;
  assign y6254 = ~n20214 ;
  assign y6255 = ~n20216 ;
  assign y6256 = ~n20219 ;
  assign y6257 = ~n20231 ;
  assign y6258 = n20233 ;
  assign y6259 = ~n20239 ;
  assign y6260 = ~n20242 ;
  assign y6261 = ~n20244 ;
  assign y6262 = n20245 ;
  assign y6263 = ~1'b0 ;
  assign y6264 = ~n20248 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = ~1'b0 ;
  assign y6267 = ~1'b0 ;
  assign y6268 = n20249 ;
  assign y6269 = ~n20264 ;
  assign y6270 = n20265 ;
  assign y6271 = n20274 ;
  assign y6272 = n20279 ;
  assign y6273 = n20288 ;
  assign y6274 = ~n20289 ;
  assign y6275 = n20291 ;
  assign y6276 = ~n20293 ;
  assign y6277 = ~n20295 ;
  assign y6278 = ~n20301 ;
  assign y6279 = ~1'b0 ;
  assign y6280 = ~1'b0 ;
  assign y6281 = ~n20308 ;
  assign y6282 = ~n20313 ;
  assign y6283 = n20316 ;
  assign y6284 = ~n20317 ;
  assign y6285 = n20321 ;
  assign y6286 = ~n20325 ;
  assign y6287 = ~n20342 ;
  assign y6288 = ~n20344 ;
  assign y6289 = ~n20345 ;
  assign y6290 = n20347 ;
  assign y6291 = ~n20357 ;
  assign y6292 = ~1'b0 ;
  assign y6293 = ~n20362 ;
  assign y6294 = n20364 ;
  assign y6295 = n20366 ;
  assign y6296 = n20367 ;
  assign y6297 = n20368 ;
  assign y6298 = n20370 ;
  assign y6299 = ~1'b0 ;
  assign y6300 = n20375 ;
  assign y6301 = ~n20382 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = ~n20387 ;
  assign y6304 = ~n20393 ;
  assign y6305 = n20398 ;
  assign y6306 = n20402 ;
  assign y6307 = ~n20406 ;
  assign y6308 = n20408 ;
  assign y6309 = ~n20411 ;
  assign y6310 = ~n20416 ;
  assign y6311 = n20428 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = ~1'b0 ;
  assign y6314 = n20432 ;
  assign y6315 = n20435 ;
  assign y6316 = ~n20440 ;
  assign y6317 = ~n20450 ;
  assign y6318 = ~1'b0 ;
  assign y6319 = ~n20458 ;
  assign y6320 = ~n20459 ;
  assign y6321 = n20469 ;
  assign y6322 = ~n20475 ;
  assign y6323 = n20477 ;
  assign y6324 = ~n20481 ;
  assign y6325 = ~n20482 ;
  assign y6326 = n20483 ;
  assign y6327 = ~n20489 ;
  assign y6328 = ~n20495 ;
  assign y6329 = ~n20497 ;
  assign y6330 = ~n20498 ;
  assign y6331 = ~n18324 ;
  assign y6332 = ~n20502 ;
  assign y6333 = n20503 ;
  assign y6334 = ~1'b0 ;
  assign y6335 = ~n20507 ;
  assign y6336 = n20509 ;
  assign y6337 = n20511 ;
  assign y6338 = ~n20512 ;
  assign y6339 = n20518 ;
  assign y6340 = n20520 ;
  assign y6341 = n20522 ;
  assign y6342 = ~n20526 ;
  assign y6343 = n20528 ;
  assign y6344 = ~n20530 ;
  assign y6345 = ~n20539 ;
  assign y6346 = ~n20540 ;
  assign y6347 = ~1'b0 ;
  assign y6348 = ~n20544 ;
  assign y6349 = n20554 ;
  assign y6350 = n20557 ;
  assign y6351 = ~n20559 ;
  assign y6352 = ~n20560 ;
  assign y6353 = n12000 ;
  assign y6354 = n20562 ;
  assign y6355 = ~1'b0 ;
  assign y6356 = n20563 ;
  assign y6357 = n20565 ;
  assign y6358 = n20570 ;
  assign y6359 = ~n20572 ;
  assign y6360 = ~n20576 ;
  assign y6361 = ~n20577 ;
  assign y6362 = n20584 ;
  assign y6363 = ~n20586 ;
  assign y6364 = n20587 ;
  assign y6365 = ~1'b0 ;
  assign y6366 = ~n20589 ;
  assign y6367 = n20593 ;
  assign y6368 = ~n20595 ;
  assign y6369 = ~n20596 ;
  assign y6370 = ~1'b0 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = ~n20600 ;
  assign y6373 = n20602 ;
  assign y6374 = n20610 ;
  assign y6375 = ~n20611 ;
  assign y6376 = n20623 ;
  assign y6377 = n20624 ;
  assign y6378 = n20631 ;
  assign y6379 = n20634 ;
  assign y6380 = n20636 ;
  assign y6381 = n20639 ;
  assign y6382 = ~n20641 ;
  assign y6383 = n20642 ;
  assign y6384 = ~n20645 ;
  assign y6385 = ~n20646 ;
  assign y6386 = ~n20647 ;
  assign y6387 = ~n20648 ;
  assign y6388 = ~n20649 ;
  assign y6389 = ~n20653 ;
  assign y6390 = ~n20661 ;
  assign y6391 = n17810 ;
  assign y6392 = ~n20665 ;
  assign y6393 = n5223 ;
  assign y6394 = n20668 ;
  assign y6395 = n20672 ;
  assign y6396 = ~1'b0 ;
  assign y6397 = n20675 ;
  assign y6398 = ~n20680 ;
  assign y6399 = n20682 ;
  assign y6400 = ~n20684 ;
  assign y6401 = ~n20687 ;
  assign y6402 = ~n20690 ;
  assign y6403 = ~n20693 ;
  assign y6404 = n20694 ;
  assign y6405 = ~n20696 ;
  assign y6406 = ~n20698 ;
  assign y6407 = ~n20700 ;
  assign y6408 = ~n20701 ;
  assign y6409 = ~n20703 ;
  assign y6410 = n20709 ;
  assign y6411 = ~n20715 ;
  assign y6412 = ~1'b0 ;
  assign y6413 = ~n20716 ;
  assign y6414 = n20719 ;
  assign y6415 = n20723 ;
  assign y6416 = ~1'b0 ;
  assign y6417 = ~n20730 ;
  assign y6418 = n20734 ;
  assign y6419 = ~n20737 ;
  assign y6420 = n20740 ;
  assign y6421 = ~n20743 ;
  assign y6422 = ~n6015 ;
  assign y6423 = n20746 ;
  assign y6424 = ~1'b0 ;
  assign y6425 = n20748 ;
  assign y6426 = ~1'b0 ;
  assign y6427 = ~1'b0 ;
  assign y6428 = ~1'b0 ;
  assign y6429 = ~1'b0 ;
  assign y6430 = ~n20751 ;
  assign y6431 = ~n20756 ;
  assign y6432 = ~n20758 ;
  assign y6433 = n20759 ;
  assign y6434 = n20761 ;
  assign y6435 = ~1'b0 ;
  assign y6436 = n20768 ;
  assign y6437 = ~n20773 ;
  assign y6438 = ~1'b0 ;
  assign y6439 = n20775 ;
  assign y6440 = ~n20778 ;
  assign y6441 = n20786 ;
  assign y6442 = n20795 ;
  assign y6443 = n20800 ;
  assign y6444 = ~n20810 ;
  assign y6445 = n20812 ;
  assign y6446 = n20815 ;
  assign y6447 = ~n20816 ;
  assign y6448 = n20823 ;
  assign y6449 = ~n20829 ;
  assign y6450 = n20835 ;
  assign y6451 = n20837 ;
  assign y6452 = n20839 ;
  assign y6453 = n20841 ;
  assign y6454 = n20844 ;
  assign y6455 = ~n20853 ;
  assign y6456 = n20854 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = n20861 ;
  assign y6459 = ~n20868 ;
  assign y6460 = ~n20882 ;
  assign y6461 = ~1'b0 ;
  assign y6462 = ~n20891 ;
  assign y6463 = n20892 ;
  assign y6464 = ~n20900 ;
  assign y6465 = ~n20902 ;
  assign y6466 = n20903 ;
  assign y6467 = ~n6115 ;
  assign y6468 = ~n20909 ;
  assign y6469 = ~n20914 ;
  assign y6470 = ~n20917 ;
  assign y6471 = ~n20920 ;
  assign y6472 = ~n20924 ;
  assign y6473 = ~n20926 ;
  assign y6474 = ~1'b0 ;
  assign y6475 = ~1'b0 ;
  assign y6476 = ~n20928 ;
  assign y6477 = ~n20929 ;
  assign y6478 = ~n20935 ;
  assign y6479 = n14618 ;
  assign y6480 = ~n20945 ;
  assign y6481 = ~n20946 ;
  assign y6482 = n20949 ;
  assign y6483 = ~n20954 ;
  assign y6484 = n20957 ;
  assign y6485 = ~n20959 ;
  assign y6486 = n14636 ;
  assign y6487 = n20966 ;
  assign y6488 = ~n20973 ;
  assign y6489 = n20976 ;
  assign y6490 = n20981 ;
  assign y6491 = ~n20984 ;
  assign y6492 = ~n20989 ;
  assign y6493 = n20992 ;
  assign y6494 = n20993 ;
  assign y6495 = n20994 ;
  assign y6496 = ~n20996 ;
  assign y6497 = n21001 ;
  assign y6498 = n21002 ;
  assign y6499 = ~n21021 ;
  assign y6500 = n21028 ;
  assign y6501 = n21030 ;
  assign y6502 = ~n21032 ;
  assign y6503 = ~n21035 ;
  assign y6504 = ~1'b0 ;
  assign y6505 = ~1'b0 ;
  assign y6506 = ~n21038 ;
  assign y6507 = ~n21039 ;
  assign y6508 = ~n21041 ;
  assign y6509 = ~n21044 ;
  assign y6510 = n21053 ;
  assign y6511 = n19819 ;
  assign y6512 = ~1'b0 ;
  assign y6513 = ~n21057 ;
  assign y6514 = n21058 ;
  assign y6515 = ~n21061 ;
  assign y6516 = ~1'b0 ;
  assign y6517 = ~n21064 ;
  assign y6518 = n21068 ;
  assign y6519 = ~n21070 ;
  assign y6520 = ~1'b0 ;
  assign y6521 = ~n21073 ;
  assign y6522 = n21079 ;
  assign y6523 = n21082 ;
  assign y6524 = ~n21089 ;
  assign y6525 = n21093 ;
  assign y6526 = n21100 ;
  assign y6527 = ~n21101 ;
  assign y6528 = n21106 ;
  assign y6529 = n21110 ;
  assign y6530 = n21111 ;
  assign y6531 = n21112 ;
  assign y6532 = ~1'b0 ;
  assign y6533 = ~1'b0 ;
  assign y6534 = n21116 ;
  assign y6535 = n21121 ;
  assign y6536 = n21122 ;
  assign y6537 = n21123 ;
  assign y6538 = ~n21126 ;
  assign y6539 = ~n15572 ;
  assign y6540 = ~n21129 ;
  assign y6541 = ~1'b0 ;
  assign y6542 = n21130 ;
  assign y6543 = ~n21135 ;
  assign y6544 = n21137 ;
  assign y6545 = ~n21140 ;
  assign y6546 = ~n21143 ;
  assign y6547 = ~n21146 ;
  assign y6548 = ~n21147 ;
  assign y6549 = n21149 ;
  assign y6550 = ~1'b0 ;
  assign y6551 = ~n21150 ;
  assign y6552 = ~n21156 ;
  assign y6553 = n21158 ;
  assign y6554 = ~n21164 ;
  assign y6555 = n21166 ;
  assign y6556 = ~1'b0 ;
  assign y6557 = ~1'b0 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = n21167 ;
  assign y6560 = n21170 ;
  assign y6561 = ~n21171 ;
  assign y6562 = ~n21172 ;
  assign y6563 = n21173 ;
  assign y6564 = ~n21175 ;
  assign y6565 = ~n21180 ;
  assign y6566 = n21181 ;
  assign y6567 = n21190 ;
  assign y6568 = ~n21192 ;
  assign y6569 = n21193 ;
  assign y6570 = ~n21195 ;
  assign y6571 = ~n21197 ;
  assign y6572 = n21200 ;
  assign y6573 = n21204 ;
  assign y6574 = ~n21205 ;
  assign y6575 = ~n21213 ;
  assign y6576 = ~1'b0 ;
  assign y6577 = n21214 ;
  assign y6578 = ~n21218 ;
  assign y6579 = ~1'b0 ;
  assign y6580 = ~n21222 ;
  assign y6581 = ~1'b0 ;
  assign y6582 = ~n21227 ;
  assign y6583 = n21229 ;
  assign y6584 = ~n21231 ;
  assign y6585 = ~1'b0 ;
  assign y6586 = n21234 ;
  assign y6587 = ~n21238 ;
  assign y6588 = n21239 ;
  assign y6589 = ~n21246 ;
  assign y6590 = ~n21250 ;
  assign y6591 = ~n21256 ;
  assign y6592 = n21258 ;
  assign y6593 = n21263 ;
  assign y6594 = n21264 ;
  assign y6595 = n21266 ;
  assign y6596 = 1'b0 ;
  assign y6597 = ~n21269 ;
  assign y6598 = n21271 ;
  assign y6599 = n21280 ;
  assign y6600 = ~n21288 ;
  assign y6601 = n21289 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = ~n21291 ;
  assign y6605 = n21292 ;
  assign y6606 = ~n21293 ;
  assign y6607 = ~1'b0 ;
  assign y6608 = ~1'b0 ;
  assign y6609 = n21301 ;
  assign y6610 = ~n21308 ;
  assign y6611 = n21311 ;
  assign y6612 = n21316 ;
  assign y6613 = ~n21318 ;
  assign y6614 = n21324 ;
  assign y6615 = ~n21325 ;
  assign y6616 = n21333 ;
  assign y6617 = ~n21337 ;
  assign y6618 = ~n21339 ;
  assign y6619 = 1'b0 ;
  assign y6620 = ~n21342 ;
  assign y6621 = ~n21346 ;
  assign y6622 = n21351 ;
  assign y6623 = n21363 ;
  assign y6624 = ~n21364 ;
  assign y6625 = ~1'b0 ;
  assign y6626 = n21368 ;
  assign y6627 = n21370 ;
  assign y6628 = n21374 ;
  assign y6629 = ~n21377 ;
  assign y6630 = ~1'b0 ;
  assign y6631 = ~n21380 ;
  assign y6632 = ~n21387 ;
  assign y6633 = ~n21388 ;
  assign y6634 = n21391 ;
  assign y6635 = n21396 ;
  assign y6636 = ~n21397 ;
  assign y6637 = ~n21407 ;
  assign y6638 = n21411 ;
  assign y6639 = ~n21415 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = ~n21417 ;
  assign y6642 = 1'b0 ;
  assign y6643 = n21421 ;
  assign y6644 = ~n21425 ;
  assign y6645 = ~n21433 ;
  assign y6646 = n21439 ;
  assign y6647 = ~n21442 ;
  assign y6648 = n21443 ;
  assign y6649 = n21447 ;
  assign y6650 = n21458 ;
  assign y6651 = n21477 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = ~1'b0 ;
  assign y6654 = ~n21480 ;
  assign y6655 = n21484 ;
  assign y6656 = ~1'b0 ;
  assign y6657 = ~1'b0 ;
  assign y6658 = n21485 ;
  assign y6659 = ~n21491 ;
  assign y6660 = ~n21493 ;
  assign y6661 = ~1'b0 ;
  assign y6662 = ~1'b0 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = ~n21495 ;
  assign y6665 = n21512 ;
  assign y6666 = n21513 ;
  assign y6667 = ~n21514 ;
  assign y6668 = n21517 ;
  assign y6669 = n21519 ;
  assign y6670 = ~1'b0 ;
  assign y6671 = n21521 ;
  assign y6672 = ~1'b0 ;
  assign y6673 = ~n21525 ;
  assign y6674 = n21528 ;
  assign y6675 = ~n21529 ;
  assign y6676 = n3694 ;
  assign y6677 = ~1'b0 ;
  assign y6678 = ~n21531 ;
  assign y6679 = ~n21534 ;
  assign y6680 = n21535 ;
  assign y6681 = ~n21540 ;
  assign y6682 = ~1'b0 ;
  assign y6683 = ~n21544 ;
  assign y6684 = n21546 ;
  assign y6685 = ~n21547 ;
  assign y6686 = ~n21548 ;
  assign y6687 = ~n21553 ;
  assign y6688 = n21557 ;
  assign y6689 = ~n21559 ;
  assign y6690 = ~n21563 ;
  assign y6691 = n21564 ;
  assign y6692 = n21567 ;
  assign y6693 = ~n21570 ;
  assign y6694 = ~n21571 ;
  assign y6695 = n21572 ;
  assign y6696 = ~n21574 ;
  assign y6697 = n21579 ;
  assign y6698 = ~1'b0 ;
  assign y6699 = ~n21584 ;
  assign y6700 = n21586 ;
  assign y6701 = ~n21587 ;
  assign y6702 = ~n21590 ;
  assign y6703 = n21592 ;
  assign y6704 = ~n21594 ;
  assign y6705 = n11332 ;
  assign y6706 = ~1'b0 ;
  assign y6707 = n21595 ;
  assign y6708 = n2985 ;
  assign y6709 = n21598 ;
  assign y6710 = ~n21599 ;
  assign y6711 = ~n21601 ;
  assign y6712 = ~n21603 ;
  assign y6713 = ~n21605 ;
  assign y6714 = n21609 ;
  assign y6715 = ~n21610 ;
  assign y6716 = ~1'b0 ;
  assign y6717 = ~n21612 ;
  assign y6718 = ~n21614 ;
  assign y6719 = n21615 ;
  assign y6720 = n21618 ;
  assign y6721 = ~n21619 ;
  assign y6722 = n21620 ;
  assign y6723 = n21626 ;
  assign y6724 = n21627 ;
  assign y6725 = ~1'b0 ;
  assign y6726 = n21631 ;
  assign y6727 = ~n21636 ;
  assign y6728 = ~1'b0 ;
  assign y6729 = n21640 ;
  assign y6730 = ~n21641 ;
  assign y6731 = n21650 ;
  assign y6732 = ~n21651 ;
  assign y6733 = ~n21654 ;
  assign y6734 = ~n21656 ;
  assign y6735 = ~n21657 ;
  assign y6736 = ~1'b0 ;
  assign y6737 = n21659 ;
  assign y6738 = ~n21665 ;
  assign y6739 = ~n21667 ;
  assign y6740 = ~1'b0 ;
  assign y6741 = ~1'b0 ;
  assign y6742 = ~n21668 ;
  assign y6743 = ~n21673 ;
  assign y6744 = ~n21675 ;
  assign y6745 = ~n21676 ;
  assign y6746 = ~n21677 ;
  assign y6747 = ~1'b0 ;
  assign y6748 = ~n21684 ;
  assign y6749 = n21688 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = n21691 ;
  assign y6752 = ~n21694 ;
  assign y6753 = n21696 ;
  assign y6754 = n21702 ;
  assign y6755 = ~n21703 ;
  assign y6756 = n21708 ;
  assign y6757 = n21715 ;
  assign y6758 = n21717 ;
  assign y6759 = n21719 ;
  assign y6760 = ~n21724 ;
  assign y6761 = n4062 ;
  assign y6762 = ~n12041 ;
  assign y6763 = ~1'b0 ;
  assign y6764 = ~n21734 ;
  assign y6765 = ~n21735 ;
  assign y6766 = n21747 ;
  assign y6767 = ~n21749 ;
  assign y6768 = n21758 ;
  assign y6769 = n21772 ;
  assign y6770 = n21774 ;
  assign y6771 = ~n21777 ;
  assign y6772 = n21782 ;
  assign y6773 = ~1'b0 ;
  assign y6774 = ~n21785 ;
  assign y6775 = ~n21786 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~n21788 ;
  assign y6778 = ~n21793 ;
  assign y6779 = n21796 ;
  assign y6780 = ~n21802 ;
  assign y6781 = ~1'b0 ;
  assign y6782 = ~1'b0 ;
  assign y6783 = ~n21805 ;
  assign y6784 = n21806 ;
  assign y6785 = n21809 ;
  assign y6786 = ~1'b0 ;
  assign y6787 = ~n21812 ;
  assign y6788 = n21814 ;
  assign y6789 = n21816 ;
  assign y6790 = n21820 ;
  assign y6791 = ~1'b0 ;
  assign y6792 = n21821 ;
  assign y6793 = ~n21824 ;
  assign y6794 = n21827 ;
  assign y6795 = n21829 ;
  assign y6796 = n21839 ;
  assign y6797 = ~n21841 ;
  assign y6798 = ~n21842 ;
  assign y6799 = n21851 ;
  assign y6800 = ~n5608 ;
  assign y6801 = ~n21853 ;
  assign y6802 = ~n21854 ;
  assign y6803 = ~n21867 ;
  assign y6804 = n21874 ;
  assign y6805 = n21881 ;
  assign y6806 = ~1'b0 ;
  assign y6807 = n21882 ;
  assign y6808 = n21884 ;
  assign y6809 = ~n21885 ;
  assign y6810 = ~n21887 ;
  assign y6811 = n21896 ;
  assign y6812 = n21898 ;
  assign y6813 = n21899 ;
  assign y6814 = ~n21901 ;
  assign y6815 = n21902 ;
  assign y6816 = n21903 ;
  assign y6817 = ~n21905 ;
  assign y6818 = n21910 ;
  assign y6819 = ~n21912 ;
  assign y6820 = ~n21915 ;
  assign y6821 = ~n14636 ;
  assign y6822 = n21920 ;
  assign y6823 = ~n21925 ;
  assign y6824 = n21930 ;
  assign y6825 = ~1'b0 ;
  assign y6826 = n21934 ;
  assign y6827 = n21937 ;
  assign y6828 = ~n21938 ;
  assign y6829 = n21939 ;
  assign y6830 = n21940 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = ~n21948 ;
  assign y6833 = ~n21953 ;
  assign y6834 = n21955 ;
  assign y6835 = ~n21957 ;
  assign y6836 = ~n21960 ;
  assign y6837 = ~1'b0 ;
  assign y6838 = n21963 ;
  assign y6839 = ~n21977 ;
  assign y6840 = ~1'b0 ;
  assign y6841 = n21979 ;
  assign y6842 = n21988 ;
  assign y6843 = n21995 ;
  assign y6844 = n21996 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = ~n21997 ;
  assign y6847 = ~n22000 ;
  assign y6848 = n22005 ;
  assign y6849 = ~1'b0 ;
  assign y6850 = n22010 ;
  assign y6851 = ~1'b0 ;
  assign y6852 = ~n22011 ;
  assign y6853 = ~1'b0 ;
  assign y6854 = n22017 ;
  assign y6855 = ~n22023 ;
  assign y6856 = n22027 ;
  assign y6857 = n22030 ;
  assign y6858 = ~n22036 ;
  assign y6859 = ~n22044 ;
  assign y6860 = ~n22045 ;
  assign y6861 = ~n22051 ;
  assign y6862 = n22052 ;
  assign y6863 = n22054 ;
  assign y6864 = ~n22066 ;
  assign y6865 = ~n22070 ;
  assign y6866 = ~1'b0 ;
  assign y6867 = ~n7563 ;
  assign y6868 = ~n22072 ;
  assign y6869 = ~n22073 ;
  assign y6870 = n22074 ;
  assign y6871 = ~1'b0 ;
  assign y6872 = ~1'b0 ;
  assign y6873 = ~n22078 ;
  assign y6874 = ~n22080 ;
  assign y6875 = ~n22084 ;
  assign y6876 = ~n22086 ;
  assign y6877 = ~n22094 ;
  assign y6878 = ~1'b0 ;
  assign y6879 = ~n22102 ;
  assign y6880 = n22103 ;
  assign y6881 = ~1'b0 ;
  assign y6882 = ~n22112 ;
  assign y6883 = ~n22115 ;
  assign y6884 = ~n22122 ;
  assign y6885 = ~n22123 ;
  assign y6886 = ~n22128 ;
  assign y6887 = ~n22137 ;
  assign y6888 = n22140 ;
  assign y6889 = n22144 ;
  assign y6890 = ~1'b0 ;
  assign y6891 = ~1'b0 ;
  assign y6892 = ~1'b0 ;
  assign y6893 = n22146 ;
  assign y6894 = ~n22148 ;
  assign y6895 = ~n22156 ;
  assign y6896 = n22157 ;
  assign y6897 = n22166 ;
  assign y6898 = ~n22169 ;
  assign y6899 = ~n22175 ;
  assign y6900 = n22176 ;
  assign y6901 = ~n22177 ;
  assign y6902 = ~n22183 ;
  assign y6903 = ~1'b0 ;
  assign y6904 = ~n22186 ;
  assign y6905 = ~1'b0 ;
  assign y6906 = ~n22189 ;
  assign y6907 = n22196 ;
  assign y6908 = ~n22197 ;
  assign y6909 = ~n19077 ;
  assign y6910 = ~n22198 ;
  assign y6911 = n22200 ;
  assign y6912 = ~n22204 ;
  assign y6913 = n22205 ;
  assign y6914 = ~n22209 ;
  assign y6915 = n22218 ;
  assign y6916 = ~n22224 ;
  assign y6917 = ~n22228 ;
  assign y6918 = ~n22232 ;
  assign y6919 = ~n22236 ;
  assign y6920 = n22242 ;
  assign y6921 = ~n22243 ;
  assign y6922 = ~n22244 ;
  assign y6923 = n22247 ;
  assign y6924 = ~n22248 ;
  assign y6925 = ~1'b0 ;
  assign y6926 = n22254 ;
  assign y6927 = ~n19657 ;
  assign y6928 = n22255 ;
  assign y6929 = n22261 ;
  assign y6930 = ~n22263 ;
  assign y6931 = n22265 ;
  assign y6932 = ~n22267 ;
  assign y6933 = n22268 ;
  assign y6934 = n22270 ;
  assign y6935 = ~n22276 ;
  assign y6936 = ~1'b0 ;
  assign y6937 = n22279 ;
  assign y6938 = ~n22289 ;
  assign y6939 = ~n22295 ;
  assign y6940 = ~n22296 ;
  assign y6941 = ~n22307 ;
  assign y6942 = n22315 ;
  assign y6943 = n22317 ;
  assign y6944 = ~n22319 ;
  assign y6945 = ~1'b0 ;
  assign y6946 = n22322 ;
  assign y6947 = n22324 ;
  assign y6948 = ~1'b0 ;
  assign y6949 = ~n22328 ;
  assign y6950 = n22329 ;
  assign y6951 = n22330 ;
  assign y6952 = ~1'b0 ;
  assign y6953 = n22331 ;
  assign y6954 = ~n22339 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = ~1'b0 ;
  assign y6957 = ~1'b0 ;
  assign y6958 = n12624 ;
  assign y6959 = n22341 ;
  assign y6960 = ~n22347 ;
  assign y6961 = n12200 ;
  assign y6962 = ~n22349 ;
  assign y6963 = n22350 ;
  assign y6964 = n22352 ;
  assign y6965 = ~n22354 ;
  assign y6966 = ~n22355 ;
  assign y6967 = 1'b0 ;
  assign y6968 = n22357 ;
  assign y6969 = ~n22359 ;
  assign y6970 = ~1'b0 ;
  assign y6971 = ~n22364 ;
  assign y6972 = ~n22368 ;
  assign y6973 = ~n22370 ;
  assign y6974 = ~n22373 ;
  assign y6975 = n22376 ;
  assign y6976 = ~n22379 ;
  assign y6977 = ~1'b0 ;
  assign y6978 = n22386 ;
  assign y6979 = ~n22388 ;
  assign y6980 = ~1'b0 ;
  assign y6981 = ~n22391 ;
  assign y6982 = ~n22393 ;
  assign y6983 = n22396 ;
  assign y6984 = ~n22400 ;
  assign y6985 = n22402 ;
  assign y6986 = ~n22403 ;
  assign y6987 = ~n22405 ;
  assign y6988 = n22408 ;
  assign y6989 = n22410 ;
  assign y6990 = n22412 ;
  assign y6991 = n22417 ;
  assign y6992 = n22421 ;
  assign y6993 = n22423 ;
  assign y6994 = ~n22425 ;
  assign y6995 = ~1'b0 ;
  assign y6996 = ~1'b0 ;
  assign y6997 = ~n22427 ;
  assign y6998 = n22428 ;
  assign y6999 = n22429 ;
  assign y7000 = ~n22430 ;
  assign y7001 = ~n22432 ;
  assign y7002 = ~n22435 ;
  assign y7003 = ~n22440 ;
  assign y7004 = n22442 ;
  assign y7005 = ~1'b0 ;
  assign y7006 = ~n22445 ;
  assign y7007 = ~n22455 ;
  assign y7008 = n22459 ;
  assign y7009 = n22461 ;
  assign y7010 = ~1'b0 ;
  assign y7011 = ~1'b0 ;
  assign y7012 = n22466 ;
  assign y7013 = n22476 ;
  assign y7014 = ~n22479 ;
  assign y7015 = ~1'b0 ;
  assign y7016 = ~n22485 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = ~n22489 ;
  assign y7019 = n22492 ;
  assign y7020 = ~n22500 ;
  assign y7021 = n22502 ;
  assign y7022 = ~1'b0 ;
  assign y7023 = n22503 ;
  assign y7024 = ~n22506 ;
  assign y7025 = ~n22511 ;
  assign y7026 = ~n22513 ;
  assign y7027 = n10729 ;
  assign y7028 = n22515 ;
  assign y7029 = n22521 ;
  assign y7030 = n22526 ;
  assign y7031 = ~n22530 ;
  assign y7032 = ~n22534 ;
  assign y7033 = n22539 ;
  assign y7034 = n22543 ;
  assign y7035 = ~n22544 ;
  assign y7036 = ~n22547 ;
  assign y7037 = n22549 ;
  assign y7038 = ~n22552 ;
  assign y7039 = ~n22554 ;
  assign y7040 = n22562 ;
  assign y7041 = ~n22570 ;
  assign y7042 = ~1'b0 ;
  assign y7043 = ~n22574 ;
  assign y7044 = n22576 ;
  assign y7045 = ~n22580 ;
  assign y7046 = ~n22582 ;
  assign y7047 = n22584 ;
  assign y7048 = ~n22587 ;
  assign y7049 = n22588 ;
  assign y7050 = ~n22591 ;
  assign y7051 = n22599 ;
  assign y7052 = n22603 ;
  assign y7053 = ~1'b0 ;
  assign y7054 = ~n22606 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = n22610 ;
  assign y7058 = ~n22611 ;
  assign y7059 = n22615 ;
  assign y7060 = n22617 ;
  assign y7061 = ~n22626 ;
  assign y7062 = ~n22627 ;
  assign y7063 = n8881 ;
  assign y7064 = ~n22630 ;
  assign y7065 = n22637 ;
  assign y7066 = n22642 ;
  assign y7067 = ~1'b0 ;
  assign y7068 = ~n22643 ;
  assign y7069 = ~1'b0 ;
  assign y7070 = ~1'b0 ;
  assign y7071 = n22654 ;
  assign y7072 = ~n22655 ;
  assign y7073 = n22656 ;
  assign y7074 = ~1'b0 ;
  assign y7075 = n22657 ;
  assign y7076 = n22661 ;
  assign y7077 = ~n22663 ;
  assign y7078 = n22665 ;
  assign y7079 = ~1'b0 ;
  assign y7080 = ~1'b0 ;
  assign y7081 = n22670 ;
  assign y7082 = n22672 ;
  assign y7083 = n22681 ;
  assign y7084 = ~1'b0 ;
  assign y7085 = ~n22684 ;
  assign y7086 = ~n22691 ;
  assign y7087 = ~1'b0 ;
  assign y7088 = ~n22694 ;
  assign y7089 = n22697 ;
  assign y7090 = n22699 ;
  assign y7091 = ~n22701 ;
  assign y7092 = ~1'b0 ;
  assign y7093 = ~n22705 ;
  assign y7094 = n22710 ;
  assign y7095 = ~n22715 ;
  assign y7096 = ~1'b0 ;
  assign y7097 = ~n22721 ;
  assign y7098 = ~n22723 ;
  assign y7099 = ~n22727 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = n22729 ;
  assign y7102 = n22730 ;
  assign y7103 = ~n22731 ;
  assign y7104 = ~n22735 ;
  assign y7105 = n22737 ;
  assign y7106 = ~1'b0 ;
  assign y7107 = n1352 ;
  assign y7108 = n22740 ;
  assign y7109 = n22744 ;
  assign y7110 = ~1'b0 ;
  assign y7111 = ~n22749 ;
  assign y7112 = ~n22755 ;
  assign y7113 = n22757 ;
  assign y7114 = ~n22762 ;
  assign y7115 = ~n22766 ;
  assign y7116 = n22768 ;
  assign y7117 = n22770 ;
  assign y7118 = n22771 ;
  assign y7119 = n22775 ;
  assign y7120 = ~n22776 ;
  assign y7121 = ~1'b0 ;
  assign y7122 = ~n22778 ;
  assign y7123 = ~1'b0 ;
  assign y7124 = ~n22780 ;
  assign y7125 = ~n22781 ;
  assign y7126 = ~n22782 ;
  assign y7127 = ~1'b0 ;
  assign y7128 = ~n22784 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~1'b0 ;
  assign y7131 = ~n22053 ;
  assign y7132 = ~n22786 ;
  assign y7133 = n22787 ;
  assign y7134 = n22791 ;
  assign y7135 = n22810 ;
  assign y7136 = n22813 ;
  assign y7137 = ~n22815 ;
  assign y7138 = n22819 ;
  assign y7139 = ~n22823 ;
  assign y7140 = ~n22830 ;
  assign y7141 = n22832 ;
  assign y7142 = ~1'b0 ;
  assign y7143 = ~n22834 ;
  assign y7144 = n22839 ;
  assign y7145 = ~n22842 ;
  assign y7146 = n22849 ;
  assign y7147 = ~n22860 ;
  assign y7148 = ~n22863 ;
  assign y7149 = ~n22869 ;
  assign y7150 = n22874 ;
  assign y7151 = n22876 ;
  assign y7152 = ~1'b0 ;
  assign y7153 = ~n22878 ;
  assign y7154 = n22880 ;
  assign y7155 = ~n22883 ;
  assign y7156 = ~n22884 ;
  assign y7157 = n22886 ;
  assign y7158 = n22889 ;
  assign y7159 = n22890 ;
  assign y7160 = n22895 ;
  assign y7161 = ~1'b0 ;
  assign y7162 = n22897 ;
  assign y7163 = ~n22900 ;
  assign y7164 = ~n22901 ;
  assign y7165 = n22906 ;
  assign y7166 = n22909 ;
  assign y7167 = n22917 ;
  assign y7168 = ~1'b0 ;
  assign y7169 = ~n22920 ;
  assign y7170 = n22924 ;
  assign y7171 = n22930 ;
  assign y7172 = n22933 ;
  assign y7173 = ~n22935 ;
  assign y7174 = ~1'b0 ;
  assign y7175 = n22940 ;
  assign y7176 = ~1'b0 ;
  assign y7177 = n22942 ;
  assign y7178 = ~n22946 ;
  assign y7179 = ~1'b0 ;
  assign y7180 = ~n22949 ;
  assign y7181 = n22951 ;
  assign y7182 = ~n22953 ;
  assign y7183 = ~n22957 ;
  assign y7184 = n22960 ;
  assign y7185 = n22972 ;
  assign y7186 = ~n22976 ;
  assign y7187 = ~n22977 ;
  assign y7188 = ~n22978 ;
  assign y7189 = ~n22985 ;
  assign y7190 = n22991 ;
  assign y7191 = n22993 ;
  assign y7192 = n22994 ;
  assign y7193 = n22997 ;
  assign y7194 = ~n22999 ;
  assign y7195 = ~1'b0 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = n23000 ;
  assign y7198 = n23012 ;
  assign y7199 = n23013 ;
  assign y7200 = ~1'b0 ;
  assign y7201 = ~n23015 ;
  assign y7202 = n23019 ;
  assign y7203 = ~1'b0 ;
  assign y7204 = ~n23025 ;
  assign y7205 = ~1'b0 ;
  assign y7206 = ~1'b0 ;
  assign y7207 = ~n23026 ;
  assign y7208 = ~1'b0 ;
  assign y7209 = ~1'b0 ;
  assign y7210 = ~n23027 ;
  assign y7211 = n23043 ;
  assign y7212 = ~n23048 ;
  assign y7213 = n23060 ;
  assign y7214 = ~n10579 ;
  assign y7215 = n23062 ;
  assign y7216 = n23065 ;
  assign y7217 = n23068 ;
  assign y7218 = n23069 ;
  assign y7219 = n23070 ;
  assign y7220 = n23071 ;
  assign y7221 = n23074 ;
  assign y7222 = n23078 ;
  assign y7223 = ~n23082 ;
  assign y7224 = n13749 ;
  assign y7225 = n23090 ;
  assign y7226 = ~n23093 ;
  assign y7227 = n23094 ;
  assign y7228 = ~n23096 ;
  assign y7229 = ~1'b0 ;
  assign y7230 = ~n23101 ;
  assign y7231 = n23104 ;
  assign y7232 = n23107 ;
  assign y7233 = ~1'b0 ;
  assign y7234 = ~n23112 ;
  assign y7235 = ~n23117 ;
  assign y7236 = ~n23120 ;
  assign y7237 = n23121 ;
  assign y7238 = n23127 ;
  assign y7239 = n23130 ;
  assign y7240 = ~1'b0 ;
  assign y7241 = ~n23132 ;
  assign y7242 = ~n23133 ;
  assign y7243 = n23134 ;
  assign y7244 = ~n23138 ;
  assign y7245 = ~n23139 ;
  assign y7246 = ~1'b0 ;
  assign y7247 = n23146 ;
  assign y7248 = n23147 ;
  assign y7249 = n23150 ;
  assign y7250 = ~n23154 ;
  assign y7251 = ~1'b0 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = ~1'b0 ;
  assign y7254 = ~n23157 ;
  assign y7255 = ~n23164 ;
  assign y7256 = ~n23169 ;
  assign y7257 = n23172 ;
  assign y7258 = ~n23174 ;
  assign y7259 = ~n23176 ;
  assign y7260 = n23180 ;
  assign y7261 = ~n23182 ;
  assign y7262 = ~n23184 ;
  assign y7263 = n23187 ;
  assign y7264 = ~n23188 ;
  assign y7265 = n23190 ;
  assign y7266 = ~n23196 ;
  assign y7267 = ~n23198 ;
  assign y7268 = ~n23201 ;
  assign y7269 = ~n23205 ;
  assign y7270 = ~n23206 ;
  assign y7271 = n23209 ;
  assign y7272 = ~n23214 ;
  assign y7273 = n23216 ;
  assign y7274 = ~n23221 ;
  assign y7275 = ~1'b0 ;
  assign y7276 = n23223 ;
  assign y7277 = n23224 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = ~n23227 ;
  assign y7280 = n23229 ;
  assign y7281 = n23231 ;
  assign y7282 = n23233 ;
  assign y7283 = n23236 ;
  assign y7284 = n23250 ;
  assign y7285 = n23252 ;
  assign y7286 = ~1'b0 ;
  assign y7287 = n23256 ;
  assign y7288 = n23257 ;
  assign y7289 = n23261 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~1'b0 ;
  assign y7292 = n23272 ;
  assign y7293 = 1'b0 ;
  assign y7294 = n23275 ;
  assign y7295 = ~n23278 ;
  assign y7296 = ~n23282 ;
  assign y7297 = n11768 ;
  assign y7298 = ~n23284 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = n23287 ;
  assign y7301 = ~n23290 ;
  assign y7302 = n23293 ;
  assign y7303 = ~n23295 ;
  assign y7304 = ~1'b0 ;
  assign y7305 = n23297 ;
  assign y7306 = ~1'b0 ;
  assign y7307 = n23299 ;
  assign y7308 = ~n23303 ;
  assign y7309 = ~n23306 ;
  assign y7310 = ~1'b0 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = n23308 ;
  assign y7313 = ~n23310 ;
  assign y7314 = n23312 ;
  assign y7315 = n23320 ;
  assign y7316 = ~1'b0 ;
  assign y7317 = ~1'b0 ;
  assign y7318 = n23323 ;
  assign y7319 = n23325 ;
  assign y7320 = n23328 ;
  assign y7321 = n23330 ;
  assign y7322 = n23334 ;
  assign y7323 = n23338 ;
  assign y7324 = n23340 ;
  assign y7325 = n23342 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = n23347 ;
  assign y7328 = ~n23351 ;
  assign y7329 = n23355 ;
  assign y7330 = ~n23361 ;
  assign y7331 = n23364 ;
  assign y7332 = ~n23368 ;
  assign y7333 = n23373 ;
  assign y7334 = ~1'b0 ;
  assign y7335 = n23374 ;
  assign y7336 = n23377 ;
  assign y7337 = n23379 ;
  assign y7338 = ~n23381 ;
  assign y7339 = n23385 ;
  assign y7340 = ~n23388 ;
  assign y7341 = ~n23390 ;
  assign y7342 = ~1'b0 ;
  assign y7343 = ~1'b0 ;
  assign y7344 = n23391 ;
  assign y7345 = ~1'b0 ;
  assign y7346 = n23393 ;
  assign y7347 = ~n23394 ;
  assign y7348 = ~n23395 ;
  assign y7349 = n23404 ;
  assign y7350 = ~1'b0 ;
  assign y7351 = ~1'b0 ;
  assign y7352 = n23405 ;
  assign y7353 = n23411 ;
  assign y7354 = n23412 ;
  assign y7355 = ~1'b0 ;
  assign y7356 = n23413 ;
  assign y7357 = ~1'b0 ;
  assign y7358 = n23414 ;
  assign y7359 = n23420 ;
  assign y7360 = n23422 ;
  assign y7361 = n23429 ;
  assign y7362 = ~n23436 ;
  assign y7363 = ~n23440 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = n23441 ;
  assign y7366 = ~n23442 ;
  assign y7367 = ~1'b0 ;
  assign y7368 = ~1'b0 ;
  assign y7369 = n23443 ;
  assign y7370 = ~1'b0 ;
  assign y7371 = ~n23445 ;
  assign y7372 = n23447 ;
  assign y7373 = ~n23452 ;
  assign y7374 = n23462 ;
  assign y7375 = ~n23463 ;
  assign y7376 = n23466 ;
  assign y7377 = n23471 ;
  assign y7378 = ~n23481 ;
  assign y7379 = n23488 ;
  assign y7380 = n23491 ;
  assign y7381 = ~n2553 ;
  assign y7382 = ~n23492 ;
  assign y7383 = n23497 ;
  assign y7384 = ~n23499 ;
  assign y7385 = ~n23503 ;
  assign y7386 = n23507 ;
  assign y7387 = ~n23508 ;
  assign y7388 = ~n23509 ;
  assign y7389 = n23514 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = n23516 ;
  assign y7392 = ~n23520 ;
  assign y7393 = ~n23525 ;
  assign y7394 = ~n23530 ;
  assign y7395 = n23534 ;
  assign y7396 = n23536 ;
  assign y7397 = ~1'b0 ;
  assign y7398 = n23539 ;
  assign y7399 = n23540 ;
  assign y7400 = ~1'b0 ;
  assign y7401 = ~1'b0 ;
  assign y7402 = ~n23541 ;
  assign y7403 = ~n23546 ;
  assign y7404 = n23548 ;
  assign y7405 = ~1'b0 ;
  assign y7406 = n23553 ;
  assign y7407 = ~n23554 ;
  assign y7408 = ~n23560 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = ~1'b0 ;
  assign y7411 = ~1'b0 ;
  assign y7412 = ~n23563 ;
  assign y7413 = ~n23566 ;
  assign y7414 = n23567 ;
  assign y7415 = n23571 ;
  assign y7416 = n23572 ;
  assign y7417 = ~1'b0 ;
  assign y7418 = ~n23584 ;
  assign y7419 = n23585 ;
  assign y7420 = n23588 ;
  assign y7421 = ~1'b0 ;
  assign y7422 = ~n23595 ;
  assign y7423 = ~n23600 ;
  assign y7424 = ~n23601 ;
  assign y7425 = ~n23603 ;
  assign y7426 = n23613 ;
  assign y7427 = ~n23615 ;
  assign y7428 = ~n23617 ;
  assign y7429 = ~1'b0 ;
  assign y7430 = n23621 ;
  assign y7431 = ~n23624 ;
  assign y7432 = n23630 ;
  assign y7433 = n23634 ;
  assign y7434 = ~n23639 ;
  assign y7435 = ~n23643 ;
  assign y7436 = n23647 ;
  assign y7437 = n23649 ;
  assign y7438 = ~n23653 ;
  assign y7439 = ~n23656 ;
  assign y7440 = ~n23657 ;
  assign y7441 = ~n23661 ;
  assign y7442 = n23663 ;
  assign y7443 = ~n23665 ;
  assign y7444 = ~n23673 ;
  assign y7445 = ~n841 ;
  assign y7446 = n23681 ;
  assign y7447 = ~1'b0 ;
  assign y7448 = n23682 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = ~n23683 ;
  assign y7451 = ~1'b0 ;
  assign y7452 = ~n23691 ;
  assign y7453 = ~n23692 ;
  assign y7454 = ~n7466 ;
  assign y7455 = ~n23698 ;
  assign y7456 = ~n23702 ;
  assign y7457 = ~n23706 ;
  assign y7458 = ~n23710 ;
  assign y7459 = n23712 ;
  assign y7460 = ~n23713 ;
  assign y7461 = ~1'b0 ;
  assign y7462 = ~n23715 ;
  assign y7463 = ~1'b0 ;
  assign y7464 = ~n23717 ;
  assign y7465 = n23719 ;
  assign y7466 = ~1'b0 ;
  assign y7467 = ~n23720 ;
  assign y7468 = n23721 ;
  assign y7469 = n23723 ;
  assign y7470 = ~n23726 ;
  assign y7471 = ~1'b0 ;
  assign y7472 = ~n23727 ;
  assign y7473 = n23729 ;
  assign y7474 = ~n23730 ;
  assign y7475 = n23732 ;
  assign y7476 = ~n23734 ;
  assign y7477 = ~n23742 ;
  assign y7478 = ~1'b0 ;
  assign y7479 = n23743 ;
  assign y7480 = ~1'b0 ;
  assign y7481 = ~n23752 ;
  assign y7482 = n23753 ;
  assign y7483 = n23755 ;
  assign y7484 = n23756 ;
  assign y7485 = n23757 ;
  assign y7486 = ~n23764 ;
  assign y7487 = ~n23765 ;
  assign y7488 = n23768 ;
  assign y7489 = ~n23770 ;
  assign y7490 = ~n23773 ;
  assign y7491 = n23775 ;
  assign y7492 = ~1'b0 ;
  assign y7493 = n23779 ;
  assign y7494 = ~1'b0 ;
  assign y7495 = ~n23785 ;
  assign y7496 = n23786 ;
  assign y7497 = n23787 ;
  assign y7498 = n23792 ;
  assign y7499 = ~n23794 ;
  assign y7500 = ~n23802 ;
  assign y7501 = n23810 ;
  assign y7502 = ~n23811 ;
  assign y7503 = n23813 ;
  assign y7504 = ~n23819 ;
  assign y7505 = ~n23828 ;
  assign y7506 = n23831 ;
  assign y7507 = ~n23834 ;
  assign y7508 = ~1'b0 ;
  assign y7509 = ~n23840 ;
  assign y7510 = n23843 ;
  assign y7511 = ~1'b0 ;
  assign y7512 = n23847 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = ~1'b0 ;
  assign y7515 = ~n23856 ;
  assign y7516 = ~1'b0 ;
  assign y7517 = ~n23861 ;
  assign y7518 = n23870 ;
  assign y7519 = ~n23872 ;
  assign y7520 = n23876 ;
  assign y7521 = ~n23877 ;
  assign y7522 = n23878 ;
  assign y7523 = n23880 ;
  assign y7524 = ~n23883 ;
  assign y7525 = ~n23884 ;
  assign y7526 = n23887 ;
  assign y7527 = ~n23888 ;
  assign y7528 = n23892 ;
  assign y7529 = ~n23893 ;
  assign y7530 = n23897 ;
  assign y7531 = n23899 ;
  assign y7532 = ~n23902 ;
  assign y7533 = n23908 ;
  assign y7534 = n23909 ;
  assign y7535 = ~n23911 ;
  assign y7536 = ~1'b0 ;
  assign y7537 = ~n23914 ;
  assign y7538 = ~1'b0 ;
  assign y7539 = n23915 ;
  assign y7540 = ~1'b0 ;
  assign y7541 = n23916 ;
  assign y7542 = n23917 ;
  assign y7543 = n23918 ;
  assign y7544 = ~n23919 ;
  assign y7545 = n23927 ;
  assign y7546 = ~1'b0 ;
  assign y7547 = ~n18929 ;
  assign y7548 = n23934 ;
  assign y7549 = n10765 ;
  assign y7550 = n23938 ;
  assign y7551 = n23939 ;
  assign y7552 = n23943 ;
  assign y7553 = ~1'b0 ;
  assign y7554 = ~n23951 ;
  assign y7555 = ~n23954 ;
  assign y7556 = ~n23959 ;
  assign y7557 = ~n23962 ;
  assign y7558 = ~n23964 ;
  assign y7559 = ~1'b0 ;
  assign y7560 = ~n23967 ;
  assign y7561 = ~n23973 ;
  assign y7562 = ~n23974 ;
  assign y7563 = ~n23975 ;
  assign y7564 = n23976 ;
  assign y7565 = ~n23984 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = ~n23987 ;
  assign y7568 = n23990 ;
  assign y7569 = ~n23993 ;
  assign y7570 = n23998 ;
  assign y7571 = n24000 ;
  assign y7572 = n24008 ;
  assign y7573 = n24010 ;
  assign y7574 = ~n24012 ;
  assign y7575 = ~1'b0 ;
  assign y7576 = ~n24013 ;
  assign y7577 = ~1'b0 ;
  assign y7578 = ~n24015 ;
  assign y7579 = n24017 ;
  assign y7580 = ~n24019 ;
  assign y7581 = n24020 ;
  assign y7582 = n24022 ;
  assign y7583 = ~1'b0 ;
  assign y7584 = ~1'b0 ;
  assign y7585 = ~1'b0 ;
  assign y7586 = n24025 ;
  assign y7587 = n24032 ;
  assign y7588 = ~n24034 ;
  assign y7589 = ~1'b0 ;
  assign y7590 = ~n24046 ;
  assign y7591 = ~1'b0 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = ~n24047 ;
  assign y7594 = ~n7790 ;
  assign y7595 = n24061 ;
  assign y7596 = ~1'b0 ;
  assign y7597 = n24069 ;
  assign y7598 = n24070 ;
  assign y7599 = ~n24072 ;
  assign y7600 = ~1'b0 ;
  assign y7601 = ~n24073 ;
  assign y7602 = n24075 ;
  assign y7603 = ~n24077 ;
  assign y7604 = ~1'b0 ;
  assign y7605 = ~n24081 ;
  assign y7606 = ~n24082 ;
  assign y7607 = ~n24084 ;
  assign y7608 = ~n24090 ;
  assign y7609 = ~1'b0 ;
  assign y7610 = n24093 ;
  assign y7611 = ~1'b0 ;
  assign y7612 = ~1'b0 ;
  assign y7613 = n24101 ;
  assign y7614 = ~n24104 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = ~1'b0 ;
  assign y7617 = n24105 ;
  assign y7618 = 1'b0 ;
  assign y7619 = ~n24107 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = n22473 ;
  assign y7622 = ~n24113 ;
  assign y7623 = ~n24116 ;
  assign y7624 = n24119 ;
  assign y7625 = ~n24123 ;
  assign y7626 = n24127 ;
  assign y7627 = ~n24128 ;
  assign y7628 = ~1'b0 ;
  assign y7629 = ~n24133 ;
  assign y7630 = n24136 ;
  assign y7631 = n24141 ;
  assign y7632 = ~n24143 ;
  assign y7633 = n24148 ;
  assign y7634 = n24151 ;
  assign y7635 = ~n24152 ;
  assign y7636 = ~n24159 ;
  assign y7637 = ~n24160 ;
  assign y7638 = ~n24167 ;
  assign y7639 = ~1'b0 ;
  assign y7640 = ~n24171 ;
  assign y7641 = ~n24173 ;
  assign y7642 = ~n24174 ;
  assign y7643 = ~n24176 ;
  assign y7644 = n24181 ;
  assign y7645 = ~1'b0 ;
  assign y7646 = ~n24182 ;
  assign y7647 = ~n24186 ;
  assign y7648 = n24199 ;
  assign y7649 = n24202 ;
  assign y7650 = ~n20125 ;
  assign y7651 = ~n24203 ;
  assign y7652 = ~n24210 ;
  assign y7653 = ~n24211 ;
  assign y7654 = ~n24217 ;
  assign y7655 = n24219 ;
  assign y7656 = n24223 ;
  assign y7657 = ~n24230 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = n24232 ;
  assign y7660 = ~n24236 ;
  assign y7661 = ~n24238 ;
  assign y7662 = n24241 ;
  assign y7663 = ~n16048 ;
  assign y7664 = n24242 ;
  assign y7665 = ~n24245 ;
  assign y7666 = ~n24250 ;
  assign y7667 = ~1'b0 ;
  assign y7668 = n24251 ;
  assign y7669 = ~n24254 ;
  assign y7670 = n24256 ;
  assign y7671 = ~n24257 ;
  assign y7672 = ~1'b0 ;
  assign y7673 = ~n24258 ;
  assign y7674 = n24262 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~n24263 ;
  assign y7677 = n24264 ;
  assign y7678 = ~n24276 ;
  assign y7679 = ~n24278 ;
  assign y7680 = ~n24282 ;
  assign y7681 = n24283 ;
  assign y7682 = ~n24292 ;
  assign y7683 = n24293 ;
  assign y7684 = ~n24295 ;
  assign y7685 = ~1'b0 ;
  assign y7686 = n24297 ;
  assign y7687 = n24301 ;
  assign y7688 = ~1'b0 ;
  assign y7689 = ~n24304 ;
  assign y7690 = n24308 ;
  assign y7691 = ~n24315 ;
  assign y7692 = n24316 ;
  assign y7693 = n24317 ;
  assign y7694 = n24319 ;
  assign y7695 = n24320 ;
  assign y7696 = n24321 ;
  assign y7697 = n24322 ;
  assign y7698 = n24323 ;
  assign y7699 = n24329 ;
  assign y7700 = ~1'b0 ;
  assign y7701 = ~1'b0 ;
  assign y7702 = ~n24332 ;
  assign y7703 = ~n24333 ;
  assign y7704 = n24340 ;
  assign y7705 = n24341 ;
  assign y7706 = n24349 ;
  assign y7707 = n24351 ;
  assign y7708 = n24364 ;
  assign y7709 = n24365 ;
  assign y7710 = ~n24367 ;
  assign y7711 = n24373 ;
  assign y7712 = ~n24375 ;
  assign y7713 = ~1'b0 ;
  assign y7714 = n24382 ;
  assign y7715 = n24384 ;
  assign y7716 = n24385 ;
  assign y7717 = ~n24393 ;
  assign y7718 = n24394 ;
  assign y7719 = n24403 ;
  assign y7720 = n24404 ;
  assign y7721 = n24406 ;
  assign y7722 = ~1'b0 ;
  assign y7723 = ~n24407 ;
  assign y7724 = ~n24408 ;
  assign y7725 = ~n10131 ;
  assign y7726 = n24409 ;
  assign y7727 = n14208 ;
  assign y7728 = n24412 ;
  assign y7729 = ~n24413 ;
  assign y7730 = n24415 ;
  assign y7731 = ~n24419 ;
  assign y7732 = n24424 ;
  assign y7733 = n24428 ;
  assign y7734 = n24429 ;
  assign y7735 = ~n24437 ;
  assign y7736 = ~n24438 ;
  assign y7737 = n24440 ;
  assign y7738 = ~n24441 ;
  assign y7739 = ~1'b0 ;
  assign y7740 = n24442 ;
  assign y7741 = ~n24444 ;
  assign y7742 = ~n24449 ;
  assign y7743 = ~n24452 ;
  assign y7744 = n24453 ;
  assign y7745 = n24455 ;
  assign y7746 = ~n24459 ;
  assign y7747 = n24461 ;
  assign y7748 = n24465 ;
  assign y7749 = n4770 ;
  assign y7750 = ~n24467 ;
  assign y7751 = n24474 ;
  assign y7752 = n24476 ;
  assign y7753 = ~1'b0 ;
  assign y7754 = ~1'b0 ;
  assign y7755 = n24478 ;
  assign y7756 = n24480 ;
  assign y7757 = n24484 ;
  assign y7758 = ~1'b0 ;
  assign y7759 = ~n24492 ;
  assign y7760 = ~n24494 ;
  assign y7761 = n24495 ;
  assign y7762 = ~n24496 ;
  assign y7763 = ~n24503 ;
  assign y7764 = n24510 ;
  assign y7765 = ~1'b0 ;
  assign y7766 = n24512 ;
  assign y7767 = n24515 ;
  assign y7768 = n24517 ;
  assign y7769 = n24521 ;
  assign y7770 = n24522 ;
  assign y7771 = ~1'b0 ;
  assign y7772 = ~n24523 ;
  assign y7773 = ~n24531 ;
  assign y7774 = n24534 ;
  assign y7775 = ~1'b0 ;
  assign y7776 = n24536 ;
  assign y7777 = ~n24539 ;
  assign y7778 = n24544 ;
  assign y7779 = ~n24545 ;
  assign y7780 = n24548 ;
  assign y7781 = ~1'b0 ;
  assign y7782 = ~n24552 ;
  assign y7783 = ~n24554 ;
  assign y7784 = ~n24556 ;
  assign y7785 = n24561 ;
  assign y7786 = ~n24564 ;
  assign y7787 = ~1'b0 ;
  assign y7788 = n10502 ;
  assign y7789 = ~n24568 ;
  assign y7790 = n24571 ;
  assign y7791 = ~n24573 ;
  assign y7792 = ~n24574 ;
  assign y7793 = n24577 ;
  assign y7794 = n24588 ;
  assign y7795 = n24591 ;
  assign y7796 = n24594 ;
  assign y7797 = n24598 ;
  assign y7798 = n24601 ;
  assign y7799 = n24604 ;
  assign y7800 = ~1'b0 ;
  assign y7801 = ~1'b0 ;
  assign y7802 = ~1'b0 ;
  assign y7803 = ~1'b0 ;
  assign y7804 = n24608 ;
  assign y7805 = ~1'b0 ;
  assign y7806 = ~n24615 ;
  assign y7807 = n24616 ;
  assign y7808 = 1'b0 ;
  assign y7809 = ~n24617 ;
  assign y7810 = n24620 ;
  assign y7811 = ~n24622 ;
  assign y7812 = ~n24623 ;
  assign y7813 = ~1'b0 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = n24625 ;
  assign y7816 = ~n24632 ;
  assign y7817 = n24637 ;
  assign y7818 = n24641 ;
  assign y7819 = n24645 ;
  assign y7820 = ~n24647 ;
  assign y7821 = ~1'b0 ;
  assign y7822 = ~1'b0 ;
  assign y7823 = ~n24650 ;
  assign y7824 = n24653 ;
  assign y7825 = n24655 ;
  assign y7826 = ~n24660 ;
  assign y7827 = n24665 ;
  assign y7828 = n24667 ;
  assign y7829 = ~1'b0 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = n24669 ;
  assign y7832 = ~1'b0 ;
  assign y7833 = ~1'b0 ;
  assign y7834 = ~n24670 ;
  assign y7835 = n24674 ;
  assign y7836 = n24675 ;
  assign y7837 = n24677 ;
  assign y7838 = n24678 ;
  assign y7839 = ~1'b0 ;
  assign y7840 = ~n24680 ;
  assign y7841 = ~n14910 ;
  assign y7842 = ~n24682 ;
  assign y7843 = ~n24687 ;
  assign y7844 = ~n24689 ;
  assign y7845 = ~1'b0 ;
  assign y7846 = ~n24692 ;
  assign y7847 = n24697 ;
  assign y7848 = ~n24699 ;
  assign y7849 = n24703 ;
  assign y7850 = n24709 ;
  assign y7851 = n24710 ;
  assign y7852 = ~n24712 ;
  assign y7853 = ~n24719 ;
  assign y7854 = ~n24721 ;
  assign y7855 = n24722 ;
  assign y7856 = n24726 ;
  assign y7857 = ~n24731 ;
  assign y7858 = ~n24733 ;
  assign y7859 = n24735 ;
  assign y7860 = n24744 ;
  assign y7861 = ~1'b0 ;
  assign y7862 = ~n24754 ;
  assign y7863 = ~n24755 ;
  assign y7864 = ~n24761 ;
  assign y7865 = n24764 ;
  assign y7866 = n24766 ;
  assign y7867 = ~1'b0 ;
  assign y7868 = n24770 ;
  assign y7869 = ~n24772 ;
  assign y7870 = n24774 ;
  assign y7871 = ~n24777 ;
  assign y7872 = n24779 ;
  assign y7873 = n24791 ;
  assign y7874 = ~1'b0 ;
  assign y7875 = ~1'b0 ;
  assign y7876 = n24794 ;
  assign y7877 = n24796 ;
  assign y7878 = n24798 ;
  assign y7879 = ~1'b0 ;
  assign y7880 = ~n24800 ;
  assign y7881 = n24803 ;
  assign y7882 = n24806 ;
  assign y7883 = ~n24810 ;
  assign y7884 = n24811 ;
  assign y7885 = ~n24813 ;
  assign y7886 = ~n24821 ;
  assign y7887 = ~n24824 ;
  assign y7888 = n24829 ;
  assign y7889 = ~n24830 ;
  assign y7890 = ~n24831 ;
  assign y7891 = ~n24835 ;
  assign y7892 = ~n24840 ;
  assign y7893 = ~n24847 ;
  assign y7894 = n24849 ;
  assign y7895 = n24855 ;
  assign y7896 = ~n24860 ;
  assign y7897 = ~n24862 ;
  assign y7898 = ~n24863 ;
  assign y7899 = ~n24867 ;
  assign y7900 = n24870 ;
  assign y7901 = ~n24871 ;
  assign y7902 = n24872 ;
  assign y7903 = ~n24874 ;
  assign y7904 = ~1'b0 ;
  assign y7905 = n24882 ;
  assign y7906 = ~n24885 ;
  assign y7907 = n24891 ;
  assign y7908 = n24899 ;
  assign y7909 = ~1'b0 ;
  assign y7910 = ~1'b0 ;
  assign y7911 = n24901 ;
  assign y7912 = ~n24902 ;
  assign y7913 = n24911 ;
  assign y7914 = ~n24914 ;
  assign y7915 = n24918 ;
  assign y7916 = ~n20937 ;
  assign y7917 = ~1'b0 ;
  assign y7918 = ~n24925 ;
  assign y7919 = n24926 ;
  assign y7920 = ~1'b0 ;
  assign y7921 = n24933 ;
  assign y7922 = n14905 ;
  assign y7923 = n24935 ;
  assign y7924 = ~1'b0 ;
  assign y7925 = ~n24939 ;
  assign y7926 = ~n24940 ;
  assign y7927 = n24943 ;
  assign y7928 = ~n24945 ;
  assign y7929 = ~n24946 ;
  assign y7930 = ~n24947 ;
  assign y7931 = n24951 ;
  assign y7932 = ~n24954 ;
  assign y7933 = ~n24965 ;
  assign y7934 = ~n24966 ;
  assign y7935 = n24967 ;
  assign y7936 = n24969 ;
  assign y7937 = ~1'b0 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = n24970 ;
  assign y7940 = n24974 ;
  assign y7941 = ~n24976 ;
  assign y7942 = n24981 ;
  assign y7943 = ~n24988 ;
  assign y7944 = ~1'b0 ;
  assign y7945 = n24994 ;
  assign y7946 = ~1'b0 ;
  assign y7947 = n24996 ;
  assign y7948 = ~n25004 ;
  assign y7949 = ~1'b0 ;
  assign y7950 = ~n25008 ;
  assign y7951 = ~1'b0 ;
  assign y7952 = ~n25009 ;
  assign y7953 = n25013 ;
  assign y7954 = n25015 ;
  assign y7955 = ~n25023 ;
  assign y7956 = ~n25028 ;
  assign y7957 = ~n25029 ;
  assign y7958 = n25036 ;
  assign y7959 = n25038 ;
  assign y7960 = ~n25039 ;
  assign y7961 = ~1'b0 ;
  assign y7962 = ~1'b0 ;
  assign y7963 = ~n25041 ;
  assign y7964 = n25046 ;
  assign y7965 = n25047 ;
  assign y7966 = ~1'b0 ;
  assign y7967 = ~n25051 ;
  assign y7968 = n25052 ;
  assign y7969 = ~n25053 ;
  assign y7970 = ~n25054 ;
  assign y7971 = ~n25055 ;
  assign y7972 = ~1'b0 ;
  assign y7973 = ~n25056 ;
  assign y7974 = ~n25062 ;
  assign y7975 = n25066 ;
  assign y7976 = n25067 ;
  assign y7977 = ~n25077 ;
  assign y7978 = ~n25081 ;
  assign y7979 = ~n25082 ;
  assign y7980 = ~n25085 ;
  assign y7981 = n25086 ;
  assign y7982 = ~1'b0 ;
  assign y7983 = n25087 ;
  assign y7984 = n25088 ;
  assign y7985 = n25093 ;
  assign y7986 = ~n25095 ;
  assign y7987 = 1'b0 ;
  assign y7988 = ~n25099 ;
  assign y7989 = ~n25100 ;
  assign y7990 = n25106 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = ~n25107 ;
  assign y7993 = n25110 ;
  assign y7994 = n25117 ;
  assign y7995 = n25118 ;
  assign y7996 = ~n25119 ;
  assign y7997 = ~n25123 ;
  assign y7998 = ~n25124 ;
  assign y7999 = ~n25126 ;
  assign y8000 = n25132 ;
  assign y8001 = ~n25141 ;
  assign y8002 = n25149 ;
  assign y8003 = ~n25152 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = n25153 ;
  assign y8006 = n25164 ;
  assign y8007 = ~n25168 ;
  assign y8008 = n25182 ;
  assign y8009 = n25186 ;
  assign y8010 = n25187 ;
  assign y8011 = n25189 ;
  assign y8012 = ~n25191 ;
  assign y8013 = ~n25193 ;
  assign y8014 = n25194 ;
  assign y8015 = ~n25196 ;
  assign y8016 = ~1'b0 ;
  assign y8017 = ~1'b0 ;
  assign y8018 = ~1'b0 ;
  assign y8019 = n25197 ;
  assign y8020 = ~n25198 ;
  assign y8021 = n25206 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = ~n25210 ;
  assign y8024 = ~n25212 ;
  assign y8025 = n25213 ;
  assign y8026 = n25216 ;
  assign y8027 = n25217 ;
  assign y8028 = ~n25219 ;
  assign y8029 = ~n25220 ;
  assign y8030 = ~n25221 ;
  assign y8031 = n25223 ;
  assign y8032 = ~n25224 ;
  assign y8033 = n25231 ;
  assign y8034 = ~1'b0 ;
  assign y8035 = ~n25232 ;
  assign y8036 = ~n25237 ;
  assign y8037 = ~n25240 ;
  assign y8038 = n25241 ;
  assign y8039 = n25244 ;
  assign y8040 = ~n25246 ;
  assign y8041 = ~n25248 ;
  assign y8042 = ~n25254 ;
  assign y8043 = n25255 ;
  assign y8044 = n25260 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = ~n25263 ;
  assign y8047 = n25272 ;
  assign y8048 = ~1'b0 ;
  assign y8049 = ~n25279 ;
  assign y8050 = n25280 ;
  assign y8051 = ~n25282 ;
  assign y8052 = ~n25286 ;
  assign y8053 = ~1'b0 ;
  assign y8054 = ~n25288 ;
  assign y8055 = ~n25289 ;
  assign y8056 = ~1'b0 ;
  assign y8057 = ~n25291 ;
  assign y8058 = ~n25292 ;
  assign y8059 = ~n25297 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = ~1'b0 ;
  assign y8062 = ~1'b0 ;
  assign y8063 = ~n25298 ;
  assign y8064 = ~n25303 ;
  assign y8065 = n25306 ;
  assign y8066 = ~1'b0 ;
  assign y8067 = ~n25309 ;
  assign y8068 = ~n25311 ;
  assign y8069 = ~n25312 ;
  assign y8070 = ~n25319 ;
  assign y8071 = ~n25322 ;
  assign y8072 = n25326 ;
  assign y8073 = n25330 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = 1'b0 ;
  assign y8076 = 1'b0 ;
  assign y8077 = n25332 ;
  assign y8078 = ~n25334 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = n25336 ;
  assign y8081 = n25341 ;
  assign y8082 = ~1'b0 ;
  assign y8083 = n25344 ;
  assign y8084 = n25345 ;
  assign y8085 = n25348 ;
  assign y8086 = ~n25351 ;
  assign y8087 = ~n25354 ;
  assign y8088 = n25356 ;
  assign y8089 = n25360 ;
  assign y8090 = n25362 ;
  assign y8091 = ~n25365 ;
  assign y8092 = ~n25377 ;
  assign y8093 = n25379 ;
  assign y8094 = ~n25380 ;
  assign y8095 = ~n25387 ;
  assign y8096 = n25389 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~n25391 ;
  assign y8099 = n25394 ;
  assign y8100 = n25396 ;
  assign y8101 = n25403 ;
  assign y8102 = n25406 ;
  assign y8103 = ~n25411 ;
  assign y8104 = n25412 ;
  assign y8105 = n18262 ;
  assign y8106 = ~n9978 ;
  assign y8107 = ~n25415 ;
  assign y8108 = ~1'b0 ;
  assign y8109 = ~1'b0 ;
  assign y8110 = n25420 ;
  assign y8111 = n25423 ;
  assign y8112 = ~n25424 ;
  assign y8113 = ~1'b0 ;
  assign y8114 = ~n25425 ;
  assign y8115 = ~n25426 ;
  assign y8116 = ~n25427 ;
  assign y8117 = ~1'b0 ;
  assign y8118 = ~n25428 ;
  assign y8119 = ~1'b0 ;
  assign y8120 = n25436 ;
  assign y8121 = ~n25438 ;
  assign y8122 = n25439 ;
  assign y8123 = ~1'b0 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = ~n25441 ;
  assign y8126 = ~n25446 ;
  assign y8127 = ~1'b0 ;
  assign y8128 = n25449 ;
  assign y8129 = n25451 ;
  assign y8130 = ~n25457 ;
  assign y8131 = ~n25463 ;
  assign y8132 = ~n4704 ;
  assign y8133 = n25467 ;
  assign y8134 = n25477 ;
  assign y8135 = n25478 ;
  assign y8136 = ~n25481 ;
  assign y8137 = n25484 ;
  assign y8138 = n25494 ;
  assign y8139 = ~1'b0 ;
  assign y8140 = n25495 ;
  assign y8141 = ~1'b0 ;
  assign y8142 = ~1'b0 ;
  assign y8143 = ~n25496 ;
  assign y8144 = ~n25499 ;
  assign y8145 = n25507 ;
  assign y8146 = ~n25511 ;
  assign y8147 = ~n25529 ;
  assign y8148 = 1'b0 ;
  assign y8149 = n25539 ;
  assign y8150 = n25540 ;
  assign y8151 = ~n25548 ;
  assign y8152 = n25554 ;
  assign y8153 = n25558 ;
  assign y8154 = n25560 ;
  assign y8155 = ~n25565 ;
  assign y8156 = ~n25568 ;
  assign y8157 = n25571 ;
  assign y8158 = n25572 ;
  assign y8159 = ~n25575 ;
  assign y8160 = ~n25581 ;
  assign y8161 = ~n25583 ;
  assign y8162 = ~n25591 ;
  assign y8163 = ~n25594 ;
  assign y8164 = ~n25596 ;
  assign y8165 = n25598 ;
  assign y8166 = ~n25601 ;
  assign y8167 = ~n25603 ;
  assign y8168 = ~n25605 ;
  assign y8169 = n25608 ;
  assign y8170 = ~n25610 ;
  assign y8171 = n25612 ;
  assign y8172 = n25615 ;
  assign y8173 = ~n25621 ;
  assign y8174 = ~n25622 ;
  assign y8175 = n25623 ;
  assign y8176 = ~n25625 ;
  assign y8177 = ~1'b0 ;
  assign y8178 = ~1'b0 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = ~1'b0 ;
  assign y8181 = ~n25629 ;
  assign y8182 = ~n25631 ;
  assign y8183 = n25636 ;
  assign y8184 = ~n25641 ;
  assign y8185 = ~n25644 ;
  assign y8186 = n25646 ;
  assign y8187 = ~n25650 ;
  assign y8188 = ~n25653 ;
  assign y8189 = ~1'b0 ;
  assign y8190 = ~1'b0 ;
  assign y8191 = ~n25655 ;
  assign y8192 = n25656 ;
  assign y8193 = n25657 ;
  assign y8194 = n25659 ;
  assign y8195 = ~n25665 ;
  assign y8196 = n25671 ;
  assign y8197 = n25678 ;
  assign y8198 = ~n25681 ;
  assign y8199 = n25693 ;
  assign y8200 = ~1'b0 ;
  assign y8201 = ~1'b0 ;
  assign y8202 = ~n25697 ;
  assign y8203 = ~n25698 ;
  assign y8204 = ~n25703 ;
  assign y8205 = n25706 ;
  assign y8206 = ~n25711 ;
  assign y8207 = ~n25719 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = n25720 ;
  assign y8210 = n25721 ;
  assign y8211 = ~n25731 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~n25732 ;
  assign y8214 = ~1'b0 ;
  assign y8215 = n25734 ;
  assign y8216 = ~n25735 ;
  assign y8217 = n25739 ;
  assign y8218 = ~n25742 ;
  assign y8219 = n25749 ;
  assign y8220 = ~n25754 ;
  assign y8221 = n25756 ;
  assign y8222 = ~n25757 ;
  assign y8223 = n25760 ;
  assign y8224 = n25761 ;
  assign y8225 = ~n25768 ;
  assign y8226 = ~n25776 ;
  assign y8227 = ~n25779 ;
  assign y8228 = ~n25782 ;
  assign y8229 = 1'b0 ;
  assign y8230 = ~1'b0 ;
  assign y8231 = ~n25785 ;
  assign y8232 = n25790 ;
  assign y8233 = ~n25792 ;
  assign y8234 = n25795 ;
  assign y8235 = ~n25796 ;
  assign y8236 = ~1'b0 ;
  assign y8237 = ~n25798 ;
  assign y8238 = n25799 ;
  assign y8239 = ~n25802 ;
  assign y8240 = ~n25803 ;
  assign y8241 = n25809 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = ~n25812 ;
  assign y8244 = ~n25813 ;
  assign y8245 = n25818 ;
  assign y8246 = ~n25819 ;
  assign y8247 = ~n25820 ;
  assign y8248 = ~n25824 ;
  assign y8249 = ~n25826 ;
  assign y8250 = ~n25832 ;
  assign y8251 = n25837 ;
  assign y8252 = ~n25842 ;
  assign y8253 = n25849 ;
  assign y8254 = ~n25850 ;
  assign y8255 = ~n25851 ;
  assign y8256 = ~1'b0 ;
  assign y8257 = ~1'b0 ;
  assign y8258 = ~n25855 ;
  assign y8259 = n25866 ;
  assign y8260 = ~n25868 ;
  assign y8261 = n25870 ;
  assign y8262 = ~n25875 ;
  assign y8263 = ~1'b0 ;
  assign y8264 = n25880 ;
  assign y8265 = n25887 ;
  assign y8266 = ~n25897 ;
  assign y8267 = ~n25905 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = ~n25912 ;
  assign y8270 = ~n25919 ;
  assign y8271 = ~n25923 ;
  assign y8272 = n12397 ;
  assign y8273 = ~n25924 ;
  assign y8274 = n25926 ;
  assign y8275 = ~n25932 ;
  assign y8276 = ~n25933 ;
  assign y8277 = ~1'b0 ;
  assign y8278 = ~n25935 ;
  assign y8279 = ~n25936 ;
  assign y8280 = n7352 ;
  assign y8281 = ~n25937 ;
  assign y8282 = ~1'b0 ;
  assign y8283 = n25940 ;
  assign y8284 = ~n25943 ;
  assign y8285 = n25948 ;
  assign y8286 = ~n25953 ;
  assign y8287 = ~1'b0 ;
  assign y8288 = ~n25959 ;
  assign y8289 = ~1'b0 ;
  assign y8290 = ~1'b0 ;
  assign y8291 = ~n25960 ;
  assign y8292 = n25963 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = ~1'b0 ;
  assign y8295 = ~1'b0 ;
  assign y8296 = n25965 ;
  assign y8297 = ~n25969 ;
  assign y8298 = n25970 ;
  assign y8299 = n25972 ;
  assign y8300 = ~n25974 ;
  assign y8301 = n25975 ;
  assign y8302 = ~1'b0 ;
  assign y8303 = n25976 ;
  assign y8304 = ~n10398 ;
  assign y8305 = ~n25978 ;
  assign y8306 = ~n25979 ;
  assign y8307 = ~1'b0 ;
  assign y8308 = ~n25983 ;
  assign y8309 = ~n25990 ;
  assign y8310 = n25991 ;
  assign y8311 = n25993 ;
  assign y8312 = ~1'b0 ;
  assign y8313 = ~1'b0 ;
  assign y8314 = n25998 ;
  assign y8315 = n26001 ;
  assign y8316 = n26004 ;
  assign y8317 = n26005 ;
  assign y8318 = ~n26011 ;
  assign y8319 = ~n26015 ;
  assign y8320 = n26016 ;
  assign y8321 = ~n26023 ;
  assign y8322 = n26028 ;
  assign y8323 = ~n26029 ;
  assign y8324 = n26031 ;
  assign y8325 = n26035 ;
  assign y8326 = n26039 ;
  assign y8327 = ~n26045 ;
  assign y8328 = ~1'b0 ;
  assign y8329 = n26050 ;
  assign y8330 = ~n26054 ;
  assign y8331 = ~n26059 ;
  assign y8332 = ~1'b0 ;
  assign y8333 = n26064 ;
  assign y8334 = ~n26065 ;
  assign y8335 = n26068 ;
  assign y8336 = ~n26071 ;
  assign y8337 = n26072 ;
  assign y8338 = n26073 ;
  assign y8339 = ~1'b0 ;
  assign y8340 = ~n26081 ;
  assign y8341 = n26082 ;
  assign y8342 = n26084 ;
  assign y8343 = ~n26086 ;
  assign y8344 = n26087 ;
  assign y8345 = ~n26091 ;
  assign y8346 = ~1'b0 ;
  assign y8347 = ~1'b0 ;
  assign y8348 = ~n26092 ;
  assign y8349 = ~n26093 ;
  assign y8350 = n26099 ;
  assign y8351 = ~n26100 ;
  assign y8352 = n26102 ;
  assign y8353 = ~n26106 ;
  assign y8354 = ~1'b0 ;
  assign y8355 = ~1'b0 ;
  assign y8356 = ~n22819 ;
  assign y8357 = ~1'b0 ;
  assign y8358 = ~1'b0 ;
  assign y8359 = n26109 ;
  assign y8360 = ~n13327 ;
  assign y8361 = n26113 ;
  assign y8362 = ~n26118 ;
  assign y8363 = ~n26126 ;
  assign y8364 = n26128 ;
  assign y8365 = ~n26129 ;
  assign y8366 = ~n26131 ;
  assign y8367 = ~n26135 ;
  assign y8368 = ~n26139 ;
  assign y8369 = ~n26141 ;
  assign y8370 = n26149 ;
  assign y8371 = ~n26156 ;
  assign y8372 = n26158 ;
  assign y8373 = ~n26160 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~1'b0 ;
  assign y8376 = ~n26163 ;
  assign y8377 = ~n26166 ;
  assign y8378 = ~n9782 ;
  assign y8379 = ~n26169 ;
  assign y8380 = ~1'b0 ;
  assign y8381 = n26177 ;
  assign y8382 = ~n26179 ;
  assign y8383 = ~n26180 ;
  assign y8384 = ~n26181 ;
  assign y8385 = n26184 ;
  assign y8386 = ~1'b0 ;
  assign y8387 = n26187 ;
  assign y8388 = ~n26189 ;
  assign y8389 = n6087 ;
  assign y8390 = ~1'b0 ;
  assign y8391 = ~1'b0 ;
  assign y8392 = ~n26191 ;
  assign y8393 = n26195 ;
  assign y8394 = ~1'b0 ;
  assign y8395 = ~n26204 ;
  assign y8396 = n26205 ;
  assign y8397 = n26206 ;
  assign y8398 = ~n26210 ;
  assign y8399 = ~n26214 ;
  assign y8400 = ~n26217 ;
  assign y8401 = ~n26218 ;
  assign y8402 = n26221 ;
  assign y8403 = ~n26223 ;
  assign y8404 = n26228 ;
  assign y8405 = ~1'b0 ;
  assign y8406 = ~n26236 ;
  assign y8407 = n26237 ;
  assign y8408 = n26239 ;
  assign y8409 = n26240 ;
  assign y8410 = ~n26242 ;
  assign y8411 = ~n26243 ;
  assign y8412 = n26248 ;
  assign y8413 = ~n26252 ;
  assign y8414 = n22246 ;
  assign y8415 = n26253 ;
  assign y8416 = ~n20522 ;
  assign y8417 = n26255 ;
  assign y8418 = ~1'b0 ;
  assign y8419 = ~n26259 ;
  assign y8420 = n26260 ;
  assign y8421 = n26263 ;
  assign y8422 = ~n26265 ;
  assign y8423 = ~n26274 ;
  assign y8424 = ~n26275 ;
  assign y8425 = ~1'b0 ;
  assign y8426 = ~1'b0 ;
  assign y8427 = ~n26280 ;
  assign y8428 = ~n26281 ;
  assign y8429 = n26284 ;
  assign y8430 = n26286 ;
  assign y8431 = ~n26297 ;
  assign y8432 = n26299 ;
  assign y8433 = n26300 ;
  assign y8434 = n26308 ;
  assign y8435 = ~n26309 ;
  assign y8436 = ~n26310 ;
  assign y8437 = ~n26316 ;
  assign y8438 = n26317 ;
  assign y8439 = n26320 ;
  assign y8440 = ~n26321 ;
  assign y8441 = n26325 ;
  assign y8442 = ~n26327 ;
  assign y8443 = ~n26330 ;
  assign y8444 = n26333 ;
  assign y8445 = n26339 ;
  assign y8446 = n26340 ;
  assign y8447 = n26345 ;
  assign y8448 = n26347 ;
  assign y8449 = n26350 ;
  assign y8450 = ~n26355 ;
  assign y8451 = n26359 ;
  assign y8452 = n26360 ;
  assign y8453 = ~1'b0 ;
  assign y8454 = n26361 ;
  assign y8455 = n26364 ;
  assign y8456 = n26367 ;
  assign y8457 = ~n26368 ;
  assign y8458 = n26374 ;
  assign y8459 = ~n26383 ;
  assign y8460 = ~n26384 ;
  assign y8461 = n26386 ;
  assign y8462 = n26390 ;
  assign y8463 = n26391 ;
  assign y8464 = n26395 ;
  assign y8465 = ~n26398 ;
  assign y8466 = ~1'b0 ;
  assign y8467 = ~n26400 ;
  assign y8468 = ~n26401 ;
  assign y8469 = n26403 ;
  assign y8470 = ~n26410 ;
  assign y8471 = ~n26416 ;
  assign y8472 = ~n26418 ;
  assign y8473 = ~1'b0 ;
  assign y8474 = n26419 ;
  assign y8475 = n26420 ;
  assign y8476 = n26425 ;
  assign y8477 = ~1'b0 ;
  assign y8478 = ~n26426 ;
  assign y8479 = ~n26427 ;
  assign y8480 = ~1'b0 ;
  assign y8481 = n26428 ;
  assign y8482 = n26431 ;
  assign y8483 = n26437 ;
  assign y8484 = n26440 ;
  assign y8485 = n26442 ;
  assign y8486 = ~n26446 ;
  assign y8487 = n26449 ;
  assign y8488 = n26450 ;
  assign y8489 = ~n26451 ;
  assign y8490 = ~1'b0 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = ~1'b0 ;
  assign y8493 = n26453 ;
  assign y8494 = ~1'b0 ;
  assign y8495 = ~n26462 ;
  assign y8496 = ~n26465 ;
  assign y8497 = ~n26468 ;
  assign y8498 = ~n26473 ;
  assign y8499 = ~n26477 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = n26480 ;
  assign y8502 = n26481 ;
  assign y8503 = ~n26486 ;
  assign y8504 = ~n26490 ;
  assign y8505 = ~n26494 ;
  assign y8506 = ~n26496 ;
  assign y8507 = n26499 ;
  assign y8508 = ~n26502 ;
  assign y8509 = ~n26506 ;
  assign y8510 = ~1'b0 ;
  assign y8511 = n26508 ;
  assign y8512 = n26513 ;
  assign y8513 = ~n15494 ;
  assign y8514 = ~1'b0 ;
  assign y8515 = ~n26517 ;
  assign y8516 = ~n26520 ;
  assign y8517 = n26533 ;
  assign y8518 = ~1'b0 ;
  assign y8519 = n26538 ;
  assign y8520 = ~n26539 ;
  assign y8521 = n26541 ;
  assign y8522 = ~n26544 ;
  assign y8523 = ~n26546 ;
  assign y8524 = n26547 ;
  assign y8525 = n26550 ;
  assign y8526 = n26553 ;
  assign y8527 = n26554 ;
  assign y8528 = n15071 ;
  assign y8529 = n26570 ;
  assign y8530 = n26574 ;
  assign y8531 = n26576 ;
  assign y8532 = ~n26578 ;
  assign y8533 = ~1'b0 ;
  assign y8534 = ~n26579 ;
  assign y8535 = n26582 ;
  assign y8536 = n26583 ;
  assign y8537 = ~n26585 ;
  assign y8538 = ~1'b0 ;
  assign y8539 = ~n26589 ;
  assign y8540 = ~n26595 ;
  assign y8541 = n26596 ;
  assign y8542 = n26597 ;
  assign y8543 = ~n26599 ;
  assign y8544 = ~n26605 ;
  assign y8545 = ~1'b0 ;
  assign y8546 = ~n26615 ;
  assign y8547 = ~n26618 ;
  assign y8548 = n26620 ;
  assign y8549 = n26623 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = n26624 ;
  assign y8553 = ~n26627 ;
  assign y8554 = n26628 ;
  assign y8555 = n26629 ;
  assign y8556 = ~n26630 ;
  assign y8557 = ~n26632 ;
  assign y8558 = n26634 ;
  assign y8559 = ~1'b0 ;
  assign y8560 = ~n26638 ;
  assign y8561 = n26642 ;
  assign y8562 = ~1'b0 ;
  assign y8563 = ~n26646 ;
  assign y8564 = ~1'b0 ;
  assign y8565 = n26647 ;
  assign y8566 = ~1'b0 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = ~1'b0 ;
  assign y8570 = ~n26649 ;
  assign y8571 = ~n26652 ;
  assign y8572 = ~n26658 ;
  assign y8573 = ~n6409 ;
  assign y8574 = ~n26660 ;
  assign y8575 = ~n26662 ;
  assign y8576 = ~n26665 ;
  assign y8577 = ~n26667 ;
  assign y8578 = ~n26675 ;
  assign y8579 = ~n26676 ;
  assign y8580 = ~n26682 ;
  assign y8581 = ~1'b0 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n26683 ;
  assign y8584 = ~n26684 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~n26685 ;
  assign y8587 = ~1'b0 ;
  assign y8588 = n26691 ;
  assign y8589 = ~n26698 ;
  assign y8590 = ~n26700 ;
  assign y8591 = n26702 ;
  assign y8592 = n26709 ;
  assign y8593 = ~n26713 ;
  assign y8594 = n26714 ;
  assign y8595 = ~1'b0 ;
  assign y8596 = n26718 ;
  assign y8597 = n26722 ;
  assign y8598 = ~1'b0 ;
  assign y8599 = ~n26730 ;
  assign y8600 = n26738 ;
  assign y8601 = ~n26740 ;
  assign y8602 = ~n26742 ;
  assign y8603 = ~1'b0 ;
  assign y8604 = ~n26744 ;
  assign y8605 = ~n26745 ;
  assign y8606 = n26748 ;
  assign y8607 = ~n26750 ;
  assign y8608 = n26756 ;
  assign y8609 = ~n26758 ;
  assign y8610 = n26761 ;
  assign y8611 = ~1'b0 ;
  assign y8612 = ~n26770 ;
  assign y8613 = ~n26771 ;
  assign y8614 = ~n26773 ;
  assign y8615 = ~1'b0 ;
  assign y8616 = n26777 ;
  assign y8617 = n26779 ;
  assign y8618 = n26780 ;
  assign y8619 = n26783 ;
  assign y8620 = ~n26785 ;
  assign y8621 = ~n26788 ;
  assign y8622 = n26791 ;
  assign y8623 = n26798 ;
  assign y8624 = n26801 ;
  assign y8625 = ~n26804 ;
  assign y8626 = n26806 ;
  assign y8627 = ~n26808 ;
  assign y8628 = ~n26819 ;
  assign y8629 = ~1'b0 ;
  assign y8630 = ~n26822 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = n26836 ;
  assign y8633 = ~n26838 ;
  assign y8634 = n26841 ;
  assign y8635 = ~1'b0 ;
  assign y8636 = ~n26842 ;
  assign y8637 = ~n26845 ;
  assign y8638 = ~n26858 ;
  assign y8639 = n26862 ;
  assign y8640 = ~n26863 ;
  assign y8641 = n21914 ;
  assign y8642 = n26869 ;
  assign y8643 = n26870 ;
  assign y8644 = n19922 ;
  assign y8645 = ~n26872 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = n26874 ;
  assign y8648 = ~n26878 ;
  assign y8649 = n26879 ;
  assign y8650 = n26881 ;
  assign y8651 = n26882 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = ~n26892 ;
  assign y8654 = n26899 ;
  assign y8655 = ~n26901 ;
  assign y8656 = ~n26902 ;
  assign y8657 = n26910 ;
  assign y8658 = n26914 ;
  assign y8659 = n26921 ;
  assign y8660 = ~n26922 ;
  assign y8661 = ~n26925 ;
  assign y8662 = n26930 ;
  assign y8663 = n26933 ;
  assign y8664 = ~1'b0 ;
  assign y8665 = ~n26935 ;
  assign y8666 = n6306 ;
  assign y8667 = n26936 ;
  assign y8668 = ~1'b0 ;
  assign y8669 = n26938 ;
  assign y8670 = n26942 ;
  assign y8671 = n26945 ;
  assign y8672 = ~1'b0 ;
  assign y8673 = ~n26947 ;
  assign y8674 = ~1'b0 ;
  assign y8675 = ~n26949 ;
  assign y8676 = ~n26953 ;
  assign y8677 = n26957 ;
  assign y8678 = ~n26962 ;
  assign y8679 = ~1'b0 ;
  assign y8680 = ~n26963 ;
  assign y8681 = n7522 ;
  assign y8682 = n26965 ;
  assign y8683 = n26966 ;
  assign y8684 = n26967 ;
  assign y8685 = n26969 ;
  assign y8686 = ~n26970 ;
  assign y8687 = ~n26977 ;
  assign y8688 = ~n26979 ;
  assign y8689 = ~n26982 ;
  assign y8690 = ~n26988 ;
  assign y8691 = ~n26989 ;
  assign y8692 = n26991 ;
  assign y8693 = ~n26994 ;
  assign y8694 = n26997 ;
  assign y8695 = ~n27002 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = n27004 ;
  assign y8698 = n27006 ;
  assign y8699 = ~n27010 ;
  assign y8700 = ~n27014 ;
  assign y8701 = ~n27018 ;
  assign y8702 = ~n27025 ;
  assign y8703 = ~1'b0 ;
  assign y8704 = n27029 ;
  assign y8705 = n27031 ;
  assign y8706 = n27032 ;
  assign y8707 = n27034 ;
  assign y8708 = ~n27036 ;
  assign y8709 = n27039 ;
  assign y8710 = ~n27041 ;
  assign y8711 = n27047 ;
  assign y8712 = ~1'b0 ;
  assign y8713 = ~1'b0 ;
  assign y8714 = n27048 ;
  assign y8715 = n27053 ;
  assign y8716 = n27055 ;
  assign y8717 = n27061 ;
  assign y8718 = n27078 ;
  assign y8719 = n27080 ;
  assign y8720 = n27085 ;
  assign y8721 = ~1'b0 ;
  assign y8722 = n27089 ;
  assign y8723 = ~n27091 ;
  assign y8724 = ~n27096 ;
  assign y8725 = n27099 ;
  assign y8726 = n27105 ;
  assign y8727 = ~n27115 ;
  assign y8728 = ~n27117 ;
  assign y8729 = ~n27120 ;
  assign y8730 = n27124 ;
  assign y8731 = n27127 ;
  assign y8732 = ~n27132 ;
  assign y8733 = n27135 ;
  assign y8734 = ~1'b0 ;
  assign y8735 = n27136 ;
  assign y8736 = ~n27139 ;
  assign y8737 = ~n27143 ;
  assign y8738 = ~n27144 ;
  assign y8739 = ~n27147 ;
  assign y8740 = n27150 ;
  assign y8741 = ~1'b0 ;
  assign y8742 = ~1'b0 ;
  assign y8743 = n27154 ;
  assign y8744 = n27155 ;
  assign y8745 = ~1'b0 ;
  assign y8746 = n27156 ;
  assign y8747 = ~n27158 ;
  assign y8748 = n27164 ;
  assign y8749 = n27165 ;
  assign y8750 = ~n27167 ;
  assign y8751 = n27169 ;
  assign y8752 = n27170 ;
  assign y8753 = n27171 ;
  assign y8754 = n27173 ;
  assign y8755 = ~n27177 ;
  assign y8756 = ~n27178 ;
  assign y8757 = n27182 ;
  assign y8758 = n27188 ;
  assign y8759 = ~1'b0 ;
  assign y8760 = ~1'b0 ;
  assign y8761 = ~n27190 ;
  assign y8762 = n27195 ;
  assign y8763 = ~n27196 ;
  assign y8764 = n27198 ;
  assign y8765 = ~n27204 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = ~n27205 ;
  assign y8768 = ~n27208 ;
  assign y8769 = ~n27209 ;
  assign y8770 = ~1'b0 ;
  assign y8771 = ~1'b0 ;
  assign y8772 = ~n27216 ;
  assign y8773 = n6875 ;
  assign y8774 = ~n27217 ;
  assign y8775 = n27218 ;
  assign y8776 = ~1'b0 ;
  assign y8777 = n27220 ;
  assign y8778 = ~n27222 ;
  assign y8779 = n27224 ;
  assign y8780 = n27227 ;
  assign y8781 = n27233 ;
  assign y8782 = ~1'b0 ;
  assign y8783 = ~n27239 ;
  assign y8784 = n27253 ;
  assign y8785 = ~n27257 ;
  assign y8786 = ~n27270 ;
  assign y8787 = ~n27272 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~n27274 ;
  assign y8790 = ~1'b0 ;
  assign y8791 = n27277 ;
  assign y8792 = n27280 ;
  assign y8793 = ~n27283 ;
  assign y8794 = 1'b0 ;
  assign y8795 = ~n27284 ;
  assign y8796 = ~n27285 ;
  assign y8797 = n27286 ;
  assign y8798 = n27295 ;
  assign y8799 = n27297 ;
  assign y8800 = ~1'b0 ;
  assign y8801 = ~1'b0 ;
  assign y8802 = n27300 ;
  assign y8803 = ~n27302 ;
  assign y8804 = n27303 ;
  assign y8805 = ~n27305 ;
  assign y8806 = ~n27308 ;
  assign y8807 = ~n27312 ;
  assign y8808 = ~n27316 ;
  assign y8809 = n27317 ;
  assign y8810 = ~n27318 ;
  assign y8811 = n27321 ;
  assign y8812 = ~n27322 ;
  assign y8813 = ~n27328 ;
  assign y8814 = ~1'b0 ;
  assign y8815 = ~1'b0 ;
  assign y8816 = n27330 ;
  assign y8817 = ~n27331 ;
  assign y8818 = n27333 ;
  assign y8819 = ~1'b0 ;
  assign y8820 = ~1'b0 ;
  assign y8821 = ~1'b0 ;
  assign y8822 = n27337 ;
  assign y8823 = ~n27341 ;
  assign y8824 = ~n27345 ;
  assign y8825 = ~n27346 ;
  assign y8826 = n27351 ;
  assign y8827 = ~n27354 ;
  assign y8828 = ~n27355 ;
  assign y8829 = ~n27359 ;
  assign y8830 = ~n27360 ;
  assign y8831 = n27361 ;
  assign y8832 = ~n27362 ;
  assign y8833 = n27364 ;
  assign y8834 = ~n27367 ;
  assign y8835 = ~n27370 ;
  assign y8836 = n27371 ;
  assign y8837 = n27374 ;
  assign y8838 = ~n27377 ;
  assign y8839 = ~n27384 ;
  assign y8840 = n27387 ;
  assign y8841 = ~1'b0 ;
  assign y8842 = n27394 ;
  assign y8843 = ~n27397 ;
  assign y8844 = ~n27398 ;
  assign y8845 = n27399 ;
  assign y8846 = ~1'b0 ;
  assign y8847 = n27405 ;
  assign y8848 = ~n27407 ;
  assign y8849 = ~n27409 ;
  assign y8850 = n27411 ;
  assign y8851 = ~n27413 ;
  assign y8852 = ~n27422 ;
  assign y8853 = ~1'b0 ;
  assign y8854 = ~n27425 ;
  assign y8855 = n27431 ;
  assign y8856 = ~n27435 ;
  assign y8857 = ~n27438 ;
  assign y8858 = ~n27439 ;
  assign y8859 = ~n27442 ;
  assign y8860 = ~n27443 ;
  assign y8861 = n27445 ;
  assign y8862 = ~n27449 ;
  assign y8863 = ~1'b0 ;
  assign y8864 = ~1'b0 ;
  assign y8865 = ~n27450 ;
  assign y8866 = n27451 ;
  assign y8867 = ~n27454 ;
  assign y8868 = n27455 ;
  assign y8869 = ~n27458 ;
  assign y8870 = ~1'b0 ;
  assign y8871 = n27466 ;
  assign y8872 = ~n27475 ;
  assign y8873 = ~n14199 ;
  assign y8874 = ~n27480 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n27483 ;
  assign y8877 = ~n27489 ;
  assign y8878 = ~1'b0 ;
  assign y8879 = ~n27492 ;
  assign y8880 = n27495 ;
  assign y8881 = ~n27498 ;
  assign y8882 = ~n27499 ;
  assign y8883 = n27501 ;
  assign y8884 = n27502 ;
  assign y8885 = ~n27504 ;
  assign y8886 = ~n27505 ;
  assign y8887 = ~n27507 ;
  assign y8888 = ~1'b0 ;
  assign y8889 = ~n27508 ;
  assign y8890 = ~n27512 ;
  assign y8891 = ~n27514 ;
  assign y8892 = n27517 ;
  assign y8893 = ~n27524 ;
  assign y8894 = ~n27526 ;
  assign y8895 = ~n27531 ;
  assign y8896 = ~n27536 ;
  assign y8897 = ~n27541 ;
  assign y8898 = n27545 ;
  assign y8899 = ~1'b0 ;
  assign y8900 = ~n27552 ;
  assign y8901 = ~1'b0 ;
  assign y8902 = n27555 ;
  assign y8903 = n27558 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = n27559 ;
  assign y8906 = ~n27561 ;
  assign y8907 = ~n27565 ;
  assign y8908 = ~n27569 ;
  assign y8909 = ~n27573 ;
  assign y8910 = n27578 ;
  assign y8911 = ~1'b0 ;
  assign y8912 = n27580 ;
  assign y8913 = ~n27583 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = ~n27585 ;
  assign y8916 = ~n27587 ;
  assign y8917 = n27588 ;
  assign y8918 = ~1'b0 ;
  assign y8919 = ~1'b0 ;
  assign y8920 = ~n27591 ;
  assign y8921 = n27592 ;
  assign y8922 = ~n1554 ;
  assign y8923 = ~n27596 ;
  assign y8924 = ~n27598 ;
  assign y8925 = ~n27601 ;
  assign y8926 = ~1'b0 ;
  assign y8927 = n27603 ;
  assign y8928 = ~n27609 ;
  assign y8929 = ~n27611 ;
  assign y8930 = ~n27617 ;
  assign y8931 = ~n27625 ;
  assign y8932 = ~n27626 ;
  assign y8933 = n27633 ;
  assign y8934 = ~1'b0 ;
  assign y8935 = ~n27634 ;
  assign y8936 = ~n27635 ;
  assign y8937 = ~n27637 ;
  assign y8938 = ~1'b0 ;
  assign y8939 = n27638 ;
  assign y8940 = ~n27646 ;
  assign y8941 = n27650 ;
  assign y8942 = ~n27652 ;
  assign y8943 = ~1'b0 ;
  assign y8944 = n27657 ;
  assign y8945 = n27660 ;
  assign y8946 = n27661 ;
  assign y8947 = ~n27666 ;
  assign y8948 = n27668 ;
  assign y8949 = ~n27671 ;
  assign y8950 = ~n27680 ;
  assign y8951 = n27686 ;
  assign y8952 = ~1'b0 ;
  assign y8953 = ~n27689 ;
  assign y8954 = ~1'b0 ;
  assign y8955 = ~n27692 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = ~1'b0 ;
  assign y8959 = ~n27694 ;
  assign y8960 = ~1'b0 ;
  assign y8961 = n27698 ;
  assign y8962 = n27705 ;
  assign y8963 = n1468 ;
  assign y8964 = n27711 ;
  assign y8965 = n27714 ;
  assign y8966 = ~n27719 ;
  assign y8967 = ~n27725 ;
  assign y8968 = n27727 ;
  assign y8969 = n27728 ;
  assign y8970 = n27730 ;
  assign y8971 = ~n27731 ;
  assign y8972 = ~n27733 ;
  assign y8973 = ~n27737 ;
  assign y8974 = ~n27742 ;
  assign y8975 = n27743 ;
  assign y8976 = ~n27749 ;
  assign y8977 = ~n27755 ;
  assign y8978 = n27756 ;
  assign y8979 = n27762 ;
  assign y8980 = n27763 ;
  assign y8981 = ~n27768 ;
  assign y8982 = ~1'b0 ;
  assign y8983 = ~n27769 ;
  assign y8984 = ~1'b0 ;
  assign y8985 = n27770 ;
  assign y8986 = ~n27772 ;
  assign y8987 = n27779 ;
  assign y8988 = ~n27780 ;
  assign y8989 = ~n27782 ;
  assign y8990 = ~n27785 ;
  assign y8991 = n27786 ;
  assign y8992 = ~n27795 ;
  assign y8993 = ~n27797 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = ~n27804 ;
  assign y8996 = n27809 ;
  assign y8997 = ~n20550 ;
  assign y8998 = ~n27811 ;
  assign y8999 = ~n27814 ;
  assign y9000 = ~n27816 ;
  assign y9001 = n27818 ;
  assign y9002 = ~n27822 ;
  assign y9003 = ~n27824 ;
  assign y9004 = n27829 ;
  assign y9005 = ~1'b0 ;
  assign y9006 = n27830 ;
  assign y9007 = ~n27831 ;
  assign y9008 = ~n27834 ;
  assign y9009 = ~n27836 ;
  assign y9010 = ~1'b0 ;
  assign y9011 = ~n27838 ;
  assign y9012 = n27839 ;
  assign y9013 = n27841 ;
  assign y9014 = n27843 ;
  assign y9015 = ~n27845 ;
  assign y9016 = ~n27847 ;
  assign y9017 = n27852 ;
  assign y9018 = ~1'b0 ;
  assign y9019 = ~1'b0 ;
  assign y9020 = ~n27853 ;
  assign y9021 = n27856 ;
  assign y9022 = ~n27859 ;
  assign y9023 = ~n27861 ;
  assign y9024 = n27866 ;
  assign y9025 = n27867 ;
  assign y9026 = n27870 ;
  assign y9027 = ~n27871 ;
  assign y9028 = ~n27873 ;
  assign y9029 = n27887 ;
  assign y9030 = ~1'b0 ;
  assign y9031 = n27890 ;
  assign y9032 = n27892 ;
  assign y9033 = n27896 ;
  assign y9034 = n27897 ;
  assign y9035 = ~1'b0 ;
  assign y9036 = n27898 ;
  assign y9037 = ~n27902 ;
  assign y9038 = ~n27905 ;
  assign y9039 = n27911 ;
  assign y9040 = ~1'b0 ;
  assign y9041 = n27914 ;
  assign y9042 = n27917 ;
  assign y9043 = ~n14991 ;
  assign y9044 = ~1'b0 ;
  assign y9045 = ~n27918 ;
  assign y9046 = ~n27919 ;
  assign y9047 = n27920 ;
  assign y9048 = ~n27923 ;
  assign y9049 = ~1'b0 ;
  assign y9050 = n27925 ;
  assign y9051 = n27926 ;
  assign y9052 = ~n27931 ;
  assign y9053 = n27932 ;
  assign y9054 = ~n27934 ;
  assign y9055 = ~1'b0 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = n27942 ;
  assign y9058 = n27943 ;
  assign y9059 = n27945 ;
  assign y9060 = 1'b0 ;
  assign y9061 = ~n27949 ;
  assign y9062 = ~n27950 ;
  assign y9063 = ~1'b0 ;
  assign y9064 = n27954 ;
  assign y9065 = ~n27956 ;
  assign y9066 = n27957 ;
  assign y9067 = n27958 ;
  assign y9068 = ~n27960 ;
  assign y9069 = ~1'b0 ;
  assign y9070 = n27964 ;
  assign y9071 = ~n27975 ;
  assign y9072 = ~n27976 ;
  assign y9073 = n27977 ;
  assign y9074 = ~n27980 ;
  assign y9075 = ~1'b0 ;
  assign y9076 = n27992 ;
  assign y9077 = ~n27994 ;
  assign y9078 = ~n28000 ;
  assign y9079 = ~1'b0 ;
  assign y9080 = n28001 ;
  assign y9081 = ~n28002 ;
  assign y9082 = n28008 ;
  assign y9083 = n28013 ;
  assign y9084 = ~1'b0 ;
  assign y9085 = ~1'b0 ;
  assign y9086 = n28018 ;
  assign y9087 = ~1'b0 ;
  assign y9088 = ~1'b0 ;
  assign y9089 = ~n28019 ;
  assign y9090 = ~n28020 ;
  assign y9091 = n6341 ;
  assign y9092 = n28021 ;
  assign y9093 = n28031 ;
  assign y9094 = n28032 ;
  assign y9095 = n28033 ;
  assign y9096 = ~n28039 ;
  assign y9097 = ~n28043 ;
  assign y9098 = ~n28045 ;
  assign y9099 = n28046 ;
  assign y9100 = n28049 ;
  assign y9101 = ~n28051 ;
  assign y9102 = n28059 ;
  assign y9103 = ~n28062 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = ~n28064 ;
  assign y9106 = ~n28069 ;
  assign y9107 = n28070 ;
  assign y9108 = n28071 ;
  assign y9109 = ~n28073 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~1'b0 ;
  assign y9112 = n28075 ;
  assign y9113 = ~n28076 ;
  assign y9114 = ~n28077 ;
  assign y9115 = ~n28078 ;
  assign y9116 = n28084 ;
  assign y9117 = n28085 ;
  assign y9118 = n28093 ;
  assign y9119 = n28096 ;
  assign y9120 = ~n28100 ;
  assign y9121 = n28102 ;
  assign y9122 = ~1'b0 ;
  assign y9123 = n28105 ;
  assign y9124 = ~n28112 ;
  assign y9125 = ~n28114 ;
  assign y9126 = ~1'b0 ;
  assign y9127 = ~n28117 ;
  assign y9128 = ~n28120 ;
  assign y9129 = ~1'b0 ;
  assign y9130 = ~n28122 ;
  assign y9131 = ~n28124 ;
  assign y9132 = ~n28125 ;
  assign y9133 = n28130 ;
  assign y9134 = ~n28134 ;
  assign y9135 = ~n28137 ;
  assign y9136 = n28139 ;
  assign y9137 = ~1'b0 ;
  assign y9138 = ~n28141 ;
  assign y9139 = n28145 ;
  assign y9140 = ~n28147 ;
  assign y9141 = ~n28149 ;
  assign y9142 = n28154 ;
  assign y9143 = ~1'b0 ;
  assign y9144 = ~1'b0 ;
  assign y9145 = ~n28157 ;
  assign y9146 = ~n28160 ;
  assign y9147 = n28174 ;
  assign y9148 = n28190 ;
  assign y9149 = n28194 ;
  assign y9150 = ~n28195 ;
  assign y9151 = n28208 ;
  assign y9152 = ~n28211 ;
  assign y9153 = ~n28213 ;
  assign y9154 = ~n28215 ;
  assign y9155 = n28216 ;
  assign y9156 = ~1'b0 ;
  assign y9157 = n28217 ;
  assign y9158 = n28227 ;
  assign y9159 = ~n28232 ;
  assign y9160 = ~1'b0 ;
  assign y9161 = 1'b0 ;
  assign y9162 = n28233 ;
  assign y9163 = n28234 ;
  assign y9164 = ~n28241 ;
  assign y9165 = ~1'b0 ;
  assign y9166 = ~1'b0 ;
  assign y9167 = n28249 ;
  assign y9168 = n28253 ;
  assign y9169 = ~1'b0 ;
  assign y9170 = ~1'b0 ;
  assign y9171 = n28257 ;
  assign y9172 = ~n28259 ;
  assign y9173 = ~1'b0 ;
  assign y9174 = n28264 ;
  assign y9175 = ~1'b0 ;
  assign y9176 = ~1'b0 ;
  assign y9177 = ~n28266 ;
  assign y9178 = n28267 ;
  assign y9179 = n28269 ;
  assign y9180 = ~n28272 ;
  assign y9181 = ~1'b0 ;
  assign y9182 = ~n28276 ;
  assign y9183 = ~n28281 ;
  assign y9184 = n28282 ;
  assign y9185 = ~n28285 ;
  assign y9186 = ~n28288 ;
  assign y9187 = ~n28290 ;
  assign y9188 = ~n28292 ;
  assign y9189 = ~n28293 ;
  assign y9190 = ~n28294 ;
  assign y9191 = n28298 ;
  assign y9192 = ~1'b0 ;
  assign y9193 = ~n28300 ;
  assign y9194 = n28302 ;
  assign y9195 = ~n28308 ;
  assign y9196 = ~1'b0 ;
  assign y9197 = n28309 ;
  assign y9198 = n28312 ;
  assign y9199 = ~n28314 ;
  assign y9200 = n28316 ;
  assign y9201 = 1'b0 ;
  assign y9202 = n28319 ;
  assign y9203 = n28322 ;
  assign y9204 = n28326 ;
  assign y9205 = ~n28328 ;
  assign y9206 = ~n28336 ;
  assign y9207 = n28346 ;
  assign y9208 = n28349 ;
  assign y9209 = n28353 ;
  assign y9210 = ~n28357 ;
  assign y9211 = n28359 ;
  assign y9212 = n28367 ;
  assign y9213 = ~n28369 ;
  assign y9214 = ~n28370 ;
  assign y9215 = ~n28385 ;
  assign y9216 = ~n28389 ;
  assign y9217 = n28390 ;
  assign y9218 = ~n28393 ;
  assign y9219 = ~n28398 ;
  assign y9220 = ~n28399 ;
  assign y9221 = ~n28402 ;
  assign y9222 = n28404 ;
  assign y9223 = ~1'b0 ;
  assign y9224 = ~n28406 ;
  assign y9225 = ~n28409 ;
  assign y9226 = ~1'b0 ;
  assign y9227 = ~n28410 ;
  assign y9228 = ~n28412 ;
  assign y9229 = n28418 ;
  assign y9230 = n28423 ;
  assign y9231 = n28424 ;
  assign y9232 = n28425 ;
  assign y9233 = ~n28426 ;
  assign y9234 = ~n28434 ;
  assign y9235 = n28436 ;
  assign y9236 = ~n28445 ;
  assign y9237 = ~n28449 ;
  assign y9238 = ~n28454 ;
  assign y9239 = n28455 ;
  assign y9240 = n28459 ;
  assign y9241 = ~1'b0 ;
  assign y9242 = n28462 ;
  assign y9243 = n28465 ;
  assign y9244 = ~n28471 ;
  assign y9245 = ~1'b0 ;
  assign y9246 = n28475 ;
  assign y9247 = ~1'b0 ;
  assign y9248 = ~n28477 ;
  assign y9249 = n28480 ;
  assign y9250 = n28483 ;
  assign y9251 = ~1'b0 ;
  assign y9252 = n28484 ;
  assign y9253 = 1'b0 ;
  assign y9254 = ~1'b0 ;
  assign y9255 = ~n28490 ;
  assign y9256 = ~1'b0 ;
  assign y9257 = n28496 ;
  assign y9258 = ~n28497 ;
  assign y9259 = n28498 ;
  assign y9260 = ~1'b0 ;
  assign y9261 = ~n28501 ;
  assign y9262 = ~n28503 ;
  assign y9263 = ~1'b0 ;
  assign y9264 = n28506 ;
  assign y9265 = ~n28513 ;
  assign y9266 = ~n28516 ;
  assign y9267 = ~n28530 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = ~1'b0 ;
  assign y9270 = n28531 ;
  assign y9271 = ~n28537 ;
  assign y9272 = ~n28539 ;
  assign y9273 = ~1'b0 ;
  assign y9274 = n28549 ;
  assign y9275 = ~n28550 ;
  assign y9276 = ~n28553 ;
  assign y9277 = ~1'b0 ;
  assign y9278 = ~n28556 ;
  assign y9279 = n28560 ;
  assign y9280 = n28564 ;
  assign y9281 = ~n2241 ;
  assign y9282 = n28566 ;
  assign y9283 = ~n28567 ;
  assign y9284 = n28568 ;
  assign y9285 = n28570 ;
  assign y9286 = ~n28572 ;
  assign y9287 = n28575 ;
  assign y9288 = n3805 ;
  assign y9289 = ~1'b0 ;
  assign y9290 = n28580 ;
  assign y9291 = ~n28586 ;
  assign y9292 = ~1'b0 ;
  assign y9293 = ~1'b0 ;
  assign y9294 = ~n28587 ;
  assign y9295 = n28590 ;
  assign y9296 = ~n28591 ;
  assign y9297 = n28593 ;
  assign y9298 = n28598 ;
  assign y9299 = n28600 ;
  assign y9300 = n28602 ;
  assign y9301 = n28605 ;
  assign y9302 = ~n28610 ;
  assign y9303 = n9290 ;
  assign y9304 = n28613 ;
  assign y9305 = n28617 ;
  assign y9306 = n28624 ;
  assign y9307 = ~n28627 ;
  assign y9308 = ~n28629 ;
  assign y9309 = n28631 ;
  assign y9310 = n28634 ;
  assign y9311 = n7615 ;
  assign y9312 = ~n28635 ;
  assign y9313 = n28645 ;
  assign y9314 = n28648 ;
  assign y9315 = ~n28654 ;
  assign y9316 = n28657 ;
  assign y9317 = n5610 ;
  assign y9318 = ~1'b0 ;
  assign y9319 = ~n28662 ;
  assign y9320 = n28663 ;
  assign y9321 = n28669 ;
  assign y9322 = ~n28670 ;
  assign y9323 = n28672 ;
  assign y9324 = ~n28675 ;
  assign y9325 = n28681 ;
  assign y9326 = n28682 ;
  assign y9327 = n28683 ;
  assign y9328 = ~1'b0 ;
  assign y9329 = ~1'b0 ;
  assign y9330 = ~n28684 ;
  assign y9331 = ~1'b0 ;
  assign y9332 = ~n28689 ;
  assign y9333 = n28691 ;
  assign y9334 = n28698 ;
  assign y9335 = n28707 ;
  assign y9336 = ~1'b0 ;
  assign y9337 = ~n28709 ;
  assign y9338 = ~n17123 ;
  assign y9339 = ~n28714 ;
  assign y9340 = n28715 ;
  assign y9341 = n28718 ;
  assign y9342 = ~n28720 ;
  assign y9343 = ~n28724 ;
  assign y9344 = n28729 ;
  assign y9345 = ~n28731 ;
  assign y9346 = n28736 ;
  assign y9347 = ~1'b0 ;
  assign y9348 = ~n28739 ;
  assign y9349 = n28742 ;
  assign y9350 = ~n28744 ;
  assign y9351 = ~n28745 ;
  assign y9352 = ~n28752 ;
  assign y9353 = n28755 ;
  assign y9354 = n28763 ;
  assign y9355 = ~n28774 ;
  assign y9356 = ~n28779 ;
  assign y9357 = n28780 ;
  assign y9358 = n28784 ;
  assign y9359 = ~n28785 ;
  assign y9360 = ~n28789 ;
  assign y9361 = n28793 ;
  assign y9362 = n28794 ;
  assign y9363 = ~n28802 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = n28805 ;
  assign y9366 = n28807 ;
  assign y9367 = ~n28809 ;
  assign y9368 = ~n28811 ;
  assign y9369 = ~n28812 ;
  assign y9370 = ~n28814 ;
  assign y9371 = n28817 ;
  assign y9372 = ~1'b0 ;
  assign y9373 = ~1'b0 ;
  assign y9374 = ~n28820 ;
  assign y9375 = ~n28821 ;
  assign y9376 = ~n28824 ;
  assign y9377 = ~n28828 ;
  assign y9378 = ~n28830 ;
  assign y9379 = ~n28835 ;
  assign y9380 = ~n28836 ;
  assign y9381 = ~n28837 ;
  assign y9382 = n28838 ;
  assign y9383 = ~n28840 ;
  assign y9384 = n28843 ;
  assign y9385 = ~n28844 ;
  assign y9386 = n28849 ;
  assign y9387 = n28856 ;
  assign y9388 = ~n28860 ;
  assign y9389 = n28869 ;
  assign y9390 = ~n28872 ;
  assign y9391 = ~1'b0 ;
  assign y9392 = n28873 ;
  assign y9393 = n28882 ;
  assign y9394 = ~n18187 ;
  assign y9395 = n28883 ;
  assign y9396 = n28886 ;
  assign y9397 = ~n28889 ;
  assign y9398 = n28891 ;
  assign y9399 = ~n28893 ;
  assign y9400 = n28898 ;
  assign y9401 = ~n28901 ;
  assign y9402 = ~n28903 ;
  assign y9403 = n28906 ;
  assign y9404 = ~n28909 ;
  assign y9405 = ~1'b0 ;
  assign y9406 = n28910 ;
  assign y9407 = n28911 ;
  assign y9408 = n28922 ;
  assign y9409 = ~n28927 ;
  assign y9410 = n28929 ;
  assign y9411 = ~1'b0 ;
  assign y9412 = n28934 ;
  assign y9413 = ~1'b0 ;
  assign y9414 = n28936 ;
  assign y9415 = ~1'b0 ;
  assign y9416 = ~n28938 ;
  assign y9417 = ~n28939 ;
  assign y9418 = n28940 ;
  assign y9419 = ~n28941 ;
  assign y9420 = ~1'b0 ;
  assign y9421 = ~1'b0 ;
  assign y9422 = n28943 ;
  assign y9423 = n28945 ;
  assign y9424 = ~n28952 ;
  assign y9425 = ~1'b0 ;
  assign y9426 = n28953 ;
  assign y9427 = n28955 ;
  assign y9428 = n28956 ;
  assign y9429 = n28958 ;
  assign y9430 = n24952 ;
  assign y9431 = ~n28964 ;
  assign y9432 = n28965 ;
  assign y9433 = n28975 ;
  assign y9434 = n28981 ;
  assign y9435 = ~n28984 ;
  assign y9436 = ~n28995 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = ~n28996 ;
  assign y9439 = ~1'b0 ;
  assign y9440 = n28999 ;
  assign y9441 = n18082 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = n29001 ;
  assign y9444 = ~n29010 ;
  assign y9445 = n29012 ;
  assign y9446 = n29013 ;
  assign y9447 = n29014 ;
  assign y9448 = ~1'b0 ;
  assign y9449 = ~n29016 ;
  assign y9450 = ~n29019 ;
  assign y9451 = ~n29021 ;
  assign y9452 = n29022 ;
  assign y9453 = ~n29027 ;
  assign y9454 = ~n29028 ;
  assign y9455 = ~n29031 ;
  assign y9456 = ~n29037 ;
  assign y9457 = ~n29038 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = ~n29039 ;
  assign y9460 = ~n29042 ;
  assign y9461 = n29043 ;
  assign y9462 = ~1'b0 ;
  assign y9463 = ~1'b0 ;
  assign y9464 = n29044 ;
  assign y9465 = ~1'b0 ;
  assign y9466 = n29047 ;
  assign y9467 = n29048 ;
  assign y9468 = ~n29054 ;
  assign y9469 = n29057 ;
  assign y9470 = ~n29059 ;
  assign y9471 = n29062 ;
  assign y9472 = n29069 ;
  assign y9473 = ~1'b0 ;
  assign y9474 = ~n29072 ;
  assign y9475 = ~n29073 ;
  assign y9476 = ~n29082 ;
  assign y9477 = ~1'b0 ;
  assign y9478 = ~n29086 ;
  assign y9479 = n29091 ;
  assign y9480 = n29099 ;
  assign y9481 = ~1'b0 ;
  assign y9482 = n29101 ;
  assign y9483 = n29102 ;
  assign y9484 = n29107 ;
  assign y9485 = ~n29109 ;
  assign y9486 = ~n29116 ;
  assign y9487 = ~n29120 ;
  assign y9488 = n29122 ;
  assign y9489 = ~1'b0 ;
  assign y9490 = ~1'b0 ;
  assign y9491 = ~n29127 ;
  assign y9492 = n11196 ;
  assign y9493 = ~n29128 ;
  assign y9494 = n29131 ;
  assign y9495 = ~n29133 ;
  assign y9496 = ~1'b0 ;
  assign y9497 = ~1'b0 ;
  assign y9498 = ~1'b0 ;
  assign y9499 = ~n29134 ;
  assign y9500 = ~n29135 ;
  assign y9501 = n29140 ;
  assign y9502 = ~1'b0 ;
  assign y9503 = n29141 ;
  assign y9504 = ~n29142 ;
  assign y9505 = ~n29145 ;
  assign y9506 = n29146 ;
  assign y9507 = n29147 ;
  assign y9508 = n29150 ;
  assign y9509 = n29152 ;
  assign y9510 = n29159 ;
  assign y9511 = n29168 ;
  assign y9512 = ~n29174 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = ~n29179 ;
  assign y9515 = n29184 ;
  assign y9516 = ~n29188 ;
  assign y9517 = n29191 ;
  assign y9518 = ~n29192 ;
  assign y9519 = n29193 ;
  assign y9520 = ~n29199 ;
  assign y9521 = n1330 ;
  assign y9522 = n29200 ;
  assign y9523 = ~n29201 ;
  assign y9524 = n29202 ;
  assign y9525 = ~n29204 ;
  assign y9526 = n29214 ;
  assign y9527 = n29221 ;
  assign y9528 = n29222 ;
  assign y9529 = ~n29227 ;
  assign y9530 = ~n29228 ;
  assign y9531 = ~1'b0 ;
  assign y9532 = ~n29232 ;
  assign y9533 = n29233 ;
  assign y9534 = ~n29234 ;
  assign y9535 = n29235 ;
  assign y9536 = ~n29238 ;
  assign y9537 = 1'b0 ;
  assign y9538 = n29241 ;
  assign y9539 = ~1'b0 ;
  assign y9540 = n29243 ;
  assign y9541 = ~n29248 ;
  assign y9542 = ~n29251 ;
  assign y9543 = n29253 ;
  assign y9544 = n29256 ;
  assign y9545 = ~1'b0 ;
  assign y9546 = ~1'b0 ;
  assign y9547 = ~n29260 ;
  assign y9548 = n29271 ;
  assign y9549 = ~n29272 ;
  assign y9550 = ~n29274 ;
  assign y9551 = ~n29275 ;
  assign y9552 = ~n29277 ;
  assign y9553 = ~n29281 ;
  assign y9554 = ~n29282 ;
  assign y9555 = ~1'b0 ;
  assign y9556 = ~n29283 ;
  assign y9557 = n29284 ;
  assign y9558 = n29287 ;
  assign y9559 = n29288 ;
  assign y9560 = ~1'b0 ;
  assign y9561 = ~n29292 ;
  assign y9562 = ~1'b0 ;
  assign y9563 = n29299 ;
  assign y9564 = n29300 ;
  assign y9565 = n29302 ;
  assign y9566 = ~n29314 ;
  assign y9567 = ~1'b0 ;
  assign y9568 = ~n29316 ;
  assign y9569 = ~n15414 ;
  assign y9570 = n29318 ;
  assign y9571 = n29319 ;
  assign y9572 = ~n29327 ;
  assign y9573 = n29336 ;
  assign y9574 = ~1'b0 ;
  assign y9575 = n29338 ;
  assign y9576 = n29341 ;
  assign y9577 = n29342 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = ~n29345 ;
  assign y9580 = ~n29350 ;
  assign y9581 = n29352 ;
  assign y9582 = n29361 ;
  assign y9583 = n29364 ;
  assign y9584 = ~n29366 ;
  assign y9585 = n29369 ;
  assign y9586 = ~n29373 ;
  assign y9587 = ~1'b0 ;
  assign y9588 = ~1'b0 ;
  assign y9589 = n29379 ;
  assign y9590 = ~n29384 ;
  assign y9591 = n29386 ;
  assign y9592 = ~n29393 ;
  assign y9593 = ~n29394 ;
  assign y9594 = n29398 ;
  assign y9595 = n29399 ;
  assign y9596 = n29401 ;
  assign y9597 = n29402 ;
  assign y9598 = ~n29404 ;
  assign y9599 = ~n29406 ;
  assign y9600 = n29411 ;
  assign y9601 = ~1'b0 ;
  assign y9602 = n29418 ;
  assign y9603 = ~n29419 ;
  assign y9604 = n29420 ;
  assign y9605 = ~n29424 ;
  assign y9606 = n29429 ;
  assign y9607 = ~n29434 ;
  assign y9608 = n29435 ;
  assign y9609 = n29438 ;
  assign y9610 = ~n29440 ;
  assign y9611 = ~1'b0 ;
  assign y9612 = n29445 ;
  assign y9613 = n29453 ;
  assign y9614 = ~1'b0 ;
  assign y9615 = ~1'b0 ;
  assign y9616 = n29458 ;
  assign y9617 = n29464 ;
  assign y9618 = n29467 ;
  assign y9619 = ~n29468 ;
  assign y9620 = ~n29469 ;
  assign y9621 = ~1'b0 ;
  assign y9622 = n29470 ;
  assign y9623 = ~1'b0 ;
  assign y9624 = ~n29477 ;
  assign y9625 = n29479 ;
  assign y9626 = ~n29481 ;
  assign y9627 = n29487 ;
  assign y9628 = ~n29490 ;
  assign y9629 = ~n29492 ;
  assign y9630 = n29497 ;
  assign y9631 = n29499 ;
  assign y9632 = ~n29500 ;
  assign y9633 = ~1'b0 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~1'b0 ;
  assign y9636 = ~1'b0 ;
  assign y9637 = n29503 ;
  assign y9638 = ~n29505 ;
  assign y9639 = ~n29509 ;
  assign y9640 = ~n29512 ;
  assign y9641 = ~n29517 ;
  assign y9642 = ~n29522 ;
  assign y9643 = n4773 ;
  assign y9644 = 1'b0 ;
  assign y9645 = ~n29523 ;
  assign y9646 = n29525 ;
  assign y9647 = ~1'b0 ;
  assign y9648 = ~1'b0 ;
  assign y9649 = ~n29526 ;
  assign y9650 = ~n29532 ;
  assign y9651 = ~n29538 ;
  assign y9652 = n29542 ;
  assign y9653 = ~n29544 ;
  assign y9654 = ~n29549 ;
  assign y9655 = n29551 ;
  assign y9656 = ~n29554 ;
  assign y9657 = n29559 ;
  assign y9658 = ~1'b0 ;
  assign y9659 = ~1'b0 ;
  assign y9660 = ~n26832 ;
  assign y9661 = 1'b0 ;
  assign y9662 = n29564 ;
  assign y9663 = ~1'b0 ;
  assign y9664 = n29574 ;
  assign y9665 = n29575 ;
  assign y9666 = n29578 ;
  assign y9667 = n29582 ;
  assign y9668 = ~n29585 ;
  assign y9669 = ~1'b0 ;
  assign y9670 = ~1'b0 ;
  assign y9671 = n29591 ;
  assign y9672 = n29597 ;
  assign y9673 = ~n29601 ;
  assign y9674 = ~n29602 ;
  assign y9675 = n29608 ;
  assign y9676 = ~n29609 ;
  assign y9677 = ~n29610 ;
  assign y9678 = n29613 ;
  assign y9679 = n29614 ;
  assign y9680 = ~1'b0 ;
  assign y9681 = ~1'b0 ;
  assign y9682 = ~n29617 ;
  assign y9683 = ~n29620 ;
  assign y9684 = ~n29622 ;
  assign y9685 = ~n29623 ;
  assign y9686 = ~n29626 ;
  assign y9687 = ~n29632 ;
  assign y9688 = ~1'b0 ;
  assign y9689 = ~n29638 ;
  assign y9690 = ~1'b0 ;
  assign y9691 = ~1'b0 ;
  assign y9692 = ~1'b0 ;
  assign y9693 = n29640 ;
  assign y9694 = ~n29644 ;
  assign y9695 = ~n29648 ;
  assign y9696 = n29649 ;
  assign y9697 = ~1'b0 ;
  assign y9698 = ~1'b0 ;
  assign y9699 = ~1'b0 ;
  assign y9700 = n29650 ;
  assign y9701 = n29659 ;
  assign y9702 = ~n29662 ;
  assign y9703 = ~n29666 ;
  assign y9704 = n29668 ;
  assign y9705 = ~n29670 ;
  assign y9706 = ~n29671 ;
  assign y9707 = ~n29673 ;
  assign y9708 = ~n29676 ;
  assign y9709 = ~n29683 ;
  assign y9710 = ~1'b0 ;
  assign y9711 = 1'b0 ;
  assign y9712 = ~n29692 ;
  assign y9713 = ~n29694 ;
  assign y9714 = ~1'b0 ;
  assign y9715 = n25745 ;
  assign y9716 = ~n29695 ;
  assign y9717 = n22413 ;
  assign y9718 = n29697 ;
  assign y9719 = n29698 ;
  assign y9720 = ~1'b0 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~n29701 ;
  assign y9723 = ~n29705 ;
  assign y9724 = ~1'b0 ;
  assign y9725 = ~n29711 ;
  assign y9726 = n29715 ;
  assign y9727 = n29716 ;
  assign y9728 = ~n29717 ;
  assign y9729 = ~1'b0 ;
  assign y9730 = n29718 ;
  assign y9731 = ~n29720 ;
  assign y9732 = ~1'b0 ;
  assign y9733 = n29721 ;
  assign y9734 = ~1'b0 ;
  assign y9735 = n29722 ;
  assign y9736 = n29723 ;
  assign y9737 = ~n29725 ;
  assign y9738 = ~n29729 ;
  assign y9739 = ~1'b0 ;
  assign y9740 = n29730 ;
  assign y9741 = n29733 ;
  assign y9742 = n29735 ;
  assign y9743 = ~n21105 ;
  assign y9744 = ~n29737 ;
  assign y9745 = n29740 ;
  assign y9746 = n29741 ;
  assign y9747 = ~1'b0 ;
  assign y9748 = n29744 ;
  assign y9749 = n29745 ;
  assign y9750 = ~n29747 ;
  assign y9751 = ~n29750 ;
  assign y9752 = n29751 ;
  assign y9753 = n29755 ;
  assign y9754 = ~1'b0 ;
  assign y9755 = ~n29756 ;
  assign y9756 = ~n29757 ;
  assign y9757 = ~1'b0 ;
  assign y9758 = n29758 ;
  assign y9759 = ~1'b0 ;
  assign y9760 = ~n29762 ;
  assign y9761 = n29763 ;
  assign y9762 = n29764 ;
  assign y9763 = n29767 ;
  assign y9764 = n29771 ;
  assign y9765 = ~1'b0 ;
  assign y9766 = ~n29775 ;
  assign y9767 = n29777 ;
  assign y9768 = ~n29781 ;
  assign y9769 = ~n29783 ;
  assign y9770 = ~n29786 ;
  assign y9771 = ~n29794 ;
  assign y9772 = ~n29796 ;
  assign y9773 = ~1'b0 ;
  assign y9774 = ~1'b0 ;
  assign y9775 = ~n12988 ;
  assign y9776 = n29797 ;
  assign y9777 = ~1'b0 ;
  assign y9778 = n29808 ;
  assign y9779 = n29811 ;
  assign y9780 = ~n29813 ;
  assign y9781 = ~n29817 ;
  assign y9782 = n29818 ;
  assign y9783 = ~1'b0 ;
  assign y9784 = n29826 ;
  assign y9785 = ~1'b0 ;
  assign y9786 = n29829 ;
  assign y9787 = ~n29838 ;
  assign y9788 = ~n29841 ;
  assign y9789 = ~n29846 ;
  assign y9790 = ~1'b0 ;
  assign y9791 = ~n29847 ;
  assign y9792 = ~n29850 ;
  assign y9793 = ~n29853 ;
  assign y9794 = ~1'b0 ;
  assign y9795 = ~n29854 ;
  assign y9796 = ~n29855 ;
  assign y9797 = ~n29861 ;
  assign y9798 = n29865 ;
  assign y9799 = n29870 ;
  assign y9800 = ~n29875 ;
  assign y9801 = ~n29876 ;
  assign y9802 = n29878 ;
  assign y9803 = ~n29879 ;
  assign y9804 = n29880 ;
  assign y9805 = n29881 ;
  assign y9806 = ~n29883 ;
  assign y9807 = ~1'b0 ;
  assign y9808 = ~n29885 ;
  assign y9809 = n29886 ;
  assign y9810 = ~n29889 ;
  assign y9811 = ~1'b0 ;
  assign y9812 = ~1'b0 ;
  assign y9813 = ~n29892 ;
  assign y9814 = ~n29895 ;
  assign y9815 = n29904 ;
  assign y9816 = n29907 ;
  assign y9817 = n29909 ;
  assign y9818 = n29913 ;
  assign y9819 = ~n29917 ;
  assign y9820 = ~n29920 ;
  assign y9821 = n29928 ;
  assign y9822 = ~n29931 ;
  assign y9823 = n29934 ;
  assign y9824 = ~n29936 ;
  assign y9825 = ~n29942 ;
  assign y9826 = ~n29945 ;
  assign y9827 = ~n29948 ;
  assign y9828 = n29951 ;
  assign y9829 = n29952 ;
  assign y9830 = n29955 ;
  assign y9831 = n29960 ;
  assign y9832 = ~n29962 ;
  assign y9833 = ~n29968 ;
  assign y9834 = ~1'b0 ;
  assign y9835 = ~n29970 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = ~n29978 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = ~1'b0 ;
  assign y9840 = n29980 ;
  assign y9841 = n29981 ;
  assign y9842 = ~n29982 ;
  assign y9843 = ~n29989 ;
  assign y9844 = ~1'b0 ;
  assign y9845 = ~n29991 ;
  assign y9846 = ~1'b0 ;
  assign y9847 = ~n29992 ;
  assign y9848 = ~n29993 ;
  assign y9849 = ~n29996 ;
  assign y9850 = n29997 ;
  assign y9851 = ~1'b0 ;
  assign y9852 = n29998 ;
  assign y9853 = ~n30004 ;
  assign y9854 = ~n30007 ;
  assign y9855 = ~n30011 ;
  assign y9856 = ~n30012 ;
  assign y9857 = ~n30013 ;
  assign y9858 = ~1'b0 ;
  assign y9859 = ~1'b0 ;
  assign y9860 = n30014 ;
  assign y9861 = ~n30017 ;
  assign y9862 = n30018 ;
  assign y9863 = ~n30024 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = n30033 ;
  assign y9866 = ~1'b0 ;
  assign y9867 = n30034 ;
  assign y9868 = ~n30035 ;
  assign y9869 = n30036 ;
  assign y9870 = ~n30038 ;
  assign y9871 = ~1'b0 ;
  assign y9872 = ~1'b0 ;
  assign y9873 = n30039 ;
  assign y9874 = n30041 ;
  assign y9875 = ~1'b0 ;
  assign y9876 = ~1'b0 ;
  assign y9877 = ~1'b0 ;
  assign y9878 = ~n30043 ;
  assign y9879 = ~n30047 ;
  assign y9880 = n30056 ;
  assign y9881 = ~1'b0 ;
  assign y9882 = ~1'b0 ;
  assign y9883 = ~1'b0 ;
  assign y9884 = n30059 ;
  assign y9885 = ~1'b0 ;
  assign y9886 = ~1'b0 ;
  assign y9887 = n30060 ;
  assign y9888 = ~n30061 ;
  assign y9889 = ~n30063 ;
  assign y9890 = ~n30064 ;
  assign y9891 = ~n30066 ;
  assign y9892 = n30070 ;
  assign y9893 = ~n30073 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = n30081 ;
  assign y9896 = ~n30082 ;
  assign y9897 = n30090 ;
  assign y9898 = n30092 ;
  assign y9899 = ~n625 ;
  assign y9900 = ~n30094 ;
  assign y9901 = ~n30097 ;
  assign y9902 = ~n30099 ;
  assign y9903 = ~1'b0 ;
  assign y9904 = ~n30109 ;
  assign y9905 = ~n30111 ;
  assign y9906 = n30113 ;
  assign y9907 = ~n30114 ;
  assign y9908 = ~1'b0 ;
  assign y9909 = ~1'b0 ;
  assign y9910 = ~1'b0 ;
  assign y9911 = ~n30121 ;
  assign y9912 = ~n30123 ;
  assign y9913 = ~n30125 ;
  assign y9914 = ~1'b0 ;
  assign y9915 = ~1'b0 ;
  assign y9916 = ~n30128 ;
  assign y9917 = ~1'b0 ;
  assign y9918 = n30132 ;
  assign y9919 = ~n30134 ;
  assign y9920 = n12978 ;
  assign y9921 = ~n30138 ;
  assign y9922 = ~1'b0 ;
  assign y9923 = ~n30139 ;
  assign y9924 = ~n30142 ;
  assign y9925 = ~1'b0 ;
  assign y9926 = ~1'b0 ;
  assign y9927 = ~n30145 ;
  assign y9928 = n30147 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = ~n30152 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = n30156 ;
  assign y9933 = n30158 ;
  assign y9934 = ~n30159 ;
  assign y9935 = ~1'b0 ;
  assign y9936 = ~n30165 ;
  assign y9937 = ~n30169 ;
  assign y9938 = ~1'b0 ;
  assign y9939 = ~n30171 ;
  assign y9940 = n30175 ;
  assign y9941 = ~n30178 ;
  assign y9942 = n30180 ;
  assign y9943 = ~n30183 ;
  assign y9944 = ~n30184 ;
  assign y9945 = n30185 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = n30186 ;
  assign y9948 = ~1'b0 ;
  assign y9949 = n30193 ;
  assign y9950 = ~n30196 ;
  assign y9951 = ~n5231 ;
  assign y9952 = ~1'b0 ;
  assign y9953 = n1264 ;
  assign y9954 = n30200 ;
  assign y9955 = ~n30208 ;
  assign y9956 = ~n30211 ;
  assign y9957 = ~n30212 ;
  assign y9958 = ~n30215 ;
  assign y9959 = n30219 ;
  assign y9960 = n30221 ;
  assign y9961 = n30223 ;
  assign y9962 = ~n30233 ;
  assign y9963 = ~1'b0 ;
  assign y9964 = n30235 ;
  assign y9965 = n30236 ;
  assign y9966 = ~n30239 ;
  assign y9967 = n30244 ;
  assign y9968 = ~1'b0 ;
  assign y9969 = n30246 ;
  assign y9970 = n30248 ;
  assign y9971 = ~n30249 ;
  assign y9972 = ~n30251 ;
  assign y9973 = n30252 ;
  assign y9974 = ~n30259 ;
  assign y9975 = n30261 ;
  assign y9976 = n30262 ;
  assign y9977 = ~n30266 ;
  assign y9978 = ~1'b0 ;
  assign y9979 = n30267 ;
  assign y9980 = n30272 ;
  assign y9981 = ~n30273 ;
  assign y9982 = n30274 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = ~n30277 ;
  assign y9985 = ~n30281 ;
  assign y9986 = n30282 ;
  assign y9987 = n30284 ;
  assign y9988 = ~1'b0 ;
  assign y9989 = ~1'b0 ;
  assign y9990 = ~1'b0 ;
  assign y9991 = ~n30287 ;
  assign y9992 = n30291 ;
  assign y9993 = n30298 ;
  assign y9994 = ~n30301 ;
  assign y9995 = ~n30302 ;
  assign y9996 = n21314 ;
  assign y9997 = ~n30307 ;
  assign y9998 = ~n30314 ;
  assign y9999 = ~n30319 ;
  assign y10000 = ~1'b0 ;
  assign y10001 = n30320 ;
  assign y10002 = ~n30321 ;
  assign y10003 = ~n30325 ;
  assign y10004 = n30331 ;
  assign y10005 = ~n30333 ;
  assign y10006 = ~1'b0 ;
  assign y10007 = n30334 ;
  assign y10008 = ~n30341 ;
  assign y10009 = ~n30344 ;
  assign y10010 = n30349 ;
  assign y10011 = ~1'b0 ;
  assign y10012 = ~n30354 ;
  assign y10013 = ~n30356 ;
  assign y10014 = ~1'b0 ;
  assign y10015 = n30360 ;
  assign y10016 = ~1'b0 ;
  assign y10017 = ~n30364 ;
  assign y10018 = ~1'b0 ;
  assign y10019 = ~n30373 ;
  assign y10020 = ~n30375 ;
  assign y10021 = n30377 ;
  assign y10022 = ~n30378 ;
  assign y10023 = ~1'b0 ;
  assign y10024 = n30386 ;
  assign y10025 = ~n30388 ;
  assign y10026 = ~n30390 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = ~1'b0 ;
  assign y10029 = n30395 ;
  assign y10030 = n30396 ;
  assign y10031 = n30401 ;
  assign y10032 = n30406 ;
  assign y10033 = n30410 ;
  assign y10034 = ~n30415 ;
  assign y10035 = n30416 ;
  assign y10036 = n30417 ;
  assign y10037 = ~n30421 ;
  assign y10038 = ~n30422 ;
  assign y10039 = n30424 ;
  assign y10040 = n30429 ;
  assign y10041 = n30434 ;
  assign y10042 = n30441 ;
  assign y10043 = n30443 ;
  assign y10044 = ~n30448 ;
  assign y10045 = ~1'b0 ;
  assign y10046 = ~1'b0 ;
  assign y10047 = ~1'b0 ;
  assign y10048 = ~n30450 ;
  assign y10049 = n30452 ;
  assign y10050 = ~n30457 ;
  assign y10051 = n30459 ;
  assign y10052 = n30464 ;
  assign y10053 = n30465 ;
  assign y10054 = ~1'b0 ;
  assign y10055 = ~1'b0 ;
  assign y10056 = n30469 ;
  assign y10057 = ~n30471 ;
  assign y10058 = n30472 ;
  assign y10059 = ~n30473 ;
  assign y10060 = ~n30476 ;
  assign y10061 = ~n30479 ;
  assign y10062 = 1'b0 ;
  assign y10063 = ~n30480 ;
  assign y10064 = n30481 ;
  assign y10065 = n30484 ;
  assign y10066 = ~n30486 ;
  assign y10067 = ~1'b0 ;
  assign y10068 = n30487 ;
  assign y10069 = n30489 ;
  assign y10070 = ~n30494 ;
  assign y10071 = ~1'b0 ;
  assign y10072 = n30495 ;
  assign y10073 = ~n30496 ;
  assign y10074 = ~n30498 ;
  assign y10075 = n30500 ;
  assign y10076 = ~n30504 ;
  assign y10077 = n30506 ;
  assign y10078 = n30508 ;
  assign y10079 = ~n30512 ;
  assign y10080 = n30513 ;
  assign y10081 = ~n30522 ;
  assign y10082 = ~n30528 ;
  assign y10083 = n14625 ;
  assign y10084 = ~n30530 ;
  assign y10085 = ~n30539 ;
  assign y10086 = n30540 ;
  assign y10087 = ~n30543 ;
  assign y10088 = ~1'b0 ;
  assign y10089 = ~n30544 ;
  assign y10090 = ~1'b0 ;
  assign y10091 = n30550 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = ~n30552 ;
  assign y10094 = ~1'b0 ;
  assign y10095 = n30554 ;
  assign y10096 = ~n30555 ;
  assign y10097 = ~n30557 ;
  assign y10098 = ~n30558 ;
  assign y10099 = n30560 ;
  assign y10100 = n30561 ;
  assign y10101 = ~n30565 ;
  assign y10102 = ~n30566 ;
  assign y10103 = n30568 ;
  assign y10104 = ~n30570 ;
  assign y10105 = 1'b0 ;
  assign y10106 = ~n30572 ;
  assign y10107 = ~n30576 ;
  assign y10108 = n30577 ;
  assign y10109 = ~n30582 ;
  assign y10110 = n30586 ;
  assign y10111 = ~n30588 ;
  assign y10112 = ~n30590 ;
  assign y10113 = ~n30597 ;
  assign y10114 = ~n30598 ;
  assign y10115 = ~n30599 ;
  assign y10116 = n30606 ;
  assign y10117 = ~1'b0 ;
  assign y10118 = n30608 ;
  assign y10119 = n30610 ;
  assign y10120 = n30612 ;
  assign y10121 = n30613 ;
  assign y10122 = n30615 ;
  assign y10123 = n30621 ;
  assign y10124 = ~n30622 ;
  assign y10125 = ~n30624 ;
  assign y10126 = ~n30628 ;
  assign y10127 = ~n30633 ;
  assign y10128 = n30638 ;
  assign y10129 = ~n30639 ;
  assign y10130 = n30640 ;
  assign y10131 = ~n30641 ;
  assign y10132 = ~n30642 ;
  assign y10133 = n30644 ;
  assign y10134 = ~n30649 ;
  assign y10135 = ~n30650 ;
  assign y10136 = ~1'b0 ;
  assign y10137 = ~1'b0 ;
  assign y10138 = ~n30652 ;
  assign y10139 = ~n30653 ;
  assign y10140 = ~1'b0 ;
  assign y10141 = ~n30655 ;
  assign y10142 = ~n30656 ;
  assign y10143 = ~n30663 ;
  assign y10144 = ~1'b0 ;
  assign y10145 = ~n30670 ;
  assign y10146 = ~1'b0 ;
  assign y10147 = ~n30674 ;
  assign y10148 = n30676 ;
  assign y10149 = n30678 ;
  assign y10150 = ~1'b0 ;
  assign y10151 = n30681 ;
  assign y10152 = ~n30683 ;
  assign y10153 = ~n30684 ;
  assign y10154 = ~n30685 ;
  assign y10155 = n30686 ;
  assign y10156 = n30690 ;
  assign y10157 = ~n30706 ;
  assign y10158 = ~1'b0 ;
  assign y10159 = ~n30711 ;
  assign y10160 = n30713 ;
  assign y10161 = n30718 ;
  assign y10162 = ~n30720 ;
  assign y10163 = ~n30721 ;
  assign y10164 = n30724 ;
  assign y10165 = ~n30725 ;
  assign y10166 = n30726 ;
  assign y10167 = n30727 ;
  assign y10168 = n30730 ;
  assign y10169 = ~1'b0 ;
  assign y10170 = 1'b0 ;
  assign y10171 = n30734 ;
  assign y10172 = n7531 ;
  assign y10173 = n30740 ;
  assign y10174 = ~1'b0 ;
  assign y10175 = ~n30743 ;
  assign y10176 = ~n30744 ;
  assign y10177 = ~n30745 ;
  assign y10178 = ~n30746 ;
  assign y10179 = ~n30748 ;
  assign y10180 = ~n30749 ;
  assign y10181 = n30750 ;
  assign y10182 = n30751 ;
  assign y10183 = ~1'b0 ;
  assign y10184 = ~n30755 ;
  assign y10185 = ~1'b0 ;
  assign y10186 = ~n30756 ;
  assign y10187 = ~n30758 ;
  assign y10188 = ~n30760 ;
  assign y10189 = ~n30762 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = n30764 ;
  assign y10192 = ~n30766 ;
  assign y10193 = ~n30767 ;
  assign y10194 = ~n30769 ;
  assign y10195 = ~1'b0 ;
  assign y10196 = ~1'b0 ;
  assign y10197 = ~n30779 ;
  assign y10198 = n30782 ;
  assign y10199 = ~n30783 ;
  assign y10200 = n30787 ;
  assign y10201 = n30789 ;
  assign y10202 = ~n30796 ;
  assign y10203 = ~1'b0 ;
  assign y10204 = ~n30797 ;
  assign y10205 = ~1'b0 ;
  assign y10206 = ~1'b0 ;
  assign y10207 = ~1'b0 ;
  assign y10208 = ~n30802 ;
  assign y10209 = ~1'b0 ;
  assign y10210 = ~n30803 ;
  assign y10211 = ~1'b0 ;
  assign y10212 = ~n30806 ;
  assign y10213 = ~n30810 ;
  assign y10214 = n30811 ;
  assign y10215 = ~n30813 ;
  assign y10216 = n30821 ;
  assign y10217 = n352 ;
  assign y10218 = ~n30822 ;
  assign y10219 = n30823 ;
  assign y10220 = n20192 ;
  assign y10221 = n30826 ;
  assign y10222 = ~1'b0 ;
  assign y10223 = ~n30827 ;
  assign y10224 = ~n30828 ;
  assign y10225 = ~n30829 ;
  assign y10226 = n30831 ;
  assign y10227 = ~1'b0 ;
  assign y10228 = n30836 ;
  assign y10229 = n30837 ;
  assign y10230 = ~n30841 ;
  assign y10231 = ~n30847 ;
  assign y10232 = ~n30849 ;
  assign y10233 = n30853 ;
  assign y10234 = n30854 ;
  assign y10235 = ~n30859 ;
  assign y10236 = ~n30862 ;
  assign y10237 = n30865 ;
  assign y10238 = ~1'b0 ;
  assign y10239 = ~1'b0 ;
  assign y10240 = ~1'b0 ;
  assign y10241 = ~n30869 ;
  assign y10242 = n30872 ;
  assign y10243 = n30874 ;
  assign y10244 = n30875 ;
  assign y10245 = n30880 ;
  assign y10246 = ~n30887 ;
  assign y10247 = ~1'b0 ;
  assign y10248 = ~n30888 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = ~n30889 ;
  assign y10251 = ~n30893 ;
  assign y10252 = ~n30895 ;
  assign y10253 = n30898 ;
  assign y10254 = ~n30904 ;
  assign y10255 = ~1'b0 ;
  assign y10256 = ~n30905 ;
  assign y10257 = n30912 ;
  assign y10258 = ~n30919 ;
  assign y10259 = ~n30921 ;
  assign y10260 = ~1'b0 ;
  assign y10261 = ~n30924 ;
  assign y10262 = n30932 ;
  assign y10263 = ~n30933 ;
  assign y10264 = n30934 ;
  assign y10265 = n30937 ;
  assign y10266 = ~n30942 ;
  assign y10267 = ~n30945 ;
  assign y10268 = ~n30946 ;
  assign y10269 = ~1'b0 ;
  assign y10270 = ~n30950 ;
  assign y10271 = ~n30952 ;
  assign y10272 = ~n30953 ;
  assign y10273 = ~n30955 ;
  assign y10274 = n5681 ;
  assign y10275 = n27150 ;
  assign y10276 = n30957 ;
  assign y10277 = ~1'b0 ;
  assign y10278 = ~n30967 ;
  assign y10279 = ~1'b0 ;
  assign y10280 = n28823 ;
  assign y10281 = n30968 ;
  assign y10282 = ~n30969 ;
  assign y10283 = ~n30970 ;
  assign y10284 = n30978 ;
  assign y10285 = ~n30980 ;
  assign y10286 = ~n30981 ;
  assign y10287 = n30983 ;
  assign y10288 = ~1'b0 ;
  assign y10289 = ~n30985 ;
  assign y10290 = ~n30991 ;
  assign y10291 = n30992 ;
  assign y10292 = n30997 ;
  assign y10293 = n30998 ;
  assign y10294 = ~n30999 ;
  assign y10295 = ~n31001 ;
  assign y10296 = ~n31002 ;
  assign y10297 = ~n31005 ;
  assign y10298 = ~n31007 ;
  assign y10299 = ~1'b0 ;
  assign y10300 = n31013 ;
  assign y10301 = n31017 ;
  assign y10302 = ~n31019 ;
  assign y10303 = ~n31027 ;
  assign y10304 = ~n31030 ;
  assign y10305 = n31034 ;
  assign y10306 = ~n31039 ;
  assign y10307 = ~1'b0 ;
  assign y10308 = ~n31045 ;
  assign y10309 = ~n31051 ;
  assign y10310 = n31056 ;
  assign y10311 = ~n31059 ;
  assign y10312 = ~n31063 ;
  assign y10313 = ~1'b0 ;
  assign y10314 = ~1'b0 ;
  assign y10315 = ~n31066 ;
  assign y10316 = n31067 ;
  assign y10317 = ~n31070 ;
  assign y10318 = ~n17513 ;
  assign y10319 = ~n31072 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = ~1'b0 ;
  assign y10322 = n31074 ;
  assign y10323 = n31075 ;
  assign y10324 = ~n31078 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~n31080 ;
  assign y10327 = n31081 ;
  assign y10328 = n31089 ;
  assign y10329 = ~n31092 ;
  assign y10330 = n31094 ;
  assign y10331 = n31095 ;
  assign y10332 = ~n31100 ;
  assign y10333 = ~n31102 ;
  assign y10334 = n31105 ;
  assign y10335 = n31112 ;
  assign y10336 = ~n31114 ;
  assign y10337 = ~1'b0 ;
  assign y10338 = ~1'b0 ;
  assign y10339 = n31116 ;
  assign y10340 = ~n31121 ;
  assign y10341 = n31127 ;
  assign y10342 = ~n31129 ;
  assign y10343 = ~n31130 ;
  assign y10344 = ~1'b0 ;
  assign y10345 = n31131 ;
  assign y10346 = n31136 ;
  assign y10347 = ~n31137 ;
  assign y10348 = ~n31144 ;
  assign y10349 = ~1'b0 ;
  assign y10350 = n31147 ;
  assign y10351 = n31153 ;
  assign y10352 = n31156 ;
  assign y10353 = ~n31157 ;
  assign y10354 = n31159 ;
  assign y10355 = n31162 ;
  assign y10356 = ~1'b0 ;
  assign y10357 = ~n31171 ;
  assign y10358 = ~1'b0 ;
  assign y10359 = ~n31172 ;
  assign y10360 = ~n31173 ;
  assign y10361 = ~n31177 ;
  assign y10362 = ~n31182 ;
  assign y10363 = ~n31190 ;
  assign y10364 = ~n31191 ;
  assign y10365 = n10113 ;
  assign y10366 = ~1'b0 ;
  assign y10367 = ~n31195 ;
  assign y10368 = ~n31196 ;
  assign y10369 = n31197 ;
  assign y10370 = n31206 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = n31208 ;
  assign y10373 = n31210 ;
  assign y10374 = ~n31212 ;
  assign y10375 = ~n31218 ;
  assign y10376 = n31222 ;
  assign y10377 = ~1'b0 ;
  assign y10378 = ~1'b0 ;
  assign y10379 = n31223 ;
  assign y10380 = ~n31225 ;
  assign y10381 = n31232 ;
  assign y10382 = n31235 ;
  assign y10383 = ~n31246 ;
  assign y10384 = n31247 ;
  assign y10385 = n31250 ;
  assign y10386 = n31256 ;
  assign y10387 = ~1'b0 ;
  assign y10388 = ~n31257 ;
  assign y10389 = n31262 ;
  assign y10390 = n31265 ;
  assign y10391 = n31267 ;
  assign y10392 = n31272 ;
  assign y10393 = ~n31274 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = n31279 ;
  assign y10396 = n31280 ;
  assign y10397 = ~n31288 ;
  assign y10398 = ~n31293 ;
  assign y10399 = ~1'b0 ;
  assign y10400 = ~1'b0 ;
  assign y10401 = n31294 ;
  assign y10402 = ~n31302 ;
  assign y10403 = n31305 ;
  assign y10404 = n31306 ;
  assign y10405 = ~n31308 ;
  assign y10406 = ~1'b0 ;
  assign y10407 = ~1'b0 ;
  assign y10408 = ~n31310 ;
  assign y10409 = n31312 ;
  assign y10410 = ~n31313 ;
  assign y10411 = ~n31317 ;
  assign y10412 = ~n31324 ;
  assign y10413 = ~1'b0 ;
  assign y10414 = ~1'b0 ;
  assign y10415 = n31328 ;
  assign y10416 = ~n31329 ;
  assign y10417 = ~1'b0 ;
  assign y10418 = ~n31333 ;
  assign y10419 = ~1'b0 ;
  assign y10420 = ~n31335 ;
  assign y10421 = ~n31340 ;
  assign y10422 = ~n31342 ;
  assign y10423 = ~n31345 ;
  assign y10424 = n31349 ;
  assign y10425 = ~1'b0 ;
  assign y10426 = ~n31356 ;
  assign y10427 = ~n31358 ;
  assign y10428 = n31364 ;
  assign y10429 = ~1'b0 ;
  assign y10430 = ~n31367 ;
  assign y10431 = n31372 ;
  assign y10432 = ~n31377 ;
  assign y10433 = ~n31378 ;
  assign y10434 = ~n31381 ;
  assign y10435 = ~n31392 ;
  assign y10436 = ~n31396 ;
  assign y10437 = ~n31397 ;
  assign y10438 = ~n31399 ;
  assign y10439 = ~n31405 ;
  assign y10440 = n31408 ;
  assign y10441 = ~n31414 ;
  assign y10442 = n31416 ;
  assign y10443 = n31419 ;
  assign y10444 = n31421 ;
  assign y10445 = ~n31422 ;
  assign y10446 = ~1'b0 ;
  assign y10447 = n31423 ;
  assign y10448 = n31427 ;
  assign y10449 = ~1'b0 ;
  assign y10450 = ~n31429 ;
  assign y10451 = n31431 ;
  assign y10452 = n31432 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = n20169 ;
  assign y10455 = n31438 ;
  assign y10456 = ~n31443 ;
  assign y10457 = n31444 ;
  assign y10458 = n31451 ;
  assign y10459 = n31452 ;
  assign y10460 = ~n31453 ;
  assign y10461 = ~1'b0 ;
  assign y10462 = ~n31455 ;
  assign y10463 = n31460 ;
  assign y10464 = ~n31462 ;
  assign y10465 = ~n31464 ;
  assign y10466 = n31465 ;
  assign y10467 = n31467 ;
  assign y10468 = ~n31469 ;
  assign y10469 = n13431 ;
  assign y10470 = n31470 ;
  assign y10471 = ~n31472 ;
  assign y10472 = n31477 ;
  assign y10473 = ~n31481 ;
  assign y10474 = ~n31483 ;
  assign y10475 = n31486 ;
  assign y10476 = ~1'b0 ;
  assign y10477 = ~n31495 ;
  assign y10478 = n31498 ;
  assign y10479 = n31503 ;
  assign y10480 = n31507 ;
  assign y10481 = ~n31513 ;
  assign y10482 = ~n31517 ;
  assign y10483 = n31522 ;
  assign y10484 = n31525 ;
  assign y10485 = n31527 ;
  assign y10486 = ~1'b0 ;
  assign y10487 = ~n31535 ;
  assign y10488 = ~n13183 ;
  assign y10489 = ~n31537 ;
  assign y10490 = ~n30572 ;
  assign y10491 = ~n31547 ;
  assign y10492 = n31549 ;
  assign y10493 = ~n31550 ;
  assign y10494 = n31558 ;
  assign y10495 = ~1'b0 ;
  assign y10496 = ~n31561 ;
  assign y10497 = n31566 ;
  assign y10498 = n31572 ;
  assign y10499 = ~n31576 ;
  assign y10500 = ~n31581 ;
  assign y10501 = ~n31583 ;
  assign y10502 = ~1'b0 ;
  assign y10503 = ~1'b0 ;
  assign y10504 = ~n31593 ;
  assign y10505 = ~n31595 ;
  assign y10506 = ~1'b0 ;
  assign y10507 = n31602 ;
  assign y10508 = ~n31604 ;
  assign y10509 = ~n31605 ;
  assign y10510 = ~n31615 ;
  assign y10511 = ~n31617 ;
  assign y10512 = ~n31627 ;
  assign y10513 = n31629 ;
  assign y10514 = ~n31635 ;
  assign y10515 = ~n31639 ;
  assign y10516 = ~n31640 ;
  assign y10517 = ~n30571 ;
  assign y10518 = ~n31641 ;
  assign y10519 = ~n31646 ;
  assign y10520 = n31649 ;
  assign y10521 = n31655 ;
  assign y10522 = ~n31656 ;
  assign y10523 = ~n31658 ;
  assign y10524 = n31663 ;
  assign y10525 = n31671 ;
  assign y10526 = ~n31673 ;
  assign y10527 = ~n31679 ;
  assign y10528 = n31680 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = n31687 ;
  assign y10532 = n31691 ;
  assign y10533 = ~n31699 ;
  assign y10534 = n31701 ;
  assign y10535 = ~n31711 ;
  assign y10536 = ~n31712 ;
  assign y10537 = ~n31716 ;
  assign y10538 = ~n31718 ;
  assign y10539 = n31720 ;
  assign y10540 = n31721 ;
  assign y10541 = ~n31723 ;
  assign y10542 = ~n31725 ;
  assign y10543 = n31730 ;
  assign y10544 = n31733 ;
  assign y10545 = ~n31738 ;
  assign y10546 = ~n31740 ;
  assign y10547 = ~n31741 ;
  assign y10548 = n31742 ;
  assign y10549 = ~1'b0 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = ~n31744 ;
  assign y10552 = ~n31747 ;
  assign y10553 = ~n31750 ;
  assign y10554 = n31752 ;
  assign y10555 = n31762 ;
  assign y10556 = ~1'b0 ;
  assign y10557 = n31763 ;
  assign y10558 = n31769 ;
  assign y10559 = ~n31774 ;
  assign y10560 = ~n31776 ;
  assign y10561 = ~n31784 ;
  assign y10562 = ~n31787 ;
  assign y10563 = n31798 ;
  assign y10564 = n31802 ;
  assign y10565 = n31806 ;
  assign y10566 = ~n31808 ;
  assign y10567 = 1'b0 ;
  assign y10568 = ~n31809 ;
  assign y10569 = ~n31810 ;
  assign y10570 = ~n31814 ;
  assign y10571 = n31821 ;
  assign y10572 = n31825 ;
  assign y10573 = ~1'b0 ;
  assign y10574 = ~1'b0 ;
  assign y10575 = ~n31827 ;
  assign y10576 = ~n31828 ;
  assign y10577 = ~n31836 ;
  assign y10578 = ~n31840 ;
  assign y10579 = ~1'b0 ;
  assign y10580 = ~n31844 ;
  assign y10581 = ~n31846 ;
  assign y10582 = ~n31847 ;
  assign y10583 = ~n31848 ;
  assign y10584 = ~1'b0 ;
  assign y10585 = ~n31849 ;
  assign y10586 = ~n31852 ;
  assign y10587 = ~1'b0 ;
  assign y10588 = ~n31853 ;
  assign y10589 = n31854 ;
  assign y10590 = ~n31858 ;
  assign y10591 = ~1'b0 ;
  assign y10592 = ~1'b0 ;
  assign y10593 = ~1'b0 ;
  assign y10594 = ~1'b0 ;
  assign y10595 = ~1'b0 ;
  assign y10596 = n4839 ;
  assign y10597 = n31874 ;
  assign y10598 = n31876 ;
  assign y10599 = n31877 ;
  assign y10600 = n31878 ;
  assign y10601 = ~n31884 ;
  assign y10602 = ~n31885 ;
  assign y10603 = ~1'b0 ;
  assign y10604 = n31890 ;
  assign y10605 = ~n31891 ;
  assign y10606 = n31895 ;
  assign y10607 = ~1'b0 ;
  assign y10608 = ~n31896 ;
  assign y10609 = ~n31901 ;
  assign y10610 = n31902 ;
  assign y10611 = ~n31903 ;
  assign y10612 = n31907 ;
  assign y10613 = n31913 ;
  assign y10614 = n31914 ;
  assign y10615 = ~1'b0 ;
  assign y10616 = n31922 ;
  assign y10617 = ~n31927 ;
  assign y10618 = ~n31928 ;
  assign y10619 = ~n31935 ;
  assign y10620 = ~n31937 ;
  assign y10621 = n31939 ;
  assign y10622 = ~n31942 ;
  assign y10623 = n31944 ;
  assign y10624 = n31945 ;
  assign y10625 = ~n31954 ;
  assign y10626 = ~n31958 ;
  assign y10627 = ~n31960 ;
  assign y10628 = n31965 ;
  assign y10629 = ~n31967 ;
  assign y10630 = ~n31968 ;
  assign y10631 = ~n31976 ;
  assign y10632 = n31977 ;
  assign y10633 = ~n31979 ;
  assign y10634 = ~n31981 ;
  assign y10635 = ~n31986 ;
  assign y10636 = ~n31989 ;
  assign y10637 = n31993 ;
  assign y10638 = ~n31995 ;
  assign y10639 = n31998 ;
  assign y10640 = ~1'b0 ;
  assign y10641 = ~n31999 ;
  assign y10642 = n32001 ;
  assign y10643 = n32004 ;
  assign y10644 = n32008 ;
  assign y10645 = ~n32011 ;
  assign y10646 = n32012 ;
  assign y10647 = ~n32016 ;
  assign y10648 = n32017 ;
  assign y10649 = ~1'b0 ;
  assign y10650 = n32019 ;
  assign y10651 = ~n32021 ;
  assign y10652 = ~1'b0 ;
  assign y10653 = n32026 ;
  assign y10654 = ~n32029 ;
  assign y10655 = ~n32035 ;
  assign y10656 = ~n32037 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = ~1'b0 ;
  assign y10659 = ~n32039 ;
  assign y10660 = ~n32046 ;
  assign y10661 = n32048 ;
  assign y10662 = n32052 ;
  assign y10663 = ~n32053 ;
  assign y10664 = ~1'b0 ;
  assign y10665 = n32056 ;
  assign y10666 = n32058 ;
  assign y10667 = n32059 ;
  assign y10668 = ~1'b0 ;
  assign y10669 = n32061 ;
  assign y10670 = n32062 ;
  assign y10671 = n10363 ;
  assign y10672 = n32064 ;
  assign y10673 = ~n32069 ;
  assign y10674 = ~n32073 ;
  assign y10675 = ~n32076 ;
  assign y10676 = ~n32077 ;
  assign y10677 = ~n32081 ;
  assign y10678 = ~n32086 ;
  assign y10679 = n32087 ;
  assign y10680 = n32088 ;
  assign y10681 = n32094 ;
  assign y10682 = n32095 ;
  assign y10683 = ~1'b0 ;
  assign y10684 = ~n32100 ;
  assign y10685 = ~1'b0 ;
  assign y10686 = ~n32102 ;
  assign y10687 = ~1'b0 ;
  assign y10688 = n32103 ;
  assign y10689 = ~n32114 ;
  assign y10690 = ~n32118 ;
  assign y10691 = ~n32125 ;
  assign y10692 = ~1'b0 ;
  assign y10693 = ~1'b0 ;
  assign y10694 = ~1'b0 ;
  assign y10695 = n32135 ;
  assign y10696 = ~n32136 ;
  assign y10697 = ~n32139 ;
  assign y10698 = n32140 ;
  assign y10699 = n32145 ;
  assign y10700 = ~n32147 ;
  assign y10701 = ~1'b0 ;
  assign y10702 = n32152 ;
  assign y10703 = n32158 ;
  assign y10704 = ~n32160 ;
  assign y10705 = n32165 ;
  assign y10706 = n32166 ;
  assign y10707 = ~1'b0 ;
  assign y10708 = ~1'b0 ;
  assign y10709 = ~n32169 ;
  assign y10710 = ~n32171 ;
  assign y10711 = ~n32184 ;
  assign y10712 = n32188 ;
  assign y10713 = ~1'b0 ;
  assign y10714 = n32192 ;
  assign y10715 = ~n32193 ;
  assign y10716 = n32198 ;
  assign y10717 = n32200 ;
  assign y10718 = n32202 ;
  assign y10719 = n32204 ;
  assign y10720 = 1'b0 ;
  assign y10721 = ~n32205 ;
  assign y10722 = n32207 ;
  assign y10723 = n32214 ;
  assign y10724 = n32215 ;
  assign y10725 = ~n32217 ;
  assign y10726 = n32221 ;
  assign y10727 = n32222 ;
  assign y10728 = n32224 ;
  assign y10729 = ~1'b0 ;
  assign y10730 = n32233 ;
  assign y10731 = n32234 ;
  assign y10732 = ~n32244 ;
  assign y10733 = n32247 ;
  assign y10734 = ~n32248 ;
  assign y10735 = ~n32252 ;
  assign y10736 = n32257 ;
  assign y10737 = ~n32258 ;
  assign y10738 = ~n32264 ;
  assign y10739 = ~n32265 ;
  assign y10740 = n32266 ;
  assign y10741 = n32271 ;
  assign y10742 = ~n32273 ;
  assign y10743 = n32278 ;
  assign y10744 = ~n32280 ;
  assign y10745 = n32281 ;
  assign y10746 = n32285 ;
  assign y10747 = n32286 ;
  assign y10748 = ~n32289 ;
  assign y10749 = n32291 ;
  assign y10750 = n25287 ;
  assign y10751 = ~1'b0 ;
  assign y10752 = ~n32294 ;
  assign y10753 = n32295 ;
  assign y10754 = n4476 ;
  assign y10755 = ~n32297 ;
  assign y10756 = n32301 ;
  assign y10757 = ~n32311 ;
  assign y10758 = ~n32313 ;
  assign y10759 = n32314 ;
  assign y10760 = ~n32315 ;
  assign y10761 = ~1'b0 ;
  assign y10762 = ~1'b0 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = n32317 ;
  assign y10765 = ~n32321 ;
  assign y10766 = ~n32323 ;
  assign y10767 = n32327 ;
  assign y10768 = n32328 ;
  assign y10769 = ~n30351 ;
  assign y10770 = ~n32331 ;
  assign y10771 = ~n32334 ;
  assign y10772 = ~n32339 ;
  assign y10773 = ~n32340 ;
  assign y10774 = n32342 ;
  assign y10775 = n32345 ;
  assign y10776 = ~n32347 ;
  assign y10777 = ~n32349 ;
  assign y10778 = n32352 ;
  assign y10779 = n32353 ;
  assign y10780 = n32361 ;
  assign y10781 = n32362 ;
  assign y10782 = n32363 ;
  assign y10783 = n32364 ;
  assign y10784 = ~n32369 ;
  assign y10785 = ~n32372 ;
  assign y10786 = ~n3523 ;
  assign y10787 = ~n32376 ;
  assign y10788 = n32378 ;
  assign y10789 = ~n32380 ;
  assign y10790 = n32382 ;
  assign y10791 = ~n32383 ;
  assign y10792 = n32393 ;
  assign y10793 = ~n32394 ;
  assign y10794 = ~n32395 ;
  assign y10795 = n32396 ;
  assign y10796 = ~n32401 ;
  assign y10797 = ~n32402 ;
  assign y10798 = n32414 ;
  assign y10799 = n32416 ;
  assign y10800 = ~1'b0 ;
  assign y10801 = ~1'b0 ;
  assign y10802 = n32418 ;
  assign y10803 = ~n32421 ;
  assign y10804 = ~n32422 ;
  assign y10805 = ~n32427 ;
  assign y10806 = ~n32428 ;
  assign y10807 = n32430 ;
  assign y10808 = n32436 ;
  assign y10809 = n32437 ;
  assign y10810 = n32441 ;
  assign y10811 = n32442 ;
  assign y10812 = n32443 ;
  assign y10813 = n32444 ;
  assign y10814 = n32451 ;
  assign y10815 = ~n32457 ;
  assign y10816 = ~n32464 ;
  assign y10817 = ~n32475 ;
  assign y10818 = ~n32477 ;
  assign y10819 = n32479 ;
  assign y10820 = ~1'b0 ;
  assign y10821 = ~n32481 ;
  assign y10822 = ~n32482 ;
  assign y10823 = ~n32484 ;
  assign y10824 = n32485 ;
  assign y10825 = ~n32487 ;
  assign y10826 = ~n32488 ;
  assign y10827 = ~n32491 ;
  assign y10828 = ~n32494 ;
  assign y10829 = ~1'b0 ;
  assign y10830 = ~n32504 ;
  assign y10831 = ~n32508 ;
  assign y10832 = n16471 ;
  assign y10833 = n32510 ;
  assign y10834 = ~n32511 ;
  assign y10835 = ~n32512 ;
  assign y10836 = ~n32515 ;
  assign y10837 = n32518 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = n32519 ;
  assign y10840 = ~n32521 ;
  assign y10841 = n32523 ;
  assign y10842 = ~n11766 ;
  assign y10843 = ~n32530 ;
  assign y10844 = ~1'b0 ;
  assign y10845 = ~n32532 ;
  assign y10846 = n32533 ;
  assign y10847 = ~1'b0 ;
  assign y10848 = ~n32535 ;
  assign y10849 = ~n32537 ;
  assign y10850 = n32540 ;
  assign y10851 = ~1'b0 ;
  assign y10852 = n32541 ;
  assign y10853 = n32543 ;
  assign y10854 = ~n32549 ;
  assign y10855 = ~n32554 ;
  assign y10856 = n32555 ;
  assign y10857 = n32557 ;
  assign y10858 = ~n32560 ;
  assign y10859 = ~1'b0 ;
  assign y10860 = ~n32561 ;
  assign y10861 = ~1'b0 ;
  assign y10862 = n32563 ;
  assign y10863 = ~n32528 ;
  assign y10864 = n32564 ;
  assign y10865 = ~n32566 ;
  assign y10866 = ~n32570 ;
  assign y10867 = ~n32572 ;
  assign y10868 = ~n32575 ;
  assign y10869 = n32576 ;
  assign y10870 = n32580 ;
  assign y10871 = ~n32582 ;
  assign y10872 = ~1'b0 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = ~n32587 ;
  assign y10875 = ~n2333 ;
  assign y10876 = ~1'b0 ;
  assign y10877 = ~n32598 ;
  assign y10878 = ~n32601 ;
  assign y10879 = n32602 ;
  assign y10880 = ~n32604 ;
  assign y10881 = n32608 ;
  assign y10882 = ~n32612 ;
  assign y10883 = ~n32615 ;
  assign y10884 = n32619 ;
  assign y10885 = ~n32620 ;
  assign y10886 = n32622 ;
  assign y10887 = ~n32624 ;
  assign y10888 = n32628 ;
  assign y10889 = ~1'b0 ;
  assign y10890 = ~n32634 ;
  assign y10891 = n32639 ;
  assign y10892 = ~n32640 ;
  assign y10893 = n32641 ;
  assign y10894 = ~n32646 ;
  assign y10895 = n32648 ;
  assign y10896 = ~n32649 ;
  assign y10897 = ~n32653 ;
  assign y10898 = n32657 ;
  assign y10899 = n32658 ;
  assign y10900 = ~1'b0 ;
  assign y10901 = ~1'b0 ;
  assign y10902 = n32659 ;
  assign y10903 = ~n32660 ;
  assign y10904 = n32661 ;
  assign y10905 = ~n32667 ;
  assign y10906 = ~n32670 ;
  assign y10907 = ~n32671 ;
  assign y10908 = ~n32674 ;
  assign y10909 = ~1'b0 ;
  assign y10910 = ~n32675 ;
  assign y10911 = n32677 ;
  assign y10912 = ~n32681 ;
  assign y10913 = ~n32683 ;
  assign y10914 = n32684 ;
  assign y10915 = n32685 ;
  assign y10916 = n32686 ;
  assign y10917 = n32693 ;
  assign y10918 = ~n32695 ;
  assign y10919 = ~n14336 ;
  assign y10920 = n32698 ;
  assign y10921 = ~n32702 ;
  assign y10922 = ~n32704 ;
  assign y10923 = ~n32707 ;
  assign y10924 = ~n32709 ;
  assign y10925 = ~n32710 ;
  assign y10926 = n32715 ;
  assign y10927 = n32722 ;
  assign y10928 = ~n32725 ;
  assign y10929 = ~n32732 ;
  assign y10930 = ~n32734 ;
  assign y10931 = ~1'b0 ;
  assign y10932 = ~1'b0 ;
  assign y10933 = n32735 ;
  assign y10934 = ~1'b0 ;
  assign y10935 = ~n32737 ;
  assign y10936 = n28819 ;
  assign y10937 = ~n32740 ;
  assign y10938 = n32742 ;
  assign y10939 = n32744 ;
  assign y10940 = ~n32747 ;
  assign y10941 = ~n32751 ;
  assign y10942 = n32755 ;
  assign y10943 = ~n32757 ;
  assign y10944 = n32765 ;
  assign y10945 = n32766 ;
  assign y10946 = ~n32777 ;
  assign y10947 = ~1'b0 ;
  assign y10948 = ~1'b0 ;
  assign y10949 = n32778 ;
  assign y10950 = ~n32781 ;
  assign y10951 = ~n32783 ;
  assign y10952 = n32784 ;
  assign y10953 = ~n32788 ;
  assign y10954 = ~1'b0 ;
  assign y10955 = n8384 ;
  assign y10956 = n31285 ;
  assign y10957 = n32793 ;
  assign y10958 = ~n32794 ;
  assign y10959 = n32795 ;
  assign y10960 = ~n32798 ;
  assign y10961 = ~n13121 ;
  assign y10962 = ~n32802 ;
  assign y10963 = ~n32804 ;
  assign y10964 = n32808 ;
  assign y10965 = n3174 ;
  assign y10966 = n32810 ;
  assign y10967 = ~n32817 ;
  assign y10968 = n32818 ;
  assign y10969 = n32821 ;
  assign y10970 = ~n32824 ;
  assign y10971 = n32825 ;
  assign y10972 = ~n32827 ;
  assign y10973 = n32828 ;
  assign y10974 = ~1'b0 ;
  assign y10975 = ~1'b0 ;
  assign y10976 = n32834 ;
  assign y10977 = ~n32838 ;
  assign y10978 = n32842 ;
  assign y10979 = ~1'b0 ;
  assign y10980 = n32845 ;
  assign y10981 = ~n32847 ;
  assign y10982 = n32849 ;
  assign y10983 = n32851 ;
  assign y10984 = ~n32852 ;
  assign y10985 = n32854 ;
  assign y10986 = ~1'b0 ;
  assign y10987 = ~1'b0 ;
  assign y10988 = n32856 ;
  assign y10989 = n32861 ;
  assign y10990 = n32869 ;
  assign y10991 = n32876 ;
  assign y10992 = n32883 ;
  assign y10993 = ~1'b0 ;
  assign y10994 = n32888 ;
  assign y10995 = n32890 ;
  assign y10996 = ~n32897 ;
  assign y10997 = ~n32898 ;
  assign y10998 = ~n32899 ;
  assign y10999 = ~1'b0 ;
  assign y11000 = n32901 ;
  assign y11001 = n32904 ;
  assign y11002 = ~1'b0 ;
  assign y11003 = n32906 ;
  assign y11004 = n32911 ;
  assign y11005 = n32912 ;
  assign y11006 = n25592 ;
  assign y11007 = ~n32914 ;
  assign y11008 = ~n32916 ;
  assign y11009 = ~n32920 ;
  assign y11010 = n32925 ;
  assign y11011 = n32928 ;
  assign y11012 = ~1'b0 ;
  assign y11013 = ~1'b0 ;
  assign y11014 = ~n32936 ;
  assign y11015 = ~n32937 ;
  assign y11016 = n24197 ;
  assign y11017 = ~n32940 ;
  assign y11018 = n32942 ;
  assign y11019 = n32944 ;
  assign y11020 = ~1'b0 ;
  assign y11021 = n32950 ;
  assign y11022 = n32952 ;
  assign y11023 = n32954 ;
  assign y11024 = n32957 ;
  assign y11025 = ~n32959 ;
  assign y11026 = ~n32962 ;
  assign y11027 = ~1'b0 ;
  assign y11028 = ~1'b0 ;
  assign y11029 = n32964 ;
  assign y11030 = n32968 ;
  assign y11031 = ~n32970 ;
  assign y11032 = ~n32973 ;
  assign y11033 = ~1'b0 ;
  assign y11034 = ~1'b0 ;
  assign y11035 = ~n32976 ;
  assign y11036 = n32977 ;
  assign y11037 = n32979 ;
  assign y11038 = ~n32981 ;
  assign y11039 = n32983 ;
  assign y11040 = ~n32989 ;
  assign y11041 = ~1'b0 ;
  assign y11042 = n32993 ;
  assign y11043 = ~n32996 ;
  assign y11044 = ~n32998 ;
  assign y11045 = n32999 ;
  assign y11046 = n33001 ;
  assign y11047 = ~n33002 ;
  assign y11048 = ~n33003 ;
  assign y11049 = n33005 ;
  assign y11050 = n33006 ;
  assign y11051 = n33008 ;
  assign y11052 = n33009 ;
  assign y11053 = ~1'b0 ;
  assign y11054 = n33010 ;
  assign y11055 = ~n33011 ;
  assign y11056 = n33012 ;
  assign y11057 = ~1'b0 ;
  assign y11058 = ~n33014 ;
  assign y11059 = ~n33018 ;
  assign y11060 = n33020 ;
  assign y11061 = ~n33021 ;
  assign y11062 = n33022 ;
  assign y11063 = ~1'b0 ;
  assign y11064 = n33026 ;
  assign y11065 = ~n33028 ;
  assign y11066 = ~1'b0 ;
  assign y11067 = n33031 ;
  assign y11068 = n33035 ;
  assign y11069 = ~n33037 ;
  assign y11070 = ~n33038 ;
  assign y11071 = ~n33040 ;
  assign y11072 = n33046 ;
  assign y11073 = n33051 ;
  assign y11074 = ~n33053 ;
  assign y11075 = ~1'b0 ;
  assign y11076 = ~n33054 ;
  assign y11077 = n33055 ;
  assign y11078 = ~n23402 ;
  assign y11079 = n33058 ;
  assign y11080 = ~n33059 ;
  assign y11081 = ~1'b0 ;
  assign y11082 = n5394 ;
  assign y11083 = n33065 ;
  assign y11084 = n33066 ;
  assign y11085 = n33071 ;
  assign y11086 = ~1'b0 ;
  assign y11087 = ~n33077 ;
  assign y11088 = ~1'b0 ;
  assign y11089 = ~1'b0 ;
  assign y11090 = ~1'b0 ;
  assign y11091 = ~n33081 ;
  assign y11092 = ~n33082 ;
  assign y11093 = n33084 ;
  assign y11094 = n33085 ;
  assign y11095 = ~1'b0 ;
  assign y11096 = n33088 ;
  assign y11097 = ~n33090 ;
  assign y11098 = ~n33091 ;
  assign y11099 = n33094 ;
  assign y11100 = ~n33095 ;
  assign y11101 = ~1'b0 ;
  assign y11102 = ~n33097 ;
  assign y11103 = ~n33099 ;
  assign y11104 = ~1'b0 ;
  assign y11105 = ~n33102 ;
  assign y11106 = ~n33105 ;
  assign y11107 = ~n21387 ;
  assign y11108 = n33106 ;
  assign y11109 = ~n33107 ;
  assign y11110 = n33109 ;
  assign y11111 = ~n33111 ;
  assign y11112 = ~n33113 ;
  assign y11113 = ~n33119 ;
  assign y11114 = n33129 ;
  assign y11115 = n33135 ;
  assign y11116 = ~n33141 ;
  assign y11117 = ~1'b0 ;
  assign y11118 = ~n33143 ;
  assign y11119 = n33144 ;
  assign y11120 = ~1'b0 ;
  assign y11121 = n33146 ;
  assign y11122 = ~n33149 ;
  assign y11123 = ~n33151 ;
  assign y11124 = n33153 ;
  assign y11125 = ~n33154 ;
  assign y11126 = ~n33159 ;
  assign y11127 = n33161 ;
  assign y11128 = ~n17060 ;
  assign y11129 = ~n33162 ;
  assign y11130 = n33165 ;
  assign y11131 = n33169 ;
  assign y11132 = ~n33174 ;
  assign y11133 = n33176 ;
  assign y11134 = ~1'b0 ;
  assign y11135 = ~n33177 ;
  assign y11136 = n33178 ;
  assign y11137 = ~1'b0 ;
  assign y11138 = 1'b0 ;
  assign y11139 = ~1'b0 ;
  assign y11140 = ~n33180 ;
  assign y11141 = n33187 ;
  assign y11142 = n33190 ;
  assign y11143 = n33191 ;
  assign y11144 = ~n33192 ;
  assign y11145 = ~n33200 ;
  assign y11146 = ~n33207 ;
  assign y11147 = ~n33210 ;
  assign y11148 = n33212 ;
  assign y11149 = ~n33215 ;
  assign y11150 = ~n33222 ;
  assign y11151 = ~n33226 ;
  assign y11152 = ~n33227 ;
  assign y11153 = ~1'b0 ;
  assign y11154 = n33234 ;
  assign y11155 = ~1'b0 ;
  assign y11156 = n33238 ;
  assign y11157 = n33240 ;
  assign y11158 = ~n33244 ;
  assign y11159 = n33247 ;
  assign y11160 = ~n33251 ;
  assign y11161 = ~n33252 ;
  assign y11162 = n21300 ;
  assign y11163 = ~n33254 ;
  assign y11164 = ~n33255 ;
  assign y11165 = n33258 ;
  assign y11166 = ~n33260 ;
  assign y11167 = ~n33263 ;
  assign y11168 = ~1'b0 ;
  assign y11169 = n33264 ;
  assign y11170 = n33266 ;
  assign y11171 = ~n33269 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = ~n33274 ;
  assign y11174 = ~n33275 ;
  assign y11175 = ~n33276 ;
  assign y11176 = n33277 ;
  assign y11177 = n33280 ;
  assign y11178 = ~n33282 ;
  assign y11179 = n3100 ;
  assign y11180 = ~1'b0 ;
  assign y11181 = ~n33283 ;
  assign y11182 = n33285 ;
  assign y11183 = n33286 ;
  assign y11184 = n33287 ;
  assign y11185 = ~n33289 ;
  assign y11186 = ~1'b0 ;
  assign y11187 = ~n33291 ;
  assign y11188 = n33294 ;
  assign y11189 = n33295 ;
  assign y11190 = ~n33300 ;
  assign y11191 = n33309 ;
  assign y11192 = n33311 ;
  assign y11193 = ~1'b0 ;
  assign y11194 = n7349 ;
  assign y11195 = ~1'b0 ;
  assign y11196 = ~n33315 ;
  assign y11197 = ~1'b0 ;
  assign y11198 = n33317 ;
  assign y11199 = ~n33320 ;
  assign y11200 = ~n33321 ;
  assign y11201 = n33322 ;
  assign y11202 = ~n33324 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = ~1'b0 ;
  assign y11205 = ~n33329 ;
  assign y11206 = n33332 ;
  assign y11207 = n33333 ;
  assign y11208 = ~n33334 ;
  assign y11209 = ~1'b0 ;
  assign y11210 = n33336 ;
  assign y11211 = n33338 ;
  assign y11212 = n33345 ;
  assign y11213 = ~n33349 ;
  assign y11214 = ~n33353 ;
  assign y11215 = n33357 ;
  assign y11216 = n33362 ;
  assign y11217 = n33368 ;
  assign y11218 = ~n33373 ;
  assign y11219 = ~n33379 ;
  assign y11220 = n33384 ;
  assign y11221 = n33385 ;
  assign y11222 = ~n33387 ;
  assign y11223 = n33392 ;
  assign y11224 = ~n33393 ;
  assign y11225 = n33394 ;
  assign y11226 = ~n33396 ;
  assign y11227 = ~1'b0 ;
  assign y11228 = n33400 ;
  assign y11229 = ~n33402 ;
  assign y11230 = ~n33407 ;
  assign y11231 = ~n33409 ;
  assign y11232 = n27391 ;
  assign y11233 = ~1'b0 ;
  assign y11234 = ~1'b0 ;
  assign y11235 = ~n33411 ;
  assign y11236 = ~1'b0 ;
  assign y11237 = n3498 ;
  assign y11238 = ~n30543 ;
  assign y11239 = n33412 ;
  assign y11240 = ~n33413 ;
  assign y11241 = ~n33416 ;
  assign y11242 = ~n33417 ;
  assign y11243 = ~1'b0 ;
  assign y11244 = ~1'b0 ;
  assign y11245 = n33421 ;
  assign y11246 = ~n33422 ;
  assign y11247 = ~n14783 ;
  assign y11248 = n33429 ;
  assign y11249 = n33431 ;
  assign y11250 = n33432 ;
  assign y11251 = ~n33433 ;
  assign y11252 = ~n33435 ;
  assign y11253 = ~n10652 ;
  assign y11254 = n33437 ;
  assign y11255 = n30795 ;
  assign y11256 = n33438 ;
  assign y11257 = ~n33439 ;
  assign y11258 = n33441 ;
  assign y11259 = ~n33449 ;
  assign y11260 = ~n33451 ;
  assign y11261 = ~1'b0 ;
  assign y11262 = ~n33457 ;
  assign y11263 = n33458 ;
  assign y11264 = ~1'b0 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = ~1'b0 ;
  assign y11267 = ~1'b0 ;
  assign y11268 = ~n33464 ;
  assign y11269 = n33465 ;
  assign y11270 = ~1'b0 ;
  assign y11271 = n33481 ;
  assign y11272 = n33482 ;
  assign y11273 = n33489 ;
  assign y11274 = ~n33491 ;
  assign y11275 = n33494 ;
  assign y11276 = ~n33496 ;
  assign y11277 = ~n33497 ;
  assign y11278 = n33499 ;
  assign y11279 = n33501 ;
  assign y11280 = ~n33504 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~n33507 ;
  assign y11283 = ~n33510 ;
  assign y11284 = n33512 ;
  assign y11285 = n33515 ;
  assign y11286 = ~n31093 ;
  assign y11287 = ~1'b0 ;
  assign y11288 = ~n33517 ;
  assign y11289 = ~1'b0 ;
  assign y11290 = ~n33518 ;
  assign y11291 = ~n33520 ;
  assign y11292 = ~n33521 ;
  assign y11293 = ~1'b0 ;
  assign y11294 = n33522 ;
  assign y11295 = n33523 ;
  assign y11296 = ~n33528 ;
  assign y11297 = n33529 ;
  assign y11298 = n33532 ;
  assign y11299 = n33535 ;
  assign y11300 = n33536 ;
  assign y11301 = ~n33540 ;
  assign y11302 = n33549 ;
  assign y11303 = ~n33550 ;
  assign y11304 = ~n33551 ;
  assign y11305 = ~n33553 ;
  assign y11306 = n33555 ;
  assign y11307 = n33556 ;
  assign y11308 = n33557 ;
  assign y11309 = ~1'b0 ;
  assign y11310 = ~n6082 ;
  assign y11311 = ~n33560 ;
  assign y11312 = ~1'b0 ;
  assign y11313 = ~n33565 ;
  assign y11314 = ~n33567 ;
  assign y11315 = ~n33570 ;
  assign y11316 = ~n33571 ;
  assign y11317 = n33579 ;
  assign y11318 = ~1'b0 ;
  assign y11319 = n33580 ;
  assign y11320 = ~1'b0 ;
  assign y11321 = ~n33581 ;
  assign y11322 = ~n33583 ;
  assign y11323 = ~1'b0 ;
  assign y11324 = n33585 ;
  assign y11325 = n33590 ;
  assign y11326 = ~n33595 ;
  assign y11327 = ~n33600 ;
  assign y11328 = ~1'b0 ;
  assign y11329 = ~n33609 ;
  assign y11330 = ~n33610 ;
  assign y11331 = n33611 ;
  assign y11332 = ~n33616 ;
  assign y11333 = n33617 ;
  assign y11334 = n33618 ;
  assign y11335 = ~n33619 ;
  assign y11336 = ~1'b0 ;
  assign y11337 = ~n33621 ;
  assign y11338 = ~n33625 ;
  assign y11339 = ~1'b0 ;
  assign y11340 = ~n33627 ;
  assign y11341 = n33630 ;
  assign y11342 = ~n33631 ;
  assign y11343 = ~n33640 ;
  assign y11344 = ~1'b0 ;
  assign y11345 = ~n33646 ;
  assign y11346 = ~n33654 ;
  assign y11347 = n33657 ;
  assign y11348 = n33660 ;
  assign y11349 = n33665 ;
  assign y11350 = n33666 ;
  assign y11351 = n33671 ;
  assign y11352 = ~n33673 ;
  assign y11353 = n33678 ;
  assign y11354 = n33681 ;
  assign y11355 = n33685 ;
  assign y11356 = ~n33690 ;
  assign y11357 = ~n33691 ;
  assign y11358 = n33693 ;
  assign y11359 = n33697 ;
  assign y11360 = ~n33699 ;
  assign y11361 = n33707 ;
  assign y11362 = ~n33709 ;
  assign y11363 = n21241 ;
  assign y11364 = ~n33714 ;
  assign y11365 = ~n33716 ;
  assign y11366 = ~1'b0 ;
  assign y11367 = ~n33721 ;
  assign y11368 = n33722 ;
  assign y11369 = ~n33725 ;
  assign y11370 = n33727 ;
  assign y11371 = ~1'b0 ;
  assign y11372 = ~1'b0 ;
  assign y11373 = n33729 ;
  assign y11374 = ~n33731 ;
  assign y11375 = ~n33733 ;
  assign y11376 = n33736 ;
  assign y11377 = ~n5370 ;
  assign y11378 = ~n33737 ;
  assign y11379 = n33739 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = ~1'b0 ;
  assign y11382 = ~n33741 ;
  assign y11383 = ~n33744 ;
  assign y11384 = n33747 ;
  assign y11385 = 1'b0 ;
  assign y11386 = n33751 ;
  assign y11387 = ~n33755 ;
  assign y11388 = ~n33758 ;
  assign y11389 = n33759 ;
  assign y11390 = n33761 ;
  assign y11391 = ~1'b0 ;
  assign y11392 = ~1'b0 ;
  assign y11393 = n33765 ;
  assign y11394 = ~n33766 ;
  assign y11395 = ~n33769 ;
  assign y11396 = n33772 ;
  assign y11397 = n33779 ;
  assign y11398 = n33783 ;
  assign y11399 = ~n33785 ;
  assign y11400 = n33787 ;
  assign y11401 = n33791 ;
  assign y11402 = n33794 ;
  assign y11403 = ~n33795 ;
  assign y11404 = n33797 ;
  assign y11405 = ~1'b0 ;
  assign y11406 = ~n33804 ;
  assign y11407 = n33806 ;
  assign y11408 = ~1'b0 ;
  assign y11409 = n33808 ;
  assign y11410 = ~n33809 ;
  assign y11411 = ~n33813 ;
  assign y11412 = n33815 ;
  assign y11413 = ~n33817 ;
  assign y11414 = n33818 ;
  assign y11415 = ~n33819 ;
  assign y11416 = ~n33823 ;
  assign y11417 = n33829 ;
  assign y11418 = ~n259 ;
  assign y11419 = n19942 ;
  assign y11420 = ~1'b0 ;
  assign y11421 = ~n33833 ;
  assign y11422 = ~n33838 ;
  assign y11423 = ~n33841 ;
  assign y11424 = ~1'b0 ;
  assign y11425 = n33842 ;
  assign y11426 = ~1'b0 ;
  assign y11427 = n33845 ;
  assign y11428 = ~n33846 ;
  assign y11429 = ~n33851 ;
  assign y11430 = n33852 ;
  assign y11431 = n25460 ;
  assign y11432 = ~n33855 ;
  assign y11433 = ~n33858 ;
  assign y11434 = ~n33863 ;
  assign y11435 = ~1'b0 ;
  assign y11436 = n33867 ;
  assign y11437 = ~n33868 ;
  assign y11438 = ~1'b0 ;
  assign y11439 = ~1'b0 ;
  assign y11440 = ~n33870 ;
  assign y11441 = n33876 ;
  assign y11442 = ~n33878 ;
  assign y11443 = ~n33881 ;
  assign y11444 = ~n33882 ;
  assign y11445 = ~n33883 ;
  assign y11446 = ~n33886 ;
  assign y11447 = ~n33887 ;
  assign y11448 = ~n33890 ;
  assign y11449 = n33892 ;
  assign y11450 = ~n33900 ;
  assign y11451 = ~1'b0 ;
  assign y11452 = n33903 ;
  assign y11453 = ~n33905 ;
  assign y11454 = n33908 ;
  assign y11455 = n33911 ;
  assign y11456 = n33912 ;
  assign y11457 = ~n33916 ;
  assign y11458 = ~1'b0 ;
  assign y11459 = n33925 ;
  assign y11460 = n33926 ;
  assign y11461 = ~n33928 ;
  assign y11462 = ~n33930 ;
  assign y11463 = ~n33941 ;
  assign y11464 = ~n33946 ;
  assign y11465 = n33947 ;
  assign y11466 = ~n33949 ;
  assign y11467 = ~n33950 ;
  assign y11468 = n33952 ;
  assign y11469 = ~n33955 ;
  assign y11470 = ~n33956 ;
  assign y11471 = ~n33959 ;
  assign y11472 = n33961 ;
  assign y11473 = ~n33962 ;
  assign y11474 = ~n33964 ;
  assign y11475 = ~n33968 ;
  assign y11476 = n33974 ;
  assign y11477 = ~n33976 ;
  assign y11478 = ~n33977 ;
  assign y11479 = n33979 ;
  assign y11480 = n33980 ;
  assign y11481 = ~n33981 ;
  assign y11482 = n33983 ;
  assign y11483 = n33987 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = ~n33991 ;
  assign y11486 = ~n33999 ;
  assign y11487 = n34003 ;
  assign y11488 = n34004 ;
  assign y11489 = n34008 ;
  assign y11490 = 1'b0 ;
  assign y11491 = ~1'b0 ;
  assign y11492 = ~1'b0 ;
  assign y11493 = n9289 ;
  assign y11494 = ~n34012 ;
  assign y11495 = ~1'b0 ;
  assign y11496 = ~n34015 ;
  assign y11497 = ~n34016 ;
  assign y11498 = ~n34020 ;
  assign y11499 = n34024 ;
  assign y11500 = n34032 ;
  assign y11501 = ~n34035 ;
  assign y11502 = ~n34039 ;
  assign y11503 = n34042 ;
  assign y11504 = n34044 ;
  assign y11505 = ~n34045 ;
  assign y11506 = ~n34046 ;
  assign y11507 = ~n34049 ;
  assign y11508 = ~n34052 ;
  assign y11509 = n34054 ;
  assign y11510 = ~n34055 ;
  assign y11511 = ~n34057 ;
  assign y11512 = n34060 ;
  assign y11513 = n34061 ;
  assign y11514 = ~n34062 ;
  assign y11515 = n34063 ;
  assign y11516 = ~n34066 ;
  assign y11517 = n34068 ;
  assign y11518 = n34073 ;
  assign y11519 = n34075 ;
  assign y11520 = ~n34082 ;
  assign y11521 = n34083 ;
  assign y11522 = n34090 ;
  assign y11523 = n34098 ;
  assign y11524 = n34099 ;
  assign y11525 = n34100 ;
  assign y11526 = n4838 ;
  assign y11527 = ~n34102 ;
  assign y11528 = ~n34104 ;
  assign y11529 = n34107 ;
  assign y11530 = n34110 ;
  assign y11531 = ~n34113 ;
  assign y11532 = n34119 ;
  assign y11533 = n34120 ;
  assign y11534 = ~n34122 ;
  assign y11535 = ~n34123 ;
  assign y11536 = ~n34127 ;
  assign y11537 = ~n34134 ;
  assign y11538 = n34136 ;
  assign y11539 = n34138 ;
  assign y11540 = ~n34140 ;
  assign y11541 = ~n34141 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = n34142 ;
  assign y11544 = n34144 ;
  assign y11545 = ~n34148 ;
  assign y11546 = ~n34151 ;
  assign y11547 = n34152 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = n34156 ;
  assign y11550 = ~n34157 ;
  assign y11551 = n34158 ;
  assign y11552 = ~1'b0 ;
  assign y11553 = ~n34159 ;
  assign y11554 = n34163 ;
  assign y11555 = ~n34170 ;
  assign y11556 = n34171 ;
  assign y11557 = n20420 ;
  assign y11558 = ~n34172 ;
  assign y11559 = ~n34173 ;
  assign y11560 = ~n34174 ;
  assign y11561 = ~n34184 ;
  assign y11562 = n34186 ;
  assign y11563 = n34188 ;
  assign y11564 = ~n27523 ;
  assign y11565 = ~n34195 ;
  assign y11566 = n34196 ;
  assign y11567 = ~n34202 ;
  assign y11568 = ~n34203 ;
  assign y11569 = ~1'b0 ;
  assign y11570 = ~1'b0 ;
  assign y11571 = n34204 ;
  assign y11572 = ~1'b0 ;
  assign y11573 = ~1'b0 ;
  assign y11574 = n34208 ;
  assign y11575 = n34211 ;
  assign y11576 = ~n34212 ;
  assign y11577 = ~n34215 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~n34228 ;
  assign y11580 = n34230 ;
  assign y11581 = n34248 ;
  assign y11582 = ~n34252 ;
  assign y11583 = ~n34255 ;
  assign y11584 = n34258 ;
  assign y11585 = n34261 ;
  assign y11586 = ~n34263 ;
  assign y11587 = ~n34264 ;
  assign y11588 = ~n34267 ;
  assign y11589 = ~n34270 ;
  assign y11590 = ~1'b0 ;
  assign y11591 = ~n34274 ;
  assign y11592 = ~n34279 ;
  assign y11593 = n34280 ;
  assign y11594 = ~n34281 ;
  assign y11595 = ~n34284 ;
  assign y11596 = n34286 ;
  assign y11597 = ~1'b0 ;
  assign y11598 = ~n34297 ;
  assign y11599 = n34298 ;
  assign y11600 = ~1'b0 ;
  assign y11601 = ~n34299 ;
  assign y11602 = n2110 ;
  assign y11603 = ~n34303 ;
  assign y11604 = n34310 ;
  assign y11605 = ~1'b0 ;
  assign y11606 = ~1'b0 ;
  assign y11607 = ~n34311 ;
  assign y11608 = ~n34312 ;
  assign y11609 = ~n34317 ;
  assign y11610 = n34319 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = ~1'b0 ;
  assign y11613 = ~n34323 ;
  assign y11614 = ~1'b0 ;
  assign y11615 = n34326 ;
  assign y11616 = n34328 ;
  assign y11617 = ~n34330 ;
  assign y11618 = n34336 ;
  assign y11619 = n34337 ;
  assign y11620 = ~1'b0 ;
  assign y11621 = ~n34344 ;
  assign y11622 = n34345 ;
  assign y11623 = ~n34347 ;
  assign y11624 = ~1'b0 ;
  assign y11625 = n34352 ;
  assign y11626 = ~n34353 ;
  assign y11627 = n34360 ;
  assign y11628 = ~n34368 ;
  assign y11629 = n34369 ;
  assign y11630 = n34374 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = n34375 ;
  assign y11633 = n34377 ;
  assign y11634 = ~n34378 ;
  assign y11635 = n34383 ;
  assign y11636 = ~n34385 ;
  assign y11637 = ~n34387 ;
  assign y11638 = ~n34388 ;
  assign y11639 = n34393 ;
  assign y11640 = n34399 ;
  assign y11641 = ~n34401 ;
  assign y11642 = n34403 ;
  assign y11643 = ~1'b0 ;
  assign y11644 = ~1'b0 ;
  assign y11645 = ~n34405 ;
  assign y11646 = ~n34411 ;
  assign y11647 = n34414 ;
  assign y11648 = n34415 ;
  assign y11649 = n34417 ;
  assign y11650 = n34418 ;
  assign y11651 = n34420 ;
  assign y11652 = ~n34427 ;
  assign y11653 = ~n34429 ;
  assign y11654 = ~n34430 ;
  assign y11655 = n34441 ;
  assign y11656 = ~1'b0 ;
  assign y11657 = n34449 ;
  assign y11658 = ~1'b0 ;
  assign y11659 = n34450 ;
  assign y11660 = ~n34454 ;
  assign y11661 = ~n34459 ;
  assign y11662 = ~n34460 ;
  assign y11663 = n34466 ;
  assign y11664 = ~1'b0 ;
  assign y11665 = n30217 ;
  assign y11666 = ~n34470 ;
  assign y11667 = ~n34472 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = n34479 ;
  assign y11670 = ~1'b0 ;
  assign y11671 = n34481 ;
  assign y11672 = n34482 ;
  assign y11673 = ~n34487 ;
  assign y11674 = ~n34489 ;
  assign y11675 = ~n34495 ;
  assign y11676 = n34497 ;
  assign y11677 = ~n2461 ;
  assign y11678 = n34500 ;
  assign y11679 = n34503 ;
  assign y11680 = ~1'b0 ;
  assign y11681 = n34505 ;
  assign y11682 = ~1'b0 ;
  assign y11683 = n34507 ;
  assign y11684 = ~1'b0 ;
  assign y11685 = ~n34513 ;
  assign y11686 = ~n34514 ;
  assign y11687 = n21736 ;
  assign y11688 = n34518 ;
  assign y11689 = ~n34520 ;
  assign y11690 = ~n34523 ;
  assign y11691 = ~n34527 ;
  assign y11692 = n34536 ;
  assign y11693 = ~n34539 ;
  assign y11694 = n34541 ;
  assign y11695 = n34543 ;
  assign y11696 = ~n34545 ;
  assign y11697 = ~n34546 ;
  assign y11698 = n34547 ;
  assign y11699 = n34548 ;
  assign y11700 = 1'b0 ;
  assign y11701 = n34550 ;
  assign y11702 = n34555 ;
  assign y11703 = ~1'b0 ;
  assign y11704 = ~n34561 ;
  assign y11705 = n34562 ;
  assign y11706 = ~n34563 ;
  assign y11707 = ~n34565 ;
  assign y11708 = ~1'b0 ;
  assign y11709 = ~n34569 ;
  assign y11710 = n34570 ;
  assign y11711 = ~n34572 ;
  assign y11712 = n34573 ;
  assign y11713 = n34577 ;
  assign y11714 = ~n34581 ;
  assign y11715 = ~n34583 ;
  assign y11716 = ~n34585 ;
  assign y11717 = ~n34588 ;
  assign y11718 = n34591 ;
  assign y11719 = n34593 ;
  assign y11720 = ~1'b0 ;
  assign y11721 = n34597 ;
  assign y11722 = n34602 ;
  assign y11723 = ~n34603 ;
  assign y11724 = n34606 ;
  assign y11725 = n34607 ;
  assign y11726 = 1'b0 ;
  assign y11727 = ~1'b0 ;
  assign y11728 = ~1'b0 ;
  assign y11729 = n34609 ;
  assign y11730 = n34622 ;
  assign y11731 = ~n34629 ;
  assign y11732 = n34631 ;
  assign y11733 = n34636 ;
  assign y11734 = n34638 ;
  assign y11735 = n34639 ;
  assign y11736 = ~1'b0 ;
  assign y11737 = ~n34644 ;
  assign y11738 = ~n34649 ;
  assign y11739 = n34651 ;
  assign y11740 = n34655 ;
  assign y11741 = ~1'b0 ;
  assign y11742 = ~n34656 ;
  assign y11743 = ~n34657 ;
  assign y11744 = ~1'b0 ;
  assign y11745 = ~n3175 ;
  assign y11746 = ~n34658 ;
  assign y11747 = ~n34661 ;
  assign y11748 = n34662 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = ~n34664 ;
  assign y11751 = n34665 ;
  assign y11752 = ~1'b0 ;
  assign y11753 = ~n34667 ;
  assign y11754 = ~n34668 ;
  assign y11755 = ~1'b0 ;
  assign y11756 = n18214 ;
  assign y11757 = ~1'b0 ;
  assign y11758 = ~n34671 ;
  assign y11759 = ~n1475 ;
  assign y11760 = n34672 ;
  assign y11761 = ~1'b0 ;
  assign y11762 = n34674 ;
  assign y11763 = ~n34678 ;
  assign y11764 = n34680 ;
  assign y11765 = ~1'b0 ;
  assign y11766 = n34682 ;
  assign y11767 = n34684 ;
  assign y11768 = n34692 ;
  assign y11769 = n34695 ;
  assign y11770 = ~n34697 ;
  assign y11771 = n34699 ;
  assign y11772 = 1'b0 ;
  assign y11773 = n34704 ;
  assign y11774 = n34707 ;
  assign y11775 = n34708 ;
  assign y11776 = n34714 ;
  assign y11777 = ~1'b0 ;
  assign y11778 = n34715 ;
  assign y11779 = ~n34716 ;
  assign y11780 = ~n34717 ;
  assign y11781 = n34718 ;
  assign y11782 = n34721 ;
  assign y11783 = n34722 ;
  assign y11784 = ~n34725 ;
  assign y11785 = ~n34727 ;
  assign y11786 = n34735 ;
  assign y11787 = n34737 ;
  assign y11788 = ~n34739 ;
  assign y11789 = n34740 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = n34745 ;
  assign y11792 = ~n34746 ;
  assign y11793 = ~n34752 ;
  assign y11794 = n34755 ;
  assign y11795 = ~1'b0 ;
  assign y11796 = n34761 ;
  assign y11797 = n34765 ;
  assign y11798 = n34767 ;
  assign y11799 = ~1'b0 ;
  assign y11800 = ~n34769 ;
  assign y11801 = ~1'b0 ;
  assign y11802 = n34770 ;
  assign y11803 = n34772 ;
  assign y11804 = ~n34775 ;
  assign y11805 = n34776 ;
  assign y11806 = n34781 ;
  assign y11807 = n34784 ;
  assign y11808 = ~1'b0 ;
  assign y11809 = ~n34785 ;
  assign y11810 = n34786 ;
  assign y11811 = ~n34787 ;
  assign y11812 = n34792 ;
  assign y11813 = ~n34796 ;
  assign y11814 = ~1'b0 ;
  assign y11815 = ~1'b0 ;
  assign y11816 = ~1'b0 ;
  assign y11817 = n34798 ;
  assign y11818 = ~n34799 ;
  assign y11819 = n34800 ;
  assign y11820 = ~n34801 ;
  assign y11821 = ~n34802 ;
  assign y11822 = n34804 ;
  assign y11823 = ~n34805 ;
  assign y11824 = n34807 ;
  assign y11825 = n34809 ;
  assign y11826 = n34821 ;
  assign y11827 = ~n34822 ;
  assign y11828 = ~n34823 ;
  assign y11829 = ~1'b0 ;
  assign y11830 = n34827 ;
  assign y11831 = ~n34830 ;
  assign y11832 = n34835 ;
  assign y11833 = n34836 ;
  assign y11834 = n34848 ;
  assign y11835 = n34855 ;
  assign y11836 = n34856 ;
  assign y11837 = ~n34857 ;
  assign y11838 = ~1'b0 ;
  assign y11839 = ~n34860 ;
  assign y11840 = ~n34865 ;
  assign y11841 = ~n34869 ;
  assign y11842 = ~n34872 ;
  assign y11843 = ~n34877 ;
  assign y11844 = n34881 ;
  assign y11845 = ~1'b0 ;
  assign y11846 = n34884 ;
  assign y11847 = ~n34885 ;
  assign y11848 = ~n34888 ;
  assign y11849 = n34891 ;
  assign y11850 = n34893 ;
  assign y11851 = n34896 ;
  assign y11852 = ~1'b0 ;
  assign y11853 = ~1'b0 ;
  assign y11854 = ~n34899 ;
  assign y11855 = ~n34905 ;
  assign y11856 = n34906 ;
  assign y11857 = n34916 ;
  assign y11858 = ~n34918 ;
  assign y11859 = n34920 ;
  assign y11860 = ~n34922 ;
  assign y11861 = n34924 ;
  assign y11862 = ~n34927 ;
  assign y11863 = ~n34929 ;
  assign y11864 = n34933 ;
  assign y11865 = ~n34934 ;
  assign y11866 = ~1'b0 ;
  assign y11867 = n34941 ;
  assign y11868 = ~n34945 ;
  assign y11869 = ~n34947 ;
  assign y11870 = ~n34951 ;
  assign y11871 = ~1'b0 ;
  assign y11872 = ~1'b0 ;
  assign y11873 = ~n34953 ;
  assign y11874 = n34954 ;
  assign y11875 = ~n34955 ;
  assign y11876 = n34956 ;
  assign y11877 = n34959 ;
  assign y11878 = ~1'b0 ;
  assign y11879 = ~1'b0 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = ~1'b0 ;
  assign y11882 = ~1'b0 ;
  assign y11883 = n34962 ;
  assign y11884 = ~n34963 ;
  assign y11885 = n34964 ;
  assign y11886 = ~n22061 ;
  assign y11887 = n34968 ;
  assign y11888 = n34974 ;
  assign y11889 = ~1'b0 ;
  assign y11890 = ~1'b0 ;
  assign y11891 = ~n34975 ;
  assign y11892 = ~n34978 ;
  assign y11893 = ~n34984 ;
  assign y11894 = ~n34997 ;
  assign y11895 = ~1'b0 ;
  assign y11896 = n34999 ;
  assign y11897 = n35010 ;
  assign y11898 = ~n35012 ;
  assign y11899 = ~n35016 ;
  assign y11900 = ~1'b0 ;
  assign y11901 = n35018 ;
  assign y11902 = ~n35023 ;
  assign y11903 = ~n35024 ;
  assign y11904 = ~n35030 ;
  assign y11905 = n35031 ;
  assign y11906 = ~n35032 ;
  assign y11907 = n35034 ;
  assign y11908 = ~n35036 ;
  assign y11909 = n35039 ;
  assign y11910 = ~1'b0 ;
  assign y11911 = ~n35040 ;
  assign y11912 = n21408 ;
  assign y11913 = n35042 ;
  assign y11914 = n35045 ;
  assign y11915 = n35046 ;
  assign y11916 = ~n35051 ;
  assign y11917 = ~n35052 ;
  assign y11918 = n35057 ;
  assign y11919 = ~n35061 ;
  assign y11920 = n35063 ;
  assign y11921 = n35065 ;
  assign y11922 = n35068 ;
  assign y11923 = ~n35071 ;
  assign y11924 = n35075 ;
  assign y11925 = n35078 ;
  assign y11926 = ~n35084 ;
  assign y11927 = n35085 ;
  assign y11928 = n35086 ;
  assign y11929 = ~n35087 ;
  assign y11930 = ~1'b0 ;
  assign y11931 = ~1'b0 ;
  assign y11932 = ~n8245 ;
  assign y11933 = ~n35091 ;
  assign y11934 = ~n35098 ;
  assign y11935 = n35102 ;
  assign y11936 = n35104 ;
  assign y11937 = n35107 ;
  assign y11938 = ~n35110 ;
  assign y11939 = ~1'b0 ;
  assign y11940 = ~1'b0 ;
  assign y11941 = n35111 ;
  assign y11942 = n15520 ;
  assign y11943 = n35116 ;
  assign y11944 = ~n35120 ;
  assign y11945 = n35126 ;
  assign y11946 = n35130 ;
  assign y11947 = ~n35131 ;
  assign y11948 = ~n35136 ;
  assign y11949 = n35144 ;
  assign y11950 = ~n35146 ;
  assign y11951 = ~n35153 ;
  assign y11952 = ~1'b0 ;
  assign y11953 = ~n35164 ;
  assign y11954 = ~n35165 ;
  assign y11955 = n35166 ;
  assign y11956 = n35169 ;
  assign y11957 = ~n35170 ;
  assign y11958 = ~n35177 ;
  assign y11959 = n35179 ;
  assign y11960 = n35184 ;
  assign y11961 = ~n35186 ;
  assign y11962 = n28403 ;
  assign y11963 = n35188 ;
  assign y11964 = n35191 ;
  assign y11965 = ~1'b0 ;
  assign y11966 = ~1'b0 ;
  assign y11967 = ~n35192 ;
  assign y11968 = n35193 ;
  assign y11969 = ~n35194 ;
  assign y11970 = ~n35198 ;
  assign y11971 = n35201 ;
  assign y11972 = n35203 ;
  assign y11973 = ~n35206 ;
  assign y11974 = ~1'b0 ;
  assign y11975 = n4653 ;
  assign y11976 = ~1'b0 ;
  assign y11977 = ~n35207 ;
  assign y11978 = ~n35208 ;
  assign y11979 = ~n35211 ;
  assign y11980 = ~1'b0 ;
  assign y11981 = ~n35212 ;
  assign y11982 = ~n35217 ;
  assign y11983 = ~n35220 ;
  assign y11984 = ~n35226 ;
  assign y11985 = ~n35228 ;
  assign y11986 = n35230 ;
  assign y11987 = n35233 ;
  assign y11988 = ~1'b0 ;
  assign y11989 = n35238 ;
  assign y11990 = ~n35239 ;
  assign y11991 = ~n35241 ;
  assign y11992 = n35245 ;
  assign y11993 = ~n35251 ;
  assign y11994 = n17284 ;
  assign y11995 = ~n35257 ;
  assign y11996 = n35259 ;
  assign y11997 = ~n35262 ;
  assign y11998 = n35263 ;
  assign y11999 = n35269 ;
  assign y12000 = ~n35271 ;
  assign y12001 = n35273 ;
  assign y12002 = n35278 ;
  assign y12003 = n35284 ;
  assign y12004 = ~n35286 ;
  assign y12005 = n35287 ;
  assign y12006 = n35289 ;
  assign y12007 = ~n35293 ;
  assign y12008 = ~n35295 ;
  assign y12009 = ~1'b0 ;
  assign y12010 = n35296 ;
  assign y12011 = ~n35305 ;
  assign y12012 = n32714 ;
  assign y12013 = n35310 ;
  assign y12014 = n615 ;
  assign y12015 = n35314 ;
  assign y12016 = n35315 ;
  assign y12017 = ~n35318 ;
  assign y12018 = ~n35319 ;
  assign y12019 = ~n35320 ;
  assign y12020 = n35321 ;
  assign y12021 = ~n35324 ;
  assign y12022 = ~n35326 ;
  assign y12023 = n35330 ;
  assign y12024 = ~n35331 ;
  assign y12025 = n35333 ;
  assign y12026 = n35335 ;
  assign y12027 = ~n35336 ;
  assign y12028 = ~n35337 ;
  assign y12029 = ~n35339 ;
  assign y12030 = n35340 ;
  assign y12031 = ~1'b0 ;
  assign y12032 = ~n35345 ;
  assign y12033 = ~n35349 ;
  assign y12034 = ~n35350 ;
  assign y12035 = n35351 ;
  assign y12036 = n35356 ;
  assign y12037 = ~n35357 ;
  assign y12038 = ~1'b0 ;
  assign y12039 = n35360 ;
  assign y12040 = ~1'b0 ;
  assign y12041 = n35363 ;
  assign y12042 = ~1'b0 ;
  assign y12043 = n35369 ;
  assign y12044 = ~n35370 ;
  assign y12045 = ~n35371 ;
  assign y12046 = ~1'b0 ;
  assign y12047 = ~n35372 ;
  assign y12048 = ~1'b0 ;
  assign y12049 = n35378 ;
  assign y12050 = n35379 ;
  assign y12051 = n35381 ;
  assign y12052 = ~n35383 ;
  assign y12053 = ~1'b0 ;
  assign y12054 = ~1'b0 ;
  assign y12055 = ~n35386 ;
  assign y12056 = ~n35389 ;
  assign y12057 = ~n35390 ;
  assign y12058 = ~n35391 ;
  assign y12059 = ~n35397 ;
  assign y12060 = ~n35399 ;
  assign y12061 = n35401 ;
  assign y12062 = ~n35404 ;
  assign y12063 = ~n35408 ;
  assign y12064 = ~n35411 ;
  assign y12065 = ~n35412 ;
  assign y12066 = n35416 ;
  assign y12067 = n35418 ;
  assign y12068 = n35422 ;
  assign y12069 = ~n35423 ;
  assign y12070 = ~n35427 ;
  assign y12071 = n35431 ;
  assign y12072 = ~1'b0 ;
  assign y12073 = ~n35434 ;
  assign y12074 = n35442 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = ~1'b0 ;
  assign y12077 = ~n35446 ;
  assign y12078 = n35449 ;
  assign y12079 = n18397 ;
  assign y12080 = 1'b0 ;
  assign y12081 = n35452 ;
  assign y12082 = ~n35454 ;
  assign y12083 = n35456 ;
  assign y12084 = ~n35457 ;
  assign y12085 = ~n35462 ;
  assign y12086 = ~n35463 ;
  assign y12087 = ~n35464 ;
  assign y12088 = ~1'b0 ;
  assign y12089 = ~n35467 ;
  assign y12090 = ~n35469 ;
  assign y12091 = n35471 ;
  assign y12092 = n35473 ;
  assign y12093 = n35477 ;
  assign y12094 = ~n35478 ;
  assign y12095 = ~n35479 ;
  assign y12096 = n735 ;
  assign y12097 = n35480 ;
  assign y12098 = n35481 ;
  assign y12099 = ~n35484 ;
  assign y12100 = n35486 ;
  assign y12101 = ~n35491 ;
  assign y12102 = ~n35494 ;
  assign y12103 = ~n35498 ;
  assign y12104 = ~n35499 ;
  assign y12105 = ~n35506 ;
  assign y12106 = ~1'b0 ;
  assign y12107 = ~1'b0 ;
  assign y12108 = ~1'b0 ;
  assign y12109 = n35515 ;
  assign y12110 = ~n35516 ;
  assign y12111 = ~n35517 ;
  assign y12112 = ~n35518 ;
  assign y12113 = n35530 ;
  assign y12114 = n35538 ;
  assign y12115 = ~1'b0 ;
  assign y12116 = ~1'b0 ;
  assign y12117 = ~n35544 ;
  assign y12118 = ~n35547 ;
  assign y12119 = ~n35554 ;
  assign y12120 = n35557 ;
  assign y12121 = n35558 ;
  assign y12122 = n35559 ;
  assign y12123 = n35561 ;
  assign y12124 = ~n35563 ;
  assign y12125 = ~n12446 ;
  assign y12126 = ~n35566 ;
  assign y12127 = ~n3837 ;
  assign y12128 = n35570 ;
  assign y12129 = n35574 ;
  assign y12130 = n35576 ;
  assign y12131 = ~n35578 ;
  assign y12132 = ~n35579 ;
  assign y12133 = ~1'b0 ;
  assign y12134 = ~n35584 ;
  assign y12135 = n35587 ;
  assign y12136 = ~n35590 ;
  assign y12137 = ~1'b0 ;
  assign y12138 = ~n35591 ;
  assign y12139 = ~n35596 ;
  assign y12140 = n35599 ;
  assign y12141 = ~n35601 ;
  assign y12142 = n35602 ;
  assign y12143 = n35606 ;
  assign y12144 = ~1'b0 ;
  assign y12145 = ~n35609 ;
  assign y12146 = ~n35610 ;
  assign y12147 = n35612 ;
  assign y12148 = n35619 ;
  assign y12149 = ~n35621 ;
  assign y12150 = n35622 ;
  assign y12151 = ~n35623 ;
  assign y12152 = ~n35626 ;
  assign y12153 = ~n35628 ;
  assign y12154 = ~n35629 ;
  assign y12155 = n35634 ;
  assign y12156 = ~1'b0 ;
  assign y12157 = ~n35638 ;
  assign y12158 = ~n35639 ;
  assign y12159 = ~n35641 ;
  assign y12160 = ~n35644 ;
  assign y12161 = n35645 ;
  assign y12162 = ~n35647 ;
  assign y12163 = ~n35650 ;
  assign y12164 = n35653 ;
  assign y12165 = n35655 ;
  assign y12166 = n9060 ;
  assign y12167 = ~n35660 ;
  assign y12168 = ~n2761 ;
  assign y12169 = ~1'b0 ;
  assign y12170 = ~1'b0 ;
  assign y12171 = n35666 ;
  assign y12172 = n35667 ;
  assign y12173 = n35679 ;
  assign y12174 = n1787 ;
  assign y12175 = ~n35680 ;
  assign y12176 = ~n35685 ;
  assign y12177 = ~n35696 ;
  assign y12178 = n35699 ;
  assign y12179 = n35700 ;
  assign y12180 = n35703 ;
  assign y12181 = ~n35709 ;
  assign y12182 = n35714 ;
  assign y12183 = ~1'b0 ;
  assign y12184 = ~1'b0 ;
  assign y12185 = n35719 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = n35721 ;
  assign y12188 = n35722 ;
  assign y12189 = ~n35729 ;
  assign y12190 = n17176 ;
  assign y12191 = ~n35730 ;
  assign y12192 = n35733 ;
  assign y12193 = ~1'b0 ;
  assign y12194 = ~n35735 ;
  assign y12195 = ~n35737 ;
  assign y12196 = ~n35741 ;
  assign y12197 = n35750 ;
  assign y12198 = ~n35753 ;
  assign y12199 = n35755 ;
  assign y12200 = ~1'b0 ;
  assign y12201 = ~n35757 ;
  assign y12202 = n35759 ;
  assign y12203 = ~n35760 ;
  assign y12204 = ~n35761 ;
  assign y12205 = n35762 ;
  assign y12206 = ~n35764 ;
  assign y12207 = ~1'b0 ;
  assign y12208 = ~1'b0 ;
  assign y12209 = n35765 ;
  assign y12210 = ~n35767 ;
  assign y12211 = ~1'b0 ;
  assign y12212 = n35769 ;
  assign y12213 = ~n35774 ;
  assign y12214 = ~n35776 ;
  assign y12215 = ~n18320 ;
  assign y12216 = n35781 ;
  assign y12217 = ~n35782 ;
  assign y12218 = ~n35784 ;
  assign y12219 = n35790 ;
  assign y12220 = ~n33570 ;
  assign y12221 = n35791 ;
  assign y12222 = n35792 ;
  assign y12223 = n35793 ;
  assign y12224 = n6330 ;
  assign y12225 = 1'b0 ;
  assign y12226 = n35795 ;
  assign y12227 = ~n35798 ;
  assign y12228 = ~1'b0 ;
  assign y12229 = ~n35802 ;
  assign y12230 = n35803 ;
  assign y12231 = n35804 ;
  assign y12232 = ~1'b0 ;
  assign y12233 = n35806 ;
  assign y12234 = ~n35808 ;
  assign y12235 = ~1'b0 ;
  assign y12236 = n35811 ;
  assign y12237 = ~n35814 ;
  assign y12238 = ~n35817 ;
  assign y12239 = n35818 ;
  assign y12240 = ~1'b0 ;
  assign y12241 = ~n35823 ;
  assign y12242 = n35825 ;
  assign y12243 = n35827 ;
  assign y12244 = ~n35828 ;
  assign y12245 = n35832 ;
  assign y12246 = n11048 ;
  assign y12247 = n35834 ;
  assign y12248 = ~n35839 ;
  assign y12249 = n35840 ;
  assign y12250 = n35844 ;
  assign y12251 = ~n35845 ;
  assign y12252 = n35848 ;
  assign y12253 = ~1'b0 ;
  assign y12254 = ~n35851 ;
  assign y12255 = n35852 ;
  assign y12256 = n35860 ;
  assign y12257 = ~1'b0 ;
  assign y12258 = ~n35867 ;
  assign y12259 = ~1'b0 ;
  assign y12260 = ~n35871 ;
  assign y12261 = ~n35872 ;
  assign y12262 = n35873 ;
  assign y12263 = ~1'b0 ;
  assign y12264 = n35878 ;
  assign y12265 = ~n35879 ;
  assign y12266 = ~n35884 ;
  assign y12267 = n35886 ;
  assign y12268 = n35887 ;
  assign y12269 = ~n35889 ;
  assign y12270 = n35890 ;
  assign y12271 = n35891 ;
  assign y12272 = n35895 ;
  assign y12273 = n35905 ;
  assign y12274 = ~n18901 ;
  assign y12275 = ~n35909 ;
  assign y12276 = n35910 ;
  assign y12277 = n35915 ;
  assign y12278 = ~n35918 ;
  assign y12279 = n35924 ;
  assign y12280 = 1'b0 ;
  assign y12281 = ~n35925 ;
  assign y12282 = n35926 ;
  assign y12283 = ~1'b0 ;
  assign y12284 = ~1'b0 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = n35929 ;
  assign y12287 = ~n35932 ;
  assign y12288 = ~n35942 ;
  assign y12289 = n35947 ;
  assign y12290 = ~1'b0 ;
  assign y12291 = ~n35951 ;
  assign y12292 = ~n35952 ;
  assign y12293 = ~n35953 ;
  assign y12294 = ~n35956 ;
  assign y12295 = ~n35961 ;
  assign y12296 = ~1'b0 ;
  assign y12297 = ~1'b0 ;
  assign y12298 = n35962 ;
  assign y12299 = ~n35963 ;
  assign y12300 = n35965 ;
  assign y12301 = n35968 ;
  assign y12302 = ~n35970 ;
  assign y12303 = n35971 ;
  assign y12304 = ~n9825 ;
  assign y12305 = ~n35976 ;
  assign y12306 = ~1'b0 ;
  assign y12307 = ~1'b0 ;
  assign y12308 = ~n35978 ;
  assign y12309 = ~n35983 ;
  assign y12310 = ~n35984 ;
  assign y12311 = n35986 ;
  assign y12312 = ~n35988 ;
  assign y12313 = ~n35995 ;
  assign y12314 = n35996 ;
  assign y12315 = n35998 ;
  assign y12316 = n36000 ;
  assign y12317 = ~1'b0 ;
  assign y12318 = n36002 ;
  assign y12319 = n36004 ;
  assign y12320 = ~n36005 ;
  assign y12321 = ~n36008 ;
  assign y12322 = n36011 ;
  assign y12323 = n36014 ;
  assign y12324 = n36018 ;
  assign y12325 = ~n36020 ;
  assign y12326 = ~1'b0 ;
  assign y12327 = n36028 ;
  assign y12328 = ~n36031 ;
  assign y12329 = n36038 ;
  assign y12330 = ~n36039 ;
  assign y12331 = n36042 ;
  assign y12332 = ~n36044 ;
  assign y12333 = ~1'b0 ;
  assign y12334 = ~n36046 ;
  assign y12335 = ~n36052 ;
  assign y12336 = ~n36053 ;
  assign y12337 = ~n36054 ;
  assign y12338 = ~n14607 ;
  assign y12339 = n36058 ;
  assign y12340 = ~1'b0 ;
  assign y12341 = ~n36063 ;
  assign y12342 = ~n36064 ;
  assign y12343 = n36068 ;
  assign y12344 = ~n36072 ;
  assign y12345 = n36084 ;
  assign y12346 = ~1'b0 ;
  assign y12347 = n36087 ;
  assign y12348 = n36088 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = n36090 ;
  assign y12351 = n36091 ;
  assign y12352 = n29175 ;
  assign y12353 = n36092 ;
  assign y12354 = ~n36093 ;
  assign y12355 = n36094 ;
  assign y12356 = n36098 ;
  assign y12357 = n36100 ;
  assign y12358 = 1'b0 ;
  assign y12359 = ~1'b0 ;
  assign y12360 = ~1'b0 ;
  assign y12361 = ~1'b0 ;
  assign y12362 = n36104 ;
  assign y12363 = n36105 ;
  assign y12364 = n36106 ;
  assign y12365 = n36109 ;
  assign y12366 = n36111 ;
  assign y12367 = ~n36113 ;
  assign y12368 = ~n36118 ;
  assign y12369 = ~n36122 ;
  assign y12370 = n36124 ;
  assign y12371 = n36125 ;
  assign y12372 = ~1'b0 ;
  assign y12373 = n36127 ;
  assign y12374 = ~n36129 ;
  assign y12375 = n36132 ;
  assign y12376 = ~n36134 ;
  assign y12377 = n36136 ;
  assign y12378 = ~n36137 ;
  assign y12379 = ~n36138 ;
  assign y12380 = n36141 ;
  assign y12381 = ~n36145 ;
  assign y12382 = ~n36147 ;
  assign y12383 = n36149 ;
  assign y12384 = n36150 ;
  assign y12385 = n36152 ;
  assign y12386 = n36154 ;
  assign y12387 = ~1'b0 ;
  assign y12388 = n36158 ;
  assign y12389 = ~n36160 ;
  assign y12390 = n36161 ;
  assign y12391 = ~n36162 ;
  assign y12392 = ~n36165 ;
  assign y12393 = ~n36170 ;
  assign y12394 = ~n36172 ;
  assign y12395 = ~n36175 ;
  assign y12396 = ~n36179 ;
  assign y12397 = ~n36182 ;
  assign y12398 = ~n36183 ;
  assign y12399 = ~1'b0 ;
  assign y12400 = ~n36186 ;
  assign y12401 = ~n36188 ;
  assign y12402 = n36191 ;
  assign y12403 = n36199 ;
  assign y12404 = ~n36207 ;
  assign y12405 = ~n36213 ;
  assign y12406 = ~n36214 ;
  assign y12407 = ~n36217 ;
  assign y12408 = n36222 ;
  assign y12409 = ~n36226 ;
  assign y12410 = ~1'b0 ;
  assign y12411 = n36228 ;
  assign y12412 = ~n36231 ;
  assign y12413 = ~n36233 ;
  assign y12414 = ~1'b0 ;
  assign y12415 = ~1'b0 ;
  assign y12416 = n36236 ;
  assign y12417 = n36237 ;
  assign y12418 = n36241 ;
  assign y12419 = ~n36246 ;
  assign y12420 = n36248 ;
  assign y12421 = ~n36249 ;
  assign y12422 = ~n36250 ;
  assign y12423 = ~n36251 ;
  assign y12424 = n36252 ;
  assign y12425 = ~n36256 ;
  assign y12426 = n36257 ;
  assign y12427 = n36259 ;
  assign y12428 = ~n36262 ;
  assign y12429 = ~n36265 ;
  assign y12430 = ~n36266 ;
  assign y12431 = ~n36269 ;
  assign y12432 = ~n36270 ;
  assign y12433 = ~n36271 ;
  assign y12434 = ~n36273 ;
  assign y12435 = ~n36276 ;
  assign y12436 = ~n36280 ;
  assign y12437 = ~n36282 ;
  assign y12438 = n36283 ;
  assign y12439 = ~n36285 ;
  assign y12440 = ~n36288 ;
  assign y12441 = ~1'b0 ;
  assign y12442 = n36289 ;
  assign y12443 = ~1'b0 ;
  assign y12444 = ~n36292 ;
  assign y12445 = n36294 ;
  assign y12446 = ~1'b0 ;
  assign y12447 = n36295 ;
  assign y12448 = ~n36299 ;
  assign y12449 = ~n36303 ;
  assign y12450 = ~n36305 ;
  assign y12451 = ~n7085 ;
  assign y12452 = ~n36306 ;
  assign y12453 = n36308 ;
  assign y12454 = ~n36309 ;
  assign y12455 = ~1'b0 ;
  assign y12456 = n36310 ;
  assign y12457 = n36311 ;
  assign y12458 = n36315 ;
  assign y12459 = n36317 ;
  assign y12460 = ~1'b0 ;
  assign y12461 = n36319 ;
  assign y12462 = ~n36323 ;
  assign y12463 = ~n36324 ;
  assign y12464 = n36329 ;
  assign y12465 = ~n36332 ;
  assign y12466 = n36333 ;
  assign y12467 = ~n36334 ;
  assign y12468 = ~n36337 ;
  assign y12469 = ~n36339 ;
  assign y12470 = ~n36341 ;
  assign y12471 = n36349 ;
  assign y12472 = ~n3441 ;
  assign y12473 = ~n36351 ;
  assign y12474 = ~n36357 ;
  assign y12475 = ~n36358 ;
  assign y12476 = n36365 ;
  assign y12477 = n36367 ;
  assign y12478 = ~n36372 ;
  assign y12479 = n36375 ;
  assign y12480 = n36377 ;
  assign y12481 = ~n36378 ;
  assign y12482 = ~n36379 ;
  assign y12483 = ~n12135 ;
  assign y12484 = ~1'b0 ;
  assign y12485 = ~n36380 ;
  assign y12486 = ~n36383 ;
  assign y12487 = ~n36387 ;
  assign y12488 = n36389 ;
  assign y12489 = ~1'b0 ;
  assign y12490 = n36393 ;
  assign y12491 = ~1'b0 ;
  assign y12492 = ~n36394 ;
  assign y12493 = ~n36399 ;
  assign y12494 = ~n36401 ;
  assign y12495 = ~1'b0 ;
  assign y12496 = ~1'b0 ;
  assign y12497 = ~n36403 ;
  assign y12498 = n36406 ;
  assign y12499 = ~n36409 ;
  assign y12500 = n36417 ;
  assign y12501 = ~n36418 ;
  assign y12502 = ~1'b0 ;
  assign y12503 = n36421 ;
  assign y12504 = ~1'b0 ;
  assign y12505 = n36424 ;
  assign y12506 = n36431 ;
  assign y12507 = n36432 ;
  assign y12508 = ~n36436 ;
  assign y12509 = n36438 ;
  assign y12510 = n36443 ;
  assign y12511 = ~n36445 ;
  assign y12512 = n36446 ;
  assign y12513 = n36450 ;
  assign y12514 = n14601 ;
  assign y12515 = ~n36452 ;
  assign y12516 = ~1'b0 ;
  assign y12517 = ~1'b0 ;
  assign y12518 = n36461 ;
  assign y12519 = n36463 ;
  assign y12520 = n36470 ;
  assign y12521 = ~1'b0 ;
  assign y12522 = ~n36472 ;
  assign y12523 = n36478 ;
  assign y12524 = n36480 ;
  assign y12525 = ~n36484 ;
  assign y12526 = ~n36488 ;
  assign y12527 = n36493 ;
  assign y12528 = n36495 ;
  assign y12529 = ~1'b0 ;
  assign y12530 = n36497 ;
  assign y12531 = ~n36499 ;
  assign y12532 = ~1'b0 ;
  assign y12533 = n36502 ;
  assign y12534 = n36509 ;
  assign y12535 = ~n36510 ;
  assign y12536 = n36513 ;
  assign y12537 = ~1'b0 ;
  assign y12538 = ~1'b0 ;
  assign y12539 = n36514 ;
  assign y12540 = ~n36518 ;
  assign y12541 = n36521 ;
  assign y12542 = n36522 ;
  assign y12543 = n36525 ;
  assign y12544 = ~1'b0 ;
  assign y12545 = ~n36529 ;
  assign y12546 = n10199 ;
  assign y12547 = ~n36531 ;
  assign y12548 = n36536 ;
  assign y12549 = ~n36538 ;
  assign y12550 = ~n36541 ;
  assign y12551 = n36542 ;
  assign y12552 = n36545 ;
  assign y12553 = ~n36547 ;
  assign y12554 = ~1'b0 ;
  assign y12555 = ~n36558 ;
  assign y12556 = n36560 ;
  assign y12557 = ~n36561 ;
  assign y12558 = n36562 ;
  assign y12559 = ~1'b0 ;
  assign y12560 = n36564 ;
  assign y12561 = n36567 ;
  assign y12562 = ~1'b0 ;
  assign y12563 = n36570 ;
  assign y12564 = n18243 ;
  assign y12565 = ~n36571 ;
  assign y12566 = ~n36573 ;
  assign y12567 = ~n36575 ;
  assign y12568 = n36576 ;
  assign y12569 = ~n36578 ;
  assign y12570 = ~n36584 ;
  assign y12571 = ~n36591 ;
  assign y12572 = n36594 ;
  assign y12573 = ~n36596 ;
  assign y12574 = ~1'b0 ;
  assign y12575 = ~n36597 ;
  assign y12576 = ~n36599 ;
  assign y12577 = ~1'b0 ;
  assign y12578 = n36600 ;
  assign y12579 = n36608 ;
  assign y12580 = n36609 ;
  assign y12581 = ~1'b0 ;
  assign y12582 = ~n36611 ;
  assign y12583 = n36614 ;
  assign y12584 = ~n36618 ;
  assign y12585 = ~n36619 ;
  assign y12586 = ~n36621 ;
  assign y12587 = n36629 ;
  assign y12588 = ~n36633 ;
  assign y12589 = ~1'b0 ;
  assign y12590 = ~n36636 ;
  assign y12591 = ~n36639 ;
  assign y12592 = n36644 ;
  assign y12593 = ~n834 ;
  assign y12594 = ~1'b0 ;
  assign y12595 = ~n36645 ;
  assign y12596 = ~n36646 ;
  assign y12597 = n36649 ;
  assign y12598 = ~n36650 ;
  assign y12599 = ~n36654 ;
  assign y12600 = ~1'b0 ;
  assign y12601 = ~n36655 ;
  assign y12602 = ~n36658 ;
  assign y12603 = ~n36660 ;
  assign y12604 = n36663 ;
  assign y12605 = ~1'b0 ;
  assign y12606 = n36664 ;
  assign y12607 = n36665 ;
  assign y12608 = n36676 ;
  assign y12609 = ~n36677 ;
  assign y12610 = n36681 ;
  assign y12611 = ~1'b0 ;
  assign y12612 = n36684 ;
  assign y12613 = ~n36685 ;
  assign y12614 = ~n36689 ;
  assign y12615 = n36691 ;
  assign y12616 = ~n36694 ;
  assign y12617 = n36699 ;
  assign y12618 = n36704 ;
  assign y12619 = ~n36706 ;
  assign y12620 = ~n36707 ;
  assign y12621 = n36709 ;
  assign y12622 = ~1'b0 ;
  assign y12623 = ~n36710 ;
  assign y12624 = ~1'b0 ;
  assign y12625 = n36712 ;
  assign y12626 = n36715 ;
  assign y12627 = ~n36716 ;
  assign y12628 = n36719 ;
  assign y12629 = n36720 ;
  assign y12630 = ~1'b0 ;
  assign y12631 = ~n36722 ;
  assign y12632 = ~n36724 ;
  assign y12633 = n36725 ;
  assign y12634 = ~n36726 ;
  assign y12635 = n36727 ;
  assign y12636 = n36729 ;
  assign y12637 = ~n36731 ;
  assign y12638 = ~1'b0 ;
  assign y12639 = n36733 ;
  assign y12640 = ~n36738 ;
  assign y12641 = n36743 ;
  assign y12642 = ~n36744 ;
  assign y12643 = n36745 ;
  assign y12644 = ~n36747 ;
  assign y12645 = n36748 ;
  assign y12646 = n36749 ;
  assign y12647 = n36751 ;
  assign y12648 = 1'b0 ;
  assign y12649 = ~1'b0 ;
  assign y12650 = n36752 ;
  assign y12651 = ~n36756 ;
  assign y12652 = ~n36759 ;
  assign y12653 = ~n36763 ;
  assign y12654 = ~1'b0 ;
  assign y12655 = ~n36765 ;
  assign y12656 = ~n36769 ;
  assign y12657 = n36771 ;
  assign y12658 = n25067 ;
  assign y12659 = ~n36772 ;
  assign y12660 = ~1'b0 ;
  assign y12661 = n36773 ;
  assign y12662 = ~n36776 ;
  assign y12663 = ~n36783 ;
  assign y12664 = n36788 ;
  assign y12665 = n36789 ;
  assign y12666 = ~n36792 ;
  assign y12667 = ~n36794 ;
  assign y12668 = n36795 ;
  assign y12669 = ~n36803 ;
  assign y12670 = ~1'b0 ;
  assign y12671 = ~n36804 ;
  assign y12672 = n36807 ;
  assign y12673 = n36809 ;
  assign y12674 = n36820 ;
  assign y12675 = ~1'b0 ;
  assign y12676 = n36824 ;
  assign y12677 = ~n36829 ;
  assign y12678 = n36832 ;
  assign y12679 = ~n36836 ;
  assign y12680 = n36839 ;
  assign y12681 = n36841 ;
  assign y12682 = ~n36842 ;
  assign y12683 = n2394 ;
  assign y12684 = n36845 ;
  assign y12685 = ~1'b0 ;
  assign y12686 = n36847 ;
  assign y12687 = ~1'b0 ;
  assign y12688 = n36853 ;
  assign y12689 = n36856 ;
  assign y12690 = n36862 ;
  assign y12691 = ~n36863 ;
  assign y12692 = n36864 ;
  assign y12693 = ~1'b0 ;
  assign y12694 = ~n36867 ;
  assign y12695 = n36870 ;
  assign y12696 = ~n36873 ;
  assign y12697 = n36874 ;
  assign y12698 = n36879 ;
  assign y12699 = ~1'b0 ;
  assign y12700 = ~n36881 ;
  assign y12701 = ~n36883 ;
  assign y12702 = ~1'b0 ;
  assign y12703 = n36884 ;
  assign y12704 = ~n36888 ;
  assign y12705 = ~n36891 ;
  assign y12706 = ~n36898 ;
  assign y12707 = ~n36899 ;
  assign y12708 = ~n36901 ;
  assign y12709 = ~n36902 ;
  assign y12710 = ~n36907 ;
  assign y12711 = ~n36909 ;
  assign y12712 = ~n36911 ;
  assign y12713 = ~1'b0 ;
  assign y12714 = ~n36912 ;
  assign y12715 = n36913 ;
  assign y12716 = ~n36916 ;
  assign y12717 = ~n36917 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = n36925 ;
  assign y12720 = ~n36927 ;
  assign y12721 = ~1'b0 ;
  assign y12722 = n36929 ;
  assign y12723 = ~n36935 ;
  assign y12724 = ~n36936 ;
  assign y12725 = ~1'b0 ;
  assign y12726 = ~n36938 ;
  assign y12727 = n36941 ;
  assign y12728 = ~n36944 ;
  assign y12729 = ~n36945 ;
  assign y12730 = ~n36947 ;
  assign y12731 = ~n36955 ;
  assign y12732 = ~n36958 ;
  assign y12733 = n36960 ;
  assign y12734 = n11612 ;
  assign y12735 = ~1'b0 ;
  assign y12736 = ~n36963 ;
  assign y12737 = ~n36965 ;
  assign y12738 = ~n36968 ;
  assign y12739 = n36976 ;
  assign y12740 = ~1'b0 ;
  assign y12741 = ~1'b0 ;
  assign y12742 = ~1'b0 ;
  assign y12743 = ~n36979 ;
  assign y12744 = ~1'b0 ;
  assign y12745 = ~n36981 ;
  assign y12746 = ~n36984 ;
  assign y12747 = ~n36986 ;
  assign y12748 = ~1'b0 ;
  assign y12749 = ~n36987 ;
  assign y12750 = ~n36990 ;
  assign y12751 = n36997 ;
  assign y12752 = n36998 ;
  assign y12753 = ~n37001 ;
  assign y12754 = ~1'b0 ;
  assign y12755 = n37006 ;
  assign y12756 = n37009 ;
  assign y12757 = ~n15057 ;
  assign y12758 = ~n37013 ;
  assign y12759 = ~1'b0 ;
  assign y12760 = ~n37014 ;
  assign y12761 = ~1'b0 ;
  assign y12762 = ~1'b0 ;
  assign y12763 = ~n37017 ;
  assign y12764 = n37018 ;
  assign y12765 = n37019 ;
  assign y12766 = ~1'b0 ;
  assign y12767 = n37021 ;
  assign y12768 = n37027 ;
  assign y12769 = ~n37033 ;
  assign y12770 = n11071 ;
  assign y12771 = n37040 ;
  assign y12772 = n37044 ;
  assign y12773 = ~1'b0 ;
  assign y12774 = ~n37049 ;
  assign y12775 = n37051 ;
  assign y12776 = ~1'b0 ;
  assign y12777 = ~n37056 ;
  assign y12778 = ~n37058 ;
  assign y12779 = n37059 ;
  assign y12780 = ~n37061 ;
  assign y12781 = ~n37068 ;
  assign y12782 = n37072 ;
  assign y12783 = n37078 ;
  assign y12784 = ~1'b0 ;
  assign y12785 = n37081 ;
  assign y12786 = n37088 ;
  assign y12787 = n37093 ;
  assign y12788 = n37096 ;
  assign y12789 = n37098 ;
  assign y12790 = 1'b0 ;
  assign y12791 = n37102 ;
  assign y12792 = ~1'b0 ;
  assign y12793 = ~n37104 ;
  assign y12794 = ~n37107 ;
  assign y12795 = n37110 ;
  assign y12796 = n37114 ;
  assign y12797 = n37115 ;
  assign y12798 = ~1'b0 ;
  assign y12799 = ~n37117 ;
  assign y12800 = ~n37120 ;
  assign y12801 = n37121 ;
  assign y12802 = ~n37127 ;
  assign y12803 = ~1'b0 ;
  assign y12804 = ~n37129 ;
  assign y12805 = ~n37131 ;
  assign y12806 = ~n37134 ;
  assign y12807 = ~n37135 ;
  assign y12808 = n37136 ;
  assign y12809 = ~n37139 ;
  assign y12810 = ~n37143 ;
  assign y12811 = ~n37147 ;
  assign y12812 = ~n37148 ;
  assign y12813 = ~n37151 ;
  assign y12814 = ~n37154 ;
  assign y12815 = ~1'b0 ;
  assign y12816 = ~n37159 ;
  assign y12817 = ~1'b0 ;
  assign y12818 = ~n37162 ;
  assign y12819 = n37163 ;
  assign y12820 = ~n37166 ;
  assign y12821 = n37169 ;
  assign y12822 = n37170 ;
  assign y12823 = ~n37177 ;
  assign y12824 = n37179 ;
  assign y12825 = ~n37181 ;
  assign y12826 = ~n37184 ;
  assign y12827 = ~n37187 ;
  assign y12828 = n37189 ;
  assign y12829 = n37196 ;
  assign y12830 = ~1'b0 ;
  assign y12831 = n37197 ;
  assign y12832 = ~1'b0 ;
  assign y12833 = ~1'b0 ;
  assign y12834 = ~n37198 ;
  assign y12835 = ~n37199 ;
  assign y12836 = n37202 ;
  assign y12837 = ~1'b0 ;
  assign y12838 = ~n37204 ;
  assign y12839 = ~n37205 ;
  assign y12840 = ~n37207 ;
  assign y12841 = ~n37209 ;
  assign y12842 = n37213 ;
  assign y12843 = ~n37219 ;
  assign y12844 = ~1'b0 ;
  assign y12845 = n37221 ;
  assign y12846 = ~1'b0 ;
  assign y12847 = ~n37223 ;
  assign y12848 = ~n37226 ;
  assign y12849 = ~n37229 ;
  assign y12850 = ~n12215 ;
  assign y12851 = n37233 ;
  assign y12852 = n37234 ;
  assign y12853 = ~n37236 ;
  assign y12854 = ~n37240 ;
  assign y12855 = n37242 ;
  assign y12856 = ~n37244 ;
  assign y12857 = ~n37248 ;
  assign y12858 = n37253 ;
  assign y12859 = n37254 ;
  assign y12860 = ~n37257 ;
  assign y12861 = ~1'b0 ;
  assign y12862 = ~n37259 ;
  assign y12863 = ~1'b0 ;
  assign y12864 = n37260 ;
  assign y12865 = ~n37261 ;
  assign y12866 = n37263 ;
  assign y12867 = ~n37266 ;
  assign y12868 = n37268 ;
  assign y12869 = ~n37270 ;
  assign y12870 = n37273 ;
  assign y12871 = n37274 ;
  assign y12872 = n37275 ;
  assign y12873 = n37282 ;
  assign y12874 = n31563 ;
  assign y12875 = n37283 ;
  assign y12876 = ~1'b0 ;
  assign y12877 = ~1'b0 ;
  assign y12878 = ~n37288 ;
  assign y12879 = ~1'b0 ;
  assign y12880 = ~n37291 ;
  assign y12881 = ~n37292 ;
  assign y12882 = ~n37293 ;
  assign y12883 = ~1'b0 ;
  assign y12884 = ~1'b0 ;
  assign y12885 = n37297 ;
  assign y12886 = ~n37299 ;
  assign y12887 = n37303 ;
  assign y12888 = n37308 ;
  assign y12889 = ~n37310 ;
  assign y12890 = n37316 ;
  assign y12891 = ~n37320 ;
  assign y12892 = ~1'b0 ;
  assign y12893 = 1'b0 ;
  assign y12894 = ~n37324 ;
  assign y12895 = ~n37326 ;
  assign y12896 = ~n37330 ;
  assign y12897 = n37335 ;
  assign y12898 = ~1'b0 ;
  assign y12899 = ~n37336 ;
  assign y12900 = ~n37337 ;
  assign y12901 = n37340 ;
  assign y12902 = n757 ;
  assign y12903 = n37341 ;
  assign y12904 = ~n37346 ;
  assign y12905 = ~n37347 ;
  assign y12906 = n37349 ;
  assign y12907 = ~n37350 ;
  assign y12908 = ~n37353 ;
  assign y12909 = ~n37355 ;
  assign y12910 = ~n37356 ;
  assign y12911 = ~1'b0 ;
  assign y12912 = n37359 ;
  assign y12913 = n37360 ;
  assign y12914 = n37364 ;
  assign y12915 = ~n37365 ;
  assign y12916 = ~1'b0 ;
  assign y12917 = ~n37367 ;
  assign y12918 = n37369 ;
  assign y12919 = n37372 ;
  assign y12920 = ~n37375 ;
  assign y12921 = n37376 ;
  assign y12922 = n37377 ;
  assign y12923 = n37378 ;
  assign y12924 = ~1'b0 ;
  assign y12925 = ~n37381 ;
  assign y12926 = ~n37382 ;
  assign y12927 = ~n37383 ;
  assign y12928 = ~n37384 ;
  assign y12929 = n37388 ;
  assign y12930 = ~n37393 ;
  assign y12931 = ~n37396 ;
  assign y12932 = ~1'b0 ;
  assign y12933 = ~n37397 ;
  assign y12934 = n37398 ;
  assign y12935 = n37400 ;
  assign y12936 = ~n37402 ;
  assign y12937 = ~n9495 ;
  assign y12938 = ~n37403 ;
  assign y12939 = n37408 ;
  assign y12940 = ~n37409 ;
  assign y12941 = ~n37413 ;
  assign y12942 = ~n37415 ;
  assign y12943 = ~n37416 ;
  assign y12944 = ~n37418 ;
  assign y12945 = n37420 ;
  assign y12946 = n37421 ;
  assign y12947 = ~n37425 ;
  assign y12948 = ~1'b0 ;
  assign y12949 = ~n37434 ;
  assign y12950 = ~n37436 ;
  assign y12951 = n37437 ;
  assign y12952 = ~1'b0 ;
  assign y12953 = ~n37438 ;
  assign y12954 = ~n37440 ;
  assign y12955 = n37444 ;
  assign y12956 = n37445 ;
  assign y12957 = ~n37447 ;
  assign y12958 = n37449 ;
  assign y12959 = n37450 ;
  assign y12960 = ~n37452 ;
  assign y12961 = n37456 ;
  assign y12962 = ~n37459 ;
  assign y12963 = ~n37460 ;
  assign y12964 = ~n37461 ;
  assign y12965 = ~n37463 ;
  assign y12966 = n37467 ;
  assign y12967 = ~n37468 ;
  assign y12968 = ~n37470 ;
  assign y12969 = ~n19980 ;
  assign y12970 = n37477 ;
  assign y12971 = ~n37479 ;
  assign y12972 = ~n37480 ;
  assign y12973 = ~1'b0 ;
  assign y12974 = n37481 ;
  assign y12975 = n37486 ;
  assign y12976 = ~n37490 ;
  assign y12977 = ~n37495 ;
  assign y12978 = ~1'b0 ;
  assign y12979 = ~n37498 ;
  assign y12980 = ~n37499 ;
  assign y12981 = ~n37502 ;
  assign y12982 = ~n37503 ;
  assign y12983 = ~n37507 ;
  assign y12984 = n37509 ;
  assign y12985 = ~1'b0 ;
  assign y12986 = n37512 ;
  assign y12987 = n37513 ;
  assign y12988 = n37515 ;
  assign y12989 = ~n37516 ;
  assign y12990 = ~n37518 ;
  assign y12991 = ~1'b0 ;
  assign y12992 = ~n37520 ;
  assign y12993 = ~1'b0 ;
  assign y12994 = ~n37522 ;
  assign y12995 = n37523 ;
  assign y12996 = n37527 ;
  assign y12997 = n37531 ;
  assign y12998 = ~n37532 ;
  assign y12999 = ~1'b0 ;
  assign y13000 = ~n37536 ;
  assign y13001 = ~1'b0 ;
  assign y13002 = n37538 ;
  assign y13003 = ~n3513 ;
  assign y13004 = ~n37539 ;
  assign y13005 = ~n37545 ;
  assign y13006 = ~n37547 ;
  assign y13007 = ~1'b0 ;
  assign y13008 = ~n37548 ;
  assign y13009 = n37549 ;
  assign y13010 = ~1'b0 ;
  assign y13011 = ~n37550 ;
  assign y13012 = ~n37553 ;
  assign y13013 = ~n37555 ;
  assign y13014 = n37562 ;
  assign y13015 = ~n37567 ;
  assign y13016 = ~n37573 ;
  assign y13017 = n37575 ;
  assign y13018 = ~n37576 ;
  assign y13019 = n37579 ;
  assign y13020 = n37582 ;
  assign y13021 = ~1'b0 ;
  assign y13022 = n37588 ;
  assign y13023 = ~1'b0 ;
  assign y13024 = ~n37589 ;
  assign y13025 = 1'b0 ;
  assign y13026 = ~n37591 ;
  assign y13027 = ~1'b0 ;
  assign y13028 = ~1'b0 ;
  assign y13029 = ~n37595 ;
  assign y13030 = n37597 ;
  assign y13031 = ~n37605 ;
  assign y13032 = n37610 ;
  assign y13033 = ~n23217 ;
  assign y13034 = ~n37612 ;
  assign y13035 = ~1'b0 ;
  assign y13036 = n37614 ;
  assign y13037 = ~n37620 ;
  assign y13038 = n37627 ;
  assign y13039 = ~n37628 ;
  assign y13040 = n37629 ;
  assign y13041 = n37633 ;
  assign y13042 = ~n37639 ;
  assign y13043 = n37641 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = n37642 ;
  assign y13046 = n37650 ;
  assign y13047 = ~n37653 ;
  assign y13048 = ~n37657 ;
  assign y13049 = ~n37659 ;
  assign y13050 = ~1'b0 ;
  assign y13051 = n37660 ;
  assign y13052 = ~1'b0 ;
  assign y13053 = ~n37661 ;
  assign y13054 = n37663 ;
  assign y13055 = ~n37668 ;
  assign y13056 = n37675 ;
  assign y13057 = n37676 ;
  assign y13058 = ~n37681 ;
  assign y13059 = ~n37683 ;
  assign y13060 = n37686 ;
  assign y13061 = n37689 ;
  assign y13062 = n37692 ;
  assign y13063 = n37695 ;
  assign y13064 = ~n37699 ;
  assign y13065 = ~n37703 ;
  assign y13066 = n37705 ;
  assign y13067 = ~n37706 ;
  assign y13068 = ~1'b0 ;
  assign y13069 = n37712 ;
  assign y13070 = n37715 ;
  assign y13071 = ~1'b0 ;
  assign y13072 = ~1'b0 ;
  assign y13073 = n37717 ;
  assign y13074 = ~n37718 ;
  assign y13075 = ~1'b0 ;
  assign y13076 = n37719 ;
  assign y13077 = ~1'b0 ;
  assign y13078 = n37728 ;
  assign y13079 = n37736 ;
  assign y13080 = ~n37737 ;
  assign y13081 = ~n37740 ;
  assign y13082 = n16481 ;
  assign y13083 = n37745 ;
  assign y13084 = ~n37747 ;
  assign y13085 = ~n37748 ;
  assign y13086 = ~n37750 ;
  assign y13087 = ~n37751 ;
  assign y13088 = ~n37755 ;
  assign y13089 = ~1'b0 ;
  assign y13090 = n37757 ;
  assign y13091 = ~1'b0 ;
  assign y13092 = ~n37761 ;
  assign y13093 = ~n37766 ;
  assign y13094 = n37770 ;
  assign y13095 = ~n37771 ;
  assign y13096 = ~n37774 ;
  assign y13097 = ~n37775 ;
  assign y13098 = ~n37783 ;
  assign y13099 = ~n37784 ;
  assign y13100 = ~n37791 ;
  assign y13101 = ~n37793 ;
  assign y13102 = ~n37794 ;
  assign y13103 = ~n37798 ;
  assign y13104 = n37799 ;
  assign y13105 = n37800 ;
  assign y13106 = n37803 ;
  assign y13107 = n37805 ;
  assign y13108 = n37807 ;
  assign y13109 = ~n37818 ;
  assign y13110 = ~1'b0 ;
  assign y13111 = ~n37821 ;
  assign y13112 = n37822 ;
  assign y13113 = n37823 ;
  assign y13114 = ~1'b0 ;
  assign y13115 = ~n37825 ;
  assign y13116 = ~1'b0 ;
  assign y13117 = ~1'b0 ;
  assign y13118 = ~n37829 ;
  assign y13119 = n37835 ;
  assign y13120 = ~n37838 ;
  assign y13121 = n37839 ;
  assign y13122 = n32599 ;
  assign y13123 = n37842 ;
  assign y13124 = n37844 ;
  assign y13125 = ~n37847 ;
  assign y13126 = n37851 ;
  assign y13127 = ~n37859 ;
  assign y13128 = ~1'b0 ;
  assign y13129 = n37863 ;
  assign y13130 = ~1'b0 ;
  assign y13131 = n37864 ;
  assign y13132 = ~n37867 ;
  assign y13133 = ~n37868 ;
  assign y13134 = n37869 ;
  assign y13135 = n37872 ;
  assign y13136 = 1'b0 ;
  assign y13137 = ~n37878 ;
  assign y13138 = n37879 ;
  assign y13139 = ~n37883 ;
  assign y13140 = n37885 ;
  assign y13141 = n37886 ;
  assign y13142 = ~1'b0 ;
  assign y13143 = n37887 ;
  assign y13144 = ~n37890 ;
  assign y13145 = ~n37892 ;
  assign y13146 = ~n37896 ;
  assign y13147 = ~1'b0 ;
  assign y13148 = n37897 ;
  assign y13149 = n37900 ;
  assign y13150 = ~n37902 ;
  assign y13151 = n37905 ;
  assign y13152 = ~n37906 ;
  assign y13153 = ~1'b0 ;
  assign y13154 = ~n37907 ;
  assign y13155 = ~n37909 ;
  assign y13156 = ~1'b0 ;
  assign y13157 = n37911 ;
  assign y13158 = n37914 ;
  assign y13159 = n37916 ;
  assign y13160 = n37919 ;
  assign y13161 = ~1'b0 ;
  assign y13162 = ~n37922 ;
  assign y13163 = ~n37926 ;
  assign y13164 = n37928 ;
  assign y13165 = n37931 ;
  assign y13166 = ~n37933 ;
  assign y13167 = n37934 ;
  assign y13168 = n37936 ;
  assign y13169 = ~n37939 ;
  assign y13170 = ~n37941 ;
  assign y13171 = ~1'b0 ;
  assign y13172 = n37947 ;
  assign y13173 = ~1'b0 ;
  assign y13174 = ~n37948 ;
  assign y13175 = ~n2394 ;
  assign y13176 = ~n31643 ;
  assign y13177 = ~n37949 ;
  assign y13178 = n37950 ;
  assign y13179 = n37953 ;
  assign y13180 = ~n37960 ;
  assign y13181 = n37967 ;
  assign y13182 = ~n37971 ;
  assign y13183 = ~n37973 ;
  assign y13184 = ~n37975 ;
  assign y13185 = ~n37976 ;
  assign y13186 = ~n37977 ;
  assign y13187 = ~n37978 ;
  assign y13188 = n37983 ;
  assign y13189 = n37984 ;
  assign y13190 = ~1'b0 ;
  assign y13191 = n37985 ;
  assign y13192 = n13055 ;
  assign y13193 = ~n36263 ;
  assign y13194 = n37989 ;
  assign y13195 = n37992 ;
  assign y13196 = ~n37994 ;
  assign y13197 = ~n37996 ;
  assign y13198 = n38000 ;
  assign y13199 = n38002 ;
  assign y13200 = ~n38004 ;
  assign y13201 = ~n38012 ;
  assign y13202 = ~1'b0 ;
  assign y13203 = n38014 ;
  assign y13204 = ~n38017 ;
  assign y13205 = n38024 ;
  assign y13206 = ~n38025 ;
  assign y13207 = ~n38026 ;
  assign y13208 = ~n38030 ;
  assign y13209 = ~1'b0 ;
  assign y13210 = ~1'b0 ;
  assign y13211 = ~n38031 ;
  assign y13212 = ~n38033 ;
  assign y13213 = n38034 ;
  assign y13214 = ~n38037 ;
  assign y13215 = ~n38042 ;
  assign y13216 = ~n38045 ;
  assign y13217 = ~1'b0 ;
  assign y13218 = ~n38048 ;
  assign y13219 = n38050 ;
  assign y13220 = n38051 ;
  assign y13221 = ~1'b0 ;
  assign y13222 = ~n38057 ;
  assign y13223 = ~1'b0 ;
  assign y13224 = n38059 ;
  assign y13225 = ~n38062 ;
  assign y13226 = ~n38069 ;
  assign y13227 = n38071 ;
  assign y13228 = ~1'b0 ;
  assign y13229 = n38072 ;
  assign y13230 = n38073 ;
  assign y13231 = n38077 ;
  assign y13232 = n38078 ;
  assign y13233 = n38080 ;
  assign y13234 = n3035 ;
  assign y13235 = n38082 ;
  assign y13236 = ~n38085 ;
  assign y13237 = ~n38087 ;
  assign y13238 = ~n38090 ;
  assign y13239 = n38093 ;
  assign y13240 = n38095 ;
  assign y13241 = ~1'b0 ;
  assign y13242 = n38096 ;
  assign y13243 = ~n38100 ;
  assign y13244 = n38108 ;
  assign y13245 = n38109 ;
  assign y13246 = ~1'b0 ;
  assign y13247 = ~n38113 ;
  assign y13248 = ~n38114 ;
  assign y13249 = ~n38115 ;
  assign y13250 = ~1'b0 ;
  assign y13251 = ~n38117 ;
  assign y13252 = 1'b0 ;
  assign y13253 = n38120 ;
  assign y13254 = ~n38121 ;
  assign y13255 = ~n38122 ;
  assign y13256 = n38125 ;
  assign y13257 = n20750 ;
  assign y13258 = ~1'b0 ;
  assign y13259 = n38131 ;
  assign y13260 = ~n38133 ;
  assign y13261 = ~n38137 ;
  assign y13262 = n38139 ;
  assign y13263 = ~n38141 ;
  assign y13264 = ~1'b0 ;
  assign y13265 = ~1'b0 ;
  assign y13266 = ~1'b0 ;
  assign y13267 = n590 ;
  assign y13268 = ~n38146 ;
  assign y13269 = ~1'b0 ;
  assign y13270 = ~n38150 ;
  assign y13271 = ~n38152 ;
  assign y13272 = ~n38153 ;
  assign y13273 = ~n38156 ;
  assign y13274 = ~n38164 ;
  assign y13275 = n38168 ;
  assign y13276 = ~1'b0 ;
  assign y13277 = ~n38170 ;
  assign y13278 = ~n38172 ;
  assign y13279 = ~1'b0 ;
  assign y13280 = ~1'b0 ;
  assign y13281 = 1'b0 ;
  assign y13282 = ~1'b0 ;
  assign y13283 = ~1'b0 ;
  assign y13284 = ~n38173 ;
  assign y13285 = n305 ;
  assign y13286 = ~1'b0 ;
  assign y13287 = ~n38174 ;
  assign y13288 = ~n38175 ;
  assign y13289 = n38176 ;
  assign y13290 = n38177 ;
  assign y13291 = ~1'b0 ;
  assign y13292 = ~n38178 ;
  assign y13293 = n38186 ;
  assign y13294 = ~1'b0 ;
  assign y13295 = ~n38189 ;
  assign y13296 = n38190 ;
  assign y13297 = ~1'b0 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~1'b0 ;
  assign y13300 = ~n38195 ;
  assign y13301 = ~n38197 ;
  assign y13302 = ~n38199 ;
  assign y13303 = n38201 ;
  assign y13304 = ~1'b0 ;
  assign y13305 = ~n38203 ;
  assign y13306 = ~n38204 ;
  assign y13307 = n38208 ;
  assign y13308 = n38211 ;
  assign y13309 = 1'b0 ;
  assign y13310 = n38218 ;
  assign y13311 = ~n38225 ;
  assign y13312 = ~n38226 ;
  assign y13313 = n38228 ;
  assign y13314 = n38229 ;
  assign y13315 = ~n38232 ;
  assign y13316 = n38234 ;
  assign y13317 = n38237 ;
  assign y13318 = n38238 ;
  assign y13319 = ~n38240 ;
  assign y13320 = ~n38242 ;
  assign y13321 = n38243 ;
  assign y13322 = ~n38244 ;
  assign y13323 = ~n38248 ;
  assign y13324 = ~n38256 ;
  assign y13325 = n38264 ;
  assign y13326 = n38271 ;
  assign y13327 = ~n36905 ;
  assign y13328 = ~1'b0 ;
  assign y13329 = ~n38272 ;
  assign y13330 = n38278 ;
  assign y13331 = ~n38279 ;
  assign y13332 = ~1'b0 ;
  assign y13333 = ~n38281 ;
  assign y13334 = n38284 ;
  assign y13335 = n38287 ;
  assign y13336 = ~n38289 ;
  assign y13337 = ~n38294 ;
  assign y13338 = ~n38295 ;
  assign y13339 = n38296 ;
  assign y13340 = n38298 ;
  assign y13341 = ~1'b0 ;
  assign y13342 = ~1'b0 ;
  assign y13343 = ~1'b0 ;
  assign y13344 = ~n38304 ;
  assign y13345 = n38310 ;
  assign y13346 = ~1'b0 ;
  assign y13347 = ~n38319 ;
  assign y13348 = ~1'b0 ;
  assign y13349 = ~1'b0 ;
  assign y13350 = n38323 ;
  assign y13351 = ~n38326 ;
  assign y13352 = ~n35548 ;
  assign y13353 = ~n38328 ;
  assign y13354 = n38331 ;
  assign y13355 = ~n38333 ;
  assign y13356 = ~n38334 ;
  assign y13357 = n38339 ;
  assign y13358 = ~n38341 ;
  assign y13359 = ~n2782 ;
  assign y13360 = ~1'b0 ;
  assign y13361 = ~1'b0 ;
  assign y13362 = ~n38343 ;
  assign y13363 = n38344 ;
  assign y13364 = n38347 ;
  assign y13365 = n38349 ;
  assign y13366 = n38350 ;
  assign y13367 = n38352 ;
  assign y13368 = ~n38354 ;
  assign y13369 = n38355 ;
  assign y13370 = ~n38359 ;
  assign y13371 = ~n38361 ;
  assign y13372 = n38363 ;
  assign y13373 = n38364 ;
  assign y13374 = n38369 ;
  assign y13375 = ~n38370 ;
  assign y13376 = ~1'b0 ;
  assign y13377 = ~n38373 ;
  assign y13378 = ~n38374 ;
  assign y13379 = n38375 ;
  assign y13380 = ~1'b0 ;
  assign y13381 = ~1'b0 ;
  assign y13382 = ~n38377 ;
  assign y13383 = n38378 ;
  assign y13384 = ~n38379 ;
  assign y13385 = n38386 ;
  assign y13386 = ~1'b0 ;
  assign y13387 = ~1'b0 ;
  assign y13388 = ~n38387 ;
  assign y13389 = n38390 ;
  assign y13390 = n38392 ;
  assign y13391 = ~n38395 ;
  assign y13392 = ~n38396 ;
  assign y13393 = n38398 ;
  assign y13394 = ~1'b0 ;
  assign y13395 = ~1'b0 ;
  assign y13396 = ~n38400 ;
  assign y13397 = n38405 ;
  assign y13398 = ~n29896 ;
  assign y13399 = n38410 ;
  assign y13400 = ~n38413 ;
  assign y13401 = ~1'b0 ;
  assign y13402 = ~n38414 ;
  assign y13403 = 1'b0 ;
  assign y13404 = n38417 ;
  assign y13405 = ~n38418 ;
  assign y13406 = n38430 ;
  assign y13407 = ~1'b0 ;
  assign y13408 = ~n38432 ;
  assign y13409 = ~n38435 ;
  assign y13410 = ~n38441 ;
  assign y13411 = n38443 ;
  assign y13412 = ~n38446 ;
  assign y13413 = n38447 ;
  assign y13414 = n38451 ;
  assign y13415 = ~1'b0 ;
  assign y13416 = n38453 ;
  assign y13417 = n38454 ;
  assign y13418 = ~n38458 ;
  assign y13419 = n38459 ;
  assign y13420 = ~n38462 ;
  assign y13421 = ~n38463 ;
  assign y13422 = ~n38467 ;
  assign y13423 = ~1'b0 ;
  assign y13424 = ~n38470 ;
  assign y13425 = ~1'b0 ;
  assign y13426 = ~n38471 ;
  assign y13427 = n38474 ;
  assign y13428 = ~1'b0 ;
  assign y13429 = ~n38479 ;
  assign y13430 = ~n38482 ;
  assign y13431 = n38486 ;
  assign y13432 = n38489 ;
  assign y13433 = ~1'b0 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = ~n38490 ;
  assign y13436 = n38493 ;
  assign y13437 = n38494 ;
  assign y13438 = n38495 ;
  assign y13439 = ~1'b0 ;
  assign y13440 = ~1'b0 ;
  assign y13441 = ~n38498 ;
  assign y13442 = n38501 ;
  assign y13443 = ~n38502 ;
  assign y13444 = n38503 ;
  assign y13445 = 1'b0 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = ~n38504 ;
  assign y13448 = ~1'b0 ;
  assign y13449 = ~n38512 ;
  assign y13450 = ~n38514 ;
  assign y13451 = n38515 ;
  assign y13452 = n38518 ;
  assign y13453 = ~1'b0 ;
  assign y13454 = n38524 ;
  assign y13455 = ~1'b0 ;
  assign y13456 = ~n38526 ;
  assign y13457 = ~n38528 ;
  assign y13458 = ~n38530 ;
  assign y13459 = n38531 ;
  assign y13460 = n38534 ;
  assign y13461 = n38538 ;
  assign y13462 = ~1'b0 ;
  assign y13463 = n38540 ;
  assign y13464 = ~n38548 ;
  assign y13465 = n38553 ;
  assign y13466 = ~n38555 ;
  assign y13467 = n38558 ;
  assign y13468 = ~1'b0 ;
  assign y13469 = ~1'b0 ;
  assign y13470 = n38559 ;
  assign y13471 = ~n38560 ;
  assign y13472 = n38563 ;
  assign y13473 = ~n38564 ;
  assign y13474 = n38568 ;
  assign y13475 = n38572 ;
  assign y13476 = ~n38573 ;
  assign y13477 = ~n38575 ;
  assign y13478 = n38576 ;
  assign y13479 = ~n38578 ;
  assign y13480 = ~n38579 ;
  assign y13481 = n38586 ;
  assign y13482 = ~1'b0 ;
  assign y13483 = ~n38590 ;
  assign y13484 = ~n38592 ;
  assign y13485 = ~1'b0 ;
  assign y13486 = ~1'b0 ;
  assign y13487 = n38599 ;
  assign y13488 = n38601 ;
  assign y13489 = n38604 ;
  assign y13490 = ~n38605 ;
  assign y13491 = ~1'b0 ;
  assign y13492 = ~1'b0 ;
  assign y13493 = ~n38608 ;
  assign y13494 = ~n38609 ;
  assign y13495 = ~n38612 ;
  assign y13496 = ~1'b0 ;
  assign y13497 = ~n38617 ;
  assign y13498 = n38624 ;
  assign y13499 = ~n38626 ;
  assign y13500 = ~n38629 ;
  assign y13501 = ~n38633 ;
  assign y13502 = ~n35552 ;
  assign y13503 = n38637 ;
  assign y13504 = ~n38640 ;
  assign y13505 = n38641 ;
  assign y13506 = ~1'b0 ;
  assign y13507 = ~1'b0 ;
  assign y13508 = ~1'b0 ;
  assign y13509 = ~1'b0 ;
  assign y13510 = n38643 ;
  assign y13511 = ~n38646 ;
  assign y13512 = ~n38648 ;
  assign y13513 = ~n38652 ;
  assign y13514 = n38653 ;
  assign y13515 = n38662 ;
  assign y13516 = n38671 ;
  assign y13517 = n38672 ;
  assign y13518 = ~n38674 ;
  assign y13519 = ~1'b0 ;
  assign y13520 = n38678 ;
  assign y13521 = ~1'b0 ;
  assign y13522 = ~n38682 ;
  assign y13523 = n38686 ;
  assign y13524 = n38687 ;
  assign y13525 = ~n38688 ;
  assign y13526 = ~n38690 ;
  assign y13527 = ~n38691 ;
  assign y13528 = ~n38692 ;
  assign y13529 = ~1'b0 ;
  assign y13530 = n38694 ;
  assign y13531 = ~n38695 ;
  assign y13532 = n38697 ;
  assign y13533 = ~n38704 ;
  assign y13534 = n38710 ;
  assign y13535 = n38714 ;
  assign y13536 = ~n38716 ;
  assign y13537 = n38720 ;
  assign y13538 = ~1'b0 ;
  assign y13539 = ~n38722 ;
  assign y13540 = ~n38724 ;
  assign y13541 = ~n38728 ;
  assign y13542 = n38732 ;
  assign y13543 = ~n38733 ;
  assign y13544 = ~n38737 ;
  assign y13545 = ~n38738 ;
  assign y13546 = ~n38740 ;
  assign y13547 = n38741 ;
  assign y13548 = ~n38750 ;
  assign y13549 = n38753 ;
  assign y13550 = n38756 ;
  assign y13551 = ~n38764 ;
  assign y13552 = n38765 ;
  assign y13553 = ~n38773 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = n38775 ;
  assign y13556 = ~n38776 ;
  assign y13557 = ~n38777 ;
  assign y13558 = ~n38782 ;
  assign y13559 = ~n38789 ;
  assign y13560 = ~n38791 ;
  assign y13561 = ~n38793 ;
  assign y13562 = n38798 ;
  assign y13563 = ~n38802 ;
  assign y13564 = ~n38803 ;
  assign y13565 = ~n38805 ;
  assign y13566 = ~n38807 ;
  assign y13567 = ~n38810 ;
  assign y13568 = n30660 ;
  assign y13569 = n38811 ;
  assign y13570 = n38812 ;
  assign y13571 = n38814 ;
  assign y13572 = ~n38818 ;
  assign y13573 = ~n38822 ;
  assign y13574 = ~1'b0 ;
  assign y13575 = ~1'b0 ;
  assign y13576 = n38827 ;
  assign y13577 = n38828 ;
  assign y13578 = n38831 ;
  assign y13579 = ~n38833 ;
  assign y13580 = ~n38836 ;
  assign y13581 = ~1'b0 ;
  assign y13582 = n38838 ;
  assign y13583 = ~n38840 ;
  assign y13584 = ~1'b0 ;
  assign y13585 = ~n38841 ;
  assign y13586 = ~n38844 ;
  assign y13587 = n38849 ;
  assign y13588 = ~1'b0 ;
  assign y13589 = ~1'b0 ;
  assign y13590 = ~n38853 ;
  assign y13591 = ~n38854 ;
  assign y13592 = n38856 ;
  assign y13593 = n38857 ;
  assign y13594 = n38860 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = n38863 ;
  assign y13597 = ~1'b0 ;
  assign y13598 = ~n38864 ;
  assign y13599 = ~n38867 ;
  assign y13600 = ~n4375 ;
  assign y13601 = ~n38869 ;
  assign y13602 = n38880 ;
  assign y13603 = ~n38884 ;
  assign y13604 = n38885 ;
  assign y13605 = n38888 ;
  assign y13606 = ~1'b0 ;
  assign y13607 = n38897 ;
  assign y13608 = n38900 ;
  assign y13609 = n38903 ;
  assign y13610 = ~n38906 ;
  assign y13611 = ~n38909 ;
  assign y13612 = n38911 ;
  assign y13613 = n38912 ;
  assign y13614 = ~1'b0 ;
  assign y13615 = n38914 ;
  assign y13616 = ~n38918 ;
  assign y13617 = n38919 ;
  assign y13618 = ~n38922 ;
  assign y13619 = n38923 ;
  assign y13620 = n38926 ;
  assign y13621 = ~1'b0 ;
  assign y13622 = n38929 ;
  assign y13623 = ~n38930 ;
  assign y13624 = ~n23476 ;
  assign y13625 = ~1'b0 ;
  assign y13626 = ~n38931 ;
  assign y13627 = n38937 ;
  assign y13628 = ~n38939 ;
  assign y13629 = n38941 ;
  assign y13630 = n38944 ;
  assign y13631 = ~n34395 ;
  assign y13632 = ~n38950 ;
  assign y13633 = ~n38952 ;
  assign y13634 = ~n38953 ;
  assign y13635 = ~n38956 ;
  assign y13636 = n38958 ;
  assign y13637 = ~n38965 ;
  assign y13638 = n18763 ;
  assign y13639 = n38969 ;
  assign y13640 = n38974 ;
  assign y13641 = n38975 ;
  assign y13642 = n38978 ;
  assign y13643 = ~n38979 ;
  assign y13644 = ~n38981 ;
  assign y13645 = ~n38982 ;
  assign y13646 = n38984 ;
  assign y13647 = ~n38986 ;
  assign y13648 = ~n38989 ;
  assign y13649 = n38992 ;
  assign y13650 = ~1'b0 ;
  assign y13651 = ~1'b0 ;
  assign y13652 = ~1'b0 ;
  assign y13653 = n38993 ;
  assign y13654 = n39001 ;
  assign y13655 = n39002 ;
  assign y13656 = n39005 ;
  assign y13657 = ~n39009 ;
  assign y13658 = n39010 ;
  assign y13659 = n39012 ;
  assign y13660 = ~n39014 ;
  assign y13661 = n39015 ;
  assign y13662 = n5537 ;
  assign y13663 = ~n39016 ;
  assign y13664 = ~n39017 ;
  assign y13665 = n39018 ;
  assign y13666 = n39019 ;
  assign y13667 = n39026 ;
  assign y13668 = ~1'b0 ;
  assign y13669 = n39028 ;
  assign y13670 = ~n39030 ;
  assign y13671 = n39032 ;
  assign y13672 = ~1'b0 ;
  assign y13673 = n39034 ;
  assign y13674 = n39035 ;
  assign y13675 = n39037 ;
  assign y13676 = n39038 ;
  assign y13677 = ~n39042 ;
  assign y13678 = ~1'b0 ;
  assign y13679 = n39054 ;
  assign y13680 = ~1'b0 ;
  assign y13681 = ~1'b0 ;
  assign y13682 = ~n39055 ;
  assign y13683 = n39056 ;
  assign y13684 = ~n39059 ;
  assign y13685 = n39061 ;
  assign y13686 = n39063 ;
  assign y13687 = n39067 ;
  assign y13688 = ~n39068 ;
  assign y13689 = ~n39069 ;
  assign y13690 = ~1'b0 ;
  assign y13691 = n39071 ;
  assign y13692 = n39073 ;
  assign y13693 = ~1'b0 ;
  assign y13694 = n39079 ;
  assign y13695 = ~n39083 ;
  assign y13696 = ~n39088 ;
  assign y13697 = ~n39089 ;
  assign y13698 = ~1'b0 ;
  assign y13699 = ~n39091 ;
  assign y13700 = ~n39096 ;
  assign y13701 = ~1'b0 ;
  assign y13702 = ~n39102 ;
  assign y13703 = ~n39105 ;
  assign y13704 = n39106 ;
  assign y13705 = ~1'b0 ;
  assign y13706 = ~n39108 ;
  assign y13707 = ~n39109 ;
  assign y13708 = ~n39115 ;
  assign y13709 = n28401 ;
  assign y13710 = ~n39122 ;
  assign y13711 = ~1'b0 ;
  assign y13712 = ~n39124 ;
  assign y13713 = n39126 ;
  assign y13714 = ~n39128 ;
  assign y13715 = ~n39129 ;
  assign y13716 = ~n39134 ;
  assign y13717 = ~n39139 ;
  assign y13718 = n39140 ;
  assign y13719 = ~n39143 ;
  assign y13720 = n16649 ;
  assign y13721 = n39146 ;
  assign y13722 = ~n39147 ;
  assign y13723 = ~1'b0 ;
  assign y13724 = n39150 ;
  assign y13725 = ~n39151 ;
  assign y13726 = n39154 ;
  assign y13727 = ~n39156 ;
  assign y13728 = ~1'b0 ;
  assign y13729 = ~n39160 ;
  assign y13730 = n39163 ;
  assign y13731 = n10369 ;
  assign y13732 = n39166 ;
  assign y13733 = ~n39172 ;
  assign y13734 = ~n39173 ;
  assign y13735 = ~1'b0 ;
  assign y13736 = n39180 ;
  assign y13737 = n39181 ;
  assign y13738 = ~n39182 ;
  assign y13739 = ~1'b0 ;
  assign y13740 = n39185 ;
  assign y13741 = n39188 ;
  assign y13742 = ~n39190 ;
  assign y13743 = ~n39193 ;
  assign y13744 = ~1'b0 ;
  assign y13745 = n39200 ;
  assign y13746 = n39201 ;
  assign y13747 = ~1'b0 ;
  assign y13748 = n39202 ;
  assign y13749 = ~n39203 ;
  assign y13750 = n39205 ;
  assign y13751 = ~1'b0 ;
  assign y13752 = n39209 ;
  assign y13753 = n39211 ;
  assign y13754 = n39217 ;
  assign y13755 = ~n39219 ;
  assign y13756 = n39221 ;
  assign y13757 = ~n39225 ;
  assign y13758 = n39226 ;
  assign y13759 = n39230 ;
  assign y13760 = ~n39232 ;
  assign y13761 = ~1'b0 ;
  assign y13762 = ~n39237 ;
  assign y13763 = 1'b0 ;
  assign y13764 = n39243 ;
  assign y13765 = ~n39244 ;
  assign y13766 = ~n39250 ;
  assign y13767 = n39251 ;
  assign y13768 = ~n39253 ;
  assign y13769 = ~n39257 ;
  assign y13770 = ~n39259 ;
  assign y13771 = n39261 ;
  assign y13772 = n39266 ;
  assign y13773 = n39272 ;
  assign y13774 = ~n39290 ;
  assign y13775 = n39295 ;
  assign y13776 = ~n39297 ;
  assign y13777 = n39300 ;
  assign y13778 = ~1'b0 ;
  assign y13779 = ~n39301 ;
  assign y13780 = n39302 ;
  assign y13781 = ~n39305 ;
  assign y13782 = n39307 ;
  assign y13783 = ~n39309 ;
  assign y13784 = ~n39310 ;
  assign y13785 = ~n39312 ;
  assign y13786 = ~n39318 ;
  assign y13787 = ~n39325 ;
  assign y13788 = ~n39326 ;
  assign y13789 = n39329 ;
  assign y13790 = n39331 ;
  assign y13791 = ~n39333 ;
  assign y13792 = ~1'b0 ;
  assign y13793 = ~n39335 ;
  assign y13794 = ~n39344 ;
  assign y13795 = ~n39345 ;
  assign y13796 = ~n39346 ;
  assign y13797 = ~n39347 ;
  assign y13798 = n39351 ;
  assign y13799 = ~n39355 ;
  assign y13800 = ~n39356 ;
  assign y13801 = n39361 ;
  assign y13802 = n39364 ;
  assign y13803 = n39366 ;
  assign y13804 = ~1'b0 ;
  assign y13805 = ~n39369 ;
  assign y13806 = ~n39371 ;
  assign y13807 = ~n39372 ;
  assign y13808 = n39373 ;
  assign y13809 = n39376 ;
  assign y13810 = n39377 ;
  assign y13811 = n39380 ;
  assign y13812 = ~n39382 ;
  assign y13813 = ~n39384 ;
  assign y13814 = n39386 ;
  assign y13815 = n39387 ;
  assign y13816 = ~n39388 ;
  assign y13817 = ~n39391 ;
  assign y13818 = ~1'b0 ;
  assign y13819 = n38557 ;
  assign y13820 = ~1'b0 ;
  assign y13821 = n39395 ;
  assign y13822 = ~n39396 ;
  assign y13823 = n39397 ;
  assign y13824 = ~n39399 ;
  assign y13825 = ~1'b0 ;
  assign y13826 = n39401 ;
  assign y13827 = n39410 ;
  assign y13828 = ~n39414 ;
  assign y13829 = n39418 ;
  assign y13830 = ~n39424 ;
  assign y13831 = ~n39426 ;
  assign y13832 = ~1'b0 ;
  assign y13833 = ~n39428 ;
  assign y13834 = n39432 ;
  assign y13835 = ~n39433 ;
  assign y13836 = ~n39434 ;
  assign y13837 = ~n39446 ;
  assign y13838 = n39448 ;
  assign y13839 = ~n39449 ;
  assign y13840 = ~1'b0 ;
  assign y13841 = n39454 ;
  assign y13842 = ~n39456 ;
  assign y13843 = ~n39457 ;
  assign y13844 = n37165 ;
  assign y13845 = n39459 ;
  assign y13846 = ~n39460 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = n39462 ;
  assign y13849 = n39468 ;
  assign y13850 = n39470 ;
  assign y13851 = n39471 ;
  assign y13852 = 1'b0 ;
  assign y13853 = n39472 ;
  assign y13854 = n39474 ;
  assign y13855 = ~n39477 ;
  assign y13856 = ~n17065 ;
  assign y13857 = n39478 ;
  assign y13858 = n39479 ;
  assign y13859 = ~n39484 ;
  assign y13860 = ~1'b0 ;
  assign y13861 = ~n39487 ;
  assign y13862 = ~1'b0 ;
  assign y13863 = ~n39490 ;
  assign y13864 = n39492 ;
  assign y13865 = n39493 ;
  assign y13866 = n39497 ;
  assign y13867 = n39498 ;
  assign y13868 = n666 ;
  assign y13869 = n39502 ;
  assign y13870 = n39505 ;
  assign y13871 = ~n39511 ;
  assign y13872 = n39512 ;
  assign y13873 = ~n39518 ;
  assign y13874 = ~n39520 ;
  assign y13875 = ~n39525 ;
  assign y13876 = ~n39527 ;
  assign y13877 = ~n39533 ;
  assign y13878 = ~n39539 ;
  assign y13879 = n39540 ;
  assign y13880 = ~n39542 ;
  assign y13881 = n39545 ;
  assign y13882 = n39549 ;
  assign y13883 = ~n39552 ;
  assign y13884 = ~n39553 ;
  assign y13885 = ~n39555 ;
  assign y13886 = ~n39557 ;
  assign y13887 = ~n39558 ;
  assign y13888 = n39559 ;
  assign y13889 = n39560 ;
  assign y13890 = ~1'b0 ;
  assign y13891 = ~1'b0 ;
  assign y13892 = ~n39562 ;
  assign y13893 = ~1'b0 ;
  assign y13894 = ~n39564 ;
  assign y13895 = ~n39566 ;
  assign y13896 = ~1'b0 ;
  assign y13897 = ~n39567 ;
  assign y13898 = n39575 ;
  assign y13899 = ~1'b0 ;
  assign y13900 = ~1'b0 ;
  assign y13901 = ~1'b0 ;
  assign y13902 = ~n39580 ;
  assign y13903 = ~n6267 ;
  assign y13904 = n39582 ;
  assign y13905 = n39584 ;
  assign y13906 = n39586 ;
  assign y13907 = ~n39590 ;
  assign y13908 = ~n39595 ;
  assign y13909 = n39599 ;
  assign y13910 = ~n39602 ;
  assign y13911 = n39608 ;
  assign y13912 = n39609 ;
  assign y13913 = ~n39615 ;
  assign y13914 = ~n39616 ;
  assign y13915 = n39621 ;
  assign y13916 = ~n39626 ;
  assign y13917 = ~1'b0 ;
  assign y13918 = n8234 ;
  assign y13919 = n39627 ;
  assign y13920 = ~n39628 ;
  assign y13921 = n39630 ;
  assign y13922 = ~1'b0 ;
  assign y13923 = ~1'b0 ;
  assign y13924 = n39631 ;
  assign y13925 = ~n39632 ;
  assign y13926 = n39633 ;
  assign y13927 = n39634 ;
  assign y13928 = n39635 ;
  assign y13929 = ~n39637 ;
  assign y13930 = n39643 ;
  assign y13931 = ~1'b0 ;
  assign y13932 = ~1'b0 ;
  assign y13933 = ~n39646 ;
  assign y13934 = n39647 ;
  assign y13935 = n39657 ;
  assign y13936 = ~n39661 ;
  assign y13937 = ~n39665 ;
  assign y13938 = n39668 ;
  assign y13939 = ~1'b0 ;
  assign y13940 = n39669 ;
  assign y13941 = ~n39671 ;
  assign y13942 = ~n39673 ;
  assign y13943 = ~n39674 ;
  assign y13944 = ~n39675 ;
  assign y13945 = n39677 ;
  assign y13946 = ~1'b0 ;
  assign y13947 = ~n39679 ;
  assign y13948 = ~n39685 ;
  assign y13949 = n39689 ;
  assign y13950 = ~n39693 ;
  assign y13951 = ~n39694 ;
  assign y13952 = n39695 ;
  assign y13953 = ~1'b0 ;
  assign y13954 = n39697 ;
  assign y13955 = n39701 ;
  assign y13956 = n39702 ;
  assign y13957 = ~n39704 ;
  assign y13958 = n39710 ;
  assign y13959 = ~n39714 ;
  assign y13960 = n39725 ;
  assign y13961 = n39732 ;
  assign y13962 = ~n39734 ;
  assign y13963 = ~n39735 ;
  assign y13964 = ~n39738 ;
  assign y13965 = n39741 ;
  assign y13966 = n39744 ;
  assign y13967 = ~1'b0 ;
  assign y13968 = ~1'b0 ;
  assign y13969 = n39745 ;
  assign y13970 = ~n39746 ;
  assign y13971 = n39748 ;
  assign y13972 = ~n39749 ;
  assign y13973 = n39752 ;
  assign y13974 = ~1'b0 ;
  assign y13975 = n39758 ;
  assign y13976 = ~n39759 ;
  assign y13977 = n39760 ;
  assign y13978 = ~n39765 ;
  assign y13979 = ~n39766 ;
  assign y13980 = n39770 ;
  assign y13981 = n39777 ;
  assign y13982 = n39779 ;
  assign y13983 = ~1'b0 ;
  assign y13984 = ~n39782 ;
  assign y13985 = ~n39785 ;
  assign y13986 = ~n39790 ;
  assign y13987 = n39793 ;
  assign y13988 = n39794 ;
  assign y13989 = ~n39795 ;
  assign y13990 = ~n39796 ;
  assign y13991 = ~n39798 ;
  assign y13992 = n39800 ;
  assign y13993 = ~n39801 ;
  assign y13994 = ~1'b0 ;
  assign y13995 = ~n39803 ;
  assign y13996 = n39806 ;
  assign y13997 = n39811 ;
  assign y13998 = ~1'b0 ;
  assign y13999 = ~n39812 ;
  assign y14000 = ~1'b0 ;
  assign y14001 = n39818 ;
  assign y14002 = ~n39819 ;
  assign y14003 = ~n39820 ;
  assign y14004 = n39822 ;
  assign y14005 = ~n39827 ;
  assign y14006 = ~n39831 ;
  assign y14007 = ~n35705 ;
  assign y14008 = ~1'b0 ;
  assign y14009 = n39834 ;
  assign y14010 = ~n39835 ;
  assign y14011 = ~n39841 ;
  assign y14012 = n39842 ;
  assign y14013 = ~1'b0 ;
  assign y14014 = ~1'b0 ;
  assign y14015 = n39846 ;
  assign y14016 = ~1'b0 ;
  assign y14017 = ~1'b0 ;
  assign y14018 = n39849 ;
  assign y14019 = ~n39850 ;
  assign y14020 = n39851 ;
  assign y14021 = ~n39852 ;
  assign y14022 = n39853 ;
  assign y14023 = n39854 ;
  assign y14024 = ~n39856 ;
  assign y14025 = n39857 ;
  assign y14026 = ~n39860 ;
  assign y14027 = ~n39862 ;
  assign y14028 = ~n39866 ;
  assign y14029 = ~n39867 ;
  assign y14030 = n39868 ;
  assign y14031 = n39869 ;
  assign y14032 = ~n39870 ;
  assign y14033 = ~n39871 ;
  assign y14034 = ~n39874 ;
  assign y14035 = ~1'b0 ;
  assign y14036 = n39877 ;
  assign y14037 = n39878 ;
  assign y14038 = n39879 ;
  assign y14039 = n25760 ;
  assign y14040 = ~1'b0 ;
  assign y14041 = ~n39881 ;
  assign y14042 = ~1'b0 ;
  assign y14043 = ~1'b0 ;
  assign y14044 = n39897 ;
  assign y14045 = ~n39898 ;
  assign y14046 = n39899 ;
  assign y14047 = ~n39902 ;
  assign y14048 = n39903 ;
  assign y14049 = ~1'b0 ;
  assign y14050 = ~n39908 ;
  assign y14051 = ~1'b0 ;
  assign y14052 = n19645 ;
  assign y14053 = ~n39910 ;
  assign y14054 = n39911 ;
  assign y14055 = n39912 ;
  assign y14056 = n39913 ;
  assign y14057 = n39915 ;
  assign y14058 = n39918 ;
  assign y14059 = ~1'b0 ;
  assign y14060 = ~1'b0 ;
  assign y14061 = ~n39925 ;
  assign y14062 = ~n39926 ;
  assign y14063 = ~n39935 ;
  assign y14064 = n26485 ;
  assign y14065 = n39939 ;
  assign y14066 = n39946 ;
  assign y14067 = n39951 ;
  assign y14068 = ~n27617 ;
  assign y14069 = ~n39957 ;
  assign y14070 = ~n39958 ;
  assign y14071 = n39967 ;
  assign y14072 = n39976 ;
  assign y14073 = ~n39980 ;
  assign y14074 = ~n39981 ;
  assign y14075 = n9788 ;
  assign y14076 = ~1'b0 ;
  assign y14077 = n39982 ;
  assign y14078 = ~n39985 ;
  assign y14079 = n39986 ;
  assign y14080 = n39992 ;
  assign y14081 = ~1'b0 ;
  assign y14082 = n39994 ;
  assign y14083 = ~1'b0 ;
  assign y14084 = ~n39998 ;
  assign y14085 = ~1'b0 ;
  assign y14086 = n40004 ;
  assign y14087 = ~n40006 ;
  assign y14088 = ~n40008 ;
  assign y14089 = ~n40010 ;
  assign y14090 = ~n40011 ;
  assign y14091 = ~1'b0 ;
  assign y14092 = n40012 ;
  assign y14093 = ~n40013 ;
  assign y14094 = ~n40014 ;
  assign y14095 = ~n40019 ;
  assign y14096 = ~1'b0 ;
  assign y14097 = ~1'b0 ;
  assign y14098 = n40020 ;
  assign y14099 = ~n40022 ;
  assign y14100 = ~n40028 ;
  assign y14101 = ~1'b0 ;
  assign y14102 = ~n40031 ;
  assign y14103 = ~n40033 ;
  assign y14104 = ~n40036 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = n40038 ;
  assign y14107 = n40044 ;
  assign y14108 = ~n40045 ;
  assign y14109 = n40046 ;
  assign y14110 = ~1'b0 ;
  assign y14111 = ~n40050 ;
  assign y14112 = ~n40054 ;
  assign y14113 = ~1'b0 ;
  assign y14114 = ~1'b0 ;
  assign y14115 = n40056 ;
  assign y14116 = n40060 ;
  assign y14117 = n40062 ;
  assign y14118 = ~n40066 ;
  assign y14119 = ~1'b0 ;
  assign y14120 = ~n40069 ;
  assign y14121 = ~n40072 ;
  assign y14122 = n40075 ;
  assign y14123 = ~n40077 ;
  assign y14124 = ~n40079 ;
  assign y14125 = n40081 ;
  assign y14126 = n40083 ;
  assign y14127 = n40085 ;
  assign y14128 = ~n40088 ;
  assign y14129 = ~n40089 ;
  assign y14130 = ~n40091 ;
  assign y14131 = n40093 ;
  assign y14132 = ~1'b0 ;
  assign y14133 = ~1'b0 ;
  assign y14134 = ~n40094 ;
  assign y14135 = ~n40096 ;
  assign y14136 = ~n40101 ;
  assign y14137 = n40103 ;
  assign y14138 = ~n40105 ;
  assign y14139 = ~1'b0 ;
  assign y14140 = ~1'b0 ;
  assign y14141 = n40111 ;
  assign y14142 = ~n40113 ;
  assign y14143 = n40114 ;
  assign y14144 = n40116 ;
  assign y14145 = ~n40117 ;
  assign y14146 = n40121 ;
  assign y14147 = n40122 ;
  assign y14148 = n40126 ;
  assign y14149 = ~n40129 ;
  assign y14150 = ~n40132 ;
  assign y14151 = ~n1337 ;
  assign y14152 = n40135 ;
  assign y14153 = ~1'b0 ;
  assign y14154 = n40137 ;
  assign y14155 = ~1'b0 ;
  assign y14156 = n40143 ;
  assign y14157 = ~n40144 ;
  assign y14158 = ~n40148 ;
  assign y14159 = ~n40151 ;
  assign y14160 = ~n40153 ;
  assign y14161 = ~1'b0 ;
  assign y14162 = n40155 ;
  assign y14163 = ~n40160 ;
  assign y14164 = n40162 ;
  assign y14165 = ~n40163 ;
  assign y14166 = ~n40169 ;
  assign y14167 = ~n40175 ;
  assign y14168 = n40177 ;
  assign y14169 = ~1'b0 ;
  assign y14170 = ~n40178 ;
  assign y14171 = n40183 ;
  assign y14172 = ~n40185 ;
  assign y14173 = n40190 ;
  assign y14174 = ~n40198 ;
  assign y14175 = ~n40199 ;
  assign y14176 = ~n40206 ;
  assign y14177 = ~1'b0 ;
  assign y14178 = ~n40208 ;
  assign y14179 = n40212 ;
  assign y14180 = ~1'b0 ;
  assign y14181 = n40214 ;
  assign y14182 = ~n40215 ;
  assign y14183 = ~n40217 ;
  assign y14184 = ~n40218 ;
  assign y14185 = n40221 ;
  assign y14186 = ~1'b0 ;
  assign y14187 = n40226 ;
  assign y14188 = ~1'b0 ;
  assign y14189 = ~n40228 ;
  assign y14190 = ~n40231 ;
  assign y14191 = ~n40242 ;
  assign y14192 = ~n40244 ;
  assign y14193 = n40245 ;
  assign y14194 = n40248 ;
  assign y14195 = ~n27510 ;
  assign y14196 = ~n40250 ;
  assign y14197 = n40251 ;
  assign y14198 = ~n40255 ;
  assign y14199 = ~n40259 ;
  assign y14200 = n8307 ;
  assign y14201 = n40261 ;
  assign y14202 = n40264 ;
  assign y14203 = n40266 ;
  assign y14204 = ~n40269 ;
  assign y14205 = n40273 ;
  assign y14206 = ~n40277 ;
  assign y14207 = n40279 ;
  assign y14208 = n40283 ;
  assign y14209 = ~n40290 ;
  assign y14210 = ~n40291 ;
  assign y14211 = ~1'b0 ;
  assign y14212 = ~n40296 ;
  assign y14213 = n40310 ;
  assign y14214 = n40311 ;
  assign y14215 = ~n40315 ;
  assign y14216 = ~n40323 ;
  assign y14217 = n40324 ;
  assign y14218 = ~1'b0 ;
  assign y14219 = ~1'b0 ;
  assign y14220 = ~n40325 ;
  assign y14221 = n40327 ;
  assign y14222 = n40329 ;
  assign y14223 = ~n40336 ;
  assign y14224 = n40337 ;
  assign y14225 = ~n40338 ;
  assign y14226 = ~n40340 ;
  assign y14227 = ~n40342 ;
  assign y14228 = ~n40345 ;
  assign y14229 = ~n40346 ;
  assign y14230 = n40348 ;
  assign y14231 = n23762 ;
  assign y14232 = ~n40351 ;
  assign y14233 = n7004 ;
  assign y14234 = ~n40353 ;
  assign y14235 = ~n40354 ;
  assign y14236 = ~1'b0 ;
  assign y14237 = ~n40355 ;
  assign y14238 = n40357 ;
  assign y14239 = n40359 ;
  assign y14240 = ~n40360 ;
  assign y14241 = n40365 ;
  assign y14242 = n40367 ;
  assign y14243 = ~n40370 ;
  assign y14244 = ~1'b0 ;
  assign y14245 = n40374 ;
  assign y14246 = ~n40375 ;
  assign y14247 = n40378 ;
  assign y14248 = n40380 ;
  assign y14249 = ~n40382 ;
  assign y14250 = n40387 ;
  assign y14251 = ~1'b0 ;
  assign y14252 = ~n11227 ;
  assign y14253 = ~n40388 ;
  assign y14254 = ~n40390 ;
  assign y14255 = n40391 ;
  assign y14256 = n40392 ;
  assign y14257 = n40398 ;
  assign y14258 = ~n18414 ;
  assign y14259 = ~1'b0 ;
  assign y14260 = ~1'b0 ;
  assign y14261 = ~n40400 ;
  assign y14262 = ~n40402 ;
  assign y14263 = n40403 ;
  assign y14264 = ~n40405 ;
  assign y14265 = ~n40406 ;
  assign y14266 = n40408 ;
  assign y14267 = 1'b0 ;
  assign y14268 = ~n40414 ;
  assign y14269 = ~n40417 ;
  assign y14270 = n40418 ;
  assign y14271 = ~1'b0 ;
  assign y14272 = n40421 ;
  assign y14273 = n40422 ;
  assign y14274 = n40424 ;
  assign y14275 = n40426 ;
  assign y14276 = n40427 ;
  assign y14277 = ~n40429 ;
  assign y14278 = ~1'b0 ;
  assign y14279 = ~n40433 ;
  assign y14280 = ~n40435 ;
  assign y14281 = ~n40436 ;
  assign y14282 = ~n40437 ;
  assign y14283 = ~n40438 ;
  assign y14284 = ~1'b0 ;
  assign y14285 = ~1'b0 ;
  assign y14286 = ~n40441 ;
  assign y14287 = n40446 ;
  assign y14288 = n40447 ;
  assign y14289 = ~n40450 ;
  assign y14290 = ~n40451 ;
  assign y14291 = n40452 ;
  assign y14292 = ~n40455 ;
  assign y14293 = ~n40457 ;
  assign y14294 = ~n40463 ;
  assign y14295 = n40464 ;
  assign y14296 = n40468 ;
  assign y14297 = n40469 ;
  assign y14298 = ~n40472 ;
  assign y14299 = ~n40473 ;
  assign y14300 = ~n40474 ;
  assign y14301 = ~n40480 ;
  assign y14302 = n40483 ;
  assign y14303 = ~1'b0 ;
  assign y14304 = ~1'b0 ;
  assign y14305 = ~n40487 ;
  assign y14306 = ~n40489 ;
  assign y14307 = n40491 ;
  assign y14308 = ~n40492 ;
  assign y14309 = ~n40498 ;
  assign y14310 = ~n40502 ;
  assign y14311 = ~1'b0 ;
  assign y14312 = n40503 ;
  assign y14313 = ~n40506 ;
  assign y14314 = n40509 ;
  assign y14315 = n40510 ;
  assign y14316 = n40518 ;
  assign y14317 = ~n40522 ;
  assign y14318 = n18579 ;
  assign y14319 = ~n40527 ;
  assign y14320 = ~n40529 ;
  assign y14321 = ~n40531 ;
  assign y14322 = n40534 ;
  assign y14323 = n17576 ;
  assign y14324 = ~n40539 ;
  assign y14325 = n40545 ;
  assign y14326 = ~n40548 ;
  assign y14327 = n40550 ;
  assign y14328 = ~1'b0 ;
  assign y14329 = n40551 ;
  assign y14330 = n40552 ;
  assign y14331 = ~n40554 ;
  assign y14332 = ~n40557 ;
  assign y14333 = n40559 ;
  assign y14334 = ~1'b0 ;
  assign y14335 = n40561 ;
  assign y14336 = ~n40563 ;
  assign y14337 = ~1'b0 ;
  assign y14338 = n40564 ;
  assign y14339 = ~n40574 ;
  assign y14340 = ~1'b0 ;
  assign y14341 = n40576 ;
  assign y14342 = ~n40582 ;
  assign y14343 = n40585 ;
  assign y14344 = ~n40586 ;
  assign y14345 = n40587 ;
  assign y14346 = n40588 ;
  assign y14347 = n40592 ;
  assign y14348 = ~n40595 ;
  assign y14349 = n40596 ;
  assign y14350 = ~n40601 ;
  assign y14351 = n40603 ;
  assign y14352 = n40605 ;
  assign y14353 = ~1'b0 ;
  assign y14354 = n40606 ;
  assign y14355 = n40611 ;
  assign y14356 = ~n40615 ;
  assign y14357 = ~n40622 ;
  assign y14358 = n40623 ;
  assign y14359 = n40626 ;
  assign y14360 = n40628 ;
  assign y14361 = ~1'b0 ;
  assign y14362 = ~n40631 ;
  assign y14363 = ~n40632 ;
  assign y14364 = n40634 ;
  assign y14365 = n40638 ;
  assign y14366 = ~n40645 ;
  assign y14367 = ~n40649 ;
  assign y14368 = ~n40653 ;
  assign y14369 = n40656 ;
  assign y14370 = ~n40660 ;
  assign y14371 = ~1'b0 ;
  assign y14372 = n40661 ;
  assign y14373 = n40662 ;
  assign y14374 = ~n40667 ;
  assign y14375 = ~1'b0 ;
  assign y14376 = ~n40673 ;
  assign y14377 = ~n40674 ;
  assign y14378 = ~n40676 ;
  assign y14379 = ~1'b0 ;
  assign y14380 = n40679 ;
  assign y14381 = ~n40689 ;
  assign y14382 = ~n40690 ;
  assign y14383 = ~n40691 ;
  assign y14384 = n40698 ;
  assign y14385 = ~1'b0 ;
  assign y14386 = ~n40699 ;
  assign y14387 = ~1'b0 ;
  assign y14388 = ~1'b0 ;
  assign y14389 = ~1'b0 ;
  assign y14390 = ~n40700 ;
  assign y14391 = n40702 ;
  assign y14392 = ~n40703 ;
  assign y14393 = n40715 ;
  assign y14394 = n40718 ;
  assign y14395 = n40719 ;
  assign y14396 = ~1'b0 ;
  assign y14397 = n40720 ;
  assign y14398 = ~n40723 ;
  assign y14399 = ~n40726 ;
  assign y14400 = n40736 ;
  assign y14401 = ~n40738 ;
  assign y14402 = n40742 ;
  assign y14403 = ~n40745 ;
  assign y14404 = n40746 ;
  assign y14405 = ~n40754 ;
  assign y14406 = ~n40755 ;
  assign y14407 = ~n40757 ;
  assign y14408 = ~n40765 ;
  assign y14409 = ~n40767 ;
  assign y14410 = n40768 ;
  assign y14411 = ~n40774 ;
  assign y14412 = ~1'b0 ;
  assign y14413 = n40780 ;
  assign y14414 = n40788 ;
  assign y14415 = ~n40791 ;
  assign y14416 = ~n40794 ;
  assign y14417 = ~n40798 ;
  assign y14418 = n40801 ;
  assign y14419 = n40802 ;
  assign y14420 = ~1'b0 ;
  assign y14421 = n40807 ;
  assign y14422 = ~n40812 ;
  assign y14423 = ~n40814 ;
  assign y14424 = n40816 ;
  assign y14425 = n40817 ;
  assign y14426 = ~n40820 ;
  assign y14427 = ~n40821 ;
  assign y14428 = ~n40826 ;
  assign y14429 = ~n40828 ;
  assign y14430 = ~n40830 ;
  assign y14431 = ~n40831 ;
  assign y14432 = n40832 ;
  assign y14433 = n40837 ;
  assign y14434 = n40838 ;
  assign y14435 = n40842 ;
  assign y14436 = n40843 ;
  assign y14437 = ~n40847 ;
  assign y14438 = n40852 ;
  assign y14439 = n40858 ;
  assign y14440 = n40864 ;
  assign y14441 = ~1'b0 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = ~1'b0 ;
  assign y14444 = ~n40865 ;
  assign y14445 = ~n40867 ;
  assign y14446 = ~n40871 ;
  assign y14447 = n40874 ;
  assign y14448 = n40880 ;
  assign y14449 = ~1'b0 ;
  assign y14450 = n40882 ;
  assign y14451 = ~1'b0 ;
  assign y14452 = n40890 ;
  assign y14453 = ~1'b0 ;
  assign y14454 = n40891 ;
  assign y14455 = n40892 ;
  assign y14456 = n40893 ;
  assign y14457 = ~n40894 ;
  assign y14458 = ~1'b0 ;
  assign y14459 = n40895 ;
  assign y14460 = ~1'b0 ;
  assign y14461 = ~n40897 ;
  assign y14462 = ~n40899 ;
  assign y14463 = n40900 ;
  assign y14464 = ~n40904 ;
  assign y14465 = ~n40908 ;
  assign y14466 = ~n40909 ;
  assign y14467 = n40911 ;
  assign y14468 = ~n40912 ;
  assign y14469 = ~n40916 ;
  assign y14470 = ~n40919 ;
  assign y14471 = ~n40921 ;
  assign y14472 = n40927 ;
  assign y14473 = ~1'b0 ;
  assign y14474 = ~n40930 ;
  assign y14475 = ~1'b0 ;
  assign y14476 = n40936 ;
  assign y14477 = ~n40937 ;
  assign y14478 = ~n40939 ;
  assign y14479 = ~1'b0 ;
  assign y14480 = ~1'b0 ;
  assign y14481 = n40941 ;
  assign y14482 = n40943 ;
  assign y14483 = ~n40947 ;
  assign y14484 = ~n40950 ;
  assign y14485 = n40952 ;
  assign y14486 = ~1'b0 ;
  assign y14487 = n40955 ;
  assign y14488 = ~1'b0 ;
  assign y14489 = ~1'b0 ;
  assign y14490 = n40956 ;
  assign y14491 = ~1'b0 ;
  assign y14492 = ~n40957 ;
  assign y14493 = ~n40958 ;
  assign y14494 = n40963 ;
  assign y14495 = ~n40967 ;
  assign y14496 = ~n40972 ;
  assign y14497 = n40974 ;
  assign y14498 = n40978 ;
  assign y14499 = ~n40980 ;
  assign y14500 = n40984 ;
  assign y14501 = n40986 ;
  assign y14502 = ~n40988 ;
  assign y14503 = ~n40992 ;
  assign y14504 = ~n40993 ;
  assign y14505 = ~n40995 ;
  assign y14506 = ~n40996 ;
  assign y14507 = ~n40999 ;
  assign y14508 = ~n41002 ;
  assign y14509 = ~n41006 ;
  assign y14510 = n41008 ;
  assign y14511 = ~n41009 ;
  assign y14512 = ~n41010 ;
  assign y14513 = n41011 ;
  assign y14514 = n6788 ;
  assign y14515 = n41013 ;
  assign y14516 = ~1'b0 ;
  assign y14517 = n18257 ;
  assign y14518 = ~n41015 ;
  assign y14519 = ~n41018 ;
  assign y14520 = n41020 ;
  assign y14521 = ~n41024 ;
  assign y14522 = ~n41027 ;
  assign y14523 = n41035 ;
  assign y14524 = ~n41037 ;
  assign y14525 = n41041 ;
  assign y14526 = ~n41043 ;
  assign y14527 = n41047 ;
  assign y14528 = ~n41048 ;
  assign y14529 = n41049 ;
  assign y14530 = ~n41051 ;
  assign y14531 = ~1'b0 ;
  assign y14532 = ~n41058 ;
  assign y14533 = n41061 ;
  assign y14534 = n17538 ;
  assign y14535 = n41063 ;
  assign y14536 = ~n41064 ;
  assign y14537 = ~1'b0 ;
  assign y14538 = ~n41066 ;
  assign y14539 = ~1'b0 ;
  assign y14540 = ~n41072 ;
  assign y14541 = ~n41073 ;
  assign y14542 = ~n41076 ;
  assign y14543 = ~n41078 ;
  assign y14544 = ~n41082 ;
  assign y14545 = ~n41085 ;
  assign y14546 = n41087 ;
  assign y14547 = ~n41090 ;
  assign y14548 = ~n41095 ;
  assign y14549 = n41096 ;
  assign y14550 = n41097 ;
  assign y14551 = n41102 ;
  assign y14552 = n41105 ;
  assign y14553 = ~1'b0 ;
  assign y14554 = n41108 ;
  assign y14555 = n41113 ;
  assign y14556 = n41116 ;
  assign y14557 = ~n41117 ;
  assign y14558 = n41118 ;
  assign y14559 = ~n41119 ;
  assign y14560 = ~n41121 ;
  assign y14561 = n41122 ;
  assign y14562 = ~n41123 ;
  assign y14563 = ~n41129 ;
  assign y14564 = ~n41134 ;
  assign y14565 = n41136 ;
  assign y14566 = n41137 ;
  assign y14567 = ~n41141 ;
  assign y14568 = ~n41145 ;
  assign y14569 = ~n41147 ;
  assign y14570 = ~n41154 ;
  assign y14571 = ~n41163 ;
  assign y14572 = ~n41166 ;
  assign y14573 = n41167 ;
  assign y14574 = n41170 ;
  assign y14575 = n41175 ;
  assign y14576 = n41177 ;
  assign y14577 = ~1'b0 ;
  assign y14578 = n41180 ;
  assign y14579 = ~n41185 ;
  assign y14580 = n41187 ;
  assign y14581 = n41188 ;
  assign y14582 = n41191 ;
  assign y14583 = n41193 ;
  assign y14584 = ~n41196 ;
  assign y14585 = n41201 ;
  assign y14586 = ~n41206 ;
  assign y14587 = n41207 ;
  assign y14588 = n41209 ;
  assign y14589 = ~1'b0 ;
  assign y14590 = n41216 ;
  assign y14591 = ~n41217 ;
  assign y14592 = ~1'b0 ;
  assign y14593 = n41218 ;
  assign y14594 = n41219 ;
  assign y14595 = ~1'b0 ;
  assign y14596 = ~1'b0 ;
  assign y14597 = ~1'b0 ;
  assign y14598 = ~1'b0 ;
  assign y14599 = n41220 ;
  assign y14600 = n41222 ;
  assign y14601 = ~n41223 ;
  assign y14602 = ~n41226 ;
  assign y14603 = ~n41229 ;
  assign y14604 = n41231 ;
  assign y14605 = ~1'b0 ;
  assign y14606 = n41235 ;
  assign y14607 = ~n41237 ;
  assign y14608 = n41240 ;
  assign y14609 = n41241 ;
  assign y14610 = n41243 ;
  assign y14611 = ~n41244 ;
  assign y14612 = ~n41246 ;
  assign y14613 = n41249 ;
  assign y14614 = n41254 ;
  assign y14615 = ~n35869 ;
  assign y14616 = ~n41258 ;
  assign y14617 = n41260 ;
  assign y14618 = ~n41264 ;
  assign y14619 = n41266 ;
  assign y14620 = n41267 ;
  assign y14621 = ~n41271 ;
  assign y14622 = ~1'b0 ;
  assign y14623 = ~n41275 ;
  assign y14624 = n41278 ;
  assign y14625 = n41280 ;
  assign y14626 = ~n41282 ;
  assign y14627 = ~n41283 ;
  assign y14628 = ~1'b0 ;
  assign y14629 = ~n41284 ;
  assign y14630 = ~1'b0 ;
  assign y14631 = n41286 ;
  assign y14632 = ~n41290 ;
  assign y14633 = ~n41291 ;
  assign y14634 = ~1'b0 ;
  assign y14635 = n41296 ;
  assign y14636 = ~n41297 ;
  assign y14637 = n41301 ;
  assign y14638 = ~n41304 ;
  assign y14639 = ~n41305 ;
  assign y14640 = n41307 ;
  assign y14641 = ~n41312 ;
  assign y14642 = ~1'b0 ;
  assign y14643 = n41315 ;
  assign y14644 = ~n41316 ;
  assign y14645 = n41317 ;
  assign y14646 = n41319 ;
  assign y14647 = ~n41321 ;
  assign y14648 = n41324 ;
  assign y14649 = ~1'b0 ;
  assign y14650 = ~n41329 ;
  assign y14651 = n41331 ;
  assign y14652 = ~n41333 ;
  assign y14653 = n41334 ;
  assign y14654 = n41340 ;
  assign y14655 = ~1'b0 ;
  assign y14656 = ~n41342 ;
  assign y14657 = n41345 ;
  assign y14658 = ~1'b0 ;
  assign y14659 = ~n41351 ;
  assign y14660 = n41352 ;
  assign y14661 = ~n41356 ;
  assign y14662 = n41357 ;
  assign y14663 = ~n41359 ;
  assign y14664 = n41363 ;
  assign y14665 = ~n41364 ;
  assign y14666 = n41366 ;
  assign y14667 = 1'b0 ;
  assign y14668 = n41373 ;
  assign y14669 = n41374 ;
  assign y14670 = n41376 ;
  assign y14671 = n41379 ;
  assign y14672 = ~1'b0 ;
  assign y14673 = n41380 ;
  assign y14674 = ~1'b0 ;
  assign y14675 = n41381 ;
  assign y14676 = ~n41382 ;
  assign y14677 = n41388 ;
  assign y14678 = ~n41394 ;
  assign y14679 = n41395 ;
  assign y14680 = ~n41397 ;
  assign y14681 = ~1'b0 ;
  assign y14682 = ~1'b0 ;
  assign y14683 = n41399 ;
  assign y14684 = n41400 ;
  assign y14685 = n41401 ;
  assign y14686 = ~n41405 ;
  assign y14687 = n41406 ;
  assign y14688 = ~n41411 ;
  assign y14689 = ~1'b0 ;
  assign y14690 = ~1'b0 ;
  assign y14691 = ~n41412 ;
  assign y14692 = n41413 ;
  assign y14693 = ~n41416 ;
  assign y14694 = ~n41417 ;
  assign y14695 = n41421 ;
  assign y14696 = ~n41422 ;
  assign y14697 = n41423 ;
  assign y14698 = ~n41424 ;
  assign y14699 = n41427 ;
  assign y14700 = n41429 ;
  assign y14701 = ~n41431 ;
  assign y14702 = ~1'b0 ;
  assign y14703 = ~n41434 ;
  assign y14704 = ~n41435 ;
  assign y14705 = n41438 ;
  assign y14706 = ~n41439 ;
  assign y14707 = n41441 ;
  assign y14708 = ~n41444 ;
  assign y14709 = n41446 ;
  assign y14710 = ~n41449 ;
  assign y14711 = n41451 ;
  assign y14712 = n41452 ;
  assign y14713 = ~n41455 ;
  assign y14714 = ~n41456 ;
  assign y14715 = n22354 ;
  assign y14716 = n41459 ;
  assign y14717 = ~1'b0 ;
  assign y14718 = n41462 ;
  assign y14719 = ~n41465 ;
  assign y14720 = n41466 ;
  assign y14721 = n41467 ;
  assign y14722 = ~n41468 ;
  assign y14723 = n41472 ;
  assign y14724 = ~1'b0 ;
  assign y14725 = ~n41476 ;
  assign y14726 = ~n41479 ;
  assign y14727 = n41481 ;
  assign y14728 = n41483 ;
  assign y14729 = n41488 ;
  assign y14730 = n41491 ;
  assign y14731 = n41492 ;
  assign y14732 = ~n41495 ;
  assign y14733 = n41499 ;
  assign y14734 = n19616 ;
  assign y14735 = n41501 ;
  assign y14736 = ~n41507 ;
  assign y14737 = ~n41508 ;
  assign y14738 = n41509 ;
  assign y14739 = n41513 ;
  assign y14740 = n41514 ;
  assign y14741 = ~n41515 ;
  assign y14742 = ~n41516 ;
  assign y14743 = ~n41518 ;
  assign y14744 = ~1'b0 ;
  assign y14745 = ~n41520 ;
  assign y14746 = ~1'b0 ;
  assign y14747 = ~n41523 ;
  assign y14748 = ~n41524 ;
  assign y14749 = ~n41526 ;
  assign y14750 = n41527 ;
  assign y14751 = ~n41529 ;
  assign y14752 = ~n41533 ;
  assign y14753 = n41534 ;
  assign y14754 = ~1'b0 ;
  assign y14755 = ~n41535 ;
  assign y14756 = n41538 ;
  assign y14757 = n41544 ;
  assign y14758 = ~n41546 ;
  assign y14759 = ~n41547 ;
  assign y14760 = n41550 ;
  assign y14761 = ~1'b0 ;
  assign y14762 = n41551 ;
  assign y14763 = ~n41552 ;
  assign y14764 = n41561 ;
  assign y14765 = n41565 ;
  assign y14766 = n41566 ;
  assign y14767 = ~n41568 ;
  assign y14768 = ~1'b0 ;
  assign y14769 = ~1'b0 ;
  assign y14770 = n41571 ;
  assign y14771 = ~n41572 ;
  assign y14772 = ~n41573 ;
  assign y14773 = n41576 ;
  assign y14774 = n41578 ;
  assign y14775 = n41580 ;
  assign y14776 = ~1'b0 ;
  assign y14777 = ~1'b0 ;
  assign y14778 = ~n41583 ;
  assign y14779 = n41592 ;
  assign y14780 = ~n41593 ;
  assign y14781 = n41594 ;
  assign y14782 = n41595 ;
  assign y14783 = ~n41597 ;
  assign y14784 = n41601 ;
  assign y14785 = ~1'b0 ;
  assign y14786 = ~1'b0 ;
  assign y14787 = ~1'b0 ;
  assign y14788 = ~1'b0 ;
  assign y14789 = ~n41602 ;
  assign y14790 = n41604 ;
  assign y14791 = ~n41606 ;
  assign y14792 = n41608 ;
  assign y14793 = ~n41614 ;
  assign y14794 = n41615 ;
  assign y14795 = n41617 ;
  assign y14796 = ~n41619 ;
  assign y14797 = ~n41622 ;
  assign y14798 = n41624 ;
  assign y14799 = n41628 ;
  assign y14800 = n5687 ;
  assign y14801 = n41630 ;
  assign y14802 = n12687 ;
  assign y14803 = ~n41633 ;
  assign y14804 = ~n41635 ;
  assign y14805 = n41638 ;
  assign y14806 = n41640 ;
  assign y14807 = n41641 ;
  assign y14808 = n41643 ;
  assign y14809 = ~n41647 ;
  assign y14810 = n41648 ;
  assign y14811 = n41650 ;
  assign y14812 = n41651 ;
  assign y14813 = ~n41653 ;
  assign y14814 = ~n41655 ;
  assign y14815 = ~n41657 ;
  assign y14816 = ~1'b0 ;
  assign y14817 = n41658 ;
  assign y14818 = n35819 ;
  assign y14819 = n41659 ;
  assign y14820 = n41663 ;
  assign y14821 = n41668 ;
  assign y14822 = ~n41671 ;
  assign y14823 = ~n41675 ;
  assign y14824 = n41679 ;
  assign y14825 = ~n41680 ;
  assign y14826 = n41681 ;
  assign y14827 = ~1'b0 ;
  assign y14828 = ~1'b0 ;
  assign y14829 = n41684 ;
  assign y14830 = n41689 ;
  assign y14831 = n41691 ;
  assign y14832 = n41695 ;
  assign y14833 = ~n41696 ;
  assign y14834 = ~n41697 ;
  assign y14835 = ~n41700 ;
  assign y14836 = ~n41701 ;
  assign y14837 = n41704 ;
  assign y14838 = ~1'b0 ;
  assign y14839 = n41706 ;
  assign y14840 = n41708 ;
  assign y14841 = ~1'b0 ;
  assign y14842 = ~n41710 ;
  assign y14843 = n41715 ;
  assign y14844 = n41716 ;
  assign y14845 = n41718 ;
  assign y14846 = ~n41719 ;
  assign y14847 = ~n41724 ;
  assign y14848 = ~n41726 ;
  assign y14849 = n41728 ;
  assign y14850 = ~1'b0 ;
  assign y14851 = ~n41729 ;
  assign y14852 = n41730 ;
  assign y14853 = n9947 ;
  assign y14854 = n41731 ;
  assign y14855 = n41732 ;
  assign y14856 = ~1'b0 ;
  assign y14857 = ~n41734 ;
  assign y14858 = ~1'b0 ;
  assign y14859 = n41735 ;
  assign y14860 = n41736 ;
  assign y14861 = n41739 ;
  assign y14862 = ~n41740 ;
  assign y14863 = ~n22563 ;
  assign y14864 = n41743 ;
  assign y14865 = ~n41747 ;
  assign y14866 = n41754 ;
  assign y14867 = ~n41756 ;
  assign y14868 = ~n41757 ;
  assign y14869 = ~n41759 ;
  assign y14870 = n41760 ;
  assign y14871 = n41762 ;
  assign y14872 = ~n41765 ;
  assign y14873 = ~1'b0 ;
  assign y14874 = ~n41770 ;
  assign y14875 = ~1'b0 ;
  assign y14876 = n961 ;
  assign y14877 = n41772 ;
  assign y14878 = ~n41775 ;
  assign y14879 = n41779 ;
  assign y14880 = n41780 ;
  assign y14881 = n10650 ;
  assign y14882 = n41782 ;
  assign y14883 = ~1'b0 ;
  assign y14884 = n41783 ;
  assign y14885 = ~n41787 ;
  assign y14886 = ~n41790 ;
  assign y14887 = ~n41794 ;
  assign y14888 = n41795 ;
  assign y14889 = n41796 ;
  assign y14890 = n41799 ;
  assign y14891 = ~1'b0 ;
  assign y14892 = ~1'b0 ;
  assign y14893 = ~n41805 ;
  assign y14894 = ~1'b0 ;
  assign y14895 = ~n41807 ;
  assign y14896 = n41808 ;
  assign y14897 = n41811 ;
  assign y14898 = ~x76 ;
  assign y14899 = ~n41812 ;
  assign y14900 = ~n41817 ;
  assign y14901 = ~1'b0 ;
  assign y14902 = ~1'b0 ;
  assign y14903 = ~n41819 ;
  assign y14904 = ~n41822 ;
  assign y14905 = n41825 ;
  assign y14906 = n41826 ;
  assign y14907 = ~n41830 ;
  assign y14908 = n41831 ;
  assign y14909 = ~n41833 ;
  assign y14910 = n41836 ;
  assign y14911 = ~1'b0 ;
  assign y14912 = n19285 ;
  assign y14913 = n41837 ;
  assign y14914 = ~n41839 ;
  assign y14915 = n41845 ;
  assign y14916 = ~n41848 ;
  assign y14917 = ~n41852 ;
  assign y14918 = ~1'b0 ;
  assign y14919 = n41853 ;
  assign y14920 = ~1'b0 ;
  assign y14921 = n41854 ;
  assign y14922 = ~n6856 ;
  assign y14923 = ~n41855 ;
  assign y14924 = ~n41856 ;
  assign y14925 = ~1'b0 ;
  assign y14926 = ~1'b0 ;
  assign y14927 = ~n41858 ;
  assign y14928 = n41859 ;
  assign y14929 = ~n41860 ;
  assign y14930 = n41861 ;
  assign y14931 = ~n41862 ;
  assign y14932 = ~n41863 ;
  assign y14933 = ~n41864 ;
  assign y14934 = ~n41868 ;
  assign y14935 = ~n41871 ;
  assign y14936 = ~1'b0 ;
  assign y14937 = n41873 ;
  assign y14938 = ~n41875 ;
  assign y14939 = ~n41876 ;
  assign y14940 = n41877 ;
  assign y14941 = n41883 ;
  assign y14942 = ~n41885 ;
  assign y14943 = ~1'b0 ;
  assign y14944 = ~1'b0 ;
  assign y14945 = n41889 ;
  assign y14946 = ~n41890 ;
  assign y14947 = ~n41894 ;
  assign y14948 = ~n41898 ;
  assign y14949 = ~1'b0 ;
  assign y14950 = ~n41901 ;
  assign y14951 = n41902 ;
  assign y14952 = n41903 ;
  assign y14953 = ~n41906 ;
  assign y14954 = n41908 ;
  assign y14955 = n41914 ;
  assign y14956 = ~n41917 ;
  assign y14957 = ~n41918 ;
  assign y14958 = ~n32606 ;
  assign y14959 = ~n41920 ;
  assign y14960 = ~n41921 ;
  assign y14961 = n41923 ;
  assign y14962 = n34192 ;
  assign y14963 = ~n41927 ;
  assign y14964 = ~n41928 ;
  assign y14965 = ~n41929 ;
  assign y14966 = n41933 ;
  assign y14967 = ~n20372 ;
  assign y14968 = ~1'b0 ;
  assign y14969 = ~1'b0 ;
  assign y14970 = ~n41935 ;
  assign y14971 = n41938 ;
  assign y14972 = ~n41939 ;
  assign y14973 = ~n41940 ;
  assign y14974 = ~n41941 ;
  assign y14975 = ~n41943 ;
  assign y14976 = n41946 ;
  assign y14977 = n41948 ;
  assign y14978 = ~1'b0 ;
  assign y14979 = ~n41949 ;
  assign y14980 = ~n41951 ;
  assign y14981 = n41956 ;
  assign y14982 = n41961 ;
  assign y14983 = ~n41964 ;
  assign y14984 = ~n41971 ;
  assign y14985 = n41973 ;
  assign y14986 = ~n41976 ;
  assign y14987 = n41977 ;
  assign y14988 = ~n41980 ;
  assign y14989 = ~n41985 ;
  assign y14990 = ~n41990 ;
  assign y14991 = n41993 ;
  assign y14992 = n41994 ;
  assign y14993 = ~n41995 ;
  assign y14994 = ~n41998 ;
  assign y14995 = n40227 ;
  assign y14996 = ~n42002 ;
  assign y14997 = ~n42004 ;
  assign y14998 = ~n42007 ;
  assign y14999 = n42010 ;
  assign y15000 = n42012 ;
  assign y15001 = n42013 ;
  assign y15002 = n42019 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = ~1'b0 ;
  assign y15005 = n42025 ;
  assign y15006 = ~1'b0 ;
  assign y15007 = ~n42028 ;
  assign y15008 = n42032 ;
  assign y15009 = ~n42033 ;
  assign y15010 = ~n42035 ;
  assign y15011 = ~n42037 ;
  assign y15012 = n42042 ;
  assign y15013 = ~n42044 ;
  assign y15014 = n42047 ;
  assign y15015 = ~n42052 ;
  assign y15016 = ~n42055 ;
  assign y15017 = n42056 ;
  assign y15018 = n42060 ;
  assign y15019 = n42064 ;
  assign y15020 = ~1'b0 ;
  assign y15021 = n42066 ;
  assign y15022 = ~1'b0 ;
  assign y15023 = ~1'b0 ;
  assign y15024 = n42069 ;
  assign y15025 = n42072 ;
  assign y15026 = n42073 ;
  assign y15027 = n42074 ;
  assign y15028 = n42077 ;
  assign y15029 = ~1'b0 ;
  assign y15030 = ~1'b0 ;
  assign y15031 = n42080 ;
  assign y15032 = n42085 ;
  assign y15033 = n42089 ;
  assign y15034 = ~n42091 ;
  assign y15035 = ~n42101 ;
  assign y15036 = ~n42104 ;
  assign y15037 = ~n42106 ;
  assign y15038 = n42108 ;
  assign y15039 = ~1'b0 ;
  assign y15040 = n42112 ;
  assign y15041 = ~n42114 ;
  assign y15042 = ~n42121 ;
  assign y15043 = ~n42124 ;
  assign y15044 = ~n42126 ;
  assign y15045 = n42129 ;
  assign y15046 = n42136 ;
  assign y15047 = ~1'b0 ;
  assign y15048 = ~1'b0 ;
  assign y15049 = n42138 ;
  assign y15050 = ~1'b0 ;
  assign y15051 = n42139 ;
  assign y15052 = n42142 ;
  assign y15053 = n42147 ;
  assign y15054 = n42149 ;
  assign y15055 = ~n42151 ;
  assign y15056 = n42153 ;
  assign y15057 = ~1'b0 ;
  assign y15058 = ~n42155 ;
  assign y15059 = ~n42159 ;
  assign y15060 = n42162 ;
  assign y15061 = n42163 ;
  assign y15062 = ~n42165 ;
  assign y15063 = ~1'b0 ;
  assign y15064 = ~1'b0 ;
  assign y15065 = n42167 ;
  assign y15066 = ~n42168 ;
  assign y15067 = ~n42171 ;
  assign y15068 = ~n42172 ;
  assign y15069 = n42174 ;
  assign y15070 = ~n42179 ;
  assign y15071 = ~1'b0 ;
  assign y15072 = ~n42184 ;
  assign y15073 = n42187 ;
  assign y15074 = n42189 ;
  assign y15075 = n42192 ;
  assign y15076 = ~n42203 ;
  assign y15077 = ~n42208 ;
  assign y15078 = ~n42210 ;
  assign y15079 = n42211 ;
  assign y15080 = n42213 ;
  assign y15081 = ~n42217 ;
  assign y15082 = ~n42219 ;
  assign y15083 = n42222 ;
  assign y15084 = ~n42223 ;
  assign y15085 = ~n42225 ;
  assign y15086 = ~n42230 ;
  assign y15087 = ~n42236 ;
  assign y15088 = ~1'b0 ;
  assign y15089 = ~1'b0 ;
  assign y15090 = n42240 ;
  assign y15091 = ~n42250 ;
  assign y15092 = n42251 ;
  assign y15093 = n42252 ;
  assign y15094 = ~n42254 ;
  assign y15095 = n10779 ;
  assign y15096 = ~1'b0 ;
  assign y15097 = ~n42255 ;
  assign y15098 = n42256 ;
  assign y15099 = n42257 ;
  assign y15100 = ~n42259 ;
  assign y15101 = ~n42262 ;
  assign y15102 = ~1'b0 ;
  assign y15103 = n42264 ;
  assign y15104 = ~n42270 ;
  assign y15105 = ~n42272 ;
  assign y15106 = n42275 ;
  assign y15107 = n42279 ;
  assign y15108 = ~1'b0 ;
  assign y15109 = ~n42281 ;
  assign y15110 = n42285 ;
  assign y15111 = ~1'b0 ;
  assign y15112 = ~n42288 ;
  assign y15113 = ~n42291 ;
  assign y15114 = ~n42292 ;
  assign y15115 = ~n42295 ;
  assign y15116 = n42298 ;
  assign y15117 = ~n42299 ;
  assign y15118 = ~1'b0 ;
  assign y15119 = ~n42303 ;
  assign y15120 = ~1'b0 ;
  assign y15121 = ~1'b0 ;
  assign y15122 = n42304 ;
  assign y15123 = n42305 ;
  assign y15124 = ~n42306 ;
  assign y15125 = ~n42310 ;
  assign y15126 = ~n42311 ;
  assign y15127 = ~n42313 ;
  assign y15128 = n42314 ;
  assign y15129 = n42316 ;
  assign y15130 = ~1'b0 ;
  assign y15131 = n42320 ;
  assign y15132 = ~n42321 ;
  assign y15133 = ~1'b0 ;
  assign y15134 = ~n42324 ;
  assign y15135 = ~n42329 ;
  assign y15136 = ~n42331 ;
  assign y15137 = n42333 ;
  assign y15138 = ~n42338 ;
  assign y15139 = ~n42347 ;
  assign y15140 = ~n42355 ;
  assign y15141 = ~n42357 ;
  assign y15142 = ~n6689 ;
  assign y15143 = ~1'b0 ;
  assign y15144 = ~n42366 ;
  assign y15145 = n42368 ;
  assign y15146 = ~1'b0 ;
  assign y15147 = n42373 ;
  assign y15148 = ~n42375 ;
  assign y15149 = n42377 ;
  assign y15150 = ~n42378 ;
  assign y15151 = ~n42382 ;
  assign y15152 = ~1'b0 ;
  assign y15153 = ~1'b0 ;
  assign y15154 = ~n42385 ;
  assign y15155 = ~n42387 ;
  assign y15156 = ~n42388 ;
  assign y15157 = n42391 ;
  assign y15158 = ~n26846 ;
  assign y15159 = n42399 ;
  assign y15160 = ~1'b0 ;
  assign y15161 = ~1'b0 ;
  assign y15162 = n42401 ;
  assign y15163 = ~1'b0 ;
  assign y15164 = n42402 ;
  assign y15165 = ~n41806 ;
  assign y15166 = n42403 ;
  assign y15167 = ~n42405 ;
  assign y15168 = ~n42407 ;
  assign y15169 = ~1'b0 ;
  assign y15170 = ~1'b0 ;
  assign y15171 = n42412 ;
  assign y15172 = n42417 ;
  assign y15173 = n42420 ;
  assign y15174 = ~1'b0 ;
  assign y15175 = ~n42425 ;
  assign y15176 = n42427 ;
  assign y15177 = n42429 ;
  assign y15178 = ~n42430 ;
  assign y15179 = n42431 ;
  assign y15180 = ~n42432 ;
  assign y15181 = ~n42433 ;
  assign y15182 = n42436 ;
  assign y15183 = ~1'b0 ;
  assign y15184 = ~n42444 ;
  assign y15185 = n42448 ;
  assign y15186 = ~n42459 ;
  assign y15187 = ~n2319 ;
  assign y15188 = n42460 ;
  assign y15189 = n42463 ;
  assign y15190 = ~n42465 ;
  assign y15191 = ~1'b0 ;
  assign y15192 = ~n42466 ;
  assign y15193 = n42470 ;
  assign y15194 = n42471 ;
  assign y15195 = ~n42475 ;
  assign y15196 = ~n42476 ;
  assign y15197 = n42477 ;
  assign y15198 = n42479 ;
  assign y15199 = ~1'b0 ;
  assign y15200 = n42481 ;
  assign y15201 = 1'b0 ;
  assign y15202 = ~1'b0 ;
  assign y15203 = ~n42482 ;
  assign y15204 = ~n42485 ;
  assign y15205 = ~n42486 ;
  assign y15206 = ~1'b0 ;
  assign y15207 = ~1'b0 ;
  assign y15208 = n42490 ;
  assign y15209 = ~n42492 ;
  assign y15210 = 1'b0 ;
  assign y15211 = n42493 ;
  assign y15212 = ~n42502 ;
  assign y15213 = ~n42503 ;
  assign y15214 = n42509 ;
  assign y15215 = n42510 ;
  assign y15216 = n42513 ;
  assign y15217 = ~1'b0 ;
  assign y15218 = ~1'b0 ;
  assign y15219 = ~n42514 ;
  assign y15220 = ~n42517 ;
  assign y15221 = ~n42519 ;
  assign y15222 = n42520 ;
  assign y15223 = n42523 ;
  assign y15224 = ~n42524 ;
  assign y15225 = ~n42526 ;
  assign y15226 = ~1'b0 ;
  assign y15227 = ~1'b0 ;
  assign y15228 = ~n42527 ;
  assign y15229 = n42529 ;
  assign y15230 = ~n36031 ;
  assign y15231 = ~n42531 ;
  assign y15232 = ~1'b0 ;
  assign y15233 = ~n42535 ;
  assign y15234 = ~1'b0 ;
  assign y15235 = ~n42539 ;
  assign y15236 = n42544 ;
  assign y15237 = n42546 ;
  assign y15238 = ~n42547 ;
  assign y15239 = n42551 ;
  assign y15240 = ~n42554 ;
  assign y15241 = ~n42555 ;
  assign y15242 = ~n42557 ;
  assign y15243 = ~n42559 ;
  assign y15244 = ~1'b0 ;
  assign y15245 = ~n42561 ;
  assign y15246 = ~n42564 ;
  assign y15247 = n42565 ;
  assign y15248 = ~n42567 ;
  assign y15249 = ~n42568 ;
  assign y15250 = ~n42571 ;
  assign y15251 = n42573 ;
  assign y15252 = ~n42574 ;
  assign y15253 = ~n42575 ;
  assign y15254 = ~n42579 ;
  assign y15255 = ~n42581 ;
  assign y15256 = ~n42584 ;
  assign y15257 = n42587 ;
  assign y15258 = ~1'b0 ;
  assign y15259 = ~1'b0 ;
  assign y15260 = ~1'b0 ;
  assign y15261 = n42589 ;
  assign y15262 = ~n42590 ;
  assign y15263 = n42591 ;
  assign y15264 = ~n42592 ;
  assign y15265 = ~n42598 ;
  assign y15266 = n42600 ;
  assign y15267 = n42601 ;
  assign y15268 = n42603 ;
  assign y15269 = n42606 ;
  assign y15270 = ~n42609 ;
  assign y15271 = ~1'b0 ;
  assign y15272 = ~n42611 ;
  assign y15273 = ~n42614 ;
  assign y15274 = ~n42615 ;
  assign y15275 = n42617 ;
  assign y15276 = n42618 ;
  assign y15277 = n42620 ;
  assign y15278 = ~1'b0 ;
  assign y15279 = ~n42622 ;
  assign y15280 = n6244 ;
  assign y15281 = n42624 ;
  assign y15282 = n42625 ;
  assign y15283 = n42627 ;
  assign y15284 = ~n29215 ;
  assign y15285 = n42628 ;
  assign y15286 = n42630 ;
  assign y15287 = ~n42632 ;
  assign y15288 = ~n42635 ;
  assign y15289 = n42638 ;
  assign y15290 = ~n42640 ;
  assign y15291 = n42641 ;
  assign y15292 = n42643 ;
  assign y15293 = ~n42645 ;
  assign y15294 = ~n42647 ;
  assign y15295 = ~n42650 ;
  assign y15296 = ~1'b0 ;
  assign y15297 = n42652 ;
  assign y15298 = ~n42655 ;
  assign y15299 = ~1'b0 ;
  assign y15300 = n42662 ;
  assign y15301 = ~n42666 ;
  assign y15302 = ~n42667 ;
  assign y15303 = ~n42669 ;
  assign y15304 = n42671 ;
  assign y15305 = ~1'b0 ;
  assign y15306 = n42674 ;
  assign y15307 = n42679 ;
  assign y15308 = ~n42683 ;
  assign y15309 = n42684 ;
  assign y15310 = ~n42685 ;
  assign y15311 = ~n42686 ;
  assign y15312 = n42687 ;
  assign y15313 = n42688 ;
  assign y15314 = ~1'b0 ;
  assign y15315 = ~1'b0 ;
  assign y15316 = ~n42690 ;
  assign y15317 = ~1'b0 ;
  assign y15318 = n42691 ;
  assign y15319 = n42692 ;
  assign y15320 = n42697 ;
  assign y15321 = n42702 ;
  assign y15322 = ~n42704 ;
  assign y15323 = ~n42705 ;
  assign y15324 = ~n42710 ;
  assign y15325 = ~n42714 ;
  assign y15326 = ~n42716 ;
  assign y15327 = n42719 ;
  assign y15328 = n42721 ;
  assign y15329 = ~n42722 ;
  assign y15330 = ~n42727 ;
  assign y15331 = ~n42732 ;
  assign y15332 = n42733 ;
  assign y15333 = n42734 ;
  assign y15334 = ~1'b0 ;
  assign y15335 = 1'b0 ;
  assign y15336 = n42742 ;
  assign y15337 = ~n42743 ;
  assign y15338 = ~n42746 ;
  assign y15339 = ~n42752 ;
  assign y15340 = ~n42756 ;
  assign y15341 = ~n42762 ;
  assign y15342 = ~n42765 ;
  assign y15343 = ~n42769 ;
  assign y15344 = ~n42773 ;
  assign y15345 = ~n42775 ;
  assign y15346 = n42780 ;
  assign y15347 = ~n42786 ;
  assign y15348 = ~1'b0 ;
  assign y15349 = ~n42791 ;
  assign y15350 = ~n42793 ;
  assign y15351 = ~n42795 ;
  assign y15352 = ~n42798 ;
  assign y15353 = ~1'b0 ;
  assign y15354 = n42799 ;
  assign y15355 = n42802 ;
  assign y15356 = ~n42804 ;
  assign y15357 = n42807 ;
  assign y15358 = ~n42808 ;
  assign y15359 = ~n42814 ;
  assign y15360 = ~1'b0 ;
  assign y15361 = ~1'b0 ;
  assign y15362 = n42819 ;
  assign y15363 = ~n42823 ;
  assign y15364 = n42824 ;
  assign y15365 = n42825 ;
  assign y15366 = n42834 ;
  assign y15367 = n42835 ;
  assign y15368 = n42838 ;
  assign y15369 = ~1'b0 ;
  assign y15370 = ~1'b0 ;
  assign y15371 = ~n42843 ;
  assign y15372 = ~1'b0 ;
  assign y15373 = ~n42844 ;
  assign y15374 = ~n42845 ;
  assign y15375 = ~n42848 ;
  assign y15376 = n42849 ;
  assign y15377 = n42851 ;
  assign y15378 = ~n42854 ;
  assign y15379 = n42857 ;
  assign y15380 = n42860 ;
  assign y15381 = ~1'b0 ;
  assign y15382 = ~n42865 ;
  assign y15383 = ~n42867 ;
  assign y15384 = ~n42868 ;
  assign y15385 = ~n42869 ;
  assign y15386 = ~n42872 ;
  assign y15387 = ~1'b0 ;
  assign y15388 = n42873 ;
  assign y15389 = ~n42877 ;
  assign y15390 = ~n42879 ;
  assign y15391 = n42882 ;
  assign y15392 = n42883 ;
  assign y15393 = n42887 ;
  assign y15394 = ~n42891 ;
  assign y15395 = ~n42900 ;
  assign y15396 = ~n42902 ;
  assign y15397 = ~1'b0 ;
  assign y15398 = ~n42906 ;
  assign y15399 = ~n42907 ;
  assign y15400 = ~n42908 ;
  assign y15401 = n42911 ;
  assign y15402 = ~1'b0 ;
  assign y15403 = ~n42912 ;
  assign y15404 = ~1'b0 ;
  assign y15405 = ~n42915 ;
  assign y15406 = n42916 ;
  assign y15407 = ~n42917 ;
  assign y15408 = n42921 ;
  assign y15409 = ~n42932 ;
  assign y15410 = ~n42933 ;
  assign y15411 = n42942 ;
  assign y15412 = ~1'b0 ;
  assign y15413 = ~n42943 ;
  assign y15414 = ~n42955 ;
  assign y15415 = n42956 ;
  assign y15416 = ~n42959 ;
  assign y15417 = n42960 ;
  assign y15418 = ~n42962 ;
  assign y15419 = ~1'b0 ;
  assign y15420 = ~1'b0 ;
  assign y15421 = n42964 ;
  assign y15422 = n42970 ;
  assign y15423 = ~n42972 ;
  assign y15424 = n42975 ;
  assign y15425 = ~n42976 ;
  assign y15426 = ~n42979 ;
  assign y15427 = ~n42980 ;
  assign y15428 = n42982 ;
  assign y15429 = ~n42986 ;
  assign y15430 = ~1'b0 ;
  assign y15431 = ~n42988 ;
  assign y15432 = n42992 ;
  assign y15433 = n42995 ;
  assign y15434 = n20638 ;
  assign y15435 = ~n42998 ;
  assign y15436 = n42999 ;
  assign y15437 = n43002 ;
  assign y15438 = ~n43005 ;
  assign y15439 = ~1'b0 ;
  assign y15440 = ~n43009 ;
  assign y15441 = ~1'b0 ;
  assign y15442 = ~1'b0 ;
  assign y15443 = n43012 ;
  assign y15444 = ~n43014 ;
  assign y15445 = ~n43016 ;
  assign y15446 = n43021 ;
  assign y15447 = ~1'b0 ;
  assign y15448 = ~n43023 ;
  assign y15449 = ~n43024 ;
  assign y15450 = n43025 ;
  assign y15451 = ~n43026 ;
  assign y15452 = n43029 ;
  assign y15453 = ~1'b0 ;
  assign y15454 = ~1'b0 ;
  assign y15455 = ~n43033 ;
  assign y15456 = n43035 ;
  assign y15457 = ~n43036 ;
  assign y15458 = ~n43037 ;
  assign y15459 = n43038 ;
  assign y15460 = ~n43039 ;
  assign y15461 = ~1'b0 ;
  assign y15462 = ~1'b0 ;
  assign y15463 = n43041 ;
  assign y15464 = ~n43048 ;
  assign y15465 = n43052 ;
  assign y15466 = n43055 ;
  assign y15467 = n43058 ;
  assign y15468 = ~n43061 ;
  assign y15469 = ~n43062 ;
  assign y15470 = ~n43064 ;
  assign y15471 = ~1'b0 ;
  assign y15472 = ~n43065 ;
  assign y15473 = ~1'b0 ;
  assign y15474 = n43066 ;
  assign y15475 = ~n3359 ;
  assign y15476 = ~n43068 ;
  assign y15477 = n43071 ;
  assign y15478 = ~n43073 ;
  assign y15479 = ~n43076 ;
  assign y15480 = ~n43081 ;
  assign y15481 = n43083 ;
  assign y15482 = ~n43084 ;
  assign y15483 = ~1'b0 ;
  assign y15484 = n43086 ;
  assign y15485 = n43088 ;
  assign y15486 = ~n43089 ;
  assign y15487 = ~n43090 ;
  assign y15488 = ~n43092 ;
  assign y15489 = ~n43095 ;
  assign y15490 = ~n43101 ;
  assign y15491 = ~1'b0 ;
  assign y15492 = ~1'b0 ;
  assign y15493 = n43102 ;
  assign y15494 = ~n43104 ;
  assign y15495 = n43109 ;
  assign y15496 = n43111 ;
  assign y15497 = ~n43112 ;
  assign y15498 = n43116 ;
  assign y15499 = n43118 ;
  assign y15500 = ~n43124 ;
  assign y15501 = ~1'b0 ;
  assign y15502 = n43127 ;
  assign y15503 = ~n43135 ;
  assign y15504 = ~n43136 ;
  assign y15505 = ~n43141 ;
  assign y15506 = ~1'b0 ;
  assign y15507 = ~n43149 ;
  assign y15508 = n43150 ;
  assign y15509 = ~n43153 ;
  assign y15510 = n43154 ;
  assign y15511 = ~n43158 ;
  assign y15512 = ~n43159 ;
  assign y15513 = ~1'b0 ;
  assign y15514 = ~1'b0 ;
  assign y15515 = ~1'b0 ;
  assign y15516 = ~n43163 ;
  assign y15517 = n43171 ;
  assign y15518 = ~n43174 ;
  assign y15519 = ~n43177 ;
  assign y15520 = ~n43184 ;
  assign y15521 = ~n43185 ;
  assign y15522 = n43187 ;
  assign y15523 = ~1'b0 ;
  assign y15524 = ~n43189 ;
  assign y15525 = ~n43191 ;
  assign y15526 = ~n43193 ;
  assign y15527 = n43198 ;
  assign y15528 = n43203 ;
  assign y15529 = ~n43204 ;
  assign y15530 = ~n43205 ;
  assign y15531 = ~n43209 ;
  assign y15532 = n43211 ;
  assign y15533 = ~n43214 ;
  assign y15534 = ~1'b0 ;
  assign y15535 = ~n43219 ;
  assign y15536 = ~n43224 ;
  assign y15537 = ~n28407 ;
  assign y15538 = n43225 ;
  assign y15539 = n43230 ;
  assign y15540 = n43235 ;
  assign y15541 = n43236 ;
  assign y15542 = n43241 ;
  assign y15543 = n43245 ;
  assign y15544 = ~1'b0 ;
  assign y15545 = n43249 ;
  assign y15546 = n43251 ;
  assign y15547 = ~n43252 ;
  assign y15548 = n43253 ;
  assign y15549 = n43254 ;
  assign y15550 = ~n43255 ;
  assign y15551 = n43256 ;
  assign y15552 = ~n41286 ;
  assign y15553 = ~1'b0 ;
  assign y15554 = n43257 ;
  assign y15555 = ~n43261 ;
  assign y15556 = n43262 ;
  assign y15557 = ~n43263 ;
  assign y15558 = ~n43264 ;
  assign y15559 = n43266 ;
  assign y15560 = ~1'b0 ;
  assign y15561 = ~1'b0 ;
  assign y15562 = n43267 ;
  assign y15563 = n43268 ;
  assign y15564 = n43273 ;
  assign y15565 = ~n43274 ;
  assign y15566 = n43276 ;
  assign y15567 = ~1'b0 ;
  assign y15568 = ~n43278 ;
  assign y15569 = n43283 ;
  assign y15570 = n43287 ;
  assign y15571 = ~n43290 ;
  assign y15572 = ~n43291 ;
  assign y15573 = ~n43292 ;
  assign y15574 = ~n43295 ;
  assign y15575 = n43297 ;
  assign y15576 = n43300 ;
  assign y15577 = n43303 ;
  assign y15578 = ~n43309 ;
  assign y15579 = n43310 ;
  assign y15580 = ~n43311 ;
  assign y15581 = ~n43312 ;
  assign y15582 = ~n43313 ;
  assign y15583 = ~1'b0 ;
  assign y15584 = ~1'b0 ;
  assign y15585 = n43317 ;
  assign y15586 = n43318 ;
  assign y15587 = n43325 ;
  assign y15588 = ~n43326 ;
  assign y15589 = n43327 ;
  assign y15590 = n43328 ;
  assign y15591 = ~n43329 ;
  assign y15592 = ~n43334 ;
  assign y15593 = ~n43336 ;
  assign y15594 = n43337 ;
  assign y15595 = ~1'b0 ;
  assign y15596 = n43339 ;
  assign y15597 = ~n43343 ;
  assign y15598 = ~n43344 ;
  assign y15599 = ~n43352 ;
  assign y15600 = n43360 ;
  assign y15601 = ~1'b0 ;
  assign y15602 = ~n43362 ;
  assign y15603 = n43364 ;
  assign y15604 = ~1'b0 ;
  assign y15605 = ~n43365 ;
  assign y15606 = ~n43367 ;
  assign y15607 = ~n43368 ;
  assign y15608 = ~n36931 ;
  assign y15609 = n43369 ;
  assign y15610 = ~n43370 ;
  assign y15611 = n43372 ;
  assign y15612 = ~n43374 ;
  assign y15613 = ~n43376 ;
  assign y15614 = n473 ;
  assign y15615 = ~n43378 ;
  assign y15616 = n43379 ;
  assign y15617 = n43380 ;
  assign y15618 = n43382 ;
  assign y15619 = n43384 ;
  assign y15620 = ~n43386 ;
  assign y15621 = ~1'b0 ;
  assign y15622 = ~n43389 ;
  assign y15623 = ~n43391 ;
  assign y15624 = n43392 ;
  assign y15625 = n43394 ;
  assign y15626 = n43398 ;
  assign y15627 = n43407 ;
  assign y15628 = n43409 ;
  assign y15629 = ~1'b0 ;
  assign y15630 = n43411 ;
  assign y15631 = n43415 ;
  assign y15632 = n43421 ;
  assign y15633 = ~n43423 ;
  assign y15634 = n43424 ;
  assign y15635 = ~n43426 ;
  assign y15636 = ~1'b0 ;
  assign y15637 = ~1'b0 ;
  assign y15638 = ~1'b0 ;
  assign y15639 = n43429 ;
  assign y15640 = ~1'b0 ;
  assign y15641 = ~n43430 ;
  assign y15642 = n43431 ;
  assign y15643 = n43432 ;
  assign y15644 = n43434 ;
  assign y15645 = n43435 ;
  assign y15646 = ~1'b0 ;
  assign y15647 = n43436 ;
  assign y15648 = ~n43439 ;
  assign y15649 = ~n43444 ;
  assign y15650 = ~1'b0 ;
  assign y15651 = n43446 ;
  assign y15652 = n43447 ;
  assign y15653 = ~n43450 ;
  assign y15654 = n43452 ;
  assign y15655 = n43453 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = n8595 ;
  assign y15658 = ~n43454 ;
  assign y15659 = ~1'b0 ;
  assign y15660 = n43456 ;
  assign y15661 = ~n5953 ;
  assign y15662 = ~n43458 ;
  assign y15663 = ~n43466 ;
  assign y15664 = ~n43470 ;
  assign y15665 = n43471 ;
  assign y15666 = n43475 ;
  assign y15667 = n43477 ;
  assign y15668 = ~n43479 ;
  assign y15669 = ~n43481 ;
  assign y15670 = ~n43482 ;
  assign y15671 = n43486 ;
  assign y15672 = ~1'b0 ;
  assign y15673 = ~n43491 ;
  assign y15674 = ~1'b0 ;
  assign y15675 = n43492 ;
  assign y15676 = n43495 ;
  assign y15677 = ~n43496 ;
  assign y15678 = n43497 ;
  assign y15679 = ~n43500 ;
  assign y15680 = ~n43503 ;
  assign y15681 = ~1'b0 ;
  assign y15682 = ~1'b0 ;
  assign y15683 = ~1'b0 ;
  assign y15684 = ~1'b0 ;
  assign y15685 = ~n43505 ;
  assign y15686 = ~n43506 ;
  assign y15687 = ~n43508 ;
  assign y15688 = n43509 ;
  assign y15689 = n43516 ;
  assign y15690 = ~n43518 ;
  assign y15691 = ~n43521 ;
  assign y15692 = ~n43523 ;
  assign y15693 = ~1'b0 ;
  assign y15694 = ~n43524 ;
  assign y15695 = ~n43526 ;
  assign y15696 = ~n43528 ;
  assign y15697 = n43531 ;
  assign y15698 = ~n43534 ;
  assign y15699 = ~n43539 ;
  assign y15700 = n43547 ;
  assign y15701 = n43549 ;
  assign y15702 = ~1'b0 ;
  assign y15703 = n43550 ;
  assign y15704 = n43551 ;
  assign y15705 = ~n43553 ;
  assign y15706 = n43555 ;
  assign y15707 = ~n43556 ;
  assign y15708 = ~1'b0 ;
  assign y15709 = n43558 ;
  assign y15710 = ~1'b0 ;
  assign y15711 = ~n43559 ;
  assign y15712 = ~n3958 ;
  assign y15713 = ~n43562 ;
  assign y15714 = n43564 ;
  assign y15715 = n43565 ;
  assign y15716 = ~n43567 ;
  assign y15717 = n43574 ;
  assign y15718 = ~1'b0 ;
  assign y15719 = n43579 ;
  assign y15720 = n43580 ;
  assign y15721 = ~n43582 ;
  assign y15722 = ~n43585 ;
  assign y15723 = ~n43589 ;
  assign y15724 = ~n43591 ;
  assign y15725 = n43593 ;
  assign y15726 = n43595 ;
  assign y15727 = ~n43598 ;
  assign y15728 = ~n43601 ;
  assign y15729 = ~n43602 ;
  assign y15730 = ~n43606 ;
  assign y15731 = n43607 ;
  assign y15732 = ~n43608 ;
  assign y15733 = 1'b0 ;
  assign y15734 = ~n43610 ;
  assign y15735 = ~1'b0 ;
  assign y15736 = n43612 ;
  assign y15737 = ~1'b0 ;
  assign y15738 = ~n43613 ;
  assign y15739 = ~n43615 ;
  assign y15740 = ~n43616 ;
  assign y15741 = n43618 ;
  assign y15742 = ~n43619 ;
  assign y15743 = ~n43622 ;
  assign y15744 = ~n43625 ;
  assign y15745 = n43627 ;
  assign y15746 = ~1'b0 ;
  assign y15747 = ~1'b0 ;
  assign y15748 = ~n43629 ;
  assign y15749 = n43632 ;
  assign y15750 = ~n43633 ;
  assign y15751 = n43634 ;
  assign y15752 = n43635 ;
  assign y15753 = ~n43638 ;
  assign y15754 = ~n43641 ;
  assign y15755 = ~1'b0 ;
  assign y15756 = n43644 ;
  assign y15757 = ~1'b0 ;
  assign y15758 = n43646 ;
  assign y15759 = n43648 ;
  assign y15760 = n43651 ;
  assign y15761 = ~n43653 ;
  assign y15762 = ~n43655 ;
  assign y15763 = n38286 ;
  assign y15764 = ~1'b0 ;
  assign y15765 = ~n43658 ;
  assign y15766 = ~n43660 ;
  assign y15767 = ~n43661 ;
  assign y15768 = n43667 ;
  assign y15769 = n43668 ;
  assign y15770 = n43673 ;
  assign y15771 = ~n43683 ;
  assign y15772 = ~n43686 ;
  assign y15773 = n43687 ;
  assign y15774 = n43688 ;
  assign y15775 = n43689 ;
  assign y15776 = ~n43692 ;
  assign y15777 = ~1'b0 ;
  assign y15778 = n43693 ;
  assign y15779 = ~1'b0 ;
  assign y15780 = ~1'b0 ;
  assign y15781 = ~1'b0 ;
  assign y15782 = ~n43694 ;
  assign y15783 = ~n43697 ;
  assign y15784 = ~n43700 ;
  assign y15785 = n43702 ;
  assign y15786 = ~n43708 ;
  assign y15787 = ~1'b0 ;
  assign y15788 = ~1'b0 ;
  assign y15789 = n43709 ;
  assign y15790 = ~n43710 ;
  assign y15791 = n43714 ;
  assign y15792 = n43715 ;
  assign y15793 = n43718 ;
  assign y15794 = ~n43723 ;
  assign y15795 = n43726 ;
  assign y15796 = n43733 ;
  assign y15797 = ~n43736 ;
  assign y15798 = ~n43745 ;
  assign y15799 = n43747 ;
  assign y15800 = ~n43748 ;
  assign y15801 = ~n43755 ;
  assign y15802 = n43756 ;
  assign y15803 = n43759 ;
  assign y15804 = ~n43761 ;
  assign y15805 = ~n43765 ;
  assign y15806 = ~1'b0 ;
  assign y15807 = ~n43769 ;
  assign y15808 = n43770 ;
  assign y15809 = n43773 ;
  assign y15810 = ~n43781 ;
  assign y15811 = n43783 ;
  assign y15812 = ~n31551 ;
  assign y15813 = ~1'b0 ;
  assign y15814 = ~n43787 ;
  assign y15815 = ~1'b0 ;
  assign y15816 = n43789 ;
  assign y15817 = ~n43792 ;
  assign y15818 = ~1'b0 ;
  assign y15819 = ~1'b0 ;
  assign y15820 = n43794 ;
  assign y15821 = n14177 ;
  assign y15822 = n43804 ;
  assign y15823 = n43805 ;
  assign y15824 = ~n22348 ;
  assign y15825 = ~1'b0 ;
  assign y15826 = 1'b0 ;
  assign y15827 = ~1'b0 ;
  assign y15828 = ~1'b0 ;
  assign y15829 = ~n43807 ;
  assign y15830 = ~n43809 ;
  assign y15831 = n43810 ;
  assign y15832 = ~n43813 ;
  assign y15833 = n43815 ;
  assign y15834 = ~n43817 ;
  assign y15835 = ~n43820 ;
  assign y15836 = ~n43822 ;
  assign y15837 = n43824 ;
  assign y15838 = n43831 ;
  assign y15839 = n43834 ;
  assign y15840 = n43835 ;
  assign y15841 = ~1'b0 ;
  assign y15842 = ~1'b0 ;
  assign y15843 = ~n43838 ;
  assign y15844 = ~n43839 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = n43842 ;
  assign y15847 = n43848 ;
  assign y15848 = ~n43849 ;
  assign y15849 = ~n43850 ;
  assign y15850 = ~n43851 ;
  assign y15851 = ~1'b0 ;
  assign y15852 = ~n43855 ;
  assign y15853 = n43857 ;
  assign y15854 = ~1'b0 ;
  assign y15855 = ~1'b0 ;
  assign y15856 = ~1'b0 ;
  assign y15857 = n43859 ;
  assign y15858 = ~n43864 ;
  assign y15859 = ~n43867 ;
  assign y15860 = ~n43868 ;
  assign y15861 = ~n43869 ;
  assign y15862 = ~n43873 ;
  assign y15863 = n43876 ;
  assign y15864 = ~1'b0 ;
  assign y15865 = n43879 ;
  assign y15866 = n43880 ;
  assign y15867 = ~n43884 ;
  assign y15868 = ~n43885 ;
  assign y15869 = n43886 ;
  assign y15870 = ~n43888 ;
  assign y15871 = ~n43890 ;
  assign y15872 = ~1'b0 ;
  assign y15873 = ~n43895 ;
  assign y15874 = ~1'b0 ;
  assign y15875 = n43898 ;
  assign y15876 = ~n43900 ;
  assign y15877 = n43901 ;
  assign y15878 = n43904 ;
  assign y15879 = n43907 ;
  assign y15880 = n43908 ;
  assign y15881 = ~n43909 ;
  assign y15882 = n43913 ;
  assign y15883 = ~1'b0 ;
  assign y15884 = n43914 ;
  assign y15885 = n43915 ;
  assign y15886 = ~n43920 ;
  assign y15887 = ~n4343 ;
  assign y15888 = ~n43923 ;
  assign y15889 = n43924 ;
  assign y15890 = ~n43927 ;
  assign y15891 = ~1'b0 ;
  assign y15892 = ~n43929 ;
  assign y15893 = ~n43931 ;
  assign y15894 = n43932 ;
  assign y15895 = n43933 ;
  assign y15896 = ~n43934 ;
  assign y15897 = n43935 ;
  assign y15898 = n43939 ;
  assign y15899 = ~1'b0 ;
  assign y15900 = n43941 ;
  assign y15901 = n43943 ;
  assign y15902 = n11748 ;
  assign y15903 = ~1'b0 ;
  assign y15904 = n43944 ;
  assign y15905 = ~n43947 ;
  assign y15906 = ~n43949 ;
  assign y15907 = ~1'b0 ;
  assign y15908 = n43951 ;
  assign y15909 = ~1'b0 ;
  assign y15910 = ~1'b0 ;
  assign y15911 = ~1'b0 ;
  assign y15912 = ~n43953 ;
  assign y15913 = ~1'b0 ;
  assign y15914 = ~n43954 ;
  assign y15915 = ~1'b0 ;
  assign y15916 = ~1'b0 ;
  assign y15917 = n43958 ;
  assign y15918 = ~n43961 ;
  assign y15919 = 1'b0 ;
  assign y15920 = ~1'b0 ;
  assign y15921 = n43962 ;
  assign y15922 = ~n43971 ;
  assign y15923 = n43973 ;
  assign y15924 = n43975 ;
  assign y15925 = n43980 ;
  assign y15926 = ~n43982 ;
  assign y15927 = ~n43985 ;
  assign y15928 = n43986 ;
  assign y15929 = n43988 ;
  assign y15930 = ~n43989 ;
  assign y15931 = n43993 ;
  assign y15932 = ~n43995 ;
  assign y15933 = n43998 ;
  assign y15934 = n44000 ;
  assign y15935 = ~n44001 ;
  assign y15936 = n20598 ;
  assign y15937 = ~n44003 ;
  assign y15938 = n44006 ;
  assign y15939 = n44011 ;
  assign y15940 = n44013 ;
  assign y15941 = n44015 ;
  assign y15942 = n44016 ;
  assign y15943 = ~n44017 ;
  assign y15944 = ~1'b0 ;
  assign y15945 = ~1'b0 ;
  assign y15946 = ~n44021 ;
  assign y15947 = ~n44024 ;
  assign y15948 = n44029 ;
  assign y15949 = n44032 ;
  assign y15950 = ~n44036 ;
  assign y15951 = ~n44039 ;
  assign y15952 = n44040 ;
  assign y15953 = n44047 ;
  assign y15954 = ~n44054 ;
  assign y15955 = ~1'b0 ;
  assign y15956 = n44056 ;
  assign y15957 = ~n44061 ;
  assign y15958 = ~n44065 ;
  assign y15959 = ~n44067 ;
  assign y15960 = n44070 ;
  assign y15961 = n44075 ;
  assign y15962 = ~n44079 ;
  assign y15963 = ~n44082 ;
  assign y15964 = n44083 ;
  assign y15965 = ~1'b0 ;
  assign y15966 = ~1'b0 ;
  assign y15967 = n44086 ;
  assign y15968 = n44087 ;
  assign y15969 = n44091 ;
  assign y15970 = n44094 ;
  assign y15971 = ~1'b0 ;
  assign y15972 = ~1'b0 ;
  assign y15973 = ~1'b0 ;
  assign y15974 = ~1'b0 ;
  assign y15975 = n44096 ;
  assign y15976 = n44101 ;
  assign y15977 = ~n44103 ;
  assign y15978 = n44108 ;
  assign y15979 = ~n44111 ;
  assign y15980 = n44112 ;
  assign y15981 = ~n44113 ;
  assign y15982 = ~n44124 ;
  assign y15983 = ~n44126 ;
  assign y15984 = n44127 ;
  assign y15985 = ~n44129 ;
  assign y15986 = ~n44131 ;
  assign y15987 = n44132 ;
  assign y15988 = n44135 ;
  assign y15989 = ~n44140 ;
  assign y15990 = ~1'b0 ;
  assign y15991 = ~n44142 ;
  assign y15992 = ~1'b0 ;
  assign y15993 = ~1'b0 ;
  assign y15994 = n44144 ;
  assign y15995 = ~n44146 ;
  assign y15996 = n44149 ;
  assign y15997 = ~n44150 ;
  assign y15998 = ~n44154 ;
  assign y15999 = ~n1705 ;
  assign y16000 = n44157 ;
  assign y16001 = ~n44158 ;
  assign y16002 = ~n44160 ;
  assign y16003 = ~1'b0 ;
  assign y16004 = ~1'b0 ;
  assign y16005 = n44163 ;
  assign y16006 = n44164 ;
  assign y16007 = ~n44170 ;
  assign y16008 = ~n44171 ;
  assign y16009 = ~1'b0 ;
  assign y16010 = ~n44174 ;
  assign y16011 = ~n44176 ;
  assign y16012 = ~1'b0 ;
  assign y16013 = n44177 ;
  assign y16014 = n44178 ;
  assign y16015 = n44182 ;
  assign y16016 = ~1'b0 ;
  assign y16017 = n44190 ;
  assign y16018 = ~1'b0 ;
  assign y16019 = n44192 ;
  assign y16020 = n44193 ;
  assign y16021 = n44195 ;
  assign y16022 = n8045 ;
  assign y16023 = n44197 ;
  assign y16024 = n44201 ;
  assign y16025 = ~1'b0 ;
  assign y16026 = ~n44202 ;
  assign y16027 = ~1'b0 ;
  assign y16028 = n44203 ;
  assign y16029 = ~n44205 ;
  assign y16030 = n44206 ;
  assign y16031 = ~n44208 ;
  assign y16032 = ~n44211 ;
  assign y16033 = ~1'b0 ;
  assign y16034 = ~n44215 ;
  assign y16035 = ~n44218 ;
  assign y16036 = ~n44220 ;
  assign y16037 = ~n44223 ;
  assign y16038 = n44224 ;
  assign y16039 = ~n44226 ;
  assign y16040 = ~1'b0 ;
  assign y16041 = n44227 ;
  assign y16042 = ~n44233 ;
  assign y16043 = n44234 ;
  assign y16044 = ~n44237 ;
  assign y16045 = n44238 ;
  assign y16046 = n44239 ;
  assign y16047 = ~1'b0 ;
  assign y16048 = ~n44243 ;
  assign y16049 = ~1'b0 ;
  assign y16050 = n44246 ;
  assign y16051 = n44249 ;
  assign y16052 = ~n44252 ;
  assign y16053 = n44253 ;
  assign y16054 = ~n44256 ;
  assign y16055 = n44257 ;
  assign y16056 = n44258 ;
  assign y16057 = n44260 ;
  assign y16058 = n44261 ;
  assign y16059 = ~n44265 ;
  assign y16060 = ~n44267 ;
  assign y16061 = ~n44269 ;
  assign y16062 = n44277 ;
  assign y16063 = n44279 ;
  assign y16064 = ~n44280 ;
  assign y16065 = ~n44285 ;
  assign y16066 = ~1'b0 ;
  assign y16067 = ~n44287 ;
  assign y16068 = n44289 ;
  assign y16069 = n44295 ;
  assign y16070 = n44296 ;
  assign y16071 = n44298 ;
  assign y16072 = n44301 ;
  assign y16073 = ~n44303 ;
  assign y16074 = ~1'b0 ;
  assign y16075 = ~1'b0 ;
  assign y16076 = ~1'b0 ;
  assign y16077 = n44306 ;
  assign y16078 = n44310 ;
  assign y16079 = n44313 ;
  assign y16080 = ~n44314 ;
  assign y16081 = ~1'b0 ;
  assign y16082 = ~1'b0 ;
  assign y16083 = ~1'b0 ;
  assign y16084 = ~n44318 ;
  assign y16085 = ~1'b0 ;
  assign y16086 = n44319 ;
  assign y16087 = n44320 ;
  assign y16088 = ~n44328 ;
  assign y16089 = ~n44329 ;
  assign y16090 = n44330 ;
  assign y16091 = n44332 ;
  assign y16092 = n40029 ;
  assign y16093 = ~1'b0 ;
  assign y16094 = n44336 ;
  assign y16095 = n44337 ;
  assign y16096 = ~n44338 ;
  assign y16097 = ~1'b0 ;
  assign y16098 = ~1'b0 ;
  assign y16099 = ~1'b0 ;
  assign y16100 = n44341 ;
  assign y16101 = ~n44344 ;
  assign y16102 = ~1'b0 ;
  assign y16103 = ~n44345 ;
  assign y16104 = n44348 ;
  assign y16105 = ~n44352 ;
  assign y16106 = n44363 ;
  assign y16107 = n44365 ;
  assign y16108 = ~n44369 ;
  assign y16109 = n44371 ;
  assign y16110 = ~n44373 ;
  assign y16111 = ~n44376 ;
  assign y16112 = ~n44377 ;
  assign y16113 = n44379 ;
  assign y16114 = ~n44380 ;
  assign y16115 = ~n44383 ;
  assign y16116 = n44387 ;
  assign y16117 = ~1'b0 ;
  assign y16118 = ~n44390 ;
  assign y16119 = n44391 ;
  assign y16120 = n44392 ;
  assign y16121 = ~n44393 ;
  assign y16122 = n44394 ;
  assign y16123 = ~1'b0 ;
  assign y16124 = n44397 ;
  assign y16125 = n44398 ;
  assign y16126 = n44399 ;
  assign y16127 = ~1'b0 ;
  assign y16128 = n44401 ;
  assign y16129 = n44403 ;
  assign y16130 = n44404 ;
  assign y16131 = ~n44409 ;
  assign y16132 = n44410 ;
  assign y16133 = ~1'b0 ;
  assign y16134 = ~n44413 ;
  assign y16135 = ~n44417 ;
  assign y16136 = ~1'b0 ;
  assign y16137 = ~n44419 ;
  assign y16138 = n44425 ;
  assign y16139 = n44430 ;
  assign y16140 = n44431 ;
  assign y16141 = ~n44432 ;
  assign y16142 = ~1'b0 ;
  assign y16143 = ~1'b0 ;
  assign y16144 = n44437 ;
  assign y16145 = n44440 ;
  assign y16146 = ~n44446 ;
  assign y16147 = n44451 ;
  assign y16148 = n44457 ;
  assign y16149 = ~n44458 ;
  assign y16150 = ~n44462 ;
  assign y16151 = ~1'b0 ;
  assign y16152 = n44464 ;
  assign y16153 = ~1'b0 ;
  assign y16154 = n44465 ;
  assign y16155 = n44471 ;
  assign y16156 = ~n44473 ;
  assign y16157 = ~n44475 ;
  assign y16158 = n44476 ;
  assign y16159 = n44484 ;
  assign y16160 = ~1'b0 ;
  assign y16161 = n44488 ;
  assign y16162 = ~1'b0 ;
  assign y16163 = ~n9941 ;
  assign y16164 = ~n44490 ;
  assign y16165 = ~n44493 ;
  assign y16166 = ~n44495 ;
  assign y16167 = n44496 ;
  assign y16168 = n44497 ;
  assign y16169 = ~1'b0 ;
  assign y16170 = ~n15187 ;
  assign y16171 = n44500 ;
  assign y16172 = ~n44502 ;
  assign y16173 = ~1'b0 ;
  assign y16174 = ~1'b0 ;
  assign y16175 = ~n44505 ;
  assign y16176 = n44508 ;
  assign y16177 = n44514 ;
  assign y16178 = ~n44516 ;
  assign y16179 = n44519 ;
  assign y16180 = n44520 ;
  assign y16181 = ~n44524 ;
  assign y16182 = ~1'b0 ;
  assign y16183 = ~1'b0 ;
  assign y16184 = ~1'b0 ;
  assign y16185 = n44525 ;
  assign y16186 = ~n44526 ;
  assign y16187 = n44528 ;
  assign y16188 = n44530 ;
  assign y16189 = ~n44533 ;
  assign y16190 = n44535 ;
  assign y16191 = ~n44536 ;
  assign y16192 = ~n44538 ;
  assign y16193 = ~n44541 ;
  assign y16194 = ~n44543 ;
  assign y16195 = ~n44546 ;
  assign y16196 = ~n44552 ;
  assign y16197 = ~1'b0 ;
  assign y16198 = ~n44553 ;
  assign y16199 = ~n44559 ;
  assign y16200 = n44560 ;
  assign y16201 = ~n44561 ;
  assign y16202 = ~n8374 ;
  assign y16203 = ~n44562 ;
  assign y16204 = ~1'b0 ;
  assign y16205 = ~1'b0 ;
  assign y16206 = ~1'b0 ;
  assign y16207 = n44564 ;
  assign y16208 = ~n44571 ;
  assign y16209 = n44574 ;
  assign y16210 = n44576 ;
  assign y16211 = n44583 ;
  assign y16212 = n44584 ;
  assign y16213 = n44586 ;
  assign y16214 = ~1'b0 ;
  assign y16215 = ~n44589 ;
  assign y16216 = n44593 ;
  assign y16217 = ~n44595 ;
  assign y16218 = ~n44596 ;
  assign y16219 = n44607 ;
  assign y16220 = ~n44608 ;
  assign y16221 = ~n44610 ;
  assign y16222 = n44612 ;
  assign y16223 = n44615 ;
  assign y16224 = n44616 ;
  assign y16225 = ~n44617 ;
  assign y16226 = ~n44619 ;
  assign y16227 = ~n44623 ;
  assign y16228 = ~n44625 ;
  assign y16229 = ~n44628 ;
  assign y16230 = ~n44632 ;
  assign y16231 = n44633 ;
  assign y16232 = ~1'b0 ;
  assign y16233 = n44635 ;
  assign y16234 = ~n44637 ;
  assign y16235 = ~n44642 ;
  assign y16236 = ~n44643 ;
  assign y16237 = ~n44644 ;
  assign y16238 = ~n44650 ;
  assign y16239 = n44656 ;
  assign y16240 = ~n44658 ;
  assign y16241 = ~1'b0 ;
  assign y16242 = n44662 ;
  assign y16243 = ~1'b0 ;
  assign y16244 = ~1'b0 ;
  assign y16245 = n44665 ;
  assign y16246 = ~n44666 ;
  assign y16247 = n44677 ;
  assign y16248 = n44683 ;
  assign y16249 = n44684 ;
  assign y16250 = ~1'b0 ;
  assign y16251 = ~n44686 ;
  assign y16252 = n44689 ;
  assign y16253 = n44696 ;
  assign y16254 = ~n44697 ;
  assign y16255 = ~n44699 ;
  assign y16256 = n44703 ;
  assign y16257 = ~n44708 ;
  assign y16258 = ~n44709 ;
  assign y16259 = ~n44715 ;
  assign y16260 = n44720 ;
  assign y16261 = ~1'b0 ;
  assign y16262 = ~1'b0 ;
  assign y16263 = n44723 ;
  assign y16264 = n44726 ;
  assign y16265 = ~n44727 ;
  assign y16266 = ~1'b0 ;
  assign y16267 = ~n44737 ;
  assign y16268 = n44739 ;
  assign y16269 = ~n44741 ;
  assign y16270 = n44743 ;
  assign y16271 = n44745 ;
  assign y16272 = n44749 ;
  assign y16273 = ~1'b0 ;
  assign y16274 = ~n44753 ;
  assign y16275 = n14131 ;
  assign y16276 = ~n44755 ;
  assign y16277 = ~1'b0 ;
  assign y16278 = ~n44757 ;
  assign y16279 = n44760 ;
  assign y16280 = ~n44761 ;
  assign y16281 = ~n44764 ;
  assign y16282 = ~n44775 ;
  assign y16283 = ~n44778 ;
  assign y16284 = ~1'b0 ;
  assign y16285 = n44781 ;
  assign y16286 = n44782 ;
  assign y16287 = n44786 ;
  assign y16288 = ~n44787 ;
  assign y16289 = n44794 ;
  assign y16290 = ~n44798 ;
  assign y16291 = ~1'b0 ;
  assign y16292 = ~n44799 ;
  assign y16293 = n44801 ;
  assign y16294 = ~1'b0 ;
  assign y16295 = n44802 ;
  assign y16296 = n44806 ;
  assign y16297 = ~n44811 ;
  assign y16298 = n44812 ;
  assign y16299 = n44813 ;
  assign y16300 = ~n44815 ;
  assign y16301 = n44816 ;
  assign y16302 = ~1'b0 ;
  assign y16303 = ~n44818 ;
  assign y16304 = ~n44820 ;
  assign y16305 = ~n44827 ;
  assign y16306 = n44830 ;
  assign y16307 = ~n44831 ;
  assign y16308 = n44835 ;
  assign y16309 = ~n5791 ;
  assign y16310 = ~1'b0 ;
  assign y16311 = ~n44837 ;
  assign y16312 = ~1'b0 ;
  assign y16313 = n44839 ;
  assign y16314 = ~n44843 ;
  assign y16315 = ~n44846 ;
  assign y16316 = ~n44848 ;
  assign y16317 = ~1'b0 ;
  assign y16318 = ~n44853 ;
  assign y16319 = ~n44857 ;
  assign y16320 = ~1'b0 ;
  assign y16321 = ~n44859 ;
  assign y16322 = ~n44860 ;
  assign y16323 = ~n44862 ;
  assign y16324 = n44866 ;
  assign y16325 = ~1'b0 ;
  assign y16326 = ~1'b0 ;
  assign y16327 = n44867 ;
  assign y16328 = ~1'b0 ;
  assign y16329 = n44870 ;
  assign y16330 = n44871 ;
  assign y16331 = n44874 ;
  assign y16332 = ~n5777 ;
  assign y16333 = ~n44878 ;
  assign y16334 = ~n44880 ;
  assign y16335 = n44882 ;
  assign y16336 = ~1'b0 ;
  assign y16337 = ~n44884 ;
  assign y16338 = ~1'b0 ;
  assign y16339 = n44885 ;
  assign y16340 = ~n9069 ;
  assign y16341 = n44886 ;
  assign y16342 = ~n44887 ;
  assign y16343 = n44890 ;
  assign y16344 = ~n44892 ;
  assign y16345 = ~1'b0 ;
  assign y16346 = ~n44894 ;
  assign y16347 = n44899 ;
  assign y16348 = n44903 ;
  assign y16349 = ~n44904 ;
  assign y16350 = ~n44912 ;
  assign y16351 = n44914 ;
  assign y16352 = n44915 ;
  assign y16353 = ~1'b0 ;
  assign y16354 = ~1'b0 ;
  assign y16355 = ~1'b0 ;
  assign y16356 = ~n44916 ;
  assign y16357 = ~n44917 ;
  assign y16358 = n44919 ;
  assign y16359 = ~1'b0 ;
  assign y16360 = ~1'b0 ;
  assign y16361 = n44921 ;
  assign y16362 = ~1'b0 ;
  assign y16363 = ~n44922 ;
  assign y16364 = ~n44925 ;
  assign y16365 = n44927 ;
  assign y16366 = n44928 ;
  assign y16367 = ~n44929 ;
  assign y16368 = ~n44932 ;
  assign y16369 = ~1'b0 ;
  assign y16370 = ~n44933 ;
  assign y16371 = ~1'b0 ;
  assign y16372 = ~n44935 ;
  assign y16373 = ~1'b0 ;
  assign y16374 = ~1'b0 ;
  assign y16375 = ~n44936 ;
  assign y16376 = ~n44937 ;
  assign y16377 = ~n44939 ;
  assign y16378 = ~n44942 ;
  assign y16379 = ~n44950 ;
  assign y16380 = ~n44954 ;
  assign y16381 = ~n44955 ;
  assign y16382 = n44960 ;
  assign y16383 = ~n44961 ;
  assign y16384 = n44968 ;
  assign y16385 = ~1'b0 ;
  assign y16386 = ~1'b0 ;
  assign y16387 = ~1'b0 ;
  assign y16388 = n27623 ;
  assign y16389 = n44970 ;
  assign y16390 = ~n44972 ;
  assign y16391 = ~n44975 ;
  assign y16392 = n44979 ;
  assign y16393 = ~n44981 ;
  assign y16394 = ~n44983 ;
  assign y16395 = n44984 ;
  assign y16396 = ~1'b0 ;
  assign y16397 = ~n44987 ;
  assign y16398 = ~n44989 ;
  assign y16399 = n44990 ;
  assign y16400 = n44992 ;
  assign y16401 = ~n44993 ;
  assign y16402 = n44995 ;
  assign y16403 = ~1'b0 ;
  assign y16404 = n44997 ;
  assign y16405 = n44998 ;
  assign y16406 = ~1'b0 ;
  assign y16407 = ~n44999 ;
  assign y16408 = n45003 ;
  assign y16409 = ~n45004 ;
  assign y16410 = ~n45006 ;
  assign y16411 = ~n45009 ;
  assign y16412 = n45012 ;
  assign y16413 = ~1'b0 ;
  assign y16414 = n45013 ;
  assign y16415 = ~1'b0 ;
  assign y16416 = ~n45016 ;
  assign y16417 = ~n45017 ;
  assign y16418 = n45018 ;
  assign y16419 = n45020 ;
  assign y16420 = n45022 ;
  assign y16421 = ~1'b0 ;
  assign y16422 = ~n45023 ;
  assign y16423 = n45025 ;
  assign y16424 = n45029 ;
  assign y16425 = ~n45030 ;
  assign y16426 = ~n45039 ;
  assign y16427 = n45043 ;
  assign y16428 = ~n45045 ;
  assign y16429 = ~n45048 ;
  assign y16430 = ~n45053 ;
  assign y16431 = ~1'b0 ;
  assign y16432 = ~1'b0 ;
  assign y16433 = ~n45058 ;
  assign y16434 = n45062 ;
  assign y16435 = n45065 ;
  assign y16436 = ~n45070 ;
  assign y16437 = ~n45071 ;
  assign y16438 = ~n45073 ;
  assign y16439 = ~1'b0 ;
  assign y16440 = ~n45075 ;
  assign y16441 = ~n45078 ;
  assign y16442 = ~n45080 ;
  assign y16443 = ~n45081 ;
  assign y16444 = ~n45082 ;
  assign y16445 = ~1'b0 ;
  assign y16446 = ~1'b0 ;
  assign y16447 = ~n45084 ;
  assign y16448 = n45085 ;
  assign y16449 = ~n45087 ;
  assign y16450 = ~n45088 ;
  assign y16451 = n45089 ;
  assign y16452 = n45091 ;
  assign y16453 = ~n45092 ;
  assign y16454 = ~n45096 ;
  assign y16455 = ~n45102 ;
  assign y16456 = ~n45103 ;
  assign y16457 = ~n45106 ;
  assign y16458 = n45112 ;
  assign y16459 = ~n11349 ;
  assign y16460 = ~1'b0 ;
  assign y16461 = ~n45114 ;
  assign y16462 = ~1'b0 ;
  assign y16463 = ~1'b0 ;
  assign y16464 = ~n45117 ;
  assign y16465 = n1202 ;
  assign y16466 = ~n45118 ;
  assign y16467 = ~n45121 ;
  assign y16468 = ~n45125 ;
  assign y16469 = ~1'b0 ;
  assign y16470 = n45127 ;
  assign y16471 = n45130 ;
  assign y16472 = ~n45133 ;
  assign y16473 = ~1'b0 ;
  assign y16474 = n45140 ;
  assign y16475 = ~n45141 ;
  assign y16476 = n45142 ;
  assign y16477 = n45143 ;
  assign y16478 = n45144 ;
  assign y16479 = ~n45147 ;
  assign y16480 = ~n45153 ;
  assign y16481 = ~n45156 ;
  assign y16482 = ~1'b0 ;
  assign y16483 = n45157 ;
  assign y16484 = n45158 ;
  assign y16485 = n45159 ;
  assign y16486 = ~n45161 ;
  assign y16487 = n45166 ;
  assign y16488 = ~n45167 ;
  assign y16489 = n45168 ;
  assign y16490 = ~n45170 ;
  assign y16491 = n45172 ;
  assign y16492 = n45174 ;
  assign y16493 = n45175 ;
  assign y16494 = n45180 ;
  assign y16495 = ~n45184 ;
  assign y16496 = n45185 ;
  assign y16497 = n45188 ;
  assign y16498 = ~n45190 ;
  assign y16499 = n45191 ;
  assign y16500 = ~n45193 ;
  assign y16501 = n45194 ;
  assign y16502 = n4757 ;
  assign y16503 = ~n45195 ;
  assign y16504 = ~n45198 ;
  assign y16505 = ~1'b0 ;
  assign y16506 = ~n45199 ;
  assign y16507 = ~1'b0 ;
  assign y16508 = ~n45200 ;
  assign y16509 = ~n45203 ;
  assign y16510 = ~n45207 ;
  assign y16511 = n45215 ;
  assign y16512 = ~n45218 ;
  assign y16513 = ~n45223 ;
  assign y16514 = n45226 ;
  assign y16515 = n45227 ;
  assign y16516 = ~n45233 ;
  assign y16517 = ~1'b0 ;
  assign y16518 = ~1'b0 ;
  assign y16519 = ~n45235 ;
  assign y16520 = n45238 ;
  assign y16521 = n45240 ;
  assign y16522 = ~n45243 ;
  assign y16523 = ~n45244 ;
  assign y16524 = ~n45246 ;
  assign y16525 = ~1'b0 ;
  assign y16526 = n45253 ;
  assign y16527 = n45254 ;
  assign y16528 = n45255 ;
  assign y16529 = ~n45257 ;
  assign y16530 = ~n45262 ;
  assign y16531 = n45265 ;
  assign y16532 = ~1'b0 ;
  assign y16533 = ~n28978 ;
  assign y16534 = n45266 ;
  assign y16535 = n45267 ;
  assign y16536 = ~n45268 ;
  assign y16537 = ~n45271 ;
  assign y16538 = ~n45272 ;
  assign y16539 = n45273 ;
  assign y16540 = ~1'b0 ;
  assign y16541 = ~n45275 ;
  assign y16542 = ~n45276 ;
  assign y16543 = n45277 ;
  assign y16544 = ~n45281 ;
  assign y16545 = ~n45286 ;
  assign y16546 = n45292 ;
  assign y16547 = ~n45296 ;
  assign y16548 = n45298 ;
  assign y16549 = ~1'b0 ;
  assign y16550 = ~1'b0 ;
  assign y16551 = n45299 ;
  assign y16552 = ~n45300 ;
  assign y16553 = ~n45302 ;
  assign y16554 = n45306 ;
  assign y16555 = n45307 ;
  assign y16556 = ~n45308 ;
  assign y16557 = ~n45311 ;
  assign y16558 = ~1'b0 ;
  assign y16559 = ~n45313 ;
  assign y16560 = n45314 ;
  assign y16561 = ~n45316 ;
  assign y16562 = ~1'b0 ;
  assign y16563 = n45319 ;
  assign y16564 = n45320 ;
  assign y16565 = n45321 ;
  assign y16566 = n45323 ;
  assign y16567 = ~n45326 ;
  assign y16568 = n45327 ;
  assign y16569 = ~n45330 ;
  assign y16570 = ~n45331 ;
  assign y16571 = ~n45332 ;
  assign y16572 = n45333 ;
  assign y16573 = ~n45335 ;
  assign y16574 = ~n45336 ;
  assign y16575 = n45338 ;
  assign y16576 = ~n45341 ;
  assign y16577 = n45342 ;
  assign y16578 = n45344 ;
  assign y16579 = ~n45347 ;
  assign y16580 = ~1'b0 ;
  assign y16581 = ~n45351 ;
  assign y16582 = ~n45352 ;
  assign y16583 = ~n45358 ;
  assign y16584 = n45363 ;
  assign y16585 = n45364 ;
  assign y16586 = ~n45365 ;
  assign y16587 = n45369 ;
  assign y16588 = ~n45372 ;
  assign y16589 = n45375 ;
  assign y16590 = ~1'b0 ;
  assign y16591 = n45377 ;
  assign y16592 = ~n45378 ;
  assign y16593 = ~n45384 ;
  assign y16594 = n45385 ;
  assign y16595 = n45387 ;
  assign y16596 = n45392 ;
  assign y16597 = n45394 ;
  assign y16598 = ~1'b0 ;
  assign y16599 = ~n45395 ;
  assign y16600 = n45402 ;
  assign y16601 = n45404 ;
  assign y16602 = ~n45405 ;
  assign y16603 = ~1'b0 ;
  assign y16604 = n45407 ;
  assign y16605 = ~n45412 ;
  assign y16606 = n45415 ;
  assign y16607 = ~n45417 ;
  assign y16608 = n45418 ;
  assign y16609 = ~n45422 ;
  assign y16610 = n45424 ;
  assign y16611 = n45425 ;
  assign y16612 = ~n45427 ;
  assign y16613 = ~n45430 ;
  assign y16614 = n45432 ;
  assign y16615 = ~1'b0 ;
  assign y16616 = ~n45433 ;
  assign y16617 = n45436 ;
  assign y16618 = ~n45438 ;
  assign y16619 = n45439 ;
  assign y16620 = ~n45440 ;
  assign y16621 = ~n45442 ;
  assign y16622 = n45448 ;
  assign y16623 = ~1'b0 ;
  assign y16624 = ~1'b0 ;
  assign y16625 = ~1'b0 ;
  assign y16626 = n45456 ;
  assign y16627 = ~n45457 ;
  assign y16628 = n45460 ;
  assign y16629 = n45463 ;
  assign y16630 = ~n45464 ;
  assign y16631 = ~n45465 ;
  assign y16632 = n45466 ;
  assign y16633 = ~1'b0 ;
  assign y16634 = ~1'b0 ;
  assign y16635 = ~n45467 ;
  assign y16636 = n1836 ;
  assign y16637 = ~n45468 ;
  assign y16638 = ~1'b0 ;
  assign y16639 = ~1'b0 ;
  assign y16640 = ~1'b0 ;
  assign y16641 = ~n45470 ;
  assign y16642 = ~n45475 ;
  assign y16643 = n45476 ;
  assign y16644 = n45478 ;
  assign y16645 = n45479 ;
  assign y16646 = n45480 ;
  assign y16647 = ~n45482 ;
  assign y16648 = n45484 ;
  assign y16649 = n45489 ;
  assign y16650 = ~1'b0 ;
  assign y16651 = ~1'b0 ;
  assign y16652 = n9334 ;
  assign y16653 = n11342 ;
  assign y16654 = n45493 ;
  assign y16655 = ~n45496 ;
  assign y16656 = n45498 ;
  assign y16657 = n45500 ;
  assign y16658 = ~n45501 ;
  assign y16659 = ~1'b0 ;
  assign y16660 = ~n45504 ;
  assign y16661 = ~n45509 ;
  assign y16662 = ~n45511 ;
  assign y16663 = ~n45515 ;
  assign y16664 = ~n45516 ;
  assign y16665 = ~n45518 ;
  assign y16666 = ~n45519 ;
  assign y16667 = n25701 ;
  assign y16668 = n45521 ;
  assign y16669 = ~1'b0 ;
  assign y16670 = ~n45523 ;
  assign y16671 = ~n45524 ;
  assign y16672 = ~n45526 ;
  assign y16673 = ~n45527 ;
  assign y16674 = n45528 ;
  assign y16675 = ~n45530 ;
  assign y16676 = ~n45533 ;
  assign y16677 = n45536 ;
  assign y16678 = ~n45537 ;
  assign y16679 = ~n45539 ;
  assign y16680 = n1214 ;
  assign y16681 = ~n45540 ;
  assign y16682 = ~n45543 ;
  assign y16683 = n45544 ;
  assign y16684 = n45548 ;
  assign y16685 = ~n45551 ;
  assign y16686 = ~1'b0 ;
  assign y16687 = ~n45555 ;
  assign y16688 = n45558 ;
  assign y16689 = ~1'b0 ;
  assign y16690 = n45564 ;
  assign y16691 = ~n45565 ;
  assign y16692 = n45568 ;
  assign y16693 = n45569 ;
  assign y16694 = n45571 ;
  assign y16695 = n45572 ;
  assign y16696 = n8092 ;
  assign y16697 = n45575 ;
  assign y16698 = n45576 ;
  assign y16699 = n45580 ;
  assign y16700 = ~n45582 ;
  assign y16701 = n45584 ;
  assign y16702 = n45587 ;
  assign y16703 = ~n45589 ;
  assign y16704 = n45592 ;
  assign y16705 = n45594 ;
  assign y16706 = ~1'b0 ;
  assign y16707 = n45595 ;
  assign y16708 = n45596 ;
  assign y16709 = n45597 ;
  assign y16710 = ~n45599 ;
  assign y16711 = ~1'b0 ;
  assign y16712 = ~1'b0 ;
  assign y16713 = ~1'b0 ;
  assign y16714 = ~n45602 ;
  assign y16715 = n45603 ;
  assign y16716 = ~n45605 ;
  assign y16717 = ~n45606 ;
  assign y16718 = n45607 ;
  assign y16719 = ~1'b0 ;
  assign y16720 = ~n28337 ;
  assign y16721 = ~1'b0 ;
  assign y16722 = ~1'b0 ;
  assign y16723 = n45608 ;
  assign y16724 = ~n45610 ;
  assign y16725 = n45613 ;
  assign y16726 = ~n45614 ;
  assign y16727 = ~n45615 ;
  assign y16728 = n45623 ;
  assign y16729 = n45625 ;
  assign y16730 = n45626 ;
  assign y16731 = n45628 ;
  assign y16732 = ~1'b0 ;
  assign y16733 = ~n45629 ;
  assign y16734 = n45631 ;
  assign y16735 = n45635 ;
  assign y16736 = n45636 ;
  assign y16737 = ~n45637 ;
  assign y16738 = n45639 ;
  assign y16739 = ~n45641 ;
  assign y16740 = n45644 ;
  assign y16741 = ~n45645 ;
  assign y16742 = ~n45648 ;
  assign y16743 = ~n45652 ;
  assign y16744 = n45653 ;
  assign y16745 = ~n45655 ;
  assign y16746 = n45658 ;
  assign y16747 = n45660 ;
  assign y16748 = ~1'b0 ;
  assign y16749 = ~n45663 ;
  assign y16750 = n45665 ;
  assign y16751 = n45666 ;
  assign y16752 = ~n45672 ;
  assign y16753 = ~n45674 ;
  assign y16754 = ~n45676 ;
  assign y16755 = ~n45678 ;
  assign y16756 = ~n45681 ;
  assign y16757 = n45686 ;
  assign y16758 = ~n45688 ;
  assign y16759 = ~1'b0 ;
  assign y16760 = ~n45689 ;
  assign y16761 = n45694 ;
  assign y16762 = n45700 ;
  assign y16763 = n45701 ;
  assign y16764 = ~n45707 ;
  assign y16765 = ~n45710 ;
  assign y16766 = n45712 ;
  assign y16767 = ~n45715 ;
  assign y16768 = n45716 ;
  assign y16769 = n45718 ;
  assign y16770 = n45721 ;
  assign y16771 = ~n45722 ;
  assign y16772 = ~n45729 ;
  assign y16773 = ~n45730 ;
  assign y16774 = n45731 ;
  assign y16775 = n45733 ;
  assign y16776 = ~1'b0 ;
  assign y16777 = ~n45734 ;
  assign y16778 = n45736 ;
  assign y16779 = n45739 ;
  assign y16780 = ~n45746 ;
  assign y16781 = n23309 ;
  assign y16782 = ~n45748 ;
  assign y16783 = n45750 ;
  assign y16784 = ~1'b0 ;
  assign y16785 = n45751 ;
  assign y16786 = n45752 ;
  assign y16787 = ~n45753 ;
  assign y16788 = n45759 ;
  assign y16789 = ~n45762 ;
  assign y16790 = ~n45763 ;
  assign y16791 = ~n45767 ;
  assign y16792 = n45768 ;
  assign y16793 = ~n45769 ;
  assign y16794 = ~n45770 ;
  assign y16795 = ~n45771 ;
  assign y16796 = ~1'b0 ;
  assign y16797 = n45778 ;
  assign y16798 = n45780 ;
  assign y16799 = n45786 ;
  assign y16800 = ~n45790 ;
  assign y16801 = n45791 ;
  assign y16802 = ~n45797 ;
  assign y16803 = ~n45798 ;
  assign y16804 = ~n45803 ;
  assign y16805 = ~n45805 ;
  assign y16806 = ~1'b0 ;
  assign y16807 = n45807 ;
  assign y16808 = n45808 ;
  assign y16809 = ~n45812 ;
  assign y16810 = ~n45813 ;
  assign y16811 = n45815 ;
  assign y16812 = n45816 ;
  assign y16813 = ~n45819 ;
  assign y16814 = ~1'b0 ;
  assign y16815 = ~n45820 ;
  assign y16816 = ~n45822 ;
  assign y16817 = ~n8719 ;
  assign y16818 = n45823 ;
  assign y16819 = n45830 ;
  assign y16820 = ~n45833 ;
  assign y16821 = ~n45835 ;
  assign y16822 = ~n45838 ;
  assign y16823 = ~n45841 ;
  assign y16824 = n45842 ;
  assign y16825 = ~n45846 ;
  assign y16826 = n45857 ;
  assign y16827 = ~1'b0 ;
  assign y16828 = ~n45859 ;
  assign y16829 = ~n45862 ;
  assign y16830 = ~n45863 ;
  assign y16831 = n45864 ;
  assign y16832 = ~n45868 ;
  assign y16833 = ~1'b0 ;
  assign y16834 = n45870 ;
  assign y16835 = n45874 ;
  assign y16836 = ~n45876 ;
  assign y16837 = n45881 ;
  assign y16838 = ~1'b0 ;
  assign y16839 = ~n45884 ;
  assign y16840 = n45885 ;
  assign y16841 = ~n45890 ;
  assign y16842 = ~n45892 ;
  assign y16843 = n45899 ;
  assign y16844 = n45902 ;
  assign y16845 = ~1'b0 ;
  assign y16846 = n45904 ;
  assign y16847 = ~n45905 ;
  assign y16848 = n45906 ;
  assign y16849 = n45910 ;
  assign y16850 = ~n45912 ;
  assign y16851 = n45914 ;
  assign y16852 = ~1'b0 ;
  assign y16853 = n45918 ;
  assign y16854 = ~n45920 ;
  assign y16855 = n45925 ;
  assign y16856 = n45929 ;
  assign y16857 = ~n45930 ;
  assign y16858 = ~n45933 ;
  assign y16859 = ~n45936 ;
  assign y16860 = ~n45937 ;
  assign y16861 = ~n45941 ;
  assign y16862 = n45944 ;
  assign y16863 = ~n45946 ;
  assign y16864 = ~1'b0 ;
  assign y16865 = ~1'b0 ;
  assign y16866 = ~1'b0 ;
  assign y16867 = ~n45952 ;
  assign y16868 = ~n45953 ;
  assign y16869 = ~n45954 ;
  assign y16870 = ~n45955 ;
  assign y16871 = n45958 ;
  assign y16872 = n45961 ;
  assign y16873 = ~1'b0 ;
  assign y16874 = n45969 ;
  assign y16875 = n45970 ;
  assign y16876 = ~1'b0 ;
  assign y16877 = ~n45971 ;
  assign y16878 = n2786 ;
  assign y16879 = ~n45973 ;
  assign y16880 = ~n45976 ;
  assign y16881 = n45977 ;
  assign y16882 = ~1'b0 ;
  assign y16883 = ~1'b0 ;
  assign y16884 = n45979 ;
  assign y16885 = n45981 ;
  assign y16886 = ~n45985 ;
  assign y16887 = n45992 ;
  assign y16888 = n45993 ;
  assign y16889 = n45997 ;
  assign y16890 = ~n45998 ;
  assign y16891 = n46000 ;
  assign y16892 = n46001 ;
  assign y16893 = n46007 ;
  assign y16894 = ~1'b0 ;
  assign y16895 = n46011 ;
  assign y16896 = ~n46014 ;
  assign y16897 = n46015 ;
  assign y16898 = n19665 ;
  assign y16899 = ~n46018 ;
  assign y16900 = ~1'b0 ;
  assign y16901 = ~1'b0 ;
  assign y16902 = ~1'b0 ;
  assign y16903 = ~1'b0 ;
  assign y16904 = ~1'b0 ;
  assign y16905 = ~1'b0 ;
  assign y16906 = ~n46023 ;
  assign y16907 = n46025 ;
  assign y16908 = ~n46028 ;
  assign y16909 = n46034 ;
  assign y16910 = n46037 ;
  assign y16911 = n46038 ;
  assign y16912 = ~n46039 ;
  assign y16913 = ~n46041 ;
  assign y16914 = n46042 ;
  assign y16915 = ~1'b0 ;
  assign y16916 = ~n46045 ;
  assign y16917 = ~n46047 ;
  assign y16918 = n46048 ;
  assign y16919 = ~n46056 ;
  assign y16920 = ~n46059 ;
  assign y16921 = n46060 ;
  assign y16922 = n46062 ;
  assign y16923 = n46064 ;
  assign y16924 = ~n46067 ;
  assign y16925 = n3184 ;
  assign y16926 = ~n46068 ;
  assign y16927 = ~n46069 ;
  assign y16928 = n46071 ;
  assign y16929 = ~n46073 ;
  assign y16930 = ~n46076 ;
  assign y16931 = ~1'b0 ;
  assign y16932 = ~n46082 ;
  assign y16933 = n46090 ;
  assign y16934 = 1'b0 ;
  assign y16935 = ~n46100 ;
  assign y16936 = n46103 ;
  assign y16937 = ~1'b0 ;
  assign y16938 = ~n46106 ;
  assign y16939 = ~n46108 ;
  assign y16940 = n46110 ;
  assign y16941 = n12983 ;
  assign y16942 = ~n46113 ;
  assign y16943 = ~n46114 ;
  assign y16944 = ~n46115 ;
  assign y16945 = n46116 ;
  assign y16946 = n46119 ;
  assign y16947 = ~n46122 ;
  assign y16948 = ~1'b0 ;
  assign y16949 = ~n46125 ;
  assign y16950 = ~n46128 ;
  assign y16951 = ~n46130 ;
  assign y16952 = ~n46131 ;
  assign y16953 = ~n46142 ;
  assign y16954 = n46143 ;
  assign y16955 = ~n46147 ;
  assign y16956 = ~1'b0 ;
  assign y16957 = n46149 ;
  assign y16958 = ~1'b0 ;
  assign y16959 = ~1'b0 ;
  assign y16960 = ~n46152 ;
  assign y16961 = n46153 ;
  assign y16962 = n46154 ;
  assign y16963 = n46155 ;
  assign y16964 = ~1'b0 ;
  assign y16965 = ~1'b0 ;
  assign y16966 = n46159 ;
  assign y16967 = n46161 ;
  assign y16968 = ~n46162 ;
  assign y16969 = n46172 ;
  assign y16970 = n6420 ;
  assign y16971 = n46176 ;
  assign y16972 = n46181 ;
  assign y16973 = ~1'b0 ;
  assign y16974 = ~n46186 ;
  assign y16975 = ~n46187 ;
  assign y16976 = n46190 ;
  assign y16977 = ~1'b0 ;
  assign y16978 = ~n46191 ;
  assign y16979 = n46194 ;
  assign y16980 = n46197 ;
  assign y16981 = ~n46201 ;
  assign y16982 = ~n46204 ;
  assign y16983 = n46205 ;
  assign y16984 = n46208 ;
  assign y16985 = ~1'b0 ;
  assign y16986 = n46209 ;
  assign y16987 = n46213 ;
  assign y16988 = n46215 ;
  assign y16989 = n46216 ;
  assign y16990 = ~n46218 ;
  assign y16991 = n46223 ;
  assign y16992 = ~1'b0 ;
  assign y16993 = ~1'b0 ;
  assign y16994 = n46225 ;
  assign y16995 = n46226 ;
  assign y16996 = n46231 ;
  assign y16997 = ~n46232 ;
  assign y16998 = ~n46235 ;
  assign y16999 = n46238 ;
  assign y17000 = n46240 ;
  assign y17001 = ~n15056 ;
  assign y17002 = n46242 ;
  assign y17003 = ~n46246 ;
  assign y17004 = ~1'b0 ;
  assign y17005 = ~1'b0 ;
  assign y17006 = ~1'b0 ;
  assign y17007 = n46248 ;
  assign y17008 = n46255 ;
  assign y17009 = n46259 ;
  assign y17010 = ~n46260 ;
  assign y17011 = n46266 ;
  assign y17012 = ~1'b0 ;
  assign y17013 = n46269 ;
  assign y17014 = ~1'b0 ;
  assign y17015 = ~n46274 ;
  assign y17016 = n46277 ;
  assign y17017 = ~n46279 ;
  assign y17018 = ~n46281 ;
  assign y17019 = n46284 ;
  assign y17020 = ~n46288 ;
  assign y17021 = ~n46291 ;
  assign y17022 = ~n46293 ;
  assign y17023 = ~n46295 ;
  assign y17024 = ~n46298 ;
  assign y17025 = ~n46299 ;
  assign y17026 = n46306 ;
  assign y17027 = ~n46307 ;
  assign y17028 = n46309 ;
  assign y17029 = ~1'b0 ;
  assign y17030 = ~1'b0 ;
  assign y17031 = ~n46312 ;
  assign y17032 = n46319 ;
  assign y17033 = ~n46323 ;
  assign y17034 = ~1'b0 ;
  assign y17035 = ~n46324 ;
  assign y17036 = ~n46326 ;
  assign y17037 = n46327 ;
  assign y17038 = n46328 ;
  assign y17039 = n46332 ;
  assign y17040 = ~1'b0 ;
  assign y17041 = ~n46333 ;
  assign y17042 = ~n46334 ;
  assign y17043 = 1'b0 ;
  assign y17044 = n46340 ;
  assign y17045 = ~n46345 ;
  assign y17046 = n46349 ;
  assign y17047 = ~n46350 ;
  assign y17048 = n46353 ;
  assign y17049 = ~n46354 ;
  assign y17050 = ~n46356 ;
  assign y17051 = ~n46362 ;
  assign y17052 = ~n46363 ;
  assign y17053 = n46365 ;
  assign y17054 = ~n46366 ;
  assign y17055 = n46368 ;
  assign y17056 = ~n46372 ;
  assign y17057 = n46373 ;
  assign y17058 = n46374 ;
  assign y17059 = n46383 ;
  assign y17060 = ~1'b0 ;
  assign y17061 = ~n46388 ;
  assign y17062 = n46389 ;
  assign y17063 = ~n46390 ;
  assign y17064 = n46393 ;
  assign y17065 = n46394 ;
  assign y17066 = ~n46395 ;
  assign y17067 = n46396 ;
  assign y17068 = ~n46398 ;
  assign y17069 = ~n46399 ;
  assign y17070 = ~n46401 ;
  assign y17071 = ~1'b0 ;
  assign y17072 = n46402 ;
  assign y17073 = n46404 ;
  assign y17074 = ~1'b0 ;
  assign y17075 = ~n46405 ;
  assign y17076 = n46411 ;
  assign y17077 = n46412 ;
  assign y17078 = ~n46414 ;
  assign y17079 = ~n46415 ;
  assign y17080 = ~n46416 ;
  assign y17081 = n46418 ;
  assign y17082 = ~1'b0 ;
  assign y17083 = ~n46421 ;
  assign y17084 = ~n46422 ;
  assign y17085 = n46426 ;
  assign y17086 = n46427 ;
  assign y17087 = ~n46429 ;
  assign y17088 = ~n46431 ;
  assign y17089 = n46434 ;
  assign y17090 = ~n46437 ;
  assign y17091 = ~1'b0 ;
  assign y17092 = ~1'b0 ;
  assign y17093 = ~1'b0 ;
  assign y17094 = ~n46439 ;
  assign y17095 = n46444 ;
  assign y17096 = ~n46446 ;
  assign y17097 = n46447 ;
  assign y17098 = ~n46450 ;
  assign y17099 = ~n46454 ;
  assign y17100 = n46455 ;
  assign y17101 = ~1'b0 ;
  assign y17102 = ~n46459 ;
  assign y17103 = ~1'b0 ;
  assign y17104 = ~n46461 ;
  assign y17105 = ~1'b0 ;
  assign y17106 = ~n46463 ;
  assign y17107 = n46464 ;
  assign y17108 = ~n11439 ;
  assign y17109 = ~1'b0 ;
  assign y17110 = ~1'b0 ;
  assign y17111 = ~1'b0 ;
  assign y17112 = ~1'b0 ;
  assign y17113 = n46468 ;
  assign y17114 = ~n46469 ;
  assign y17115 = ~n46473 ;
  assign y17116 = ~n46474 ;
  assign y17117 = n46475 ;
  assign y17118 = ~n38466 ;
  assign y17119 = ~n46476 ;
  assign y17120 = ~n46478 ;
  assign y17121 = n46482 ;
  assign y17122 = ~n46485 ;
  assign y17123 = n46490 ;
  assign y17124 = ~n46491 ;
  assign y17125 = ~n46498 ;
  assign y17126 = n46501 ;
  assign y17127 = n46503 ;
  assign y17128 = n46506 ;
  assign y17129 = ~n46508 ;
  assign y17130 = ~1'b0 ;
  assign y17131 = n46510 ;
  assign y17132 = ~1'b0 ;
  assign y17133 = n46512 ;
  assign y17134 = ~n46517 ;
  assign y17135 = n46518 ;
  assign y17136 = n46519 ;
  assign y17137 = n46522 ;
  assign y17138 = n46524 ;
  assign y17139 = ~n46527 ;
  assign y17140 = n46531 ;
  assign y17141 = ~1'b0 ;
  assign y17142 = ~n46532 ;
  assign y17143 = ~1'b0 ;
  assign y17144 = n46533 ;
  assign y17145 = ~n46536 ;
  assign y17146 = ~n46539 ;
  assign y17147 = n46542 ;
  assign y17148 = ~n46543 ;
  assign y17149 = ~n46547 ;
  assign y17150 = ~n46551 ;
  assign y17151 = n46552 ;
  assign y17152 = n46553 ;
  assign y17153 = ~n46554 ;
  assign y17154 = n46559 ;
  assign y17155 = n46565 ;
  assign y17156 = n46567 ;
  assign y17157 = ~n46569 ;
  assign y17158 = ~n46573 ;
  assign y17159 = ~1'b0 ;
  assign y17160 = ~n46575 ;
  assign y17161 = ~n46576 ;
  assign y17162 = ~n46577 ;
  assign y17163 = ~n46579 ;
  assign y17164 = ~n46581 ;
  assign y17165 = ~1'b0 ;
  assign y17166 = n46583 ;
  assign y17167 = ~n46584 ;
  assign y17168 = ~n46590 ;
  assign y17169 = ~n46593 ;
  assign y17170 = ~n46595 ;
  assign y17171 = n46597 ;
  assign y17172 = ~n46600 ;
  assign y17173 = ~n46606 ;
  assign y17174 = ~n46610 ;
  assign y17175 = ~n46612 ;
  assign y17176 = ~n46614 ;
  assign y17177 = ~n46615 ;
  assign y17178 = n46618 ;
  assign y17179 = n46622 ;
  assign y17180 = ~1'b0 ;
  assign y17181 = ~n46624 ;
  assign y17182 = n46627 ;
  assign y17183 = n46628 ;
  assign y17184 = n46632 ;
  assign y17185 = n46634 ;
  assign y17186 = ~n46636 ;
  assign y17187 = n46641 ;
  assign y17188 = n46643 ;
  assign y17189 = ~1'b0 ;
  assign y17190 = ~n46648 ;
  assign y17191 = n46654 ;
  assign y17192 = n46658 ;
  assign y17193 = ~1'b0 ;
  assign y17194 = n46663 ;
  assign y17195 = ~n46664 ;
  assign y17196 = n46665 ;
  assign y17197 = ~n46666 ;
  assign y17198 = ~n46667 ;
  assign y17199 = ~n46672 ;
  assign y17200 = n46674 ;
  assign y17201 = 1'b0 ;
  assign y17202 = n46676 ;
  assign y17203 = n46678 ;
  assign y17204 = n46679 ;
  assign y17205 = ~n46681 ;
  assign y17206 = ~n46682 ;
  assign y17207 = n46685 ;
  assign y17208 = ~n46687 ;
  assign y17209 = ~n46689 ;
  assign y17210 = ~n46691 ;
  assign y17211 = ~1'b0 ;
  assign y17212 = ~n46693 ;
  assign y17213 = n46695 ;
  assign y17214 = ~n46699 ;
  assign y17215 = ~n46700 ;
  assign y17216 = n46701 ;
  assign y17217 = n46704 ;
  assign y17218 = ~1'b0 ;
  assign y17219 = ~1'b0 ;
  assign y17220 = n46706 ;
  assign y17221 = n46710 ;
  assign y17222 = n46712 ;
  assign y17223 = n46713 ;
  assign y17224 = n46715 ;
  assign y17225 = ~n46719 ;
  assign y17226 = ~n46723 ;
  assign y17227 = ~1'b0 ;
  assign y17228 = ~n46725 ;
  assign y17229 = ~n46726 ;
  assign y17230 = ~1'b0 ;
  assign y17231 = n46727 ;
  assign y17232 = ~n46728 ;
  assign y17233 = n46729 ;
  assign y17234 = n46731 ;
  assign y17235 = ~n46734 ;
  assign y17236 = ~1'b0 ;
  assign y17237 = ~1'b0 ;
  assign y17238 = n46737 ;
  assign y17239 = ~1'b0 ;
  assign y17240 = ~n46739 ;
  assign y17241 = ~n46742 ;
  assign y17242 = n46744 ;
  assign y17243 = n46745 ;
  assign y17244 = n46754 ;
  assign y17245 = n46755 ;
  assign y17246 = ~1'b0 ;
  assign y17247 = ~n46756 ;
  assign y17248 = ~n46760 ;
  assign y17249 = n46763 ;
  assign y17250 = ~n46768 ;
  assign y17251 = n46770 ;
  assign y17252 = ~n46775 ;
  assign y17253 = n46779 ;
  assign y17254 = n46780 ;
  assign y17255 = ~n46782 ;
  assign y17256 = n46783 ;
  assign y17257 = ~1'b0 ;
  assign y17258 = ~n46785 ;
  assign y17259 = ~n46786 ;
  assign y17260 = ~n46787 ;
  assign y17261 = ~n46791 ;
  assign y17262 = n46792 ;
  assign y17263 = n46798 ;
  assign y17264 = ~1'b0 ;
  assign y17265 = ~1'b0 ;
  assign y17266 = ~1'b0 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = n46799 ;
  assign y17269 = n46801 ;
  assign y17270 = n899 ;
  assign y17271 = n46802 ;
  assign y17272 = ~n46803 ;
  assign y17273 = n46805 ;
  assign y17274 = ~n46811 ;
  assign y17275 = n46812 ;
  assign y17276 = ~n46814 ;
  assign y17277 = ~n46815 ;
  assign y17278 = n46817 ;
  assign y17279 = n31314 ;
  assign y17280 = n46819 ;
  assign y17281 = ~n46821 ;
  assign y17282 = n46823 ;
  assign y17283 = n46827 ;
  assign y17284 = ~1'b0 ;
  assign y17285 = ~1'b0 ;
  assign y17286 = ~n46829 ;
  assign y17287 = ~n46830 ;
  assign y17288 = ~n46835 ;
  assign y17289 = n46839 ;
  assign y17290 = n46845 ;
  assign y17291 = ~1'b0 ;
  assign y17292 = ~1'b0 ;
  assign y17293 = n46847 ;
  assign y17294 = n46853 ;
  assign y17295 = n46854 ;
  assign y17296 = ~n46858 ;
  assign y17297 = n46862 ;
  assign y17298 = ~n46866 ;
  assign y17299 = ~1'b0 ;
  assign y17300 = ~1'b0 ;
  assign y17301 = ~n46867 ;
  assign y17302 = n46869 ;
  assign y17303 = n46876 ;
  assign y17304 = n46877 ;
  assign y17305 = n46880 ;
  assign y17306 = n46881 ;
  assign y17307 = n46882 ;
  assign y17308 = n46886 ;
  assign y17309 = n46888 ;
  assign y17310 = ~n46891 ;
  assign y17311 = n46893 ;
  assign y17312 = n46895 ;
  assign y17313 = ~n46896 ;
  assign y17314 = n46897 ;
  assign y17315 = n46905 ;
  assign y17316 = n46907 ;
  assign y17317 = ~n19496 ;
  assign y17318 = n46912 ;
  assign y17319 = 1'b0 ;
  assign y17320 = n46913 ;
  assign y17321 = ~n46918 ;
  assign y17322 = n46920 ;
  assign y17323 = n46929 ;
  assign y17324 = n46931 ;
  assign y17325 = ~1'b0 ;
  assign y17326 = ~1'b0 ;
  assign y17327 = n46935 ;
  assign y17328 = ~n46936 ;
  assign y17329 = ~n46939 ;
  assign y17330 = ~n46941 ;
  assign y17331 = ~n46943 ;
  assign y17332 = n46944 ;
  assign y17333 = n46950 ;
  assign y17334 = n46952 ;
  assign y17335 = n46953 ;
  assign y17336 = n46956 ;
  assign y17337 = ~1'b0 ;
  assign y17338 = ~n46961 ;
  assign y17339 = ~n46963 ;
  assign y17340 = ~n46965 ;
  assign y17341 = ~n46968 ;
  assign y17342 = ~1'b0 ;
  assign y17343 = ~n46972 ;
  assign y17344 = n46976 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = ~n46979 ;
  assign y17347 = n46981 ;
  assign y17348 = n46982 ;
  assign y17349 = ~n46983 ;
  assign y17350 = n46985 ;
  assign y17351 = ~1'b0 ;
  assign y17352 = n46988 ;
  assign y17353 = n46989 ;
  assign y17354 = ~1'b0 ;
  assign y17355 = ~n13226 ;
  assign y17356 = ~1'b0 ;
  assign y17357 = ~n46991 ;
  assign y17358 = ~n46998 ;
  assign y17359 = n46999 ;
  assign y17360 = ~n47002 ;
  assign y17361 = ~n47005 ;
  assign y17362 = n47007 ;
  assign y17363 = n47008 ;
  assign y17364 = ~1'b0 ;
  assign y17365 = n47010 ;
  assign y17366 = n47011 ;
  assign y17367 = n47013 ;
  assign y17368 = ~n47015 ;
  assign y17369 = n47016 ;
  assign y17370 = ~n47017 ;
  assign y17371 = n47018 ;
  assign y17372 = n47020 ;
  assign y17373 = n47024 ;
  assign y17374 = 1'b0 ;
  assign y17375 = n47025 ;
  assign y17376 = n47029 ;
  assign y17377 = n47032 ;
  assign y17378 = ~n47035 ;
  assign y17379 = ~n47039 ;
  assign y17380 = n47041 ;
  assign y17381 = n47043 ;
  assign y17382 = ~n47044 ;
  assign y17383 = ~n47046 ;
  assign y17384 = n47047 ;
  assign y17385 = ~n47048 ;
  assign y17386 = n47049 ;
  assign y17387 = n47051 ;
  assign y17388 = n47053 ;
  assign y17389 = ~n47054 ;
  assign y17390 = ~n47058 ;
  assign y17391 = 1'b0 ;
  assign y17392 = ~n40684 ;
  assign y17393 = ~n47059 ;
  assign y17394 = ~n47063 ;
  assign y17395 = n46870 ;
  assign y17396 = ~n47073 ;
  assign y17397 = ~n47074 ;
  assign y17398 = ~1'b0 ;
  assign y17399 = n47075 ;
  assign y17400 = ~n47079 ;
  assign y17401 = n47083 ;
  assign y17402 = n47084 ;
  assign y17403 = n47085 ;
  assign y17404 = n47088 ;
  assign y17405 = ~n47089 ;
  assign y17406 = n47093 ;
  assign y17407 = n47098 ;
  assign y17408 = ~1'b0 ;
  assign y17409 = ~1'b0 ;
  assign y17410 = ~n47099 ;
  assign y17411 = n47100 ;
  assign y17412 = n47103 ;
  assign y17413 = ~n47104 ;
  assign y17414 = ~n47106 ;
  assign y17415 = ~1'b0 ;
  assign y17416 = ~n47108 ;
  assign y17417 = ~1'b0 ;
  assign y17418 = n47111 ;
  assign y17419 = ~n47113 ;
  assign y17420 = ~n47114 ;
  assign y17421 = ~n47117 ;
  assign y17422 = n47118 ;
  assign y17423 = n47121 ;
  assign y17424 = n47124 ;
  assign y17425 = ~n47125 ;
  assign y17426 = ~1'b0 ;
  assign y17427 = n47128 ;
  assign y17428 = ~n47132 ;
  assign y17429 = n47135 ;
  assign y17430 = n47140 ;
  assign y17431 = n47142 ;
  assign y17432 = ~n47145 ;
  assign y17433 = n47147 ;
  assign y17434 = n47152 ;
  assign y17435 = ~n47157 ;
  assign y17436 = ~n47159 ;
  assign y17437 = n47162 ;
  assign y17438 = n47167 ;
  assign y17439 = ~n47168 ;
  assign y17440 = ~n47171 ;
  assign y17441 = ~n47172 ;
  assign y17442 = ~n47174 ;
  assign y17443 = ~n47176 ;
  assign y17444 = ~1'b0 ;
  assign y17445 = n47178 ;
  assign y17446 = n47180 ;
  assign y17447 = n47185 ;
  assign y17448 = ~n47188 ;
  assign y17449 = n47190 ;
  assign y17450 = n47191 ;
  assign y17451 = ~n47192 ;
  assign y17452 = ~1'b0 ;
  assign y17453 = n47193 ;
  assign y17454 = n47198 ;
  assign y17455 = ~n47204 ;
  assign y17456 = ~n47207 ;
  assign y17457 = ~n47208 ;
  assign y17458 = n47209 ;
  assign y17459 = ~n47210 ;
  assign y17460 = ~n47211 ;
  assign y17461 = ~1'b0 ;
  assign y17462 = ~1'b0 ;
  assign y17463 = n47214 ;
  assign y17464 = ~n47215 ;
  assign y17465 = n47216 ;
  assign y17466 = n47218 ;
  assign y17467 = n47219 ;
  assign y17468 = n47224 ;
  assign y17469 = n47225 ;
  assign y17470 = n47228 ;
  assign y17471 = n47230 ;
  assign y17472 = n47232 ;
  assign y17473 = n47237 ;
  assign y17474 = ~n47238 ;
  assign y17475 = ~n47240 ;
  assign y17476 = ~n47242 ;
  assign y17477 = ~n47244 ;
  assign y17478 = n47249 ;
  assign y17479 = n47250 ;
  assign y17480 = n47254 ;
  assign y17481 = ~1'b0 ;
  assign y17482 = ~n47257 ;
  assign y17483 = ~n47258 ;
  assign y17484 = n47264 ;
  assign y17485 = ~n47265 ;
  assign y17486 = ~n47266 ;
  assign y17487 = ~n47267 ;
  assign y17488 = n47268 ;
  assign y17489 = ~n47269 ;
  assign y17490 = ~n47272 ;
  assign y17491 = n47275 ;
  assign y17492 = ~1'b0 ;
  assign y17493 = n17212 ;
  assign y17494 = n47282 ;
  assign y17495 = n47287 ;
  assign y17496 = n47288 ;
  assign y17497 = ~n47290 ;
  assign y17498 = ~n47291 ;
  assign y17499 = ~n47292 ;
  assign y17500 = ~n47299 ;
  assign y17501 = n47301 ;
  assign y17502 = ~1'b0 ;
  assign y17503 = n47303 ;
  assign y17504 = ~n47304 ;
  assign y17505 = ~n47306 ;
  assign y17506 = n47307 ;
  assign y17507 = ~n47308 ;
  assign y17508 = ~n47313 ;
  assign y17509 = n47314 ;
  assign y17510 = ~n47317 ;
  assign y17511 = ~n47318 ;
  assign y17512 = ~1'b0 ;
  assign y17513 = ~1'b0 ;
  assign y17514 = ~n47320 ;
  assign y17515 = ~n47323 ;
  assign y17516 = n47325 ;
  assign y17517 = n47328 ;
  assign y17518 = ~n47329 ;
  assign y17519 = ~n47330 ;
  assign y17520 = n47336 ;
  assign y17521 = ~1'b0 ;
  assign y17522 = n47338 ;
  assign y17523 = ~n47340 ;
  assign y17524 = ~n47341 ;
  assign y17525 = n47342 ;
  assign y17526 = ~n47347 ;
  assign y17527 = ~n47350 ;
  assign y17528 = n9931 ;
  assign y17529 = n47354 ;
  assign y17530 = n47356 ;
  assign y17531 = n47357 ;
  assign y17532 = n47359 ;
  assign y17533 = ~n47364 ;
  assign y17534 = ~n47365 ;
  assign y17535 = n47366 ;
  assign y17536 = ~n47374 ;
  assign y17537 = n47377 ;
  assign y17538 = n47379 ;
  assign y17539 = ~n47381 ;
  assign y17540 = ~n47384 ;
  assign y17541 = ~1'b0 ;
  assign y17542 = n47388 ;
  assign y17543 = n6958 ;
  assign y17544 = ~n47391 ;
  assign y17545 = ~n47392 ;
  assign y17546 = ~n47400 ;
  assign y17547 = ~n47402 ;
  assign y17548 = n47403 ;
  assign y17549 = ~n47404 ;
  assign y17550 = ~n47409 ;
  assign y17551 = ~1'b0 ;
  assign y17552 = n47410 ;
  assign y17553 = ~n47415 ;
  assign y17554 = n47418 ;
  assign y17555 = n47420 ;
  assign y17556 = ~n47421 ;
  assign y17557 = n47422 ;
  assign y17558 = n47424 ;
  assign y17559 = n47425 ;
  assign y17560 = ~1'b0 ;
  assign y17561 = ~n47428 ;
  assign y17562 = n47429 ;
  assign y17563 = ~1'b0 ;
  assign y17564 = n47431 ;
  assign y17565 = ~n47436 ;
  assign y17566 = n47438 ;
  assign y17567 = n47439 ;
  assign y17568 = ~1'b0 ;
  assign y17569 = ~n47441 ;
  assign y17570 = ~n47445 ;
  assign y17571 = n47447 ;
  assign y17572 = ~n40209 ;
  assign y17573 = ~n47448 ;
  assign y17574 = n47449 ;
  assign y17575 = ~n47452 ;
  assign y17576 = ~n47456 ;
  assign y17577 = ~n47460 ;
  assign y17578 = ~1'b0 ;
  assign y17579 = ~n47467 ;
  assign y17580 = ~n47472 ;
  assign y17581 = ~1'b0 ;
  assign y17582 = n47473 ;
  assign y17583 = n47474 ;
  assign y17584 = ~n47475 ;
  assign y17585 = n47476 ;
  assign y17586 = n47483 ;
  assign y17587 = ~n47484 ;
  assign y17588 = n47490 ;
  assign y17589 = ~n47492 ;
  assign y17590 = ~n47493 ;
  assign y17591 = n47495 ;
  assign y17592 = ~n47497 ;
  assign y17593 = ~n47502 ;
  assign y17594 = n47503 ;
  assign y17595 = ~n47505 ;
  assign y17596 = ~n47510 ;
  assign y17597 = ~n47512 ;
  assign y17598 = ~1'b0 ;
  assign y17599 = ~1'b0 ;
  assign y17600 = ~1'b0 ;
  assign y17601 = n47514 ;
  assign y17602 = n47515 ;
  assign y17603 = ~n47522 ;
  assign y17604 = ~1'b0 ;
  assign y17605 = n47523 ;
  assign y17606 = ~n47524 ;
  assign y17607 = n47532 ;
  assign y17608 = ~n47533 ;
  assign y17609 = ~n47534 ;
  assign y17610 = n47537 ;
  assign y17611 = n47541 ;
  assign y17612 = ~n47542 ;
  assign y17613 = n10251 ;
  assign y17614 = n47545 ;
  assign y17615 = n47546 ;
  assign y17616 = ~n47548 ;
  assign y17617 = ~1'b0 ;
  assign y17618 = ~1'b0 ;
  assign y17619 = ~1'b0 ;
  assign y17620 = ~n47549 ;
  assign y17621 = ~n47551 ;
  assign y17622 = ~n47552 ;
  assign y17623 = ~n47556 ;
  assign y17624 = n47560 ;
  assign y17625 = ~n47563 ;
  assign y17626 = ~n47564 ;
  assign y17627 = ~n47566 ;
  assign y17628 = ~1'b0 ;
  assign y17629 = n3285 ;
  assign y17630 = n47568 ;
  assign y17631 = ~n47569 ;
  assign y17632 = ~n29915 ;
  assign y17633 = n47572 ;
  assign y17634 = ~1'b0 ;
  assign y17635 = ~n47573 ;
  assign y17636 = ~n47577 ;
  assign y17637 = ~n47580 ;
  assign y17638 = n47581 ;
  assign y17639 = n47585 ;
  assign y17640 = n47586 ;
  assign y17641 = n47589 ;
  assign y17642 = ~n47591 ;
  assign y17643 = 1'b0 ;
  assign y17644 = n47593 ;
  assign y17645 = n47597 ;
  assign y17646 = n47598 ;
  assign y17647 = n47599 ;
  assign y17648 = ~n47601 ;
  assign y17649 = ~n47604 ;
  assign y17650 = ~1'b0 ;
  assign y17651 = n47606 ;
  assign y17652 = n47608 ;
  assign y17653 = ~n47610 ;
  assign y17654 = ~1'b0 ;
  assign y17655 = ~n47613 ;
  assign y17656 = n47616 ;
  assign y17657 = n47617 ;
  assign y17658 = ~1'b0 ;
  assign y17659 = ~n47619 ;
  assign y17660 = n47621 ;
  assign y17661 = ~1'b0 ;
  assign y17662 = ~1'b0 ;
  assign y17663 = ~1'b0 ;
  assign y17664 = ~n47623 ;
  assign y17665 = ~1'b0 ;
  assign y17666 = ~n47626 ;
  assign y17667 = n47629 ;
  assign y17668 = ~n47631 ;
  assign y17669 = n47632 ;
  assign y17670 = ~n47633 ;
  assign y17671 = ~n47635 ;
  assign y17672 = ~1'b0 ;
  assign y17673 = ~n47638 ;
  assign y17674 = ~n47641 ;
  assign y17675 = ~n47643 ;
  assign y17676 = n47644 ;
  assign y17677 = ~n47647 ;
  assign y17678 = ~n47650 ;
  assign y17679 = ~n47652 ;
  assign y17680 = ~n47653 ;
  assign y17681 = ~n47655 ;
  assign y17682 = ~n47657 ;
  assign y17683 = n47660 ;
  assign y17684 = ~n47662 ;
  assign y17685 = ~1'b0 ;
  assign y17686 = n47663 ;
  assign y17687 = ~n47666 ;
  assign y17688 = ~n47671 ;
  assign y17689 = n47674 ;
  assign y17690 = n47677 ;
  assign y17691 = ~n47680 ;
  assign y17692 = ~1'b0 ;
  assign y17693 = n47682 ;
  assign y17694 = ~1'b0 ;
  assign y17695 = n47685 ;
  assign y17696 = ~n47687 ;
  assign y17697 = ~n47688 ;
  assign y17698 = n47690 ;
  assign y17699 = ~n47695 ;
  assign y17700 = n47696 ;
  assign y17701 = n26266 ;
  assign y17702 = ~n47697 ;
  assign y17703 = ~n47703 ;
  assign y17704 = ~1'b0 ;
  assign y17705 = ~n47705 ;
  assign y17706 = ~n47709 ;
  assign y17707 = ~n47711 ;
  assign y17708 = ~n47715 ;
  assign y17709 = ~n47717 ;
  assign y17710 = n47722 ;
  assign y17711 = ~n47725 ;
  assign y17712 = n47727 ;
  assign y17713 = ~1'b0 ;
  assign y17714 = n47728 ;
  assign y17715 = ~n47731 ;
  assign y17716 = ~n47733 ;
  assign y17717 = n47734 ;
  assign y17718 = ~n47735 ;
  assign y17719 = ~n47737 ;
  assign y17720 = ~n47739 ;
  assign y17721 = n47750 ;
  assign y17722 = n47751 ;
  assign y17723 = ~n47753 ;
  assign y17724 = n47754 ;
  assign y17725 = n47760 ;
  assign y17726 = n47761 ;
  assign y17727 = n47766 ;
  assign y17728 = ~1'b0 ;
  assign y17729 = ~n47770 ;
  assign y17730 = ~1'b0 ;
  assign y17731 = ~n47772 ;
  assign y17732 = ~1'b0 ;
  assign y17733 = n47773 ;
  assign y17734 = ~n47774 ;
  assign y17735 = n31468 ;
  assign y17736 = n47776 ;
  assign y17737 = n47777 ;
  assign y17738 = ~n47781 ;
  assign y17739 = n47783 ;
  assign y17740 = ~n47785 ;
  assign y17741 = n47787 ;
  assign y17742 = ~n47789 ;
  assign y17743 = ~n47791 ;
  assign y17744 = ~n47793 ;
  assign y17745 = ~n47796 ;
  assign y17746 = n47799 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = n47801 ;
  assign y17749 = ~n47802 ;
  assign y17750 = n47804 ;
  assign y17751 = ~n47808 ;
  assign y17752 = ~n47810 ;
  assign y17753 = ~n47815 ;
  assign y17754 = n47816 ;
  assign y17755 = n47818 ;
  assign y17756 = ~n47819 ;
  assign y17757 = n47821 ;
  assign y17758 = n47822 ;
  assign y17759 = ~1'b0 ;
  assign y17760 = n47823 ;
  assign y17761 = ~n47827 ;
  assign y17762 = n47833 ;
  assign y17763 = n47837 ;
  assign y17764 = n47840 ;
  assign y17765 = ~n47842 ;
  assign y17766 = ~n47845 ;
  assign y17767 = n23521 ;
  assign y17768 = ~1'b0 ;
  assign y17769 = n47846 ;
  assign y17770 = ~n47848 ;
  assign y17771 = ~1'b0 ;
  assign y17772 = ~n47850 ;
  assign y17773 = n47855 ;
  assign y17774 = ~n47856 ;
  assign y17775 = ~n47857 ;
  assign y17776 = ~n47858 ;
  assign y17777 = ~1'b0 ;
  assign y17778 = ~1'b0 ;
  assign y17779 = n47861 ;
  assign y17780 = n23626 ;
  assign y17781 = n47863 ;
  assign y17782 = ~n47865 ;
  assign y17783 = n47866 ;
  assign y17784 = ~n47867 ;
  assign y17785 = ~n47870 ;
  assign y17786 = ~n47872 ;
  assign y17787 = 1'b0 ;
  assign y17788 = ~n47873 ;
  assign y17789 = n47876 ;
  assign y17790 = n47878 ;
  assign y17791 = ~n47882 ;
  assign y17792 = ~1'b0 ;
  assign y17793 = ~n47883 ;
  assign y17794 = ~n47886 ;
  assign y17795 = ~n47888 ;
  assign y17796 = n47894 ;
  assign y17797 = ~n47900 ;
  assign y17798 = ~1'b0 ;
  assign y17799 = ~n47904 ;
  assign y17800 = n47908 ;
  assign y17801 = n47910 ;
  assign y17802 = ~n47911 ;
  assign y17803 = n47918 ;
  assign y17804 = n47920 ;
  assign y17805 = ~1'b0 ;
  assign y17806 = n47921 ;
  assign y17807 = ~n47922 ;
  assign y17808 = ~1'b0 ;
  assign y17809 = n47924 ;
  assign y17810 = ~n47926 ;
  assign y17811 = n47930 ;
  assign y17812 = n47933 ;
  assign y17813 = n47935 ;
  assign y17814 = ~n47940 ;
  assign y17815 = ~n47942 ;
  assign y17816 = n47944 ;
  assign y17817 = ~1'b0 ;
  assign y17818 = n31490 ;
  assign y17819 = ~n47946 ;
  assign y17820 = ~1'b0 ;
  assign y17821 = n47947 ;
  assign y17822 = ~n47951 ;
  assign y17823 = ~n47952 ;
  assign y17824 = n30886 ;
  assign y17825 = ~n47953 ;
  assign y17826 = ~1'b0 ;
  assign y17827 = ~1'b0 ;
  assign y17828 = ~n47955 ;
  assign y17829 = ~n47957 ;
  assign y17830 = ~1'b0 ;
  assign y17831 = n47963 ;
  assign y17832 = ~n47966 ;
  assign y17833 = n47967 ;
  assign y17834 = n47968 ;
  assign y17835 = n47971 ;
  assign y17836 = n47972 ;
  assign y17837 = ~n47976 ;
  assign y17838 = ~n47978 ;
  assign y17839 = ~n47986 ;
  assign y17840 = ~1'b0 ;
  assign y17841 = ~1'b0 ;
  assign y17842 = n47990 ;
  assign y17843 = n47992 ;
  assign y17844 = ~n47993 ;
  assign y17845 = ~n47996 ;
  assign y17846 = ~1'b0 ;
  assign y17847 = n47998 ;
  assign y17848 = ~1'b0 ;
  assign y17849 = ~1'b0 ;
  assign y17850 = n48003 ;
  assign y17851 = n48007 ;
  assign y17852 = ~n48008 ;
  assign y17853 = n48011 ;
  assign y17854 = ~n48013 ;
  assign y17855 = n48016 ;
  assign y17856 = ~1'b0 ;
  assign y17857 = ~1'b0 ;
  assign y17858 = n48018 ;
  assign y17859 = ~n48020 ;
  assign y17860 = ~1'b0 ;
  assign y17861 = n48026 ;
  assign y17862 = n48027 ;
  assign y17863 = ~n48033 ;
  assign y17864 = ~1'b0 ;
  assign y17865 = ~n48037 ;
  assign y17866 = ~1'b0 ;
  assign y17867 = ~1'b0 ;
  assign y17868 = ~1'b0 ;
  assign y17869 = ~n48039 ;
  assign y17870 = n48043 ;
  assign y17871 = ~1'b0 ;
  assign y17872 = ~n48047 ;
  assign y17873 = ~n48051 ;
  assign y17874 = n48052 ;
  assign y17875 = ~n48053 ;
  assign y17876 = ~n48054 ;
  assign y17877 = ~1'b0 ;
  assign y17878 = ~1'b0 ;
  assign y17879 = ~1'b0 ;
  assign y17880 = ~n48057 ;
  assign y17881 = n48058 ;
  assign y17882 = ~n48061 ;
  assign y17883 = ~n48062 ;
  assign y17884 = ~n48063 ;
  assign y17885 = ~n48064 ;
  assign y17886 = ~n48066 ;
  assign y17887 = ~n48067 ;
  assign y17888 = ~n48071 ;
  assign y17889 = ~1'b0 ;
  assign y17890 = n48075 ;
  assign y17891 = ~n48076 ;
  assign y17892 = n48077 ;
  assign y17893 = n48080 ;
  assign y17894 = n48081 ;
  assign y17895 = n48084 ;
  assign y17896 = ~n48086 ;
  assign y17897 = ~1'b0 ;
  assign y17898 = ~1'b0 ;
  assign y17899 = n48088 ;
  assign y17900 = ~n48094 ;
  assign y17901 = n48098 ;
  assign y17902 = n48103 ;
  assign y17903 = n48109 ;
  assign y17904 = ~n48113 ;
  assign y17905 = n13828 ;
  assign y17906 = ~n48115 ;
  assign y17907 = ~n48116 ;
  assign y17908 = ~n48118 ;
  assign y17909 = n48119 ;
  assign y17910 = n48122 ;
  assign y17911 = ~1'b0 ;
  assign y17912 = ~n48123 ;
  assign y17913 = n48125 ;
  assign y17914 = ~n48126 ;
  assign y17915 = n48133 ;
  assign y17916 = n48134 ;
  assign y17917 = 1'b0 ;
  assign y17918 = ~n48135 ;
  assign y17919 = n48140 ;
  assign y17920 = ~n48144 ;
  assign y17921 = ~1'b0 ;
  assign y17922 = ~n48145 ;
  assign y17923 = n48146 ;
  assign y17924 = ~n48155 ;
  assign y17925 = n48158 ;
  assign y17926 = ~n48161 ;
  assign y17927 = n48162 ;
  assign y17928 = ~n48166 ;
  assign y17929 = n48169 ;
  assign y17930 = ~1'b0 ;
  assign y17931 = ~n48170 ;
  assign y17932 = n48175 ;
  assign y17933 = n48178 ;
  assign y17934 = ~n48179 ;
  assign y17935 = ~n48185 ;
  assign y17936 = ~n48186 ;
  assign y17937 = ~1'b0 ;
  assign y17938 = ~n48188 ;
  assign y17939 = n48190 ;
  assign y17940 = ~n48194 ;
  assign y17941 = ~1'b0 ;
  assign y17942 = ~n48195 ;
  assign y17943 = n48201 ;
  assign y17944 = ~n48202 ;
  assign y17945 = n48212 ;
  assign y17946 = n48215 ;
  assign y17947 = n48217 ;
  assign y17948 = ~n48219 ;
  assign y17949 = ~1'b0 ;
  assign y17950 = ~n48220 ;
  assign y17951 = ~n48221 ;
  assign y17952 = ~n48222 ;
  assign y17953 = n48225 ;
  assign y17954 = ~n48226 ;
  assign y17955 = n48228 ;
  assign y17956 = ~1'b0 ;
  assign y17957 = ~n48232 ;
  assign y17958 = ~1'b0 ;
  assign y17959 = n48233 ;
  assign y17960 = n48239 ;
  assign y17961 = n48240 ;
  assign y17962 = n48244 ;
  assign y17963 = n48247 ;
  assign y17964 = n33958 ;
  assign y17965 = n48253 ;
  assign y17966 = n48255 ;
  assign y17967 = n48257 ;
  assign y17968 = ~n48259 ;
  assign y17969 = n48264 ;
  assign y17970 = ~n48265 ;
  assign y17971 = ~n48266 ;
  assign y17972 = ~n48267 ;
  assign y17973 = ~n48271 ;
  assign y17974 = n48272 ;
  assign y17975 = n48274 ;
  assign y17976 = ~1'b0 ;
  assign y17977 = n48280 ;
  assign y17978 = ~n48281 ;
  assign y17979 = n48285 ;
  assign y17980 = n48286 ;
  assign y17981 = ~n48287 ;
  assign y17982 = n48291 ;
  assign y17983 = ~1'b0 ;
  assign y17984 = n48294 ;
  assign y17985 = ~n48296 ;
  assign y17986 = ~1'b0 ;
  assign y17987 = ~n48298 ;
  assign y17988 = n48300 ;
  assign y17989 = n48301 ;
  assign y17990 = ~n48304 ;
  assign y17991 = n48305 ;
  assign y17992 = n48306 ;
  assign y17993 = ~n48307 ;
  assign y17994 = n48309 ;
  assign y17995 = n48315 ;
  assign y17996 = ~1'b0 ;
  assign y17997 = n48316 ;
  assign y17998 = ~1'b0 ;
  assign y17999 = ~n48318 ;
  assign y18000 = ~n48322 ;
  assign y18001 = ~n48323 ;
  assign y18002 = ~n48324 ;
  assign y18003 = n48327 ;
  assign y18004 = ~n48333 ;
  assign y18005 = ~n48335 ;
  assign y18006 = ~n48336 ;
  assign y18007 = n48338 ;
  assign y18008 = ~1'b0 ;
  assign y18009 = ~1'b0 ;
  assign y18010 = ~n48340 ;
  assign y18011 = ~n48347 ;
  assign y18012 = ~n48351 ;
  assign y18013 = ~n48352 ;
  assign y18014 = n48353 ;
  assign y18015 = ~1'b0 ;
  assign y18016 = n48355 ;
  assign y18017 = n16864 ;
  assign y18018 = n48358 ;
  assign y18019 = n48363 ;
  assign y18020 = ~1'b0 ;
  assign y18021 = ~n48364 ;
  assign y18022 = ~n48367 ;
  assign y18023 = ~n48368 ;
  assign y18024 = n48370 ;
  assign y18025 = n48376 ;
  assign y18026 = n48378 ;
  assign y18027 = n48382 ;
  assign y18028 = ~n48385 ;
  assign y18029 = ~n48387 ;
  assign y18030 = ~1'b0 ;
  assign y18031 = n48393 ;
  assign y18032 = ~n34088 ;
  assign y18033 = n48394 ;
  assign y18034 = n48397 ;
  assign y18035 = n48400 ;
  assign y18036 = n48404 ;
  assign y18037 = n48405 ;
  assign y18038 = n48406 ;
  assign y18039 = ~n48412 ;
  assign y18040 = ~n48416 ;
  assign y18041 = ~n48417 ;
  assign y18042 = n48420 ;
  assign y18043 = ~n48427 ;
  assign y18044 = ~n48430 ;
  assign y18045 = n48434 ;
  assign y18046 = ~1'b0 ;
  assign y18047 = ~n48436 ;
  assign y18048 = 1'b0 ;
  assign y18049 = ~n48440 ;
  assign y18050 = n48442 ;
  assign y18051 = n48445 ;
  assign y18052 = n48451 ;
  assign y18053 = ~1'b0 ;
  assign y18054 = n48452 ;
  assign y18055 = ~n48454 ;
  assign y18056 = ~n48456 ;
  assign y18057 = n48458 ;
  assign y18058 = n48462 ;
  assign y18059 = n48463 ;
  assign y18060 = ~n48466 ;
  assign y18061 = n48469 ;
  assign y18062 = ~n48472 ;
  assign y18063 = ~n48474 ;
  assign y18064 = n48480 ;
  assign y18065 = ~1'b0 ;
  assign y18066 = ~1'b0 ;
  assign y18067 = ~n48483 ;
  assign y18068 = n48485 ;
  assign y18069 = n48486 ;
  assign y18070 = ~n48488 ;
  assign y18071 = ~n48489 ;
  assign y18072 = n48490 ;
  assign y18073 = n48495 ;
  assign y18074 = ~1'b0 ;
  assign y18075 = ~n48502 ;
  assign y18076 = ~n48506 ;
  assign y18077 = n48507 ;
  assign y18078 = n48516 ;
  assign y18079 = n48518 ;
  assign y18080 = ~n48519 ;
  assign y18081 = n26020 ;
  assign y18082 = n48520 ;
  assign y18083 = ~n48521 ;
  assign y18084 = ~1'b0 ;
  assign y18085 = n48523 ;
  assign y18086 = n48525 ;
  assign y18087 = ~n48527 ;
  assign y18088 = ~n48528 ;
  assign y18089 = ~n48529 ;
  assign y18090 = n48533 ;
  assign y18091 = ~n48534 ;
  assign y18092 = ~1'b0 ;
  assign y18093 = ~1'b0 ;
  assign y18094 = ~n48538 ;
  assign y18095 = ~n48541 ;
  assign y18096 = ~n48542 ;
  assign y18097 = ~1'b0 ;
  assign y18098 = n48552 ;
  assign y18099 = ~n48554 ;
  assign y18100 = n48555 ;
  assign y18101 = ~n48557 ;
  assign y18102 = ~n48558 ;
  assign y18103 = ~1'b0 ;
  assign y18104 = ~1'b0 ;
  assign y18105 = n48559 ;
  assign y18106 = n48565 ;
  assign y18107 = n48566 ;
  assign y18108 = n48567 ;
  assign y18109 = ~n48569 ;
  assign y18110 = ~n48572 ;
  assign y18111 = n48574 ;
  assign y18112 = n48576 ;
  assign y18113 = ~1'b0 ;
  assign y18114 = n48579 ;
  assign y18115 = n48580 ;
  assign y18116 = n48583 ;
  assign y18117 = n48584 ;
  assign y18118 = ~n48588 ;
  assign y18119 = ~n48590 ;
  assign y18120 = n48592 ;
  assign y18121 = n48593 ;
  assign y18122 = ~1'b0 ;
  assign y18123 = ~n48594 ;
  assign y18124 = ~n48596 ;
  assign y18125 = ~1'b0 ;
  assign y18126 = ~n48599 ;
  assign y18127 = ~n48600 ;
  assign y18128 = n48601 ;
  assign y18129 = n48603 ;
  assign y18130 = ~n48613 ;
  assign y18131 = n48616 ;
  assign y18132 = n48619 ;
  assign y18133 = n48623 ;
  assign y18134 = ~n48624 ;
  assign y18135 = ~n48627 ;
  assign y18136 = ~1'b0 ;
  assign y18137 = ~1'b0 ;
  assign y18138 = ~n48628 ;
  assign y18139 = n48631 ;
  assign y18140 = n48634 ;
  assign y18141 = ~n48635 ;
  assign y18142 = n48636 ;
  assign y18143 = n48637 ;
  assign y18144 = ~n48639 ;
  assign y18145 = ~n48640 ;
  assign y18146 = ~n48642 ;
  assign y18147 = ~1'b0 ;
  assign y18148 = ~n48645 ;
  assign y18149 = ~n48646 ;
  assign y18150 = n48647 ;
  assign y18151 = n48656 ;
  assign y18152 = ~n48657 ;
  assign y18153 = n48668 ;
  assign y18154 = n48671 ;
  assign y18155 = ~n48674 ;
  assign y18156 = n48676 ;
  assign y18157 = ~n48678 ;
  assign y18158 = ~n20008 ;
  assign y18159 = ~n48679 ;
  assign y18160 = n48680 ;
  assign y18161 = ~n48681 ;
  assign y18162 = ~1'b0 ;
  assign y18163 = n48686 ;
  assign y18164 = ~1'b0 ;
  assign y18165 = ~n48690 ;
  assign y18166 = ~1'b0 ;
  assign y18167 = n48696 ;
  assign y18168 = n48704 ;
  assign y18169 = n48705 ;
  assign y18170 = ~n48708 ;
  assign y18171 = ~n48710 ;
  assign y18172 = n48711 ;
  assign y18173 = ~n27870 ;
  assign y18174 = ~n48713 ;
  assign y18175 = n48715 ;
  assign y18176 = ~1'b0 ;
  assign y18177 = n48717 ;
  assign y18178 = n48718 ;
  assign y18179 = n48721 ;
  assign y18180 = ~n48724 ;
  assign y18181 = n48725 ;
  assign y18182 = ~n48726 ;
  assign y18183 = ~n48730 ;
  assign y18184 = ~1'b0 ;
  assign y18185 = ~n48731 ;
  assign y18186 = ~n48733 ;
  assign y18187 = ~1'b0 ;
  assign y18188 = n48736 ;
  assign y18189 = n48737 ;
  assign y18190 = n48741 ;
  assign y18191 = n48743 ;
  assign y18192 = n48745 ;
  assign y18193 = ~1'b0 ;
  assign y18194 = n48747 ;
  assign y18195 = n48750 ;
  assign y18196 = ~n48751 ;
  assign y18197 = n48753 ;
  assign y18198 = n8136 ;
  assign y18199 = ~n48754 ;
  assign y18200 = n48755 ;
  assign y18201 = n48756 ;
  assign y18202 = n48759 ;
  assign y18203 = n48760 ;
  assign y18204 = n48761 ;
  assign y18205 = ~1'b0 ;
  assign y18206 = n48762 ;
  assign y18207 = n48764 ;
  assign y18208 = ~n48767 ;
  assign y18209 = ~n48768 ;
  assign y18210 = ~n48771 ;
  assign y18211 = n48773 ;
  assign y18212 = ~1'b0 ;
  assign y18213 = n48775 ;
  assign y18214 = ~1'b0 ;
  assign y18215 = n48777 ;
  assign y18216 = ~1'b0 ;
  assign y18217 = ~1'b0 ;
  assign y18218 = ~1'b0 ;
  assign y18219 = n48783 ;
  assign y18220 = n48784 ;
  assign y18221 = n48785 ;
  assign y18222 = ~1'b0 ;
  assign y18223 = n16116 ;
  assign y18224 = ~1'b0 ;
  assign y18225 = ~n48788 ;
  assign y18226 = n48795 ;
  assign y18227 = ~n48800 ;
  assign y18228 = n48805 ;
  assign y18229 = ~n48806 ;
  assign y18230 = n48813 ;
  assign y18231 = ~n48818 ;
  assign y18232 = ~n48820 ;
  assign y18233 = ~n48824 ;
  assign y18234 = ~1'b0 ;
  assign y18235 = ~n48826 ;
  assign y18236 = ~n48827 ;
  assign y18237 = ~n48829 ;
  assign y18238 = n5208 ;
  assign y18239 = ~n48831 ;
  assign y18240 = ~n48839 ;
  assign y18241 = n48841 ;
  assign y18242 = n48846 ;
  assign y18243 = n48848 ;
  assign y18244 = ~1'b0 ;
  assign y18245 = ~n48852 ;
  assign y18246 = ~n48854 ;
  assign y18247 = ~n48855 ;
  assign y18248 = n48856 ;
  assign y18249 = n48858 ;
  assign y18250 = n48860 ;
  assign y18251 = n48862 ;
  assign y18252 = ~n48864 ;
  assign y18253 = n48867 ;
  assign y18254 = n48870 ;
  assign y18255 = ~n48871 ;
  assign y18256 = ~1'b0 ;
  assign y18257 = ~n48873 ;
  assign y18258 = n48874 ;
  assign y18259 = ~n48881 ;
  assign y18260 = ~n48882 ;
  assign y18261 = n48884 ;
  assign y18262 = ~n48885 ;
  assign y18263 = n48886 ;
  assign y18264 = ~1'b0 ;
  assign y18265 = ~1'b0 ;
  assign y18266 = ~1'b0 ;
  assign y18267 = n48889 ;
  assign y18268 = n48890 ;
  assign y18269 = n48892 ;
  assign y18270 = n48899 ;
  assign y18271 = ~n15928 ;
  assign y18272 = ~n48902 ;
  assign y18273 = ~n48905 ;
  assign y18274 = ~1'b0 ;
  assign y18275 = ~n48906 ;
  assign y18276 = n48908 ;
  assign y18277 = n48910 ;
  assign y18278 = ~n48915 ;
  assign y18279 = ~n48918 ;
  assign y18280 = ~n48919 ;
  assign y18281 = ~n48922 ;
  assign y18282 = n48926 ;
  assign y18283 = ~n48930 ;
  assign y18284 = n48935 ;
  assign y18285 = n48937 ;
  assign y18286 = ~n48938 ;
  assign y18287 = ~n48940 ;
  assign y18288 = n48941 ;
  assign y18289 = ~n48943 ;
  assign y18290 = ~n48945 ;
  assign y18291 = ~n48947 ;
  assign y18292 = ~n48953 ;
  assign y18293 = ~n48956 ;
  assign y18294 = ~1'b0 ;
  assign y18295 = ~n48957 ;
  assign y18296 = n48958 ;
  assign y18297 = ~n48960 ;
  assign y18298 = n48962 ;
  assign y18299 = n48967 ;
  assign y18300 = n48970 ;
  assign y18301 = ~n48971 ;
  assign y18302 = n48972 ;
  assign y18303 = ~n48975 ;
  assign y18304 = ~n48978 ;
  assign y18305 = n48980 ;
  assign y18306 = ~1'b0 ;
  assign y18307 = ~n48981 ;
  assign y18308 = n48983 ;
  assign y18309 = ~n48985 ;
  assign y18310 = n48986 ;
  assign y18311 = n48989 ;
  assign y18312 = ~n48993 ;
  assign y18313 = ~n6438 ;
  assign y18314 = n48994 ;
  assign y18315 = n48996 ;
  assign y18316 = ~n49000 ;
  assign y18317 = ~n49001 ;
  assign y18318 = n49003 ;
  assign y18319 = n49005 ;
  assign y18320 = ~n49006 ;
  assign y18321 = ~n49007 ;
  assign y18322 = ~n49010 ;
  assign y18323 = n49012 ;
  assign y18324 = ~1'b0 ;
  assign y18325 = ~n49019 ;
  assign y18326 = ~1'b0 ;
  assign y18327 = ~n49021 ;
  assign y18328 = ~n49022 ;
  assign y18329 = ~1'b0 ;
  assign y18330 = n49024 ;
  assign y18331 = n26619 ;
  assign y18332 = ~n49025 ;
  assign y18333 = n49028 ;
  assign y18334 = n49029 ;
  assign y18335 = n49031 ;
  assign y18336 = ~1'b0 ;
  assign y18337 = ~n49036 ;
  assign y18338 = ~1'b0 ;
  assign y18339 = ~n46575 ;
  assign y18340 = n49038 ;
  assign y18341 = n49041 ;
  assign y18342 = n11913 ;
  assign y18343 = ~n49044 ;
  assign y18344 = n49045 ;
  assign y18345 = n49048 ;
  assign y18346 = n49050 ;
  assign y18347 = ~1'b0 ;
  assign y18348 = ~1'b0 ;
  assign y18349 = ~1'b0 ;
  assign y18350 = ~n49052 ;
  assign y18351 = ~n49053 ;
  assign y18352 = ~n49056 ;
  assign y18353 = n49057 ;
  assign y18354 = ~n49062 ;
  assign y18355 = ~1'b0 ;
  assign y18356 = ~n49064 ;
  assign y18357 = ~1'b0 ;
  assign y18358 = ~n49066 ;
  assign y18359 = 1'b0 ;
  assign y18360 = ~n49071 ;
  assign y18361 = ~n49072 ;
  assign y18362 = n49073 ;
  assign y18363 = n49078 ;
  assign y18364 = n49082 ;
  assign y18365 = n49083 ;
  assign y18366 = ~n49085 ;
  assign y18367 = n49087 ;
  assign y18368 = ~1'b0 ;
  assign y18369 = ~n49088 ;
  assign y18370 = ~n49090 ;
  assign y18371 = ~n49091 ;
  assign y18372 = ~n49092 ;
  assign y18373 = ~n49093 ;
  assign y18374 = ~n49095 ;
  assign y18375 = ~n49097 ;
  assign y18376 = ~n49101 ;
  assign y18377 = ~n49105 ;
  assign y18378 = ~1'b0 ;
  assign y18379 = n9596 ;
  assign y18380 = ~n49106 ;
  assign y18381 = n49108 ;
  assign y18382 = ~1'b0 ;
  assign y18383 = ~n49109 ;
  assign y18384 = ~n49110 ;
  assign y18385 = ~n49114 ;
  assign y18386 = n49117 ;
  assign y18387 = ~1'b0 ;
  assign y18388 = ~n49122 ;
  assign y18389 = n26609 ;
  assign y18390 = ~n22470 ;
  assign y18391 = ~n49123 ;
  assign y18392 = ~n49124 ;
  assign y18393 = n49125 ;
  assign y18394 = n28611 ;
  assign y18395 = ~n49131 ;
  assign y18396 = n49132 ;
  assign y18397 = n49133 ;
  assign y18398 = ~1'b0 ;
  assign y18399 = ~n49135 ;
  assign y18400 = n49136 ;
  assign y18401 = n49138 ;
  assign y18402 = n49140 ;
  assign y18403 = ~n49144 ;
  assign y18404 = ~n49146 ;
  assign y18405 = n49148 ;
  assign y18406 = ~n49153 ;
  assign y18407 = n49156 ;
  assign y18408 = ~n49158 ;
  assign y18409 = n12222 ;
  assign y18410 = ~1'b0 ;
  assign y18411 = n49161 ;
  assign y18412 = ~n49162 ;
  assign y18413 = ~n49163 ;
  assign y18414 = n49173 ;
  assign y18415 = n49174 ;
  assign y18416 = ~n49175 ;
  assign y18417 = n49183 ;
  assign y18418 = ~n49188 ;
  assign y18419 = n49191 ;
  assign y18420 = ~1'b0 ;
  assign y18421 = ~1'b0 ;
  assign y18422 = n49193 ;
  assign y18423 = ~1'b0 ;
  assign y18424 = ~n49195 ;
  assign y18425 = ~n49196 ;
  assign y18426 = ~n49199 ;
  assign y18427 = ~n49202 ;
  assign y18428 = ~n49203 ;
  assign y18429 = n49206 ;
  assign y18430 = 1'b0 ;
  assign y18431 = n49210 ;
  assign y18432 = n49217 ;
  assign y18433 = ~n49220 ;
  assign y18434 = ~n49221 ;
  assign y18435 = ~n49225 ;
  assign y18436 = n49230 ;
  assign y18437 = ~1'b0 ;
  assign y18438 = n49232 ;
  assign y18439 = n49237 ;
  assign y18440 = ~1'b0 ;
  assign y18441 = n49239 ;
  assign y18442 = ~n49242 ;
  assign y18443 = n49243 ;
  assign y18444 = ~n49245 ;
  assign y18445 = ~n49246 ;
  assign y18446 = ~n49247 ;
  assign y18447 = ~n49250 ;
  assign y18448 = n49251 ;
  assign y18449 = n49252 ;
  assign y18450 = n49255 ;
  assign y18451 = n49257 ;
  assign y18452 = ~n49261 ;
  assign y18453 = ~n49266 ;
  assign y18454 = ~n49267 ;
  assign y18455 = n49270 ;
  assign y18456 = ~n49271 ;
  assign y18457 = ~n49272 ;
  assign y18458 = ~1'b0 ;
  assign y18459 = n49274 ;
  assign y18460 = n49278 ;
  assign y18461 = ~n49280 ;
  assign y18462 = ~n49285 ;
  assign y18463 = n49287 ;
  assign y18464 = ~n49289 ;
  assign y18465 = n49297 ;
  assign y18466 = ~n49301 ;
  assign y18467 = ~n49302 ;
  assign y18468 = n49304 ;
  assign y18469 = ~1'b0 ;
  assign y18470 = n49306 ;
  assign y18471 = ~1'b0 ;
  assign y18472 = n49308 ;
  assign y18473 = ~n49311 ;
  assign y18474 = n49314 ;
  assign y18475 = n49316 ;
  assign y18476 = n49317 ;
  assign y18477 = ~n49318 ;
  assign y18478 = n49319 ;
  assign y18479 = ~n49321 ;
  assign y18480 = ~n49323 ;
  assign y18481 = ~1'b0 ;
  assign y18482 = ~n49326 ;
  assign y18483 = n49328 ;
  assign y18484 = ~n44630 ;
  assign y18485 = ~n49329 ;
  assign y18486 = ~n49332 ;
  assign y18487 = ~n49335 ;
  assign y18488 = ~n49338 ;
  assign y18489 = ~n49340 ;
  assign y18490 = n49344 ;
  assign y18491 = ~n49345 ;
  assign y18492 = n49348 ;
  assign y18493 = n2497 ;
  assign y18494 = ~n49350 ;
  assign y18495 = ~n49355 ;
  assign y18496 = n49356 ;
  assign y18497 = n49357 ;
  assign y18498 = ~1'b0 ;
  assign y18499 = ~n49359 ;
  assign y18500 = ~1'b0 ;
  assign y18501 = n49360 ;
  assign y18502 = ~n49364 ;
  assign y18503 = ~n49365 ;
  assign y18504 = ~n49367 ;
  assign y18505 = ~1'b0 ;
  assign y18506 = n49368 ;
  assign y18507 = ~1'b0 ;
  assign y18508 = ~1'b0 ;
  assign y18509 = ~n49372 ;
  assign y18510 = ~n49373 ;
  assign y18511 = n49375 ;
  assign y18512 = ~n49377 ;
  assign y18513 = n49378 ;
  assign y18514 = ~n49381 ;
  assign y18515 = ~1'b0 ;
  assign y18516 = ~n49383 ;
  assign y18517 = n49384 ;
  assign y18518 = n49385 ;
  assign y18519 = n29416 ;
  assign y18520 = ~n49392 ;
  assign y18521 = ~n49394 ;
  assign y18522 = n49396 ;
  assign y18523 = ~n49399 ;
  assign y18524 = n49401 ;
  assign y18525 = ~n49402 ;
  assign y18526 = ~n49403 ;
  assign y18527 = n49405 ;
  assign y18528 = n49408 ;
  assign y18529 = ~1'b0 ;
  assign y18530 = ~n49410 ;
  assign y18531 = n49417 ;
  assign y18532 = n49419 ;
  assign y18533 = n49420 ;
  assign y18534 = ~n49424 ;
  assign y18535 = n49427 ;
  assign y18536 = ~1'b0 ;
  assign y18537 = ~n49432 ;
  assign y18538 = ~1'b0 ;
  assign y18539 = ~1'b0 ;
  assign y18540 = n49434 ;
  assign y18541 = n49436 ;
  assign y18542 = ~n49438 ;
  assign y18543 = ~n36543 ;
  assign y18544 = n49443 ;
  assign y18545 = ~n49444 ;
  assign y18546 = ~n49447 ;
  assign y18547 = ~1'b0 ;
  assign y18548 = n49449 ;
  assign y18549 = n49451 ;
  assign y18550 = n49455 ;
  assign y18551 = ~n49457 ;
  assign y18552 = n49460 ;
  assign y18553 = n49461 ;
  assign y18554 = ~n49463 ;
  assign y18555 = ~n49465 ;
  assign y18556 = n49469 ;
  assign y18557 = n49472 ;
  assign y18558 = ~1'b0 ;
  assign y18559 = ~n49476 ;
  assign y18560 = n49477 ;
  assign y18561 = ~1'b0 ;
  assign y18562 = ~n49479 ;
  assign y18563 = n49482 ;
  assign y18564 = n49483 ;
  assign y18565 = ~n49484 ;
  assign y18566 = ~n49485 ;
  assign y18567 = n49486 ;
  assign y18568 = n49487 ;
  assign y18569 = ~1'b0 ;
  assign y18570 = n49489 ;
  assign y18571 = n49491 ;
  assign y18572 = ~1'b0 ;
  assign y18573 = ~1'b0 ;
  assign y18574 = ~n49492 ;
  assign y18575 = n49493 ;
  assign y18576 = n49495 ;
  assign y18577 = n49496 ;
  assign y18578 = n49498 ;
  assign y18579 = ~n49503 ;
  assign y18580 = ~1'b0 ;
  assign y18581 = n49504 ;
  assign y18582 = ~n49506 ;
  assign y18583 = n49513 ;
  assign y18584 = n49514 ;
  assign y18585 = ~n49515 ;
  assign y18586 = n49516 ;
  assign y18587 = n8635 ;
  assign y18588 = ~n49518 ;
  assign y18589 = ~n14601 ;
  assign y18590 = ~1'b0 ;
  assign y18591 = n49519 ;
  assign y18592 = ~1'b0 ;
  assign y18593 = n49522 ;
  assign y18594 = n49525 ;
  assign y18595 = n49526 ;
  assign y18596 = ~n49530 ;
  assign y18597 = n49531 ;
  assign y18598 = ~n49534 ;
  assign y18599 = ~1'b0 ;
  assign y18600 = ~n49537 ;
  assign y18601 = ~1'b0 ;
  assign y18602 = ~1'b0 ;
  assign y18603 = ~n49543 ;
  assign y18604 = ~n49544 ;
  assign y18605 = n49545 ;
  assign y18606 = n49551 ;
  assign y18607 = n49552 ;
  assign y18608 = ~1'b0 ;
  assign y18609 = ~1'b0 ;
  assign y18610 = ~n49557 ;
  assign y18611 = ~n49559 ;
  assign y18612 = 1'b0 ;
  assign y18613 = n49561 ;
  assign y18614 = n49562 ;
  assign y18615 = ~n49563 ;
  assign y18616 = n49566 ;
  assign y18617 = n49569 ;
  assign y18618 = ~n49570 ;
  assign y18619 = n49572 ;
  assign y18620 = ~1'b0 ;
  assign y18621 = n49578 ;
  assign y18622 = n49580 ;
  assign y18623 = n49583 ;
  assign y18624 = ~n49585 ;
  assign y18625 = n49586 ;
  assign y18626 = ~n49588 ;
  assign y18627 = n49589 ;
  assign y18628 = ~n49591 ;
  assign y18629 = ~n49599 ;
  assign y18630 = ~1'b0 ;
  assign y18631 = ~n49604 ;
  assign y18632 = ~n49610 ;
  assign y18633 = ~n49611 ;
  assign y18634 = ~n49616 ;
  assign y18635 = ~1'b0 ;
  assign y18636 = ~n49617 ;
  assign y18637 = n49620 ;
  assign y18638 = n49622 ;
  assign y18639 = ~n49624 ;
  assign y18640 = ~n49625 ;
  assign y18641 = n49627 ;
  assign y18642 = n49629 ;
  assign y18643 = ~n49630 ;
  assign y18644 = ~n49632 ;
  assign y18645 = n49637 ;
  assign y18646 = ~n49639 ;
  assign y18647 = ~n49640 ;
  assign y18648 = n49641 ;
  assign y18649 = n49642 ;
  assign y18650 = n49644 ;
  assign y18651 = ~1'b0 ;
  assign y18652 = n49647 ;
  assign y18653 = n49650 ;
  assign y18654 = ~1'b0 ;
  assign y18655 = ~1'b0 ;
  assign y18656 = ~n49654 ;
  assign y18657 = ~n4567 ;
  assign y18658 = n49655 ;
  assign y18659 = n49657 ;
  assign y18660 = n49659 ;
  assign y18661 = ~n49661 ;
  assign y18662 = 1'b0 ;
  assign y18663 = ~1'b0 ;
  assign y18664 = ~1'b0 ;
  assign y18665 = n49664 ;
  assign y18666 = ~n49668 ;
  assign y18667 = n49669 ;
  assign y18668 = ~n49670 ;
  assign y18669 = ~n49673 ;
  assign y18670 = n49675 ;
  assign y18671 = ~1'b0 ;
  assign y18672 = ~1'b0 ;
  assign y18673 = ~1'b0 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = ~n49677 ;
  assign y18676 = n49681 ;
  assign y18677 = ~n49683 ;
  assign y18678 = ~n6463 ;
  assign y18679 = n49684 ;
  assign y18680 = ~1'b0 ;
  assign y18681 = n49685 ;
  assign y18682 = ~1'b0 ;
  assign y18683 = ~1'b0 ;
  assign y18684 = n49691 ;
  assign y18685 = ~1'b0 ;
  assign y18686 = ~n49692 ;
  assign y18687 = ~n49695 ;
  assign y18688 = ~n49698 ;
  assign y18689 = n49700 ;
  assign y18690 = ~n49705 ;
  assign y18691 = ~n49709 ;
  assign y18692 = ~1'b0 ;
  assign y18693 = ~1'b0 ;
  assign y18694 = ~n49711 ;
  assign y18695 = ~n49716 ;
  assign y18696 = ~n49719 ;
  assign y18697 = n49720 ;
  assign y18698 = ~n49722 ;
  assign y18699 = n49727 ;
  assign y18700 = ~n15029 ;
  assign y18701 = ~n49728 ;
  assign y18702 = ~n49730 ;
  assign y18703 = n49736 ;
  assign y18704 = ~n49737 ;
  assign y18705 = ~1'b0 ;
  assign y18706 = ~n49738 ;
  assign y18707 = ~n49741 ;
  assign y18708 = ~n49742 ;
  assign y18709 = ~n49746 ;
  assign y18710 = ~n49750 ;
  assign y18711 = ~1'b0 ;
  assign y18712 = n49753 ;
  assign y18713 = ~n49754 ;
  assign y18714 = ~n6729 ;
  assign y18715 = n49763 ;
  assign y18716 = n49764 ;
  assign y18717 = ~n49768 ;
  assign y18718 = n49769 ;
  assign y18719 = n49770 ;
  assign y18720 = ~1'b0 ;
  assign y18721 = ~n49772 ;
  assign y18722 = ~n49775 ;
  assign y18723 = ~n49777 ;
  assign y18724 = 1'b0 ;
  assign y18725 = n49779 ;
  assign y18726 = n49780 ;
  assign y18727 = ~n49781 ;
  assign y18728 = ~n49789 ;
  assign y18729 = ~n49791 ;
  assign y18730 = n49793 ;
  assign y18731 = ~1'b0 ;
  assign y18732 = ~1'b0 ;
  assign y18733 = ~n49794 ;
  assign y18734 = ~1'b0 ;
  assign y18735 = n49795 ;
  assign y18736 = ~n49805 ;
  assign y18737 = n49806 ;
  assign y18738 = ~n49807 ;
  assign y18739 = n49812 ;
  assign y18740 = n49814 ;
  assign y18741 = ~1'b0 ;
  assign y18742 = ~n49816 ;
  assign y18743 = ~n49817 ;
  assign y18744 = ~1'b0 ;
  assign y18745 = ~1'b0 ;
  assign y18746 = ~n49819 ;
  assign y18747 = ~n49820 ;
  assign y18748 = n49823 ;
  assign y18749 = ~n49824 ;
  assign y18750 = n49825 ;
  assign y18751 = ~1'b0 ;
  assign y18752 = ~1'b0 ;
  assign y18753 = ~n49830 ;
  assign y18754 = ~n49832 ;
  assign y18755 = ~n49834 ;
  assign y18756 = ~n49837 ;
  assign y18757 = n5445 ;
  assign y18758 = n49838 ;
  assign y18759 = n49840 ;
  assign y18760 = n49844 ;
  assign y18761 = ~n49849 ;
  assign y18762 = n28538 ;
  assign y18763 = ~1'b0 ;
  assign y18764 = ~1'b0 ;
  assign y18765 = ~n18591 ;
  assign y18766 = n49850 ;
  assign y18767 = n49851 ;
  assign y18768 = n49856 ;
  assign y18769 = ~n49857 ;
  assign y18770 = ~n49860 ;
  assign y18771 = 1'b0 ;
  assign y18772 = ~n49862 ;
  assign y18773 = ~n49870 ;
  assign y18774 = ~n49872 ;
  assign y18775 = n49873 ;
  assign y18776 = n49874 ;
  assign y18777 = n49879 ;
  assign y18778 = n40797 ;
  assign y18779 = n49880 ;
  assign y18780 = ~n49881 ;
  assign y18781 = ~n49884 ;
  assign y18782 = ~1'b0 ;
  assign y18783 = ~1'b0 ;
  assign y18784 = ~1'b0 ;
  assign y18785 = n49887 ;
  assign y18786 = ~n49888 ;
  assign y18787 = n49892 ;
  assign y18788 = ~n49894 ;
  assign y18789 = ~n49895 ;
  assign y18790 = n49898 ;
  assign y18791 = n49899 ;
  assign y18792 = n49900 ;
  assign y18793 = ~1'b0 ;
  assign y18794 = ~n49902 ;
  assign y18795 = ~1'b0 ;
  assign y18796 = n49904 ;
  assign y18797 = n49905 ;
  assign y18798 = n49909 ;
  assign y18799 = ~n49910 ;
  assign y18800 = n49912 ;
  assign y18801 = ~n49916 ;
  assign y18802 = ~n49918 ;
  assign y18803 = ~1'b0 ;
  assign y18804 = ~n49920 ;
  assign y18805 = ~n49932 ;
  assign y18806 = ~n49935 ;
  assign y18807 = ~1'b0 ;
  assign y18808 = ~n49936 ;
  assign y18809 = n49938 ;
  assign y18810 = ~n49939 ;
  assign y18811 = ~n49940 ;
  assign y18812 = ~1'b0 ;
  assign y18813 = ~n49941 ;
  assign y18814 = ~n8396 ;
  assign y18815 = n49944 ;
  assign y18816 = ~1'b0 ;
  assign y18817 = n49946 ;
  assign y18818 = n49948 ;
  assign y18819 = n49952 ;
  assign y18820 = ~n49956 ;
  assign y18821 = n49957 ;
  assign y18822 = ~n49959 ;
  assign y18823 = ~1'b0 ;
  assign y18824 = ~1'b0 ;
  assign y18825 = ~n49962 ;
  assign y18826 = ~1'b0 ;
  assign y18827 = ~1'b0 ;
  assign y18828 = n49963 ;
  assign y18829 = ~n5188 ;
  assign y18830 = ~n49966 ;
  assign y18831 = ~n49967 ;
  assign y18832 = n49969 ;
  assign y18833 = ~n49971 ;
  assign y18834 = ~1'b0 ;
  assign y18835 = ~1'b0 ;
  assign y18836 = ~1'b0 ;
  assign y18837 = ~1'b0 ;
  assign y18838 = n24360 ;
  assign y18839 = n49974 ;
  assign y18840 = n49975 ;
  assign y18841 = n49976 ;
  assign y18842 = n49979 ;
  assign y18843 = ~n49981 ;
  assign y18844 = ~n49985 ;
  assign y18845 = n49986 ;
  assign y18846 = ~1'b0 ;
  assign y18847 = ~n49991 ;
  assign y18848 = ~n49992 ;
  assign y18849 = n49995 ;
  assign y18850 = ~n29272 ;
  assign y18851 = ~n49996 ;
  assign y18852 = ~n49998 ;
  assign y18853 = ~n50001 ;
  assign y18854 = ~x29 ;
  assign y18855 = n50002 ;
  assign y18856 = ~n50016 ;
  assign y18857 = ~n50017 ;
  assign y18858 = ~n50022 ;
  assign y18859 = ~n50026 ;
  assign y18860 = ~n50031 ;
  assign y18861 = n50033 ;
  assign y18862 = n50035 ;
  assign y18863 = n50037 ;
  assign y18864 = ~1'b0 ;
  assign y18865 = n50039 ;
  assign y18866 = ~n50041 ;
  assign y18867 = ~n50043 ;
  assign y18868 = n50045 ;
  assign y18869 = ~n50046 ;
  assign y18870 = ~n50047 ;
  assign y18871 = n50049 ;
  assign y18872 = ~n50051 ;
  assign y18873 = ~n50052 ;
  assign y18874 = ~1'b0 ;
  assign y18875 = ~n50053 ;
  assign y18876 = ~n50058 ;
  assign y18877 = n50060 ;
  assign y18878 = ~n50064 ;
  assign y18879 = ~n50065 ;
  assign y18880 = ~n50069 ;
  assign y18881 = n33637 ;
  assign y18882 = n50070 ;
  assign y18883 = ~1'b0 ;
  assign y18884 = ~1'b0 ;
  assign y18885 = ~n50075 ;
  assign y18886 = n50078 ;
  assign y18887 = n24883 ;
  assign y18888 = ~n50079 ;
  assign y18889 = ~1'b0 ;
  assign y18890 = ~n50080 ;
  assign y18891 = n50083 ;
  assign y18892 = n50085 ;
  assign y18893 = ~n50086 ;
  assign y18894 = n12561 ;
  assign y18895 = ~n50087 ;
  assign y18896 = n50090 ;
  assign y18897 = ~n50091 ;
  assign y18898 = n50093 ;
  assign y18899 = n50094 ;
  assign y18900 = ~1'b0 ;
  assign y18901 = ~1'b0 ;
  assign y18902 = ~n50096 ;
  assign y18903 = n50097 ;
  assign y18904 = ~n2430 ;
  assign y18905 = ~1'b0 ;
  assign y18906 = n50100 ;
  assign y18907 = n50105 ;
  assign y18908 = ~n50106 ;
  assign y18909 = n50107 ;
  assign y18910 = ~n50109 ;
  assign y18911 = n50111 ;
  assign y18912 = ~n50112 ;
  assign y18913 = n50114 ;
  assign y18914 = ~n50116 ;
  assign y18915 = ~1'b0 ;
  assign y18916 = n50123 ;
  assign y18917 = n50124 ;
  assign y18918 = ~n50129 ;
  assign y18919 = ~n50130 ;
  assign y18920 = ~n50131 ;
  assign y18921 = ~n50134 ;
  assign y18922 = ~n50136 ;
  assign y18923 = n50138 ;
  assign y18924 = n50140 ;
  assign y18925 = ~1'b0 ;
  assign y18926 = n50142 ;
  assign y18927 = n50144 ;
  assign y18928 = n50145 ;
  assign y18929 = ~n50148 ;
  assign y18930 = n50151 ;
  assign y18931 = ~n50153 ;
  assign y18932 = n50158 ;
  assign y18933 = n50160 ;
  assign y18934 = n50163 ;
  assign y18935 = n50167 ;
  assign y18936 = ~1'b0 ;
  assign y18937 = ~1'b0 ;
  assign y18938 = n50168 ;
  assign y18939 = ~n50171 ;
  assign y18940 = ~n50175 ;
  assign y18941 = ~n50181 ;
  assign y18942 = n50183 ;
  assign y18943 = n50184 ;
  assign y18944 = ~n50187 ;
  assign y18945 = ~n50189 ;
  assign y18946 = ~1'b0 ;
  assign y18947 = n50193 ;
  assign y18948 = n50196 ;
  assign y18949 = ~1'b0 ;
  assign y18950 = ~n50197 ;
  assign y18951 = n50198 ;
  assign y18952 = n50200 ;
  assign y18953 = ~1'b0 ;
  assign y18954 = n50201 ;
  assign y18955 = ~n50210 ;
  assign y18956 = ~n50212 ;
  assign y18957 = ~n50213 ;
  assign y18958 = n50215 ;
  assign y18959 = n50216 ;
  assign y18960 = n50221 ;
  assign y18961 = n50222 ;
  assign y18962 = ~n50226 ;
  assign y18963 = ~n50227 ;
  assign y18964 = n50229 ;
  assign y18965 = n50230 ;
  assign y18966 = ~n50231 ;
  assign y18967 = n50234 ;
  assign y18968 = ~n50237 ;
  assign y18969 = n50238 ;
  assign y18970 = n50247 ;
  assign y18971 = ~n50251 ;
  assign y18972 = ~n50253 ;
  assign y18973 = n50255 ;
  assign y18974 = ~n50257 ;
  assign y18975 = ~n50261 ;
  assign y18976 = ~n50263 ;
  assign y18977 = ~1'b0 ;
  assign y18978 = n50264 ;
  assign y18979 = ~n50269 ;
  assign y18980 = n50278 ;
  assign y18981 = ~n50286 ;
  assign y18982 = ~n50287 ;
  assign y18983 = ~n50288 ;
  assign y18984 = ~1'b0 ;
  assign y18985 = ~n50293 ;
  assign y18986 = n50297 ;
  assign y18987 = ~1'b0 ;
  assign y18988 = ~1'b0 ;
  assign y18989 = n50301 ;
  assign y18990 = ~n50302 ;
  assign y18991 = ~n50304 ;
  assign y18992 = n50310 ;
  assign y18993 = n50313 ;
  assign y18994 = n50314 ;
  assign y18995 = ~1'b0 ;
  assign y18996 = n50318 ;
  assign y18997 = n50319 ;
  assign y18998 = ~1'b0 ;
  assign y18999 = n50321 ;
  assign y19000 = ~n50325 ;
  assign y19001 = ~n50327 ;
  assign y19002 = ~n50329 ;
  assign y19003 = n50330 ;
  assign y19004 = ~1'b0 ;
  assign y19005 = ~n50331 ;
  assign y19006 = n50334 ;
  assign y19007 = n50336 ;
  assign y19008 = ~n50338 ;
  assign y19009 = ~1'b0 ;
  assign y19010 = n50342 ;
  assign y19011 = ~n50344 ;
  assign y19012 = ~n50347 ;
  assign y19013 = ~n50348 ;
  assign y19014 = n12237 ;
  assign y19015 = n50350 ;
  assign y19016 = ~1'b0 ;
  assign y19017 = n24570 ;
  assign y19018 = n50355 ;
  assign y19019 = ~n50359 ;
  assign y19020 = n50360 ;
  assign y19021 = ~n50361 ;
  assign y19022 = ~n50364 ;
  assign y19023 = ~n50368 ;
  assign y19024 = n50370 ;
  assign y19025 = ~n50372 ;
  assign y19026 = n50374 ;
  assign y19027 = ~1'b0 ;
  assign y19028 = n50376 ;
  assign y19029 = ~n50378 ;
  assign y19030 = ~n50379 ;
  assign y19031 = ~n50380 ;
  assign y19032 = n50383 ;
  assign y19033 = n50384 ;
  assign y19034 = n50385 ;
  assign y19035 = ~n50386 ;
  assign y19036 = n50388 ;
  assign y19037 = ~n50391 ;
  assign y19038 = ~n50392 ;
  assign y19039 = ~n50397 ;
  assign y19040 = ~1'b0 ;
  assign y19041 = ~n50399 ;
  assign y19042 = ~n50405 ;
  assign y19043 = n50406 ;
  assign y19044 = n50407 ;
  assign y19045 = n50408 ;
  assign y19046 = ~n50410 ;
  assign y19047 = ~1'b0 ;
  assign y19048 = n50411 ;
  assign y19049 = ~n50413 ;
  assign y19050 = n50418 ;
  assign y19051 = ~n50421 ;
  assign y19052 = n50422 ;
  assign y19053 = n50425 ;
  assign y19054 = ~n50426 ;
  assign y19055 = n50427 ;
  assign y19056 = ~n50433 ;
  assign y19057 = n50434 ;
  assign y19058 = ~1'b0 ;
  assign y19059 = ~1'b0 ;
  assign y19060 = ~n50438 ;
  assign y19061 = n50439 ;
  assign y19062 = ~n50441 ;
  assign y19063 = n50442 ;
  assign y19064 = n50444 ;
  assign y19065 = ~1'b0 ;
  assign y19066 = n50447 ;
  assign y19067 = ~n50449 ;
  assign y19068 = ~1'b0 ;
  assign y19069 = n50456 ;
  assign y19070 = ~n50457 ;
  assign y19071 = n50458 ;
  assign y19072 = ~n50459 ;
  assign y19073 = ~n50462 ;
  assign y19074 = ~n50463 ;
  assign y19075 = n50464 ;
  assign y19076 = ~n50466 ;
  assign y19077 = ~n50469 ;
  assign y19078 = n50473 ;
  assign y19079 = n50474 ;
  assign y19080 = ~1'b0 ;
  assign y19081 = ~n50477 ;
  assign y19082 = ~n50478 ;
  assign y19083 = n50479 ;
  assign y19084 = ~n50480 ;
  assign y19085 = ~n48369 ;
  assign y19086 = ~n50489 ;
  assign y19087 = ~1'b0 ;
  assign y19088 = ~1'b0 ;
  assign y19089 = ~n50491 ;
  assign y19090 = n50493 ;
  assign y19091 = n50497 ;
  assign y19092 = ~1'b0 ;
  assign y19093 = ~n50500 ;
  assign y19094 = ~n50501 ;
  assign y19095 = n50503 ;
  assign y19096 = n50504 ;
  assign y19097 = ~n50506 ;
  assign y19098 = ~n50509 ;
  assign y19099 = ~n50513 ;
  assign y19100 = ~1'b0 ;
  assign y19101 = ~n50515 ;
  assign y19102 = n50518 ;
  assign y19103 = n50519 ;
  assign y19104 = n50523 ;
  assign y19105 = ~n50524 ;
  assign y19106 = ~n50528 ;
  assign y19107 = ~n50529 ;
  assign y19108 = ~n50532 ;
  assign y19109 = n50534 ;
  assign y19110 = ~1'b0 ;
  assign y19111 = ~1'b0 ;
  assign y19112 = n50537 ;
  assign y19113 = ~n50542 ;
  assign y19114 = n50543 ;
  assign y19115 = ~n50544 ;
  assign y19116 = n50545 ;
  assign y19117 = ~1'b0 ;
  assign y19118 = ~n50548 ;
  assign y19119 = n50553 ;
  assign y19120 = n50558 ;
  assign y19121 = ~1'b0 ;
  assign y19122 = n50562 ;
  assign y19123 = ~n50566 ;
  assign y19124 = ~n50568 ;
  assign y19125 = ~n50570 ;
  assign y19126 = n50572 ;
  assign y19127 = ~n50573 ;
  assign y19128 = ~1'b0 ;
  assign y19129 = ~n50575 ;
  assign y19130 = ~n50576 ;
  assign y19131 = n50578 ;
  assign y19132 = n50579 ;
  assign y19133 = ~n50580 ;
  assign y19134 = n50581 ;
  assign y19135 = n50584 ;
  assign y19136 = ~n50585 ;
  assign y19137 = ~n50587 ;
  assign y19138 = ~1'b0 ;
  assign y19139 = ~n50589 ;
  assign y19140 = ~1'b0 ;
  assign y19141 = ~1'b0 ;
  assign y19142 = ~1'b0 ;
  assign y19143 = n50591 ;
  assign y19144 = ~n50598 ;
  assign y19145 = ~n50599 ;
  assign y19146 = ~n50600 ;
  assign y19147 = n50601 ;
  assign y19148 = n50606 ;
  assign y19149 = ~n50607 ;
  assign y19150 = ~n50614 ;
  assign y19151 = n50617 ;
  assign y19152 = n50620 ;
  assign y19153 = ~n50623 ;
  assign y19154 = n50626 ;
  assign y19155 = n50630 ;
  assign y19156 = n50635 ;
  assign y19157 = n50636 ;
  assign y19158 = ~n50639 ;
  assign y19159 = ~n50643 ;
  assign y19160 = ~n50645 ;
  assign y19161 = n50647 ;
  assign y19162 = ~n50649 ;
  assign y19163 = ~1'b0 ;
  assign y19164 = ~n50652 ;
  assign y19165 = ~n50656 ;
  assign y19166 = n50659 ;
  assign y19167 = ~n50660 ;
  assign y19168 = n50663 ;
  assign y19169 = ~1'b0 ;
  assign y19170 = ~n50670 ;
  assign y19171 = n50677 ;
  assign y19172 = n50681 ;
  assign y19173 = n50682 ;
  assign y19174 = n50683 ;
  assign y19175 = n50684 ;
  assign y19176 = n50689 ;
  assign y19177 = n50695 ;
  assign y19178 = n50699 ;
  assign y19179 = ~1'b0 ;
  assign y19180 = n50702 ;
  assign y19181 = ~n50705 ;
  assign y19182 = ~n50706 ;
  assign y19183 = ~n50709 ;
  assign y19184 = n50713 ;
  assign y19185 = n50714 ;
  assign y19186 = n50717 ;
  assign y19187 = ~n50721 ;
  assign y19188 = n3613 ;
  assign y19189 = ~n50722 ;
  assign y19190 = ~1'b0 ;
  assign y19191 = ~n50727 ;
  assign y19192 = ~1'b0 ;
  assign y19193 = ~n50731 ;
  assign y19194 = ~1'b0 ;
  assign y19195 = ~n50734 ;
  assign y19196 = ~n50735 ;
  assign y19197 = n50736 ;
  assign y19198 = ~n50737 ;
  assign y19199 = ~n50738 ;
  assign y19200 = ~1'b0 ;
  assign y19201 = ~n50740 ;
  assign y19202 = ~n50742 ;
  assign y19203 = ~n50743 ;
  assign y19204 = ~n50747 ;
  assign y19205 = n50748 ;
  assign y19206 = ~n50750 ;
  assign y19207 = n50753 ;
  assign y19208 = ~n50754 ;
  assign y19209 = n50755 ;
  assign y19210 = ~n50756 ;
  assign y19211 = n50758 ;
  assign y19212 = n50764 ;
  assign y19213 = n50766 ;
  assign y19214 = n50767 ;
  assign y19215 = n50768 ;
  assign y19216 = n50770 ;
  assign y19217 = ~n50773 ;
  assign y19218 = ~n50774 ;
  assign y19219 = ~1'b0 ;
  assign y19220 = ~n50776 ;
  assign y19221 = ~n50778 ;
  assign y19222 = ~1'b0 ;
  assign y19223 = ~n12164 ;
  assign y19224 = ~1'b0 ;
  assign y19225 = n50779 ;
  assign y19226 = ~n50780 ;
  assign y19227 = n50781 ;
  assign y19228 = n50782 ;
  assign y19229 = ~1'b0 ;
  assign y19230 = n50786 ;
  assign y19231 = ~n50787 ;
  assign y19232 = n50790 ;
  assign y19233 = ~1'b0 ;
  assign y19234 = ~1'b0 ;
  assign y19235 = ~n50792 ;
  assign y19236 = ~n50793 ;
  assign y19237 = n50794 ;
  assign y19238 = n50796 ;
  assign y19239 = n50797 ;
  assign y19240 = n50798 ;
  assign y19241 = n50802 ;
  assign y19242 = n50805 ;
  assign y19243 = ~1'b0 ;
  assign y19244 = n50807 ;
  assign y19245 = ~n50809 ;
  assign y19246 = ~n50810 ;
  assign y19247 = n50812 ;
  assign y19248 = ~n50819 ;
  assign y19249 = n50823 ;
  assign y19250 = ~n50826 ;
  assign y19251 = ~n46897 ;
  assign y19252 = ~n50830 ;
  assign y19253 = n50833 ;
  assign y19254 = ~1'b0 ;
  assign y19255 = n50839 ;
  assign y19256 = ~n50840 ;
  assign y19257 = ~n50846 ;
  assign y19258 = n50851 ;
  assign y19259 = n50856 ;
  assign y19260 = ~n50858 ;
  assign y19261 = ~1'b0 ;
  assign y19262 = n50859 ;
  assign y19263 = n50860 ;
  assign y19264 = n50863 ;
  assign y19265 = ~n50867 ;
  assign y19266 = ~n50869 ;
  assign y19267 = n50872 ;
  assign y19268 = n50874 ;
  assign y19269 = ~n50875 ;
  assign y19270 = n50876 ;
  assign y19271 = n50879 ;
  assign y19272 = n50881 ;
  assign y19273 = n50888 ;
  assign y19274 = ~1'b0 ;
  assign y19275 = ~n50889 ;
  assign y19276 = ~n50890 ;
  assign y19277 = n50893 ;
  assign y19278 = n50894 ;
  assign y19279 = ~n50896 ;
  assign y19280 = n50900 ;
  assign y19281 = n50903 ;
  assign y19282 = ~1'b0 ;
  assign y19283 = n50907 ;
  assign y19284 = n50909 ;
  assign y19285 = ~n50912 ;
  assign y19286 = ~1'b0 ;
  assign y19287 = ~1'b0 ;
  assign y19288 = n50916 ;
  assign y19289 = n50919 ;
  assign y19290 = ~n50922 ;
  assign y19291 = n50926 ;
  assign y19292 = n50931 ;
  assign y19293 = ~n50932 ;
  assign y19294 = ~1'b0 ;
  assign y19295 = ~n50934 ;
  assign y19296 = ~n50936 ;
  assign y19297 = ~n50938 ;
  assign y19298 = ~n50941 ;
  assign y19299 = n50942 ;
  assign y19300 = ~n50943 ;
  assign y19301 = ~n50945 ;
  assign y19302 = ~n50946 ;
  assign y19303 = n50947 ;
  assign y19304 = ~1'b0 ;
  assign y19305 = n50949 ;
  assign y19306 = n50950 ;
  assign y19307 = ~1'b0 ;
  assign y19308 = ~n50954 ;
  assign y19309 = n50955 ;
  assign y19310 = ~n50961 ;
  assign y19311 = ~n50964 ;
  assign y19312 = ~n50967 ;
  assign y19313 = n50969 ;
  assign y19314 = n50970 ;
  assign y19315 = ~n50974 ;
  assign y19316 = ~n50975 ;
  assign y19317 = n50976 ;
  assign y19318 = ~n50980 ;
  assign y19319 = ~1'b0 ;
  assign y19320 = ~n50981 ;
  assign y19321 = ~n50984 ;
  assign y19322 = ~n50986 ;
  assign y19323 = n50987 ;
  assign y19324 = 1'b0 ;
  assign y19325 = ~n50988 ;
  assign y19326 = n50989 ;
  assign y19327 = ~1'b0 ;
  assign y19328 = n50992 ;
  assign y19329 = n50994 ;
  assign y19330 = ~1'b0 ;
  assign y19331 = ~n50995 ;
  assign y19332 = ~n50996 ;
  assign y19333 = ~n51004 ;
  assign y19334 = ~n51012 ;
  assign y19335 = ~n51014 ;
  assign y19336 = ~n51017 ;
  assign y19337 = n51019 ;
  assign y19338 = n51021 ;
  assign y19339 = n51024 ;
  assign y19340 = n51030 ;
  assign y19341 = ~n51032 ;
  assign y19342 = ~n51033 ;
  assign y19343 = n51034 ;
  assign y19344 = ~n51038 ;
  assign y19345 = n51041 ;
  assign y19346 = ~n51049 ;
  assign y19347 = n51052 ;
  assign y19348 = n51053 ;
  assign y19349 = ~1'b0 ;
  assign y19350 = ~n51055 ;
  assign y19351 = ~n51061 ;
  assign y19352 = ~1'b0 ;
  assign y19353 = n51062 ;
  assign y19354 = ~n51063 ;
  assign y19355 = n51064 ;
  assign y19356 = ~n51065 ;
  assign y19357 = ~n51067 ;
  assign y19358 = ~1'b0 ;
  assign y19359 = n51069 ;
  assign y19360 = n51070 ;
  assign y19361 = ~1'b0 ;
  assign y19362 = n51073 ;
  assign y19363 = ~n51074 ;
  assign y19364 = n51077 ;
  assign y19365 = ~n51078 ;
  assign y19366 = ~n51079 ;
  assign y19367 = n51081 ;
  assign y19368 = n27400 ;
  assign y19369 = ~1'b0 ;
  assign y19370 = n51082 ;
  assign y19371 = n51085 ;
  assign y19372 = n51091 ;
  assign y19373 = ~n51093 ;
  assign y19374 = n12250 ;
  assign y19375 = n51099 ;
  assign y19376 = n51102 ;
  assign y19377 = ~n51104 ;
  assign y19378 = n51107 ;
  assign y19379 = ~n51109 ;
  assign y19380 = ~n51116 ;
  assign y19381 = n51117 ;
  assign y19382 = n51121 ;
  assign y19383 = n51127 ;
  assign y19384 = ~n51132 ;
  assign y19385 = ~n51137 ;
  assign y19386 = ~1'b0 ;
  assign y19387 = ~n51139 ;
  assign y19388 = ~1'b0 ;
  assign y19389 = ~1'b0 ;
  assign y19390 = ~n51141 ;
  assign y19391 = ~n51142 ;
  assign y19392 = n51144 ;
  assign y19393 = ~n51145 ;
  assign y19394 = ~n51148 ;
  assign y19395 = n51150 ;
  assign y19396 = ~n51152 ;
  assign y19397 = ~1'b0 ;
  assign y19398 = ~n51160 ;
  assign y19399 = ~1'b0 ;
  assign y19400 = n51167 ;
  assign y19401 = n51168 ;
  assign y19402 = ~n51170 ;
  assign y19403 = ~n51174 ;
  assign y19404 = ~n51178 ;
  assign y19405 = ~n51179 ;
  assign y19406 = n51184 ;
  assign y19407 = ~1'b0 ;
  assign y19408 = n51186 ;
  assign y19409 = n51187 ;
  assign y19410 = n51188 ;
  assign y19411 = ~1'b0 ;
  assign y19412 = n51190 ;
  assign y19413 = ~n51191 ;
  assign y19414 = ~n51195 ;
  assign y19415 = ~n51197 ;
  assign y19416 = ~n37648 ;
  assign y19417 = ~n51201 ;
  assign y19418 = n51206 ;
  assign y19419 = ~n51208 ;
  assign y19420 = n51210 ;
  assign y19421 = ~1'b0 ;
  assign y19422 = n51211 ;
  assign y19423 = ~n51212 ;
  assign y19424 = n51214 ;
  assign y19425 = n51218 ;
  assign y19426 = ~n51219 ;
  assign y19427 = n51220 ;
  assign y19428 = n51222 ;
  assign y19429 = ~n51227 ;
  assign y19430 = n51229 ;
  assign y19431 = ~n51234 ;
  assign y19432 = ~1'b0 ;
  assign y19433 = n51235 ;
  assign y19434 = ~n51239 ;
  assign y19435 = ~n51240 ;
  assign y19436 = ~n51241 ;
  assign y19437 = ~n51244 ;
  assign y19438 = ~n51246 ;
  assign y19439 = n51248 ;
  assign y19440 = ~n51250 ;
  assign y19441 = ~1'b0 ;
  assign y19442 = ~n51251 ;
  assign y19443 = ~1'b0 ;
  assign y19444 = ~n51253 ;
  assign y19445 = n51254 ;
  assign y19446 = ~n51257 ;
  assign y19447 = n51261 ;
  assign y19448 = n51264 ;
  assign y19449 = ~n51266 ;
  assign y19450 = ~n51272 ;
  assign y19451 = ~1'b0 ;
  assign y19452 = ~n51273 ;
  assign y19453 = ~n51274 ;
  assign y19454 = n51275 ;
  assign y19455 = ~n51276 ;
  assign y19456 = ~n51278 ;
  assign y19457 = ~n51282 ;
  assign y19458 = ~n51284 ;
  assign y19459 = n27199 ;
  assign y19460 = ~1'b0 ;
  assign y19461 = n51288 ;
  assign y19462 = n51290 ;
  assign y19463 = ~n51291 ;
  assign y19464 = ~1'b0 ;
  assign y19465 = ~n51294 ;
  assign y19466 = 1'b0 ;
  assign y19467 = ~n51295 ;
  assign y19468 = ~n51299 ;
  assign y19469 = ~n51300 ;
  assign y19470 = ~n51301 ;
  assign y19471 = ~n51303 ;
  assign y19472 = 1'b0 ;
  assign y19473 = ~n51304 ;
  assign y19474 = n51308 ;
  assign y19475 = ~1'b0 ;
  assign y19476 = ~1'b0 ;
  assign y19477 = n51309 ;
  assign y19478 = ~1'b0 ;
  assign y19479 = ~n51310 ;
  assign y19480 = n51311 ;
  assign y19481 = n33083 ;
  assign y19482 = ~1'b0 ;
  assign y19483 = ~1'b0 ;
  assign y19484 = n51318 ;
  assign y19485 = n51329 ;
  assign y19486 = ~n51334 ;
  assign y19487 = ~n51336 ;
  assign y19488 = n51342 ;
  assign y19489 = n51344 ;
  assign y19490 = ~n51345 ;
  assign y19491 = ~n51346 ;
  assign y19492 = n51348 ;
  assign y19493 = n51352 ;
  assign y19494 = n51354 ;
  assign y19495 = ~1'b0 ;
  assign y19496 = ~n51356 ;
  assign y19497 = ~1'b0 ;
  assign y19498 = n25831 ;
  assign y19499 = ~n51362 ;
  assign y19500 = ~n51363 ;
  assign y19501 = ~1'b0 ;
  assign y19502 = n51364 ;
  assign y19503 = n51365 ;
  assign y19504 = ~n51368 ;
  assign y19505 = ~1'b0 ;
  assign y19506 = ~n51370 ;
  assign y19507 = ~1'b0 ;
  assign y19508 = ~1'b0 ;
  assign y19509 = ~n23957 ;
  assign y19510 = n51373 ;
  assign y19511 = n51374 ;
  assign y19512 = n51376 ;
  assign y19513 = ~n51380 ;
  assign y19514 = ~n51382 ;
  assign y19515 = n51386 ;
  assign y19516 = ~1'b0 ;
  assign y19517 = n51388 ;
  assign y19518 = ~n51391 ;
  assign y19519 = ~n51396 ;
  assign y19520 = n51402 ;
  assign y19521 = ~n51403 ;
  assign y19522 = ~n51404 ;
  assign y19523 = n51406 ;
  assign y19524 = ~n51409 ;
  assign y19525 = ~1'b0 ;
  assign y19526 = ~n51410 ;
  assign y19527 = n51413 ;
  assign y19528 = ~1'b0 ;
  assign y19529 = ~1'b0 ;
  assign y19530 = n51414 ;
  assign y19531 = n51416 ;
  assign y19532 = n51418 ;
  assign y19533 = n20881 ;
  assign y19534 = n51421 ;
  assign y19535 = ~1'b0 ;
  assign y19536 = ~1'b0 ;
  assign y19537 = ~1'b0 ;
  assign y19538 = ~1'b0 ;
  assign y19539 = ~1'b0 ;
  assign y19540 = ~n51427 ;
  assign y19541 = n51429 ;
  assign y19542 = n51430 ;
  assign y19543 = n51431 ;
  assign y19544 = n51433 ;
  assign y19545 = n51435 ;
  assign y19546 = n51438 ;
  assign y19547 = n51440 ;
  assign y19548 = ~1'b0 ;
  assign y19549 = ~1'b0 ;
  assign y19550 = n51442 ;
  assign y19551 = ~1'b0 ;
  assign y19552 = ~1'b0 ;
  assign y19553 = ~n51448 ;
  assign y19554 = ~n51450 ;
  assign y19555 = ~n51452 ;
  assign y19556 = n51456 ;
  assign y19557 = ~n51471 ;
  assign y19558 = n51472 ;
  assign y19559 = ~1'b0 ;
  assign y19560 = n51473 ;
  assign y19561 = ~n51474 ;
  assign y19562 = ~1'b0 ;
  assign y19563 = n51476 ;
  assign y19564 = ~n51479 ;
  assign y19565 = n51480 ;
  assign y19566 = ~n51481 ;
  assign y19567 = ~n51489 ;
  assign y19568 = ~n51491 ;
  assign y19569 = ~n51492 ;
  assign y19570 = n51493 ;
  assign y19571 = n51495 ;
  assign y19572 = ~n51498 ;
  assign y19573 = n51502 ;
  assign y19574 = n51503 ;
  assign y19575 = n51504 ;
  assign y19576 = n51505 ;
  assign y19577 = ~n51508 ;
  assign y19578 = ~1'b0 ;
  assign y19579 = ~n51511 ;
  assign y19580 = ~1'b0 ;
  assign y19581 = n51513 ;
  assign y19582 = n51515 ;
  assign y19583 = n51516 ;
  assign y19584 = n51517 ;
  assign y19585 = n51518 ;
  assign y19586 = n51521 ;
  assign y19587 = ~n51524 ;
  assign y19588 = ~n51528 ;
  assign y19589 = n51529 ;
  assign y19590 = ~n51531 ;
  assign y19591 = ~1'b0 ;
  assign y19592 = n51533 ;
  assign y19593 = ~n51537 ;
  assign y19594 = n51539 ;
  assign y19595 = ~n51541 ;
  assign y19596 = ~n51544 ;
  assign y19597 = ~n51547 ;
  assign y19598 = ~n51550 ;
  assign y19599 = n51554 ;
  assign y19600 = ~1'b0 ;
  assign y19601 = n51557 ;
  assign y19602 = ~1'b0 ;
  assign y19603 = ~n51559 ;
  assign y19604 = ~n51565 ;
  assign y19605 = ~n51574 ;
  assign y19606 = n51576 ;
  assign y19607 = ~n51578 ;
  assign y19608 = n51579 ;
  assign y19609 = ~1'b0 ;
  assign y19610 = n51580 ;
  assign y19611 = n51582 ;
  assign y19612 = n51584 ;
  assign y19613 = n51590 ;
  assign y19614 = n51591 ;
  assign y19615 = ~n51595 ;
  assign y19616 = ~n51596 ;
  assign y19617 = ~n51597 ;
  assign y19618 = ~n51598 ;
  assign y19619 = ~n51600 ;
  assign y19620 = n51603 ;
  assign y19621 = ~1'b0 ;
  assign y19622 = n51605 ;
  assign y19623 = ~n51607 ;
  assign y19624 = n51612 ;
  assign y19625 = ~n51614 ;
  assign y19626 = ~n51618 ;
  assign y19627 = ~n51619 ;
  assign y19628 = n51621 ;
  assign y19629 = ~n51624 ;
  assign y19630 = ~1'b0 ;
  assign y19631 = ~n51628 ;
  assign y19632 = ~n51631 ;
  assign y19633 = n51632 ;
  assign y19634 = n51633 ;
  assign y19635 = n51634 ;
  assign y19636 = ~n51635 ;
  assign y19637 = n51636 ;
  assign y19638 = n51637 ;
  assign y19639 = n51638 ;
  assign y19640 = ~1'b0 ;
  assign y19641 = ~n51642 ;
  assign y19642 = ~1'b0 ;
  assign y19643 = ~1'b0 ;
  assign y19644 = ~1'b0 ;
  assign y19645 = n51647 ;
  assign y19646 = ~n51648 ;
  assign y19647 = ~n51650 ;
  assign y19648 = n51651 ;
  assign y19649 = n51652 ;
  assign y19650 = ~n51654 ;
  assign y19651 = ~1'b0 ;
  assign y19652 = n51656 ;
  assign y19653 = ~n51658 ;
  assign y19654 = ~n51660 ;
  assign y19655 = ~1'b0 ;
  assign y19656 = n51666 ;
  assign y19657 = n51670 ;
  assign y19658 = ~n51671 ;
  assign y19659 = ~n4912 ;
  assign y19660 = ~n51672 ;
  assign y19661 = ~1'b0 ;
  assign y19662 = n51678 ;
  assign y19663 = ~1'b0 ;
  assign y19664 = ~n51679 ;
  assign y19665 = n51684 ;
  assign y19666 = n51685 ;
  assign y19667 = n51686 ;
  assign y19668 = ~n51688 ;
  assign y19669 = n51689 ;
  assign y19670 = ~n51690 ;
  assign y19671 = ~n51692 ;
  assign y19672 = ~1'b0 ;
  assign y19673 = ~n51696 ;
  assign y19674 = ~1'b0 ;
  assign y19675 = ~1'b0 ;
  assign y19676 = ~1'b0 ;
  assign y19677 = n51698 ;
  assign y19678 = n51699 ;
  assign y19679 = ~n51701 ;
  assign y19680 = n51702 ;
  assign y19681 = n51704 ;
  assign y19682 = n20533 ;
  assign y19683 = ~1'b0 ;
  assign y19684 = ~1'b0 ;
  assign y19685 = ~n51705 ;
  assign y19686 = ~n51707 ;
  assign y19687 = n51710 ;
  assign y19688 = ~1'b0 ;
  assign y19689 = n51713 ;
  assign y19690 = ~n51714 ;
  assign y19691 = ~n51715 ;
  assign y19692 = n28810 ;
  assign y19693 = ~n51719 ;
  assign y19694 = ~n51721 ;
  assign y19695 = n51723 ;
  assign y19696 = n51725 ;
  assign y19697 = n51729 ;
  assign y19698 = n51734 ;
  assign y19699 = ~n51736 ;
  assign y19700 = n51740 ;
  assign y19701 = ~n51741 ;
  assign y19702 = ~n51746 ;
  assign y19703 = n51753 ;
  assign y19704 = ~n51756 ;
  assign y19705 = n51758 ;
  assign y19706 = ~1'b0 ;
  assign y19707 = n51762 ;
  assign y19708 = n51764 ;
  assign y19709 = ~1'b0 ;
  assign y19710 = ~n51767 ;
  assign y19711 = n51768 ;
  assign y19712 = ~n51771 ;
  assign y19713 = ~n51773 ;
  assign y19714 = n38946 ;
  assign y19715 = n51774 ;
  assign y19716 = ~n51780 ;
  assign y19717 = ~n51789 ;
  assign y19718 = ~1'b0 ;
  assign y19719 = n51791 ;
  assign y19720 = n51793 ;
  assign y19721 = ~n51795 ;
  assign y19722 = ~n51798 ;
  assign y19723 = n51799 ;
  assign y19724 = ~n51802 ;
  assign y19725 = ~n51805 ;
  assign y19726 = n51807 ;
  assign y19727 = n51809 ;
  assign y19728 = ~n51811 ;
  assign y19729 = ~n51813 ;
  assign y19730 = ~n51817 ;
  assign y19731 = n8387 ;
  assign y19732 = ~n51819 ;
  assign y19733 = ~n51824 ;
  assign y19734 = n51827 ;
  assign y19735 = n51829 ;
  assign y19736 = n51832 ;
  assign y19737 = ~n51833 ;
  assign y19738 = ~1'b0 ;
  assign y19739 = ~1'b0 ;
  assign y19740 = n51834 ;
  assign y19741 = n51836 ;
  assign y19742 = ~n51838 ;
  assign y19743 = ~1'b0 ;
  assign y19744 = ~n21683 ;
  assign y19745 = n51839 ;
  assign y19746 = ~n51841 ;
  assign y19747 = ~n51843 ;
  assign y19748 = ~n51845 ;
  assign y19749 = ~1'b0 ;
  assign y19750 = n51846 ;
  assign y19751 = ~n51848 ;
  assign y19752 = n51850 ;
  assign y19753 = ~n51853 ;
  assign y19754 = ~n51855 ;
  assign y19755 = n51856 ;
  assign y19756 = ~n51859 ;
  assign y19757 = ~n51863 ;
  assign y19758 = n51866 ;
  assign y19759 = ~n51872 ;
  assign y19760 = ~n51875 ;
  assign y19761 = ~n51878 ;
  assign y19762 = ~n51882 ;
  assign y19763 = n51886 ;
  assign y19764 = ~n51890 ;
  assign y19765 = ~1'b0 ;
  assign y19766 = n51892 ;
  assign y19767 = n51895 ;
  assign y19768 = n51897 ;
  assign y19769 = ~n51899 ;
  assign y19770 = n51900 ;
  assign y19771 = ~1'b0 ;
  assign y19772 = n47739 ;
  assign y19773 = n51901 ;
  assign y19774 = ~n51905 ;
  assign y19775 = ~1'b0 ;
  assign y19776 = ~n51908 ;
  assign y19777 = n51910 ;
  assign y19778 = ~n51913 ;
  assign y19779 = n51914 ;
  assign y19780 = ~n51916 ;
  assign y19781 = ~n51918 ;
  assign y19782 = n51921 ;
  assign y19783 = ~1'b0 ;
  assign y19784 = ~1'b0 ;
  assign y19785 = n51924 ;
  assign y19786 = ~n51926 ;
  assign y19787 = n51929 ;
  assign y19788 = ~n51931 ;
  assign y19789 = ~n51932 ;
  assign y19790 = n51933 ;
  assign y19791 = ~n51934 ;
  assign y19792 = n51935 ;
  assign y19793 = n51937 ;
  assign y19794 = ~n51941 ;
  assign y19795 = ~1'b0 ;
  assign y19796 = ~n51945 ;
  assign y19797 = ~n51947 ;
  assign y19798 = ~n51950 ;
  assign y19799 = n51951 ;
  assign y19800 = ~n51957 ;
  assign y19801 = ~n51958 ;
  assign y19802 = ~n51959 ;
  assign y19803 = ~n51960 ;
  assign y19804 = n51961 ;
  assign y19805 = ~1'b0 ;
  assign y19806 = ~1'b0 ;
  assign y19807 = n51964 ;
  assign y19808 = ~1'b0 ;
  assign y19809 = ~n51966 ;
  assign y19810 = ~n51968 ;
  assign y19811 = n51972 ;
  assign y19812 = n51973 ;
  assign y19813 = n51974 ;
  assign y19814 = n18121 ;
  assign y19815 = ~n51976 ;
  assign y19816 = ~n51980 ;
  assign y19817 = ~n51982 ;
  assign y19818 = ~n51984 ;
  assign y19819 = n51987 ;
  assign y19820 = 1'b0 ;
  assign y19821 = ~n51988 ;
  assign y19822 = n51991 ;
  assign y19823 = n51993 ;
  assign y19824 = n51994 ;
  assign y19825 = n51997 ;
  assign y19826 = n52000 ;
  assign y19827 = ~1'b0 ;
  assign y19828 = n52002 ;
  assign y19829 = n52004 ;
  assign y19830 = ~1'b0 ;
  assign y19831 = ~n52007 ;
  assign y19832 = n52010 ;
  assign y19833 = ~n52011 ;
  assign y19834 = ~n52014 ;
  assign y19835 = ~n52017 ;
  assign y19836 = n52018 ;
  assign y19837 = n52020 ;
  assign y19838 = 1'b0 ;
  assign y19839 = ~n52022 ;
  assign y19840 = ~n52024 ;
  assign y19841 = ~n52025 ;
  assign y19842 = ~n52028 ;
  assign y19843 = n52029 ;
  assign y19844 = ~n52034 ;
  assign y19845 = ~n52035 ;
  assign y19846 = n52041 ;
  assign y19847 = n52045 ;
  assign y19848 = ~n52046 ;
  assign y19849 = ~1'b0 ;
  assign y19850 = ~n52049 ;
  assign y19851 = n52050 ;
  assign y19852 = ~n52051 ;
  assign y19853 = ~n52052 ;
  assign y19854 = n52055 ;
  assign y19855 = n52056 ;
  assign y19856 = ~n52058 ;
  assign y19857 = ~n52059 ;
  assign y19858 = ~n52060 ;
  assign y19859 = ~1'b0 ;
  assign y19860 = ~n52062 ;
  assign y19861 = ~n52064 ;
  assign y19862 = ~n52066 ;
  assign y19863 = ~1'b0 ;
  assign y19864 = ~n52072 ;
  assign y19865 = ~n52073 ;
  assign y19866 = n52074 ;
  assign y19867 = ~n52075 ;
  assign y19868 = n52077 ;
  assign y19869 = ~n52078 ;
  assign y19870 = ~n32462 ;
  assign y19871 = ~1'b0 ;
  assign y19872 = ~1'b0 ;
  assign y19873 = ~n52079 ;
  assign y19874 = ~1'b0 ;
  assign y19875 = ~n52089 ;
  assign y19876 = ~n52091 ;
  assign y19877 = n52092 ;
  assign y19878 = ~n52095 ;
  assign y19879 = ~n52103 ;
  assign y19880 = n52110 ;
  assign y19881 = ~n52112 ;
  assign y19882 = n52114 ;
  assign y19883 = ~n52116 ;
  assign y19884 = n52121 ;
  assign y19885 = n52123 ;
  assign y19886 = n52126 ;
  assign y19887 = ~n52127 ;
  assign y19888 = ~n52131 ;
  assign y19889 = n52133 ;
  assign y19890 = n52134 ;
  assign y19891 = n52136 ;
  assign y19892 = ~1'b0 ;
  assign y19893 = ~n6458 ;
  assign y19894 = ~n52139 ;
  assign y19895 = ~n52144 ;
  assign y19896 = ~1'b0 ;
  assign y19897 = ~n12092 ;
  assign y19898 = n52145 ;
  assign y19899 = ~n52147 ;
  assign y19900 = ~n52154 ;
  assign y19901 = ~n52155 ;
  assign y19902 = ~n52160 ;
  assign y19903 = ~n52161 ;
  assign y19904 = ~n52164 ;
  assign y19905 = ~1'b0 ;
  assign y19906 = ~1'b0 ;
  assign y19907 = ~n52166 ;
  assign y19908 = ~n52168 ;
  assign y19909 = ~n52177 ;
  assign y19910 = n52182 ;
  assign y19911 = ~n52183 ;
  assign y19912 = ~n52184 ;
  assign y19913 = ~n52186 ;
  assign y19914 = n52188 ;
  assign y19915 = ~n2448 ;
  assign y19916 = n52195 ;
  assign y19917 = ~1'b0 ;
  assign y19918 = ~1'b0 ;
  assign y19919 = n52197 ;
  assign y19920 = n52208 ;
  assign y19921 = ~n52212 ;
  assign y19922 = n52217 ;
  assign y19923 = ~n52218 ;
  assign y19924 = ~n52222 ;
  assign y19925 = n52224 ;
  assign y19926 = ~n52228 ;
  assign y19927 = ~1'b0 ;
  assign y19928 = n52230 ;
  assign y19929 = ~n52231 ;
  assign y19930 = ~n52234 ;
  assign y19931 = ~1'b0 ;
  assign y19932 = n52237 ;
  assign y19933 = ~n52242 ;
  assign y19934 = n52243 ;
  assign y19935 = ~1'b0 ;
  assign y19936 = ~1'b0 ;
  assign y19937 = ~n52244 ;
  assign y19938 = n52249 ;
  assign y19939 = ~1'b0 ;
  assign y19940 = ~n52252 ;
  assign y19941 = ~n52255 ;
  assign y19942 = ~n52260 ;
  assign y19943 = n52261 ;
  assign y19944 = n52263 ;
  assign y19945 = ~n52265 ;
  assign y19946 = ~n52266 ;
  assign y19947 = ~n26355 ;
  assign y19948 = ~n52268 ;
  assign y19949 = n52270 ;
  assign y19950 = ~1'b0 ;
  assign y19951 = n583 ;
  assign y19952 = ~n52275 ;
  assign y19953 = ~n52277 ;
  assign y19954 = ~n52278 ;
  assign y19955 = n52279 ;
  assign y19956 = n52280 ;
  assign y19957 = ~1'b0 ;
  assign y19958 = ~1'b0 ;
  assign y19959 = ~n52287 ;
  assign y19960 = ~1'b0 ;
  assign y19961 = n52288 ;
  assign y19962 = n52291 ;
  assign y19963 = ~n52301 ;
  assign y19964 = n52302 ;
  assign y19965 = n52303 ;
  assign y19966 = ~n52305 ;
  assign y19967 = ~n52308 ;
  assign y19968 = n52310 ;
  assign y19969 = ~1'b0 ;
  assign y19970 = ~n52313 ;
  assign y19971 = n52315 ;
  assign y19972 = ~n52318 ;
  assign y19973 = ~n52320 ;
  assign y19974 = ~n52322 ;
  assign y19975 = n52325 ;
  assign y19976 = n52328 ;
  assign y19977 = n52329 ;
  assign y19978 = n52331 ;
  assign y19979 = ~n52332 ;
  assign y19980 = ~n52334 ;
  assign y19981 = n52336 ;
  assign y19982 = ~n52341 ;
  assign y19983 = ~n52343 ;
  assign y19984 = n52345 ;
  assign y19985 = ~n52357 ;
  assign y19986 = ~n52359 ;
  assign y19987 = n841 ;
  assign y19988 = ~n52361 ;
  assign y19989 = n52365 ;
  assign y19990 = ~1'b0 ;
  assign y19991 = 1'b0 ;
  assign y19992 = ~n52368 ;
  assign y19993 = ~1'b0 ;
  assign y19994 = n52371 ;
  assign y19995 = n52372 ;
  assign y19996 = n52373 ;
  assign y19997 = n52376 ;
  assign y19998 = ~n52377 ;
  assign y19999 = n52378 ;
  assign y20000 = ~n52381 ;
  assign y20001 = ~n52384 ;
  assign y20002 = n52385 ;
  assign y20003 = ~n52388 ;
  assign y20004 = ~1'b0 ;
  assign y20005 = ~n52391 ;
  assign y20006 = n52394 ;
  assign y20007 = ~n52395 ;
  assign y20008 = n52400 ;
  assign y20009 = n52401 ;
  assign y20010 = ~n52412 ;
  assign y20011 = ~n52416 ;
  assign y20012 = ~1'b0 ;
  assign y20013 = ~1'b0 ;
  assign y20014 = ~n52419 ;
  assign y20015 = ~n52421 ;
  assign y20016 = ~n52422 ;
  assign y20017 = n52424 ;
  assign y20018 = n52425 ;
  assign y20019 = n52427 ;
  assign y20020 = n52430 ;
  assign y20021 = n52435 ;
  assign y20022 = n52436 ;
  assign y20023 = ~1'b0 ;
  assign y20024 = ~n52442 ;
  assign y20025 = 1'b0 ;
  assign y20026 = n25261 ;
  assign y20027 = n52443 ;
  assign y20028 = ~n52444 ;
  assign y20029 = ~n52445 ;
  assign y20030 = n52446 ;
  assign y20031 = n52448 ;
  assign y20032 = ~1'b0 ;
  assign y20033 = ~1'b0 ;
  assign y20034 = ~n52450 ;
  assign y20035 = n52454 ;
  assign y20036 = ~n52456 ;
  assign y20037 = ~n48693 ;
  assign y20038 = n52457 ;
  assign y20039 = ~1'b0 ;
  assign y20040 = ~n52458 ;
  assign y20041 = n52459 ;
  assign y20042 = ~n52462 ;
  assign y20043 = ~n52464 ;
  assign y20044 = n52466 ;
  assign y20045 = ~1'b0 ;
  assign y20046 = ~1'b0 ;
  assign y20047 = n52468 ;
  assign y20048 = ~n52470 ;
  assign y20049 = ~n52474 ;
  assign y20050 = ~n52475 ;
  assign y20051 = n52477 ;
  assign y20052 = ~n52478 ;
  assign y20053 = 1'b0 ;
  assign y20054 = ~1'b0 ;
  assign y20055 = n52479 ;
  assign y20056 = n52481 ;
  assign y20057 = ~1'b0 ;
  assign y20058 = ~n52482 ;
  assign y20059 = n52483 ;
  assign y20060 = n52486 ;
  assign y20061 = ~n52487 ;
  assign y20062 = n52492 ;
  assign y20063 = ~n52495 ;
  assign y20064 = ~1'b0 ;
  assign y20065 = n52497 ;
  assign y20066 = ~1'b0 ;
  assign y20067 = ~n52501 ;
  assign y20068 = ~n52504 ;
  assign y20069 = n52506 ;
  assign y20070 = ~n52507 ;
  assign y20071 = n52510 ;
  assign y20072 = n52511 ;
  assign y20073 = n52513 ;
  assign y20074 = n52515 ;
  assign y20075 = ~1'b0 ;
  assign y20076 = n52518 ;
  assign y20077 = n52519 ;
  assign y20078 = ~n52521 ;
  assign y20079 = n52523 ;
  assign y20080 = ~1'b0 ;
  assign y20081 = ~n52526 ;
  assign y20082 = ~n52527 ;
  assign y20083 = ~n42653 ;
  assign y20084 = n52528 ;
  assign y20085 = n52532 ;
  assign y20086 = ~1'b0 ;
  assign y20087 = ~n52533 ;
  assign y20088 = ~n52537 ;
  assign y20089 = ~1'b0 ;
  assign y20090 = n52541 ;
  assign y20091 = n52544 ;
  assign y20092 = n52552 ;
  assign y20093 = n52555 ;
  assign y20094 = n52558 ;
  assign y20095 = ~n52559 ;
  assign y20096 = ~n52562 ;
  assign y20097 = n52568 ;
  assign y20098 = ~1'b0 ;
  assign y20099 = ~1'b0 ;
  assign y20100 = ~n52572 ;
  assign y20101 = n52574 ;
  assign y20102 = ~n52576 ;
  assign y20103 = n52578 ;
  assign y20104 = ~n52581 ;
  assign y20105 = ~n52582 ;
  assign y20106 = n52583 ;
  assign y20107 = ~1'b0 ;
  assign y20108 = ~1'b0 ;
  assign y20109 = n52587 ;
  assign y20110 = n4139 ;
  assign y20111 = n52589 ;
  assign y20112 = ~1'b0 ;
  assign y20113 = ~n52591 ;
  assign y20114 = n52598 ;
  assign y20115 = n52601 ;
  assign y20116 = ~n52605 ;
  assign y20117 = ~n52606 ;
  assign y20118 = n52608 ;
  assign y20119 = ~n52612 ;
  assign y20120 = ~1'b0 ;
  assign y20121 = ~n38332 ;
  assign y20122 = n52613 ;
  assign y20123 = ~n52616 ;
  assign y20124 = n52620 ;
  assign y20125 = ~n52621 ;
  assign y20126 = n52623 ;
  assign y20127 = n52624 ;
  assign y20128 = n52625 ;
  assign y20129 = ~1'b0 ;
  assign y20130 = n52627 ;
  assign y20131 = ~1'b0 ;
  assign y20132 = ~1'b0 ;
  assign y20133 = ~n52629 ;
  assign y20134 = ~n52631 ;
  assign y20135 = n52639 ;
  assign y20136 = ~n52640 ;
  assign y20137 = n52644 ;
  assign y20138 = ~n52647 ;
  assign y20139 = n52648 ;
  assign y20140 = ~n52656 ;
  assign y20141 = ~n52658 ;
  assign y20142 = ~1'b0 ;
  assign y20143 = ~n52660 ;
  assign y20144 = ~1'b0 ;
  assign y20145 = n52664 ;
  assign y20146 = n52668 ;
  assign y20147 = n52669 ;
  assign y20148 = n52674 ;
  assign y20149 = ~n52675 ;
  assign y20150 = n52680 ;
  assign y20151 = ~1'b0 ;
  assign y20152 = ~n52681 ;
  assign y20153 = n52682 ;
  assign y20154 = ~n52683 ;
  assign y20155 = ~n52687 ;
  assign y20156 = n52688 ;
  assign y20157 = n52691 ;
  assign y20158 = n52692 ;
  assign y20159 = n52694 ;
  assign y20160 = ~n52695 ;
  assign y20161 = ~n52696 ;
  assign y20162 = ~1'b0 ;
  assign y20163 = ~1'b0 ;
  assign y20164 = ~n52700 ;
  assign y20165 = n52705 ;
  assign y20166 = ~1'b0 ;
  assign y20167 = n52709 ;
  assign y20168 = n52712 ;
  assign y20169 = n52713 ;
  assign y20170 = ~n52714 ;
  assign y20171 = n52717 ;
  assign y20172 = n52723 ;
  assign y20173 = n52724 ;
  assign y20174 = n52730 ;
  assign y20175 = ~1'b0 ;
  assign y20176 = n52731 ;
  assign y20177 = ~n52733 ;
  assign y20178 = ~1'b0 ;
  assign y20179 = n52737 ;
  assign y20180 = ~n52740 ;
  assign y20181 = n52741 ;
  assign y20182 = ~n52742 ;
  assign y20183 = ~n52743 ;
  assign y20184 = ~1'b0 ;
  assign y20185 = ~n52745 ;
  assign y20186 = ~1'b0 ;
  assign y20187 = ~n52747 ;
  assign y20188 = ~1'b0 ;
  assign y20189 = ~1'b0 ;
  assign y20190 = ~n52748 ;
  assign y20191 = ~n52749 ;
  assign y20192 = ~n52750 ;
  assign y20193 = ~n52751 ;
  assign y20194 = n52755 ;
  assign y20195 = ~1'b0 ;
  assign y20196 = ~n52757 ;
  assign y20197 = n52759 ;
  assign y20198 = ~n52761 ;
  assign y20199 = ~1'b0 ;
  assign y20200 = ~n52764 ;
  assign y20201 = n52774 ;
  assign y20202 = n52775 ;
  assign y20203 = n52779 ;
  assign y20204 = ~n52780 ;
  assign y20205 = ~n52782 ;
  assign y20206 = ~n52786 ;
  assign y20207 = ~n52787 ;
  assign y20208 = ~n52790 ;
  assign y20209 = n52792 ;
  assign y20210 = ~n52793 ;
  assign y20211 = ~n52794 ;
  assign y20212 = ~n52795 ;
  assign y20213 = n52796 ;
  assign y20214 = n52797 ;
  assign y20215 = n52798 ;
  assign y20216 = ~n52799 ;
  assign y20217 = ~1'b0 ;
  assign y20218 = ~n52801 ;
  assign y20219 = ~1'b0 ;
  assign y20220 = ~n52803 ;
  assign y20221 = ~1'b0 ;
  assign y20222 = ~1'b0 ;
  assign y20223 = ~n52804 ;
  assign y20224 = ~n52807 ;
  assign y20225 = ~n52808 ;
  assign y20226 = n52812 ;
  assign y20227 = n52814 ;
  assign y20228 = ~1'b0 ;
  assign y20229 = ~n52822 ;
  assign y20230 = ~n52827 ;
  assign y20231 = ~n52830 ;
  assign y20232 = n52831 ;
  assign y20233 = ~1'b0 ;
  assign y20234 = n52834 ;
  assign y20235 = n52836 ;
  assign y20236 = ~n52839 ;
  assign y20237 = ~n52842 ;
  assign y20238 = n52843 ;
  assign y20239 = ~1'b0 ;
  assign y20240 = ~1'b0 ;
  assign y20241 = n52845 ;
endmodule
