module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7309 , n7310 , n7311 ;
  assign n136 = x77 & x128 ;
  assign n137 = x129 & n136 ;
  assign n138 = x78 & ~x128 ;
  assign n139 = x129 & n138 ;
  assign n140 = ~n137 & ~n139 ;
  assign n141 = x80 & ~x128 ;
  assign n142 = ~x129 & n141 ;
  assign n143 = x79 & x128 ;
  assign n144 = ~x129 & n143 ;
  assign n145 = ~n142 & ~n144 ;
  assign n146 = n140 & n145 ;
  assign n147 = ~x130 & ~x131 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = x73 & x128 ;
  assign n150 = x129 & n149 ;
  assign n151 = x74 & ~x128 ;
  assign n152 = x129 & n151 ;
  assign n153 = ~n150 & ~n152 ;
  assign n154 = x76 & ~x128 ;
  assign n155 = ~x129 & n154 ;
  assign n156 = x75 & x128 ;
  assign n157 = ~x129 & n156 ;
  assign n158 = ~n155 & ~n157 ;
  assign n159 = n153 & n158 ;
  assign n160 = x130 & ~x131 ;
  assign n161 = ~n159 & n160 ;
  assign n162 = ~n148 & ~n161 ;
  assign n163 = x65 & x128 ;
  assign n164 = x129 & n163 ;
  assign n165 = x66 & ~x128 ;
  assign n166 = x129 & n165 ;
  assign n167 = ~n164 & ~n166 ;
  assign n168 = x68 & ~x128 ;
  assign n169 = ~x129 & n168 ;
  assign n170 = x67 & x128 ;
  assign n171 = ~x129 & n170 ;
  assign n172 = ~n169 & ~n171 ;
  assign n173 = n167 & n172 ;
  assign n174 = x130 & x131 ;
  assign n175 = ~n173 & n174 ;
  assign n176 = x69 & x128 ;
  assign n177 = x129 & n176 ;
  assign n178 = x70 & ~x128 ;
  assign n179 = x129 & n178 ;
  assign n180 = ~n177 & ~n179 ;
  assign n181 = x72 & ~x128 ;
  assign n182 = ~x129 & n181 ;
  assign n183 = x71 & x128 ;
  assign n184 = ~x129 & n183 ;
  assign n185 = ~n182 & ~n184 ;
  assign n186 = n180 & n185 ;
  assign n187 = ~x130 & x131 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = ~n175 & ~n188 ;
  assign n190 = n162 & n189 ;
  assign n191 = x132 & x133 ;
  assign n192 = ~n190 & n191 ;
  assign n193 = x93 & x128 ;
  assign n194 = x129 & n193 ;
  assign n195 = x94 & ~x128 ;
  assign n196 = x129 & n195 ;
  assign n197 = ~n194 & ~n196 ;
  assign n198 = x96 & ~x128 ;
  assign n199 = ~x129 & n198 ;
  assign n200 = x95 & x128 ;
  assign n201 = ~x129 & n200 ;
  assign n202 = ~n199 & ~n201 ;
  assign n203 = n197 & n202 ;
  assign n204 = n147 & ~n203 ;
  assign n205 = x89 & x128 ;
  assign n206 = x129 & n205 ;
  assign n207 = x90 & ~x128 ;
  assign n208 = x129 & n207 ;
  assign n209 = ~n206 & ~n208 ;
  assign n210 = x92 & ~x128 ;
  assign n211 = ~x129 & n210 ;
  assign n212 = x91 & x128 ;
  assign n213 = ~x129 & n212 ;
  assign n214 = ~n211 & ~n213 ;
  assign n215 = n209 & n214 ;
  assign n216 = n160 & ~n215 ;
  assign n217 = ~n204 & ~n216 ;
  assign n218 = x81 & x128 ;
  assign n219 = x129 & n218 ;
  assign n220 = x82 & ~x128 ;
  assign n221 = x129 & n220 ;
  assign n222 = ~n219 & ~n221 ;
  assign n223 = x84 & ~x128 ;
  assign n224 = ~x129 & n223 ;
  assign n225 = x83 & x128 ;
  assign n226 = ~x129 & n225 ;
  assign n227 = ~n224 & ~n226 ;
  assign n228 = n222 & n227 ;
  assign n229 = n174 & ~n228 ;
  assign n230 = x85 & x128 ;
  assign n231 = x129 & n230 ;
  assign n232 = x86 & ~x128 ;
  assign n233 = x129 & n232 ;
  assign n234 = ~n231 & ~n233 ;
  assign n235 = x88 & ~x128 ;
  assign n236 = ~x129 & n235 ;
  assign n237 = x87 & x128 ;
  assign n238 = ~x129 & n237 ;
  assign n239 = ~n236 & ~n238 ;
  assign n240 = n234 & n239 ;
  assign n241 = n187 & ~n240 ;
  assign n242 = ~n229 & ~n241 ;
  assign n243 = n217 & n242 ;
  assign n244 = ~x132 & x133 ;
  assign n245 = ~n243 & n244 ;
  assign n246 = ~n192 & ~n245 ;
  assign n247 = x125 & x128 ;
  assign n248 = x129 & n247 ;
  assign n249 = x126 & ~x128 ;
  assign n250 = x129 & n249 ;
  assign n251 = ~n248 & ~n250 ;
  assign n252 = x0 & ~x128 ;
  assign n253 = ~x129 & n252 ;
  assign n254 = x127 & x128 ;
  assign n255 = ~x129 & n254 ;
  assign n256 = ~n253 & ~n255 ;
  assign n257 = n251 & n256 ;
  assign n258 = n147 & ~n257 ;
  assign n259 = x121 & x128 ;
  assign n260 = x129 & n259 ;
  assign n261 = x122 & ~x128 ;
  assign n262 = x129 & n261 ;
  assign n263 = ~n260 & ~n262 ;
  assign n264 = x124 & ~x128 ;
  assign n265 = ~x129 & n264 ;
  assign n266 = x123 & x128 ;
  assign n267 = ~x129 & n266 ;
  assign n268 = ~n265 & ~n267 ;
  assign n269 = n263 & n268 ;
  assign n270 = n160 & ~n269 ;
  assign n271 = ~n258 & ~n270 ;
  assign n272 = x113 & x128 ;
  assign n273 = x129 & n272 ;
  assign n274 = x114 & ~x128 ;
  assign n275 = x129 & n274 ;
  assign n276 = ~n273 & ~n275 ;
  assign n277 = x116 & ~x128 ;
  assign n278 = ~x129 & n277 ;
  assign n279 = x115 & x128 ;
  assign n280 = ~x129 & n279 ;
  assign n281 = ~n278 & ~n280 ;
  assign n282 = n276 & n281 ;
  assign n283 = n174 & ~n282 ;
  assign n284 = x117 & x128 ;
  assign n285 = x129 & n284 ;
  assign n286 = x118 & ~x128 ;
  assign n287 = x129 & n286 ;
  assign n288 = ~n285 & ~n287 ;
  assign n289 = x120 & ~x128 ;
  assign n290 = ~x129 & n289 ;
  assign n291 = x119 & x128 ;
  assign n292 = ~x129 & n291 ;
  assign n293 = ~n290 & ~n292 ;
  assign n294 = n288 & n293 ;
  assign n295 = n187 & ~n294 ;
  assign n296 = ~n283 & ~n295 ;
  assign n297 = n271 & n296 ;
  assign n298 = ~x132 & ~x133 ;
  assign n299 = ~n297 & n298 ;
  assign n300 = x109 & x128 ;
  assign n301 = x129 & n300 ;
  assign n302 = x110 & ~x128 ;
  assign n303 = x129 & n302 ;
  assign n304 = ~n301 & ~n303 ;
  assign n305 = x112 & ~x128 ;
  assign n306 = ~x129 & n305 ;
  assign n307 = x111 & x128 ;
  assign n308 = ~x129 & n307 ;
  assign n309 = ~n306 & ~n308 ;
  assign n310 = n304 & n309 ;
  assign n311 = n147 & ~n310 ;
  assign n312 = x105 & x128 ;
  assign n313 = x129 & n312 ;
  assign n314 = x106 & ~x128 ;
  assign n315 = x129 & n314 ;
  assign n316 = ~n313 & ~n315 ;
  assign n317 = x108 & ~x128 ;
  assign n318 = ~x129 & n317 ;
  assign n319 = x107 & x128 ;
  assign n320 = ~x129 & n319 ;
  assign n321 = ~n318 & ~n320 ;
  assign n322 = n316 & n321 ;
  assign n323 = n160 & ~n322 ;
  assign n324 = ~n311 & ~n323 ;
  assign n325 = x97 & x128 ;
  assign n326 = x129 & n325 ;
  assign n327 = x98 & ~x128 ;
  assign n328 = x129 & n327 ;
  assign n329 = ~n326 & ~n328 ;
  assign n330 = x100 & ~x128 ;
  assign n331 = ~x129 & n330 ;
  assign n332 = x99 & x128 ;
  assign n333 = ~x129 & n332 ;
  assign n334 = ~n331 & ~n333 ;
  assign n335 = n329 & n334 ;
  assign n336 = n174 & ~n335 ;
  assign n337 = x101 & x128 ;
  assign n338 = x129 & n337 ;
  assign n339 = x102 & ~x128 ;
  assign n340 = x129 & n339 ;
  assign n341 = ~n338 & ~n340 ;
  assign n342 = x104 & ~x128 ;
  assign n343 = ~x129 & n342 ;
  assign n344 = x103 & x128 ;
  assign n345 = ~x129 & n344 ;
  assign n346 = ~n343 & ~n345 ;
  assign n347 = n341 & n346 ;
  assign n348 = n187 & ~n347 ;
  assign n349 = ~n336 & ~n348 ;
  assign n350 = n324 & n349 ;
  assign n351 = x132 & ~x133 ;
  assign n352 = ~n350 & n351 ;
  assign n353 = ~n299 & ~n352 ;
  assign n354 = n246 & n353 ;
  assign n355 = ~x134 & ~n354 ;
  assign n356 = x13 & x128 ;
  assign n357 = x129 & n356 ;
  assign n358 = x14 & ~x128 ;
  assign n359 = x129 & n358 ;
  assign n360 = ~n357 & ~n359 ;
  assign n361 = x16 & ~x128 ;
  assign n362 = ~x129 & n361 ;
  assign n363 = x15 & x128 ;
  assign n364 = ~x129 & n363 ;
  assign n365 = ~n362 & ~n364 ;
  assign n366 = n360 & n365 ;
  assign n367 = n147 & ~n366 ;
  assign n368 = x9 & x128 ;
  assign n369 = x129 & n368 ;
  assign n370 = x10 & ~x128 ;
  assign n371 = x129 & n370 ;
  assign n372 = ~n369 & ~n371 ;
  assign n373 = x12 & ~x128 ;
  assign n374 = ~x129 & n373 ;
  assign n375 = x11 & x128 ;
  assign n376 = ~x129 & n375 ;
  assign n377 = ~n374 & ~n376 ;
  assign n378 = n372 & n377 ;
  assign n379 = n160 & ~n378 ;
  assign n380 = ~n367 & ~n379 ;
  assign n381 = x1 & x128 ;
  assign n382 = x129 & n381 ;
  assign n383 = x2 & ~x128 ;
  assign n384 = x129 & n383 ;
  assign n385 = ~n382 & ~n384 ;
  assign n386 = x4 & ~x128 ;
  assign n387 = ~x129 & n386 ;
  assign n388 = x3 & x128 ;
  assign n389 = ~x129 & n388 ;
  assign n390 = ~n387 & ~n389 ;
  assign n391 = n385 & n390 ;
  assign n392 = n174 & ~n391 ;
  assign n393 = x5 & x128 ;
  assign n394 = x129 & n393 ;
  assign n395 = x6 & ~x128 ;
  assign n396 = x129 & n395 ;
  assign n397 = ~n394 & ~n396 ;
  assign n398 = x8 & ~x128 ;
  assign n399 = ~x129 & n398 ;
  assign n400 = x7 & x128 ;
  assign n401 = ~x129 & n400 ;
  assign n402 = ~n399 & ~n401 ;
  assign n403 = n397 & n402 ;
  assign n404 = n187 & ~n403 ;
  assign n405 = ~n392 & ~n404 ;
  assign n406 = n380 & n405 ;
  assign n407 = n191 & ~n406 ;
  assign n408 = x29 & x128 ;
  assign n409 = x129 & n408 ;
  assign n410 = x30 & ~x128 ;
  assign n411 = x129 & n410 ;
  assign n412 = ~n409 & ~n411 ;
  assign n413 = x32 & ~x128 ;
  assign n414 = ~x129 & n413 ;
  assign n415 = x31 & x128 ;
  assign n416 = ~x129 & n415 ;
  assign n417 = ~n414 & ~n416 ;
  assign n418 = n412 & n417 ;
  assign n419 = n147 & ~n418 ;
  assign n420 = x25 & x128 ;
  assign n421 = x129 & n420 ;
  assign n422 = x26 & ~x128 ;
  assign n423 = x129 & n422 ;
  assign n424 = ~n421 & ~n423 ;
  assign n425 = x28 & ~x128 ;
  assign n426 = ~x129 & n425 ;
  assign n427 = x27 & x128 ;
  assign n428 = ~x129 & n427 ;
  assign n429 = ~n426 & ~n428 ;
  assign n430 = n424 & n429 ;
  assign n431 = n160 & ~n430 ;
  assign n432 = ~n419 & ~n431 ;
  assign n433 = x17 & x128 ;
  assign n434 = x129 & n433 ;
  assign n435 = x18 & ~x128 ;
  assign n436 = x129 & n435 ;
  assign n437 = ~n434 & ~n436 ;
  assign n438 = x20 & ~x128 ;
  assign n439 = ~x129 & n438 ;
  assign n440 = x19 & x128 ;
  assign n441 = ~x129 & n440 ;
  assign n442 = ~n439 & ~n441 ;
  assign n443 = n437 & n442 ;
  assign n444 = n174 & ~n443 ;
  assign n445 = x21 & x128 ;
  assign n446 = x129 & n445 ;
  assign n447 = x22 & ~x128 ;
  assign n448 = x129 & n447 ;
  assign n449 = ~n446 & ~n448 ;
  assign n450 = x24 & ~x128 ;
  assign n451 = ~x129 & n450 ;
  assign n452 = x23 & x128 ;
  assign n453 = ~x129 & n452 ;
  assign n454 = ~n451 & ~n453 ;
  assign n455 = n449 & n454 ;
  assign n456 = n187 & ~n455 ;
  assign n457 = ~n444 & ~n456 ;
  assign n458 = n432 & n457 ;
  assign n459 = n244 & ~n458 ;
  assign n460 = ~n407 & ~n459 ;
  assign n461 = x61 & x128 ;
  assign n462 = x129 & n461 ;
  assign n463 = x62 & ~x128 ;
  assign n464 = x129 & n463 ;
  assign n465 = ~n462 & ~n464 ;
  assign n466 = x64 & ~x128 ;
  assign n467 = ~x129 & n466 ;
  assign n468 = x63 & x128 ;
  assign n469 = ~x129 & n468 ;
  assign n470 = ~n467 & ~n469 ;
  assign n471 = n465 & n470 ;
  assign n472 = n147 & ~n471 ;
  assign n473 = x57 & x128 ;
  assign n474 = x129 & n473 ;
  assign n475 = x58 & ~x128 ;
  assign n476 = x129 & n475 ;
  assign n477 = ~n474 & ~n476 ;
  assign n478 = x60 & ~x128 ;
  assign n479 = ~x129 & n478 ;
  assign n480 = x59 & x128 ;
  assign n481 = ~x129 & n480 ;
  assign n482 = ~n479 & ~n481 ;
  assign n483 = n477 & n482 ;
  assign n484 = n160 & ~n483 ;
  assign n485 = ~n472 & ~n484 ;
  assign n486 = x49 & x128 ;
  assign n487 = x129 & n486 ;
  assign n488 = x50 & ~x128 ;
  assign n489 = x129 & n488 ;
  assign n490 = ~n487 & ~n489 ;
  assign n491 = x52 & ~x128 ;
  assign n492 = ~x129 & n491 ;
  assign n493 = x51 & x128 ;
  assign n494 = ~x129 & n493 ;
  assign n495 = ~n492 & ~n494 ;
  assign n496 = n490 & n495 ;
  assign n497 = n174 & ~n496 ;
  assign n498 = x53 & x128 ;
  assign n499 = x129 & n498 ;
  assign n500 = x54 & ~x128 ;
  assign n501 = x129 & n500 ;
  assign n502 = ~n499 & ~n501 ;
  assign n503 = x56 & ~x128 ;
  assign n504 = ~x129 & n503 ;
  assign n505 = x55 & x128 ;
  assign n506 = ~x129 & n505 ;
  assign n507 = ~n504 & ~n506 ;
  assign n508 = n502 & n507 ;
  assign n509 = n187 & ~n508 ;
  assign n510 = ~n497 & ~n509 ;
  assign n511 = n485 & n510 ;
  assign n512 = n298 & ~n511 ;
  assign n513 = x45 & x128 ;
  assign n514 = x129 & n513 ;
  assign n515 = x46 & ~x128 ;
  assign n516 = x129 & n515 ;
  assign n517 = ~n514 & ~n516 ;
  assign n518 = x48 & ~x128 ;
  assign n519 = ~x129 & n518 ;
  assign n520 = x47 & x128 ;
  assign n521 = ~x129 & n520 ;
  assign n522 = ~n519 & ~n521 ;
  assign n523 = n517 & n522 ;
  assign n524 = n147 & ~n523 ;
  assign n525 = x41 & x128 ;
  assign n526 = x129 & n525 ;
  assign n527 = x42 & ~x128 ;
  assign n528 = x129 & n527 ;
  assign n529 = ~n526 & ~n528 ;
  assign n530 = x44 & ~x128 ;
  assign n531 = ~x129 & n530 ;
  assign n532 = x43 & x128 ;
  assign n533 = ~x129 & n532 ;
  assign n534 = ~n531 & ~n533 ;
  assign n535 = n529 & n534 ;
  assign n536 = n160 & ~n535 ;
  assign n537 = ~n524 & ~n536 ;
  assign n538 = x33 & x128 ;
  assign n539 = x129 & n538 ;
  assign n540 = x34 & ~x128 ;
  assign n541 = x129 & n540 ;
  assign n542 = ~n539 & ~n541 ;
  assign n543 = x36 & ~x128 ;
  assign n544 = ~x129 & n543 ;
  assign n545 = x35 & x128 ;
  assign n546 = ~x129 & n545 ;
  assign n547 = ~n544 & ~n546 ;
  assign n548 = n542 & n547 ;
  assign n549 = n174 & ~n548 ;
  assign n550 = x40 & ~x128 ;
  assign n551 = ~x129 & n550 ;
  assign n552 = x37 & x128 ;
  assign n553 = x129 & n552 ;
  assign n554 = ~n551 & ~n553 ;
  assign n555 = x39 & x128 ;
  assign n556 = ~x129 & n555 ;
  assign n557 = x38 & ~x128 ;
  assign n558 = x129 & n557 ;
  assign n559 = ~n556 & ~n558 ;
  assign n560 = n554 & n559 ;
  assign n561 = n187 & ~n560 ;
  assign n562 = ~n549 & ~n561 ;
  assign n563 = n537 & n562 ;
  assign n564 = n351 & ~n563 ;
  assign n565 = ~n512 & ~n564 ;
  assign n566 = n460 & n565 ;
  assign n567 = x134 & ~n566 ;
  assign n568 = ~n355 & ~n567 ;
  assign n995 = ~n568 & x135 ;
  assign n569 = ~x77 & ~x128 ;
  assign n570 = ~x129 & n569 ;
  assign n571 = ~x78 & x128 ;
  assign n572 = ~x129 & n571 ;
  assign n573 = ~n570 & ~n572 ;
  assign n574 = ~x80 & x128 ;
  assign n575 = x129 & n574 ;
  assign n576 = ~x79 & ~x128 ;
  assign n577 = x129 & n576 ;
  assign n578 = ~n575 & ~n577 ;
  assign n579 = n573 & n578 ;
  assign n580 = n174 & ~n579 ;
  assign n581 = ~x73 & ~x128 ;
  assign n582 = ~x129 & n581 ;
  assign n583 = ~x74 & x128 ;
  assign n584 = ~x129 & n583 ;
  assign n585 = ~n582 & ~n584 ;
  assign n586 = ~x76 & x128 ;
  assign n587 = x129 & n586 ;
  assign n588 = ~x75 & ~x128 ;
  assign n589 = x129 & n588 ;
  assign n590 = ~n587 & ~n589 ;
  assign n591 = n585 & n590 ;
  assign n592 = n187 & ~n591 ;
  assign n593 = ~n580 & ~n592 ;
  assign n594 = ~x65 & ~x128 ;
  assign n595 = ~x129 & n594 ;
  assign n596 = ~x66 & x128 ;
  assign n597 = ~x129 & n596 ;
  assign n598 = ~n595 & ~n597 ;
  assign n599 = ~x68 & x128 ;
  assign n600 = x129 & n599 ;
  assign n601 = ~x67 & ~x128 ;
  assign n602 = x129 & n601 ;
  assign n603 = ~n600 & ~n602 ;
  assign n604 = n598 & n603 ;
  assign n605 = n147 & ~n604 ;
  assign n606 = ~x69 & ~x128 ;
  assign n607 = ~x129 & n606 ;
  assign n608 = ~x70 & x128 ;
  assign n609 = ~x129 & n608 ;
  assign n610 = ~n607 & ~n609 ;
  assign n611 = ~x72 & x128 ;
  assign n612 = x129 & n611 ;
  assign n613 = ~x71 & ~x128 ;
  assign n614 = x129 & n613 ;
  assign n615 = ~n612 & ~n614 ;
  assign n616 = n610 & n615 ;
  assign n617 = n160 & ~n616 ;
  assign n618 = ~n605 & ~n617 ;
  assign n619 = n593 & n618 ;
  assign n620 = n298 & ~n619 ;
  assign n621 = ~x93 & ~x128 ;
  assign n622 = ~x129 & n621 ;
  assign n623 = ~x94 & x128 ;
  assign n624 = ~x129 & n623 ;
  assign n625 = ~n622 & ~n624 ;
  assign n626 = ~x96 & x128 ;
  assign n627 = x129 & n626 ;
  assign n628 = ~x95 & ~x128 ;
  assign n629 = x129 & n628 ;
  assign n630 = ~n627 & ~n629 ;
  assign n631 = n625 & n630 ;
  assign n632 = n174 & ~n631 ;
  assign n633 = ~x89 & ~x128 ;
  assign n634 = ~x129 & n633 ;
  assign n635 = ~x90 & x128 ;
  assign n636 = ~x129 & n635 ;
  assign n637 = ~n634 & ~n636 ;
  assign n638 = ~x92 & x128 ;
  assign n639 = x129 & n638 ;
  assign n640 = ~x91 & ~x128 ;
  assign n641 = x129 & n640 ;
  assign n642 = ~n639 & ~n641 ;
  assign n643 = n637 & n642 ;
  assign n644 = n187 & ~n643 ;
  assign n645 = ~n632 & ~n644 ;
  assign n646 = ~x81 & ~x128 ;
  assign n647 = ~x129 & n646 ;
  assign n648 = ~x82 & x128 ;
  assign n649 = ~x129 & n648 ;
  assign n650 = ~n647 & ~n649 ;
  assign n651 = ~x84 & x128 ;
  assign n652 = x129 & n651 ;
  assign n653 = ~x83 & ~x128 ;
  assign n654 = x129 & n653 ;
  assign n655 = ~n652 & ~n654 ;
  assign n656 = n650 & n655 ;
  assign n657 = n147 & ~n656 ;
  assign n658 = ~x85 & ~x128 ;
  assign n659 = ~x129 & n658 ;
  assign n660 = ~x86 & x128 ;
  assign n661 = ~x129 & n660 ;
  assign n662 = ~n659 & ~n661 ;
  assign n663 = ~x88 & x128 ;
  assign n664 = x129 & n663 ;
  assign n665 = ~x87 & ~x128 ;
  assign n666 = x129 & n665 ;
  assign n667 = ~n664 & ~n666 ;
  assign n668 = n662 & n667 ;
  assign n669 = n160 & ~n668 ;
  assign n670 = ~n657 & ~n669 ;
  assign n671 = n645 & n670 ;
  assign n672 = n351 & ~n671 ;
  assign n673 = ~n620 & ~n672 ;
  assign n674 = ~x125 & ~x128 ;
  assign n675 = ~x129 & n674 ;
  assign n676 = ~x126 & x128 ;
  assign n677 = ~x129 & n676 ;
  assign n678 = ~n675 & ~n677 ;
  assign n679 = ~x0 & x128 ;
  assign n680 = x129 & n679 ;
  assign n681 = ~x127 & ~x128 ;
  assign n682 = x129 & n681 ;
  assign n683 = ~n680 & ~n682 ;
  assign n684 = n678 & n683 ;
  assign n685 = n174 & ~n684 ;
  assign n686 = ~x121 & ~x128 ;
  assign n687 = ~x129 & n686 ;
  assign n688 = ~x122 & x128 ;
  assign n689 = ~x129 & n688 ;
  assign n690 = ~n687 & ~n689 ;
  assign n691 = ~x124 & x128 ;
  assign n692 = x129 & n691 ;
  assign n693 = ~x123 & ~x128 ;
  assign n694 = x129 & n693 ;
  assign n695 = ~n692 & ~n694 ;
  assign n696 = n690 & n695 ;
  assign n697 = n187 & ~n696 ;
  assign n698 = ~n685 & ~n697 ;
  assign n699 = ~x113 & ~x128 ;
  assign n700 = ~x129 & n699 ;
  assign n701 = ~x114 & x128 ;
  assign n702 = ~x129 & n701 ;
  assign n703 = ~n700 & ~n702 ;
  assign n704 = ~x116 & x128 ;
  assign n705 = x129 & n704 ;
  assign n706 = ~x115 & ~x128 ;
  assign n707 = x129 & n706 ;
  assign n708 = ~n705 & ~n707 ;
  assign n709 = n703 & n708 ;
  assign n710 = n147 & ~n709 ;
  assign n711 = ~x117 & ~x128 ;
  assign n712 = ~x129 & n711 ;
  assign n713 = ~x118 & x128 ;
  assign n714 = ~x129 & n713 ;
  assign n715 = ~n712 & ~n714 ;
  assign n716 = ~x120 & x128 ;
  assign n717 = x129 & n716 ;
  assign n718 = ~x119 & ~x128 ;
  assign n719 = x129 & n718 ;
  assign n720 = ~n717 & ~n719 ;
  assign n721 = n715 & n720 ;
  assign n722 = n160 & ~n721 ;
  assign n723 = ~n710 & ~n722 ;
  assign n724 = n698 & n723 ;
  assign n725 = n191 & ~n724 ;
  assign n726 = ~x109 & ~x128 ;
  assign n727 = ~x129 & n726 ;
  assign n728 = ~x110 & x128 ;
  assign n729 = ~x129 & n728 ;
  assign n730 = ~n727 & ~n729 ;
  assign n731 = ~x112 & x128 ;
  assign n732 = x129 & n731 ;
  assign n733 = ~x111 & ~x128 ;
  assign n734 = x129 & n733 ;
  assign n735 = ~n732 & ~n734 ;
  assign n736 = n730 & n735 ;
  assign n737 = n174 & ~n736 ;
  assign n738 = ~x105 & ~x128 ;
  assign n739 = ~x129 & n738 ;
  assign n740 = ~x106 & x128 ;
  assign n741 = ~x129 & n740 ;
  assign n742 = ~n739 & ~n741 ;
  assign n743 = ~x108 & x128 ;
  assign n744 = x129 & n743 ;
  assign n745 = ~x107 & ~x128 ;
  assign n746 = x129 & n745 ;
  assign n747 = ~n744 & ~n746 ;
  assign n748 = n742 & n747 ;
  assign n749 = n187 & ~n748 ;
  assign n750 = ~n737 & ~n749 ;
  assign n751 = ~x97 & ~x128 ;
  assign n752 = ~x129 & n751 ;
  assign n753 = ~x98 & x128 ;
  assign n754 = ~x129 & n753 ;
  assign n755 = ~n752 & ~n754 ;
  assign n756 = ~x100 & x128 ;
  assign n757 = x129 & n756 ;
  assign n758 = ~x99 & ~x128 ;
  assign n759 = x129 & n758 ;
  assign n760 = ~n757 & ~n759 ;
  assign n761 = n755 & n760 ;
  assign n762 = n147 & ~n761 ;
  assign n763 = ~x101 & ~x128 ;
  assign n764 = ~x129 & n763 ;
  assign n765 = ~x102 & x128 ;
  assign n766 = ~x129 & n765 ;
  assign n767 = ~n764 & ~n766 ;
  assign n768 = ~x104 & x128 ;
  assign n769 = x129 & n768 ;
  assign n770 = ~x103 & ~x128 ;
  assign n771 = x129 & n770 ;
  assign n772 = ~n769 & ~n771 ;
  assign n773 = n767 & n772 ;
  assign n774 = n160 & ~n773 ;
  assign n775 = ~n762 & ~n774 ;
  assign n776 = n750 & n775 ;
  assign n777 = n244 & ~n776 ;
  assign n778 = ~n725 & ~n777 ;
  assign n779 = n673 & n778 ;
  assign n780 = x134 & ~n779 ;
  assign n781 = ~x13 & ~x128 ;
  assign n782 = ~x129 & n781 ;
  assign n783 = ~x14 & x128 ;
  assign n784 = ~x129 & n783 ;
  assign n785 = ~n782 & ~n784 ;
  assign n786 = ~x16 & x128 ;
  assign n787 = x129 & n786 ;
  assign n788 = ~x15 & ~x128 ;
  assign n789 = x129 & n788 ;
  assign n790 = ~n787 & ~n789 ;
  assign n791 = n785 & n790 ;
  assign n792 = n174 & ~n791 ;
  assign n793 = ~x9 & ~x128 ;
  assign n794 = ~x129 & n793 ;
  assign n795 = ~x10 & x128 ;
  assign n796 = ~x129 & n795 ;
  assign n797 = ~n794 & ~n796 ;
  assign n798 = ~x12 & x128 ;
  assign n799 = x129 & n798 ;
  assign n800 = ~x11 & ~x128 ;
  assign n801 = x129 & n800 ;
  assign n802 = ~n799 & ~n801 ;
  assign n803 = n797 & n802 ;
  assign n804 = n187 & ~n803 ;
  assign n805 = ~n792 & ~n804 ;
  assign n806 = ~x1 & ~x128 ;
  assign n807 = ~x129 & n806 ;
  assign n808 = ~x2 & x128 ;
  assign n809 = ~x129 & n808 ;
  assign n810 = ~n807 & ~n809 ;
  assign n811 = ~x4 & x128 ;
  assign n812 = x129 & n811 ;
  assign n813 = ~x3 & ~x128 ;
  assign n814 = x129 & n813 ;
  assign n815 = ~n812 & ~n814 ;
  assign n816 = n810 & n815 ;
  assign n817 = n147 & ~n816 ;
  assign n818 = ~x5 & ~x128 ;
  assign n819 = ~x129 & n818 ;
  assign n820 = ~x6 & x128 ;
  assign n821 = ~x129 & n820 ;
  assign n822 = ~n819 & ~n821 ;
  assign n823 = ~x8 & x128 ;
  assign n824 = x129 & n823 ;
  assign n825 = ~x7 & ~x128 ;
  assign n826 = x129 & n825 ;
  assign n827 = ~n824 & ~n826 ;
  assign n828 = n822 & n827 ;
  assign n829 = n160 & ~n828 ;
  assign n830 = ~n817 & ~n829 ;
  assign n831 = n805 & n830 ;
  assign n832 = n298 & ~n831 ;
  assign n833 = ~x29 & ~x128 ;
  assign n834 = ~x129 & n833 ;
  assign n835 = ~x30 & x128 ;
  assign n836 = ~x129 & n835 ;
  assign n837 = ~n834 & ~n836 ;
  assign n838 = ~x32 & x128 ;
  assign n839 = x129 & n838 ;
  assign n840 = ~x31 & ~x128 ;
  assign n841 = x129 & n840 ;
  assign n842 = ~n839 & ~n841 ;
  assign n843 = n837 & n842 ;
  assign n844 = n174 & ~n843 ;
  assign n845 = ~x25 & ~x128 ;
  assign n846 = ~x129 & n845 ;
  assign n847 = ~x26 & x128 ;
  assign n848 = ~x129 & n847 ;
  assign n849 = ~n846 & ~n848 ;
  assign n850 = ~x28 & x128 ;
  assign n851 = x129 & n850 ;
  assign n852 = ~x27 & ~x128 ;
  assign n853 = x129 & n852 ;
  assign n854 = ~n851 & ~n853 ;
  assign n855 = n849 & n854 ;
  assign n856 = n187 & ~n855 ;
  assign n857 = ~n844 & ~n856 ;
  assign n858 = ~x17 & ~x128 ;
  assign n859 = ~x129 & n858 ;
  assign n860 = ~x18 & x128 ;
  assign n861 = ~x129 & n860 ;
  assign n862 = ~n859 & ~n861 ;
  assign n863 = ~x20 & x128 ;
  assign n864 = x129 & n863 ;
  assign n865 = ~x19 & ~x128 ;
  assign n866 = x129 & n865 ;
  assign n867 = ~n864 & ~n866 ;
  assign n868 = n862 & n867 ;
  assign n869 = n147 & ~n868 ;
  assign n870 = ~x21 & ~x128 ;
  assign n871 = ~x129 & n870 ;
  assign n872 = ~x22 & x128 ;
  assign n873 = ~x129 & n872 ;
  assign n874 = ~n871 & ~n873 ;
  assign n875 = ~x24 & x128 ;
  assign n876 = x129 & n875 ;
  assign n877 = ~x23 & ~x128 ;
  assign n878 = x129 & n877 ;
  assign n879 = ~n876 & ~n878 ;
  assign n880 = n874 & n879 ;
  assign n881 = n160 & ~n880 ;
  assign n882 = ~n869 & ~n881 ;
  assign n883 = n857 & n882 ;
  assign n884 = n351 & ~n883 ;
  assign n885 = ~n832 & ~n884 ;
  assign n886 = ~x61 & ~x128 ;
  assign n887 = ~x129 & n886 ;
  assign n888 = ~x62 & x128 ;
  assign n889 = ~x129 & n888 ;
  assign n890 = ~n887 & ~n889 ;
  assign n891 = ~x64 & x128 ;
  assign n892 = x129 & n891 ;
  assign n893 = ~x63 & ~x128 ;
  assign n894 = x129 & n893 ;
  assign n895 = ~n892 & ~n894 ;
  assign n896 = n890 & n895 ;
  assign n897 = n174 & ~n896 ;
  assign n898 = ~x57 & ~x128 ;
  assign n899 = ~x129 & n898 ;
  assign n900 = ~x58 & x128 ;
  assign n901 = ~x129 & n900 ;
  assign n902 = ~n899 & ~n901 ;
  assign n903 = ~x60 & x128 ;
  assign n904 = x129 & n903 ;
  assign n905 = ~x59 & ~x128 ;
  assign n906 = x129 & n905 ;
  assign n907 = ~n904 & ~n906 ;
  assign n908 = n902 & n907 ;
  assign n909 = n187 & ~n908 ;
  assign n910 = ~n897 & ~n909 ;
  assign n911 = ~x49 & ~x128 ;
  assign n912 = ~x129 & n911 ;
  assign n913 = ~x50 & x128 ;
  assign n914 = ~x129 & n913 ;
  assign n915 = ~n912 & ~n914 ;
  assign n916 = ~x52 & x128 ;
  assign n917 = x129 & n916 ;
  assign n918 = ~x51 & ~x128 ;
  assign n919 = x129 & n918 ;
  assign n920 = ~n917 & ~n919 ;
  assign n921 = n915 & n920 ;
  assign n922 = n147 & ~n921 ;
  assign n923 = ~x53 & ~x128 ;
  assign n924 = ~x129 & n923 ;
  assign n925 = ~x54 & x128 ;
  assign n926 = ~x129 & n925 ;
  assign n927 = ~n924 & ~n926 ;
  assign n928 = ~x56 & x128 ;
  assign n929 = x129 & n928 ;
  assign n930 = ~x55 & ~x128 ;
  assign n931 = x129 & n930 ;
  assign n932 = ~n929 & ~n931 ;
  assign n933 = n927 & n932 ;
  assign n934 = n160 & ~n933 ;
  assign n935 = ~n922 & ~n934 ;
  assign n936 = n910 & n935 ;
  assign n937 = n191 & ~n936 ;
  assign n938 = ~x45 & ~x128 ;
  assign n939 = ~x129 & n938 ;
  assign n940 = ~x46 & x128 ;
  assign n941 = ~x129 & n940 ;
  assign n942 = ~n939 & ~n941 ;
  assign n943 = ~x48 & x128 ;
  assign n944 = x129 & n943 ;
  assign n945 = ~x47 & ~x128 ;
  assign n946 = x129 & n945 ;
  assign n947 = ~n944 & ~n946 ;
  assign n948 = n942 & n947 ;
  assign n949 = n174 & ~n948 ;
  assign n950 = ~x41 & ~x128 ;
  assign n951 = ~x129 & n950 ;
  assign n952 = ~x42 & x128 ;
  assign n953 = ~x129 & n952 ;
  assign n954 = ~n951 & ~n953 ;
  assign n955 = ~x44 & x128 ;
  assign n956 = x129 & n955 ;
  assign n957 = ~x43 & ~x128 ;
  assign n958 = x129 & n957 ;
  assign n959 = ~n956 & ~n958 ;
  assign n960 = n954 & n959 ;
  assign n961 = n187 & ~n960 ;
  assign n962 = ~n949 & ~n961 ;
  assign n963 = ~x33 & ~x128 ;
  assign n964 = ~x129 & n963 ;
  assign n965 = ~x34 & x128 ;
  assign n966 = ~x129 & n965 ;
  assign n967 = ~n964 & ~n966 ;
  assign n968 = ~x36 & x128 ;
  assign n969 = x129 & n968 ;
  assign n970 = ~x35 & ~x128 ;
  assign n971 = x129 & n970 ;
  assign n972 = ~n969 & ~n971 ;
  assign n973 = n967 & n972 ;
  assign n974 = n147 & ~n973 ;
  assign n975 = ~x40 & x128 ;
  assign n976 = x129 & n975 ;
  assign n977 = ~x37 & ~x128 ;
  assign n978 = ~x129 & n977 ;
  assign n979 = ~n976 & ~n978 ;
  assign n980 = ~x39 & ~x128 ;
  assign n981 = x129 & n980 ;
  assign n982 = ~x38 & x128 ;
  assign n983 = ~x129 & n982 ;
  assign n984 = ~n981 & ~n983 ;
  assign n985 = n979 & n984 ;
  assign n986 = n160 & ~n985 ;
  assign n987 = ~n974 & ~n986 ;
  assign n988 = n962 & n987 ;
  assign n989 = n244 & ~n988 ;
  assign n990 = ~n937 & ~n989 ;
  assign n991 = n885 & n990 ;
  assign n992 = ~x134 & ~n991 ;
  assign n993 = ~n780 & ~n992 ;
  assign n996 = n993 & ~x135 ;
  assign n997 = ~n995 & ~n996 ;
  assign n998 = x81 & ~x128 ;
  assign n999 = ~x129 & n998 ;
  assign n1000 = x78 & x128 ;
  assign n1001 = x129 & n1000 ;
  assign n1002 = ~n999 & ~n1001 ;
  assign n1003 = x80 & x128 ;
  assign n1004 = ~x129 & n1003 ;
  assign n1005 = x79 & ~x128 ;
  assign n1006 = x129 & n1005 ;
  assign n1007 = ~n1004 & ~n1006 ;
  assign n1008 = n1002 & n1007 ;
  assign n1009 = n147 & ~n1008 ;
  assign n1010 = x77 & ~x128 ;
  assign n1011 = ~x129 & n1010 ;
  assign n1012 = x74 & x128 ;
  assign n1013 = x129 & n1012 ;
  assign n1014 = ~n1011 & ~n1013 ;
  assign n1015 = x76 & x128 ;
  assign n1016 = ~x129 & n1015 ;
  assign n1017 = x75 & ~x128 ;
  assign n1018 = x129 & n1017 ;
  assign n1019 = ~n1016 & ~n1018 ;
  assign n1020 = n1014 & n1019 ;
  assign n1021 = n160 & ~n1020 ;
  assign n1022 = ~n1009 & ~n1021 ;
  assign n1023 = x69 & ~x128 ;
  assign n1024 = ~x129 & n1023 ;
  assign n1025 = x66 & x128 ;
  assign n1026 = x129 & n1025 ;
  assign n1027 = ~n1024 & ~n1026 ;
  assign n1028 = x68 & x128 ;
  assign n1029 = ~x129 & n1028 ;
  assign n1030 = x67 & ~x128 ;
  assign n1031 = x129 & n1030 ;
  assign n1032 = ~n1029 & ~n1031 ;
  assign n1033 = n1027 & n1032 ;
  assign n1034 = n174 & ~n1033 ;
  assign n1035 = x73 & ~x128 ;
  assign n1036 = ~x129 & n1035 ;
  assign n1037 = x70 & x128 ;
  assign n1038 = x129 & n1037 ;
  assign n1039 = ~n1036 & ~n1038 ;
  assign n1040 = x72 & x128 ;
  assign n1041 = ~x129 & n1040 ;
  assign n1042 = x71 & ~x128 ;
  assign n1043 = x129 & n1042 ;
  assign n1044 = ~n1041 & ~n1043 ;
  assign n1045 = n1039 & n1044 ;
  assign n1046 = n187 & ~n1045 ;
  assign n1047 = ~n1034 & ~n1046 ;
  assign n1048 = n1022 & n1047 ;
  assign n1049 = n191 & ~n1048 ;
  assign n1050 = x97 & ~x128 ;
  assign n1051 = ~x129 & n1050 ;
  assign n1052 = x94 & x128 ;
  assign n1053 = x129 & n1052 ;
  assign n1054 = ~n1051 & ~n1053 ;
  assign n1055 = x96 & x128 ;
  assign n1056 = ~x129 & n1055 ;
  assign n1057 = x95 & ~x128 ;
  assign n1058 = x129 & n1057 ;
  assign n1059 = ~n1056 & ~n1058 ;
  assign n1060 = n1054 & n1059 ;
  assign n1061 = n147 & ~n1060 ;
  assign n1062 = x93 & ~x128 ;
  assign n1063 = ~x129 & n1062 ;
  assign n1064 = x90 & x128 ;
  assign n1065 = x129 & n1064 ;
  assign n1066 = ~n1063 & ~n1065 ;
  assign n1067 = x92 & x128 ;
  assign n1068 = ~x129 & n1067 ;
  assign n1069 = x91 & ~x128 ;
  assign n1070 = x129 & n1069 ;
  assign n1071 = ~n1068 & ~n1070 ;
  assign n1072 = n1066 & n1071 ;
  assign n1073 = n160 & ~n1072 ;
  assign n1074 = ~n1061 & ~n1073 ;
  assign n1075 = x85 & ~x128 ;
  assign n1076 = ~x129 & n1075 ;
  assign n1077 = x82 & x128 ;
  assign n1078 = x129 & n1077 ;
  assign n1079 = ~n1076 & ~n1078 ;
  assign n1080 = x84 & x128 ;
  assign n1081 = ~x129 & n1080 ;
  assign n1082 = x83 & ~x128 ;
  assign n1083 = x129 & n1082 ;
  assign n1084 = ~n1081 & ~n1083 ;
  assign n1085 = n1079 & n1084 ;
  assign n1086 = n174 & ~n1085 ;
  assign n1087 = x89 & ~x128 ;
  assign n1088 = ~x129 & n1087 ;
  assign n1089 = x86 & x128 ;
  assign n1090 = x129 & n1089 ;
  assign n1091 = ~n1088 & ~n1090 ;
  assign n1092 = x88 & x128 ;
  assign n1093 = ~x129 & n1092 ;
  assign n1094 = x87 & ~x128 ;
  assign n1095 = x129 & n1094 ;
  assign n1096 = ~n1093 & ~n1095 ;
  assign n1097 = n1091 & n1096 ;
  assign n1098 = n187 & ~n1097 ;
  assign n1099 = ~n1086 & ~n1098 ;
  assign n1100 = n1074 & n1099 ;
  assign n1101 = n244 & ~n1100 ;
  assign n1102 = ~n1049 & ~n1101 ;
  assign n1103 = x1 & ~x128 ;
  assign n1104 = ~x129 & n1103 ;
  assign n1105 = x126 & x128 ;
  assign n1106 = x129 & n1105 ;
  assign n1107 = ~n1104 & ~n1106 ;
  assign n1108 = x0 & x128 ;
  assign n1109 = ~x129 & n1108 ;
  assign n1110 = x127 & ~x128 ;
  assign n1111 = x129 & n1110 ;
  assign n1112 = ~n1109 & ~n1111 ;
  assign n1113 = n1107 & n1112 ;
  assign n1114 = n147 & ~n1113 ;
  assign n1115 = x125 & ~x128 ;
  assign n1116 = ~x129 & n1115 ;
  assign n1117 = x122 & x128 ;
  assign n1118 = x129 & n1117 ;
  assign n1119 = ~n1116 & ~n1118 ;
  assign n1120 = x124 & x128 ;
  assign n1121 = ~x129 & n1120 ;
  assign n1122 = x123 & ~x128 ;
  assign n1123 = x129 & n1122 ;
  assign n1124 = ~n1121 & ~n1123 ;
  assign n1125 = n1119 & n1124 ;
  assign n1126 = n160 & ~n1125 ;
  assign n1127 = ~n1114 & ~n1126 ;
  assign n1128 = x117 & ~x128 ;
  assign n1129 = ~x129 & n1128 ;
  assign n1130 = x114 & x128 ;
  assign n1131 = x129 & n1130 ;
  assign n1132 = ~n1129 & ~n1131 ;
  assign n1133 = x116 & x128 ;
  assign n1134 = ~x129 & n1133 ;
  assign n1135 = x115 & ~x128 ;
  assign n1136 = x129 & n1135 ;
  assign n1137 = ~n1134 & ~n1136 ;
  assign n1138 = n1132 & n1137 ;
  assign n1139 = n174 & ~n1138 ;
  assign n1140 = x121 & ~x128 ;
  assign n1141 = ~x129 & n1140 ;
  assign n1142 = x118 & x128 ;
  assign n1143 = x129 & n1142 ;
  assign n1144 = ~n1141 & ~n1143 ;
  assign n1145 = x120 & x128 ;
  assign n1146 = ~x129 & n1145 ;
  assign n1147 = x119 & ~x128 ;
  assign n1148 = x129 & n1147 ;
  assign n1149 = ~n1146 & ~n1148 ;
  assign n1150 = n1144 & n1149 ;
  assign n1151 = n187 & ~n1150 ;
  assign n1152 = ~n1139 & ~n1151 ;
  assign n1153 = n1127 & n1152 ;
  assign n1154 = n298 & ~n1153 ;
  assign n1155 = x113 & ~x128 ;
  assign n1156 = ~x129 & n1155 ;
  assign n1157 = x110 & x128 ;
  assign n1158 = x129 & n1157 ;
  assign n1159 = ~n1156 & ~n1158 ;
  assign n1160 = x112 & x128 ;
  assign n1161 = ~x129 & n1160 ;
  assign n1162 = x111 & ~x128 ;
  assign n1163 = x129 & n1162 ;
  assign n1164 = ~n1161 & ~n1163 ;
  assign n1165 = n1159 & n1164 ;
  assign n1166 = n147 & ~n1165 ;
  assign n1167 = x109 & ~x128 ;
  assign n1168 = ~x129 & n1167 ;
  assign n1169 = x106 & x128 ;
  assign n1170 = x129 & n1169 ;
  assign n1171 = ~n1168 & ~n1170 ;
  assign n1172 = x108 & x128 ;
  assign n1173 = ~x129 & n1172 ;
  assign n1174 = x107 & ~x128 ;
  assign n1175 = x129 & n1174 ;
  assign n1176 = ~n1173 & ~n1175 ;
  assign n1177 = n1171 & n1176 ;
  assign n1178 = n160 & ~n1177 ;
  assign n1179 = ~n1166 & ~n1178 ;
  assign n1180 = x101 & ~x128 ;
  assign n1181 = ~x129 & n1180 ;
  assign n1182 = x98 & x128 ;
  assign n1183 = x129 & n1182 ;
  assign n1184 = ~n1181 & ~n1183 ;
  assign n1185 = x100 & x128 ;
  assign n1186 = ~x129 & n1185 ;
  assign n1187 = x99 & ~x128 ;
  assign n1188 = x129 & n1187 ;
  assign n1189 = ~n1186 & ~n1188 ;
  assign n1190 = n1184 & n1189 ;
  assign n1191 = n174 & ~n1190 ;
  assign n1192 = x105 & ~x128 ;
  assign n1193 = ~x129 & n1192 ;
  assign n1194 = x102 & x128 ;
  assign n1195 = x129 & n1194 ;
  assign n1196 = ~n1193 & ~n1195 ;
  assign n1197 = x104 & x128 ;
  assign n1198 = ~x129 & n1197 ;
  assign n1199 = x103 & ~x128 ;
  assign n1200 = x129 & n1199 ;
  assign n1201 = ~n1198 & ~n1200 ;
  assign n1202 = n1196 & n1201 ;
  assign n1203 = n187 & ~n1202 ;
  assign n1204 = ~n1191 & ~n1203 ;
  assign n1205 = n1179 & n1204 ;
  assign n1206 = n351 & ~n1205 ;
  assign n1207 = ~n1154 & ~n1206 ;
  assign n1208 = n1102 & n1207 ;
  assign n1209 = ~x134 & ~n1208 ;
  assign n1210 = x65 & ~x128 ;
  assign n1211 = ~x129 & n1210 ;
  assign n1212 = x62 & x128 ;
  assign n1213 = x129 & n1212 ;
  assign n1214 = ~n1211 & ~n1213 ;
  assign n1215 = x64 & x128 ;
  assign n1216 = ~x129 & n1215 ;
  assign n1217 = x63 & ~x128 ;
  assign n1218 = x129 & n1217 ;
  assign n1219 = ~n1216 & ~n1218 ;
  assign n1220 = n1214 & n1219 ;
  assign n1221 = n147 & ~n1220 ;
  assign n1222 = x61 & ~x128 ;
  assign n1223 = ~x129 & n1222 ;
  assign n1224 = x58 & x128 ;
  assign n1225 = x129 & n1224 ;
  assign n1226 = ~n1223 & ~n1225 ;
  assign n1227 = x60 & x128 ;
  assign n1228 = ~x129 & n1227 ;
  assign n1229 = x59 & ~x128 ;
  assign n1230 = x129 & n1229 ;
  assign n1231 = ~n1228 & ~n1230 ;
  assign n1232 = n1226 & n1231 ;
  assign n1233 = n160 & ~n1232 ;
  assign n1234 = ~n1221 & ~n1233 ;
  assign n1235 = x53 & ~x128 ;
  assign n1236 = ~x129 & n1235 ;
  assign n1237 = x50 & x128 ;
  assign n1238 = x129 & n1237 ;
  assign n1239 = ~n1236 & ~n1238 ;
  assign n1240 = x52 & x128 ;
  assign n1241 = ~x129 & n1240 ;
  assign n1242 = x51 & ~x128 ;
  assign n1243 = x129 & n1242 ;
  assign n1244 = ~n1241 & ~n1243 ;
  assign n1245 = n1239 & n1244 ;
  assign n1246 = n174 & ~n1245 ;
  assign n1247 = x57 & ~x128 ;
  assign n1248 = ~x129 & n1247 ;
  assign n1249 = x54 & x128 ;
  assign n1250 = x129 & n1249 ;
  assign n1251 = ~n1248 & ~n1250 ;
  assign n1252 = x56 & x128 ;
  assign n1253 = ~x129 & n1252 ;
  assign n1254 = x55 & ~x128 ;
  assign n1255 = x129 & n1254 ;
  assign n1256 = ~n1253 & ~n1255 ;
  assign n1257 = n1251 & n1256 ;
  assign n1258 = n187 & ~n1257 ;
  assign n1259 = ~n1246 & ~n1258 ;
  assign n1260 = n1234 & n1259 ;
  assign n1261 = n298 & ~n1260 ;
  assign n1262 = x17 & ~x128 ;
  assign n1263 = ~x129 & n1262 ;
  assign n1264 = x14 & x128 ;
  assign n1265 = x129 & n1264 ;
  assign n1266 = ~n1263 & ~n1265 ;
  assign n1267 = x16 & x128 ;
  assign n1268 = ~x129 & n1267 ;
  assign n1269 = x15 & ~x128 ;
  assign n1270 = x129 & n1269 ;
  assign n1271 = ~n1268 & ~n1270 ;
  assign n1272 = n1266 & n1271 ;
  assign n1273 = n147 & ~n1272 ;
  assign n1274 = x13 & ~x128 ;
  assign n1275 = ~x129 & n1274 ;
  assign n1276 = x10 & x128 ;
  assign n1277 = x129 & n1276 ;
  assign n1278 = ~n1275 & ~n1277 ;
  assign n1279 = x12 & x128 ;
  assign n1280 = ~x129 & n1279 ;
  assign n1281 = x11 & ~x128 ;
  assign n1282 = x129 & n1281 ;
  assign n1283 = ~n1280 & ~n1282 ;
  assign n1284 = n1278 & n1283 ;
  assign n1285 = n160 & ~n1284 ;
  assign n1286 = ~n1273 & ~n1285 ;
  assign n1287 = x5 & ~x128 ;
  assign n1288 = ~x129 & n1287 ;
  assign n1289 = x2 & x128 ;
  assign n1290 = x129 & n1289 ;
  assign n1291 = ~n1288 & ~n1290 ;
  assign n1292 = x4 & x128 ;
  assign n1293 = ~x129 & n1292 ;
  assign n1294 = x3 & ~x128 ;
  assign n1295 = x129 & n1294 ;
  assign n1296 = ~n1293 & ~n1295 ;
  assign n1297 = n1291 & n1296 ;
  assign n1298 = n174 & ~n1297 ;
  assign n1299 = x9 & ~x128 ;
  assign n1300 = ~x129 & n1299 ;
  assign n1301 = x6 & x128 ;
  assign n1302 = x129 & n1301 ;
  assign n1303 = ~n1300 & ~n1302 ;
  assign n1304 = x8 & x128 ;
  assign n1305 = ~x129 & n1304 ;
  assign n1306 = x7 & ~x128 ;
  assign n1307 = x129 & n1306 ;
  assign n1308 = ~n1305 & ~n1307 ;
  assign n1309 = n1303 & n1308 ;
  assign n1310 = n187 & ~n1309 ;
  assign n1311 = ~n1298 & ~n1310 ;
  assign n1312 = n1286 & n1311 ;
  assign n1313 = n191 & ~n1312 ;
  assign n1314 = ~n1261 & ~n1313 ;
  assign n1315 = x49 & ~x128 ;
  assign n1316 = ~x129 & n1315 ;
  assign n1317 = x46 & x128 ;
  assign n1318 = x129 & n1317 ;
  assign n1319 = ~n1316 & ~n1318 ;
  assign n1320 = x48 & x128 ;
  assign n1321 = ~x129 & n1320 ;
  assign n1322 = x47 & ~x128 ;
  assign n1323 = x129 & n1322 ;
  assign n1324 = ~n1321 & ~n1323 ;
  assign n1325 = n1319 & n1324 ;
  assign n1326 = n147 & ~n1325 ;
  assign n1327 = x42 & x128 ;
  assign n1328 = x129 & n1327 ;
  assign n1329 = x43 & ~x128 ;
  assign n1330 = x129 & n1329 ;
  assign n1331 = ~n1328 & ~n1330 ;
  assign n1332 = x45 & ~x128 ;
  assign n1333 = ~x129 & n1332 ;
  assign n1334 = x44 & x128 ;
  assign n1335 = ~x129 & n1334 ;
  assign n1336 = ~n1333 & ~n1335 ;
  assign n1337 = n1331 & n1336 ;
  assign n1338 = n160 & ~n1337 ;
  assign n1339 = ~n1326 & ~n1338 ;
  assign n1340 = x37 & ~x128 ;
  assign n1341 = ~x129 & n1340 ;
  assign n1342 = x34 & x128 ;
  assign n1343 = x129 & n1342 ;
  assign n1344 = ~n1341 & ~n1343 ;
  assign n1345 = x36 & x128 ;
  assign n1346 = ~x129 & n1345 ;
  assign n1347 = x35 & ~x128 ;
  assign n1348 = x129 & n1347 ;
  assign n1349 = ~n1346 & ~n1348 ;
  assign n1350 = n1344 & n1349 ;
  assign n1351 = n174 & ~n1350 ;
  assign n1352 = x41 & ~x128 ;
  assign n1353 = ~x129 & n1352 ;
  assign n1354 = x40 & x128 ;
  assign n1355 = ~x129 & n1354 ;
  assign n1356 = ~n1353 & ~n1355 ;
  assign n1357 = x39 & ~x128 ;
  assign n1358 = x129 & n1357 ;
  assign n1359 = x38 & x128 ;
  assign n1360 = x129 & n1359 ;
  assign n1361 = ~n1358 & ~n1360 ;
  assign n1362 = n1356 & n1361 ;
  assign n1363 = n187 & ~n1362 ;
  assign n1364 = ~n1351 & ~n1363 ;
  assign n1365 = n1339 & n1364 ;
  assign n1366 = n351 & ~n1365 ;
  assign n1367 = x33 & ~x128 ;
  assign n1368 = ~x129 & n1367 ;
  assign n1369 = x30 & x128 ;
  assign n1370 = x129 & n1369 ;
  assign n1371 = ~n1368 & ~n1370 ;
  assign n1372 = x32 & x128 ;
  assign n1373 = ~x129 & n1372 ;
  assign n1374 = x31 & ~x128 ;
  assign n1375 = x129 & n1374 ;
  assign n1376 = ~n1373 & ~n1375 ;
  assign n1377 = n1371 & n1376 ;
  assign n1378 = n147 & ~n1377 ;
  assign n1379 = x29 & ~x128 ;
  assign n1380 = ~x129 & n1379 ;
  assign n1381 = x26 & x128 ;
  assign n1382 = x129 & n1381 ;
  assign n1383 = ~n1380 & ~n1382 ;
  assign n1384 = x28 & x128 ;
  assign n1385 = ~x129 & n1384 ;
  assign n1386 = x27 & ~x128 ;
  assign n1387 = x129 & n1386 ;
  assign n1388 = ~n1385 & ~n1387 ;
  assign n1389 = n1383 & n1388 ;
  assign n1390 = n160 & ~n1389 ;
  assign n1391 = ~n1378 & ~n1390 ;
  assign n1392 = x21 & ~x128 ;
  assign n1393 = ~x129 & n1392 ;
  assign n1394 = x18 & x128 ;
  assign n1395 = x129 & n1394 ;
  assign n1396 = ~n1393 & ~n1395 ;
  assign n1397 = x20 & x128 ;
  assign n1398 = ~x129 & n1397 ;
  assign n1399 = x19 & ~x128 ;
  assign n1400 = x129 & n1399 ;
  assign n1401 = ~n1398 & ~n1400 ;
  assign n1402 = n1396 & n1401 ;
  assign n1403 = n174 & ~n1402 ;
  assign n1404 = x25 & ~x128 ;
  assign n1405 = ~x129 & n1404 ;
  assign n1406 = x22 & x128 ;
  assign n1407 = x129 & n1406 ;
  assign n1408 = ~n1405 & ~n1407 ;
  assign n1409 = x24 & x128 ;
  assign n1410 = ~x129 & n1409 ;
  assign n1411 = x23 & ~x128 ;
  assign n1412 = x129 & n1411 ;
  assign n1413 = ~n1410 & ~n1412 ;
  assign n1414 = n1408 & n1413 ;
  assign n1415 = n187 & ~n1414 ;
  assign n1416 = ~n1403 & ~n1415 ;
  assign n1417 = n1391 & n1416 ;
  assign n1418 = n244 & ~n1417 ;
  assign n1419 = ~n1366 & ~n1418 ;
  assign n1420 = n1314 & n1419 ;
  assign n1421 = x134 & ~n1420 ;
  assign n1422 = ~n1209 & ~n1421 ;
  assign n1849 = ~n1422 & x136 ;
  assign n1423 = ~x81 & x128 ;
  assign n1424 = x129 & n1423 ;
  assign n1425 = ~x78 & ~x128 ;
  assign n1426 = ~x129 & n1425 ;
  assign n1427 = ~n1424 & ~n1426 ;
  assign n1428 = ~x80 & ~x128 ;
  assign n1429 = x129 & n1428 ;
  assign n1430 = ~x79 & x128 ;
  assign n1431 = ~x129 & n1430 ;
  assign n1432 = ~n1429 & ~n1431 ;
  assign n1433 = n1427 & n1432 ;
  assign n1434 = n174 & ~n1433 ;
  assign n1435 = ~x77 & x128 ;
  assign n1436 = x129 & n1435 ;
  assign n1437 = ~x74 & ~x128 ;
  assign n1438 = ~x129 & n1437 ;
  assign n1439 = ~n1436 & ~n1438 ;
  assign n1440 = ~x76 & ~x128 ;
  assign n1441 = x129 & n1440 ;
  assign n1442 = ~x75 & x128 ;
  assign n1443 = ~x129 & n1442 ;
  assign n1444 = ~n1441 & ~n1443 ;
  assign n1445 = n1439 & n1444 ;
  assign n1446 = n187 & ~n1445 ;
  assign n1447 = ~n1434 & ~n1446 ;
  assign n1448 = ~x69 & x128 ;
  assign n1449 = x129 & n1448 ;
  assign n1450 = ~x66 & ~x128 ;
  assign n1451 = ~x129 & n1450 ;
  assign n1452 = ~n1449 & ~n1451 ;
  assign n1453 = ~x68 & ~x128 ;
  assign n1454 = x129 & n1453 ;
  assign n1455 = ~x67 & x128 ;
  assign n1456 = ~x129 & n1455 ;
  assign n1457 = ~n1454 & ~n1456 ;
  assign n1458 = n1452 & n1457 ;
  assign n1459 = n147 & ~n1458 ;
  assign n1460 = ~x73 & x128 ;
  assign n1461 = x129 & n1460 ;
  assign n1462 = ~x70 & ~x128 ;
  assign n1463 = ~x129 & n1462 ;
  assign n1464 = ~n1461 & ~n1463 ;
  assign n1465 = ~x72 & ~x128 ;
  assign n1466 = x129 & n1465 ;
  assign n1467 = ~x71 & x128 ;
  assign n1468 = ~x129 & n1467 ;
  assign n1469 = ~n1466 & ~n1468 ;
  assign n1470 = n1464 & n1469 ;
  assign n1471 = n160 & ~n1470 ;
  assign n1472 = ~n1459 & ~n1471 ;
  assign n1473 = n1447 & n1472 ;
  assign n1474 = n298 & ~n1473 ;
  assign n1475 = ~x97 & x128 ;
  assign n1476 = x129 & n1475 ;
  assign n1477 = ~x94 & ~x128 ;
  assign n1478 = ~x129 & n1477 ;
  assign n1479 = ~n1476 & ~n1478 ;
  assign n1480 = ~x96 & ~x128 ;
  assign n1481 = x129 & n1480 ;
  assign n1482 = ~x95 & x128 ;
  assign n1483 = ~x129 & n1482 ;
  assign n1484 = ~n1481 & ~n1483 ;
  assign n1485 = n1479 & n1484 ;
  assign n1486 = n174 & ~n1485 ;
  assign n1487 = ~x93 & x128 ;
  assign n1488 = x129 & n1487 ;
  assign n1489 = ~x90 & ~x128 ;
  assign n1490 = ~x129 & n1489 ;
  assign n1491 = ~n1488 & ~n1490 ;
  assign n1492 = ~x92 & ~x128 ;
  assign n1493 = x129 & n1492 ;
  assign n1494 = ~x91 & x128 ;
  assign n1495 = ~x129 & n1494 ;
  assign n1496 = ~n1493 & ~n1495 ;
  assign n1497 = n1491 & n1496 ;
  assign n1498 = n187 & ~n1497 ;
  assign n1499 = ~n1486 & ~n1498 ;
  assign n1500 = ~x85 & x128 ;
  assign n1501 = x129 & n1500 ;
  assign n1502 = ~x82 & ~x128 ;
  assign n1503 = ~x129 & n1502 ;
  assign n1504 = ~n1501 & ~n1503 ;
  assign n1505 = ~x84 & ~x128 ;
  assign n1506 = x129 & n1505 ;
  assign n1507 = ~x83 & x128 ;
  assign n1508 = ~x129 & n1507 ;
  assign n1509 = ~n1506 & ~n1508 ;
  assign n1510 = n1504 & n1509 ;
  assign n1511 = n147 & ~n1510 ;
  assign n1512 = ~x89 & x128 ;
  assign n1513 = x129 & n1512 ;
  assign n1514 = ~x86 & ~x128 ;
  assign n1515 = ~x129 & n1514 ;
  assign n1516 = ~n1513 & ~n1515 ;
  assign n1517 = ~x88 & ~x128 ;
  assign n1518 = x129 & n1517 ;
  assign n1519 = ~x87 & x128 ;
  assign n1520 = ~x129 & n1519 ;
  assign n1521 = ~n1518 & ~n1520 ;
  assign n1522 = n1516 & n1521 ;
  assign n1523 = n160 & ~n1522 ;
  assign n1524 = ~n1511 & ~n1523 ;
  assign n1525 = n1499 & n1524 ;
  assign n1526 = n351 & ~n1525 ;
  assign n1527 = ~n1474 & ~n1526 ;
  assign n1528 = ~x1 & x128 ;
  assign n1529 = x129 & n1528 ;
  assign n1530 = ~x126 & ~x128 ;
  assign n1531 = ~x129 & n1530 ;
  assign n1532 = ~n1529 & ~n1531 ;
  assign n1533 = ~x0 & ~x128 ;
  assign n1534 = x129 & n1533 ;
  assign n1535 = ~x127 & x128 ;
  assign n1536 = ~x129 & n1535 ;
  assign n1537 = ~n1534 & ~n1536 ;
  assign n1538 = n1532 & n1537 ;
  assign n1539 = n174 & ~n1538 ;
  assign n1540 = ~x125 & x128 ;
  assign n1541 = x129 & n1540 ;
  assign n1542 = ~x122 & ~x128 ;
  assign n1543 = ~x129 & n1542 ;
  assign n1544 = ~n1541 & ~n1543 ;
  assign n1545 = ~x124 & ~x128 ;
  assign n1546 = x129 & n1545 ;
  assign n1547 = ~x123 & x128 ;
  assign n1548 = ~x129 & n1547 ;
  assign n1549 = ~n1546 & ~n1548 ;
  assign n1550 = n1544 & n1549 ;
  assign n1551 = n187 & ~n1550 ;
  assign n1552 = ~n1539 & ~n1551 ;
  assign n1553 = ~x117 & x128 ;
  assign n1554 = x129 & n1553 ;
  assign n1555 = ~x114 & ~x128 ;
  assign n1556 = ~x129 & n1555 ;
  assign n1557 = ~n1554 & ~n1556 ;
  assign n1558 = ~x116 & ~x128 ;
  assign n1559 = x129 & n1558 ;
  assign n1560 = ~x115 & x128 ;
  assign n1561 = ~x129 & n1560 ;
  assign n1562 = ~n1559 & ~n1561 ;
  assign n1563 = n1557 & n1562 ;
  assign n1564 = n147 & ~n1563 ;
  assign n1565 = ~x121 & x128 ;
  assign n1566 = x129 & n1565 ;
  assign n1567 = ~x118 & ~x128 ;
  assign n1568 = ~x129 & n1567 ;
  assign n1569 = ~n1566 & ~n1568 ;
  assign n1570 = ~x120 & ~x128 ;
  assign n1571 = x129 & n1570 ;
  assign n1572 = ~x119 & x128 ;
  assign n1573 = ~x129 & n1572 ;
  assign n1574 = ~n1571 & ~n1573 ;
  assign n1575 = n1569 & n1574 ;
  assign n1576 = n160 & ~n1575 ;
  assign n1577 = ~n1564 & ~n1576 ;
  assign n1578 = n1552 & n1577 ;
  assign n1579 = n191 & ~n1578 ;
  assign n1580 = ~x113 & x128 ;
  assign n1581 = x129 & n1580 ;
  assign n1582 = ~x110 & ~x128 ;
  assign n1583 = ~x129 & n1582 ;
  assign n1584 = ~n1581 & ~n1583 ;
  assign n1585 = ~x112 & ~x128 ;
  assign n1586 = x129 & n1585 ;
  assign n1587 = ~x111 & x128 ;
  assign n1588 = ~x129 & n1587 ;
  assign n1589 = ~n1586 & ~n1588 ;
  assign n1590 = n1584 & n1589 ;
  assign n1591 = n174 & ~n1590 ;
  assign n1592 = ~x109 & x128 ;
  assign n1593 = x129 & n1592 ;
  assign n1594 = ~x106 & ~x128 ;
  assign n1595 = ~x129 & n1594 ;
  assign n1596 = ~n1593 & ~n1595 ;
  assign n1597 = ~x108 & ~x128 ;
  assign n1598 = x129 & n1597 ;
  assign n1599 = ~x107 & x128 ;
  assign n1600 = ~x129 & n1599 ;
  assign n1601 = ~n1598 & ~n1600 ;
  assign n1602 = n1596 & n1601 ;
  assign n1603 = n187 & ~n1602 ;
  assign n1604 = ~n1591 & ~n1603 ;
  assign n1605 = ~x101 & x128 ;
  assign n1606 = x129 & n1605 ;
  assign n1607 = ~x98 & ~x128 ;
  assign n1608 = ~x129 & n1607 ;
  assign n1609 = ~n1606 & ~n1608 ;
  assign n1610 = ~x100 & ~x128 ;
  assign n1611 = x129 & n1610 ;
  assign n1612 = ~x99 & x128 ;
  assign n1613 = ~x129 & n1612 ;
  assign n1614 = ~n1611 & ~n1613 ;
  assign n1615 = n1609 & n1614 ;
  assign n1616 = n147 & ~n1615 ;
  assign n1617 = ~x105 & x128 ;
  assign n1618 = x129 & n1617 ;
  assign n1619 = ~x102 & ~x128 ;
  assign n1620 = ~x129 & n1619 ;
  assign n1621 = ~n1618 & ~n1620 ;
  assign n1622 = ~x104 & ~x128 ;
  assign n1623 = x129 & n1622 ;
  assign n1624 = ~x103 & x128 ;
  assign n1625 = ~x129 & n1624 ;
  assign n1626 = ~n1623 & ~n1625 ;
  assign n1627 = n1621 & n1626 ;
  assign n1628 = n160 & ~n1627 ;
  assign n1629 = ~n1616 & ~n1628 ;
  assign n1630 = n1604 & n1629 ;
  assign n1631 = n244 & ~n1630 ;
  assign n1632 = ~n1579 & ~n1631 ;
  assign n1633 = n1527 & n1632 ;
  assign n1634 = x134 & ~n1633 ;
  assign n1635 = ~x65 & x128 ;
  assign n1636 = x129 & n1635 ;
  assign n1637 = ~x62 & ~x128 ;
  assign n1638 = ~x129 & n1637 ;
  assign n1639 = ~n1636 & ~n1638 ;
  assign n1640 = ~x64 & ~x128 ;
  assign n1641 = x129 & n1640 ;
  assign n1642 = ~x63 & x128 ;
  assign n1643 = ~x129 & n1642 ;
  assign n1644 = ~n1641 & ~n1643 ;
  assign n1645 = n1639 & n1644 ;
  assign n1646 = n174 & ~n1645 ;
  assign n1647 = ~x61 & x128 ;
  assign n1648 = x129 & n1647 ;
  assign n1649 = ~x58 & ~x128 ;
  assign n1650 = ~x129 & n1649 ;
  assign n1651 = ~n1648 & ~n1650 ;
  assign n1652 = ~x60 & ~x128 ;
  assign n1653 = x129 & n1652 ;
  assign n1654 = ~x59 & x128 ;
  assign n1655 = ~x129 & n1654 ;
  assign n1656 = ~n1653 & ~n1655 ;
  assign n1657 = n1651 & n1656 ;
  assign n1658 = n187 & ~n1657 ;
  assign n1659 = ~n1646 & ~n1658 ;
  assign n1660 = ~x53 & x128 ;
  assign n1661 = x129 & n1660 ;
  assign n1662 = ~x50 & ~x128 ;
  assign n1663 = ~x129 & n1662 ;
  assign n1664 = ~n1661 & ~n1663 ;
  assign n1665 = ~x52 & ~x128 ;
  assign n1666 = x129 & n1665 ;
  assign n1667 = ~x51 & x128 ;
  assign n1668 = ~x129 & n1667 ;
  assign n1669 = ~n1666 & ~n1668 ;
  assign n1670 = n1664 & n1669 ;
  assign n1671 = n147 & ~n1670 ;
  assign n1672 = ~x57 & x128 ;
  assign n1673 = x129 & n1672 ;
  assign n1674 = ~x54 & ~x128 ;
  assign n1675 = ~x129 & n1674 ;
  assign n1676 = ~n1673 & ~n1675 ;
  assign n1677 = ~x56 & ~x128 ;
  assign n1678 = x129 & n1677 ;
  assign n1679 = ~x55 & x128 ;
  assign n1680 = ~x129 & n1679 ;
  assign n1681 = ~n1678 & ~n1680 ;
  assign n1682 = n1676 & n1681 ;
  assign n1683 = n160 & ~n1682 ;
  assign n1684 = ~n1671 & ~n1683 ;
  assign n1685 = n1659 & n1684 ;
  assign n1686 = n191 & ~n1685 ;
  assign n1687 = ~x17 & x128 ;
  assign n1688 = x129 & n1687 ;
  assign n1689 = ~x14 & ~x128 ;
  assign n1690 = ~x129 & n1689 ;
  assign n1691 = ~n1688 & ~n1690 ;
  assign n1692 = ~x16 & ~x128 ;
  assign n1693 = x129 & n1692 ;
  assign n1694 = ~x15 & x128 ;
  assign n1695 = ~x129 & n1694 ;
  assign n1696 = ~n1693 & ~n1695 ;
  assign n1697 = n1691 & n1696 ;
  assign n1698 = n174 & ~n1697 ;
  assign n1699 = ~x13 & x128 ;
  assign n1700 = x129 & n1699 ;
  assign n1701 = ~x10 & ~x128 ;
  assign n1702 = ~x129 & n1701 ;
  assign n1703 = ~n1700 & ~n1702 ;
  assign n1704 = ~x12 & ~x128 ;
  assign n1705 = x129 & n1704 ;
  assign n1706 = ~x11 & x128 ;
  assign n1707 = ~x129 & n1706 ;
  assign n1708 = ~n1705 & ~n1707 ;
  assign n1709 = n1703 & n1708 ;
  assign n1710 = n187 & ~n1709 ;
  assign n1711 = ~n1698 & ~n1710 ;
  assign n1712 = ~x5 & x128 ;
  assign n1713 = x129 & n1712 ;
  assign n1714 = ~x2 & ~x128 ;
  assign n1715 = ~x129 & n1714 ;
  assign n1716 = ~n1713 & ~n1715 ;
  assign n1717 = ~x4 & ~x128 ;
  assign n1718 = x129 & n1717 ;
  assign n1719 = ~x3 & x128 ;
  assign n1720 = ~x129 & n1719 ;
  assign n1721 = ~n1718 & ~n1720 ;
  assign n1722 = n1716 & n1721 ;
  assign n1723 = n147 & ~n1722 ;
  assign n1724 = ~x9 & x128 ;
  assign n1725 = x129 & n1724 ;
  assign n1726 = ~x6 & ~x128 ;
  assign n1727 = ~x129 & n1726 ;
  assign n1728 = ~n1725 & ~n1727 ;
  assign n1729 = ~x8 & ~x128 ;
  assign n1730 = x129 & n1729 ;
  assign n1731 = ~x7 & x128 ;
  assign n1732 = ~x129 & n1731 ;
  assign n1733 = ~n1730 & ~n1732 ;
  assign n1734 = n1728 & n1733 ;
  assign n1735 = n160 & ~n1734 ;
  assign n1736 = ~n1723 & ~n1735 ;
  assign n1737 = n1711 & n1736 ;
  assign n1738 = n298 & ~n1737 ;
  assign n1739 = ~n1686 & ~n1738 ;
  assign n1740 = ~x49 & x128 ;
  assign n1741 = x129 & n1740 ;
  assign n1742 = ~x46 & ~x128 ;
  assign n1743 = ~x129 & n1742 ;
  assign n1744 = ~n1741 & ~n1743 ;
  assign n1745 = ~x48 & ~x128 ;
  assign n1746 = x129 & n1745 ;
  assign n1747 = ~x47 & x128 ;
  assign n1748 = ~x129 & n1747 ;
  assign n1749 = ~n1746 & ~n1748 ;
  assign n1750 = n1744 & n1749 ;
  assign n1751 = n174 & ~n1750 ;
  assign n1752 = ~x42 & ~x128 ;
  assign n1753 = ~x129 & n1752 ;
  assign n1754 = ~x43 & x128 ;
  assign n1755 = ~x129 & n1754 ;
  assign n1756 = ~n1753 & ~n1755 ;
  assign n1757 = ~x45 & x128 ;
  assign n1758 = x129 & n1757 ;
  assign n1759 = ~x44 & ~x128 ;
  assign n1760 = x129 & n1759 ;
  assign n1761 = ~n1758 & ~n1760 ;
  assign n1762 = n1756 & n1761 ;
  assign n1763 = n187 & ~n1762 ;
  assign n1764 = ~n1751 & ~n1763 ;
  assign n1765 = ~x37 & x128 ;
  assign n1766 = x129 & n1765 ;
  assign n1767 = ~x34 & ~x128 ;
  assign n1768 = ~x129 & n1767 ;
  assign n1769 = ~n1766 & ~n1768 ;
  assign n1770 = ~x36 & ~x128 ;
  assign n1771 = x129 & n1770 ;
  assign n1772 = ~x35 & x128 ;
  assign n1773 = ~x129 & n1772 ;
  assign n1774 = ~n1771 & ~n1773 ;
  assign n1775 = n1769 & n1774 ;
  assign n1776 = n147 & ~n1775 ;
  assign n1777 = ~x41 & x128 ;
  assign n1778 = x129 & n1777 ;
  assign n1779 = ~x40 & ~x128 ;
  assign n1780 = x129 & n1779 ;
  assign n1781 = ~n1778 & ~n1780 ;
  assign n1782 = ~x39 & x128 ;
  assign n1783 = ~x129 & n1782 ;
  assign n1784 = ~x38 & ~x128 ;
  assign n1785 = ~x129 & n1784 ;
  assign n1786 = ~n1783 & ~n1785 ;
  assign n1787 = n1781 & n1786 ;
  assign n1788 = n160 & ~n1787 ;
  assign n1789 = ~n1776 & ~n1788 ;
  assign n1790 = n1764 & n1789 ;
  assign n1791 = n244 & ~n1790 ;
  assign n1792 = ~x33 & x128 ;
  assign n1793 = x129 & n1792 ;
  assign n1794 = ~x30 & ~x128 ;
  assign n1795 = ~x129 & n1794 ;
  assign n1796 = ~n1793 & ~n1795 ;
  assign n1797 = ~x32 & ~x128 ;
  assign n1798 = x129 & n1797 ;
  assign n1799 = ~x31 & x128 ;
  assign n1800 = ~x129 & n1799 ;
  assign n1801 = ~n1798 & ~n1800 ;
  assign n1802 = n1796 & n1801 ;
  assign n1803 = n174 & ~n1802 ;
  assign n1804 = ~x29 & x128 ;
  assign n1805 = x129 & n1804 ;
  assign n1806 = ~x26 & ~x128 ;
  assign n1807 = ~x129 & n1806 ;
  assign n1808 = ~n1805 & ~n1807 ;
  assign n1809 = ~x28 & ~x128 ;
  assign n1810 = x129 & n1809 ;
  assign n1811 = ~x27 & x128 ;
  assign n1812 = ~x129 & n1811 ;
  assign n1813 = ~n1810 & ~n1812 ;
  assign n1814 = n1808 & n1813 ;
  assign n1815 = n187 & ~n1814 ;
  assign n1816 = ~n1803 & ~n1815 ;
  assign n1817 = ~x21 & x128 ;
  assign n1818 = x129 & n1817 ;
  assign n1819 = ~x18 & ~x128 ;
  assign n1820 = ~x129 & n1819 ;
  assign n1821 = ~n1818 & ~n1820 ;
  assign n1822 = ~x20 & ~x128 ;
  assign n1823 = x129 & n1822 ;
  assign n1824 = ~x19 & x128 ;
  assign n1825 = ~x129 & n1824 ;
  assign n1826 = ~n1823 & ~n1825 ;
  assign n1827 = n1821 & n1826 ;
  assign n1828 = n147 & ~n1827 ;
  assign n1829 = ~x25 & x128 ;
  assign n1830 = x129 & n1829 ;
  assign n1831 = ~x22 & ~x128 ;
  assign n1832 = ~x129 & n1831 ;
  assign n1833 = ~n1830 & ~n1832 ;
  assign n1834 = ~x24 & ~x128 ;
  assign n1835 = x129 & n1834 ;
  assign n1836 = ~x23 & x128 ;
  assign n1837 = ~x129 & n1836 ;
  assign n1838 = ~n1835 & ~n1837 ;
  assign n1839 = n1833 & n1838 ;
  assign n1840 = n160 & ~n1839 ;
  assign n1841 = ~n1828 & ~n1840 ;
  assign n1842 = n1816 & n1841 ;
  assign n1843 = n351 & ~n1842 ;
  assign n1844 = ~n1791 & ~n1843 ;
  assign n1845 = n1739 & n1844 ;
  assign n1846 = ~x134 & ~n1845 ;
  assign n1847 = ~n1634 & ~n1846 ;
  assign n1850 = n1847 & ~x136 ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = ~x129 & n218 ;
  assign n1853 = ~x129 & n220 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = x129 & n141 ;
  assign n1856 = x129 & n143 ;
  assign n1857 = ~n1855 & ~n1856 ;
  assign n1858 = n1854 & n1857 ;
  assign n1859 = n147 & ~n1858 ;
  assign n1860 = ~x129 & n136 ;
  assign n1861 = ~x129 & n138 ;
  assign n1862 = ~n1860 & ~n1861 ;
  assign n1863 = x129 & n154 ;
  assign n1864 = x129 & n156 ;
  assign n1865 = ~n1863 & ~n1864 ;
  assign n1866 = n1862 & n1865 ;
  assign n1867 = n160 & ~n1866 ;
  assign n1868 = ~n1859 & ~n1867 ;
  assign n1869 = ~x129 & n176 ;
  assign n1870 = ~x129 & n178 ;
  assign n1871 = ~n1869 & ~n1870 ;
  assign n1872 = x129 & n168 ;
  assign n1873 = x129 & n170 ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = n1871 & n1874 ;
  assign n1876 = n174 & ~n1875 ;
  assign n1877 = ~x129 & n149 ;
  assign n1878 = ~x129 & n151 ;
  assign n1879 = ~n1877 & ~n1878 ;
  assign n1880 = x129 & n181 ;
  assign n1881 = x129 & n183 ;
  assign n1882 = ~n1880 & ~n1881 ;
  assign n1883 = n1879 & n1882 ;
  assign n1884 = n187 & ~n1883 ;
  assign n1885 = ~n1876 & ~n1884 ;
  assign n1886 = n1868 & n1885 ;
  assign n1887 = n191 & ~n1886 ;
  assign n1888 = ~x129 & n325 ;
  assign n1889 = ~x129 & n327 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = x129 & n198 ;
  assign n1892 = x129 & n200 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = n1890 & n1893 ;
  assign n1895 = n147 & ~n1894 ;
  assign n1896 = ~x129 & n193 ;
  assign n1897 = ~x129 & n195 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1899 = x129 & n210 ;
  assign n1900 = x129 & n212 ;
  assign n1901 = ~n1899 & ~n1900 ;
  assign n1902 = n1898 & n1901 ;
  assign n1903 = n160 & ~n1902 ;
  assign n1904 = ~n1895 & ~n1903 ;
  assign n1905 = ~x129 & n230 ;
  assign n1906 = ~x129 & n232 ;
  assign n1907 = ~n1905 & ~n1906 ;
  assign n1908 = x129 & n223 ;
  assign n1909 = x129 & n225 ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1911 = n1907 & n1910 ;
  assign n1912 = n174 & ~n1911 ;
  assign n1913 = ~x129 & n205 ;
  assign n1914 = ~x129 & n207 ;
  assign n1915 = ~n1913 & ~n1914 ;
  assign n1916 = x129 & n235 ;
  assign n1917 = x129 & n237 ;
  assign n1918 = ~n1916 & ~n1917 ;
  assign n1919 = n1915 & n1918 ;
  assign n1920 = n187 & ~n1919 ;
  assign n1921 = ~n1912 & ~n1920 ;
  assign n1922 = n1904 & n1921 ;
  assign n1923 = n244 & ~n1922 ;
  assign n1924 = ~n1887 & ~n1923 ;
  assign n1925 = ~x129 & n381 ;
  assign n1926 = ~x129 & n383 ;
  assign n1927 = ~n1925 & ~n1926 ;
  assign n1928 = x129 & n252 ;
  assign n1929 = x129 & n254 ;
  assign n1930 = ~n1928 & ~n1929 ;
  assign n1931 = n1927 & n1930 ;
  assign n1932 = n147 & ~n1931 ;
  assign n1933 = ~x129 & n247 ;
  assign n1934 = ~x129 & n249 ;
  assign n1935 = ~n1933 & ~n1934 ;
  assign n1936 = x129 & n264 ;
  assign n1937 = x129 & n266 ;
  assign n1938 = ~n1936 & ~n1937 ;
  assign n1939 = n1935 & n1938 ;
  assign n1940 = n160 & ~n1939 ;
  assign n1941 = ~n1932 & ~n1940 ;
  assign n1942 = ~x129 & n284 ;
  assign n1943 = ~x129 & n286 ;
  assign n1944 = ~n1942 & ~n1943 ;
  assign n1945 = x129 & n277 ;
  assign n1946 = x129 & n279 ;
  assign n1947 = ~n1945 & ~n1946 ;
  assign n1948 = n1944 & n1947 ;
  assign n1949 = n174 & ~n1948 ;
  assign n1950 = ~x129 & n259 ;
  assign n1951 = ~x129 & n261 ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1953 = x129 & n289 ;
  assign n1954 = x129 & n291 ;
  assign n1955 = ~n1953 & ~n1954 ;
  assign n1956 = n1952 & n1955 ;
  assign n1957 = n187 & ~n1956 ;
  assign n1958 = ~n1949 & ~n1957 ;
  assign n1959 = n1941 & n1958 ;
  assign n1960 = n298 & ~n1959 ;
  assign n1961 = ~x129 & n272 ;
  assign n1962 = ~x129 & n274 ;
  assign n1963 = ~n1961 & ~n1962 ;
  assign n1964 = x129 & n305 ;
  assign n1965 = x129 & n307 ;
  assign n1966 = ~n1964 & ~n1965 ;
  assign n1967 = n1963 & n1966 ;
  assign n1968 = n147 & ~n1967 ;
  assign n1969 = ~x129 & n300 ;
  assign n1970 = ~x129 & n302 ;
  assign n1971 = ~n1969 & ~n1970 ;
  assign n1972 = x129 & n317 ;
  assign n1973 = x129 & n319 ;
  assign n1974 = ~n1972 & ~n1973 ;
  assign n1975 = n1971 & n1974 ;
  assign n1976 = n160 & ~n1975 ;
  assign n1977 = ~n1968 & ~n1976 ;
  assign n1978 = ~x129 & n337 ;
  assign n1979 = ~x129 & n339 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = x129 & n330 ;
  assign n1982 = x129 & n332 ;
  assign n1983 = ~n1981 & ~n1982 ;
  assign n1984 = n1980 & n1983 ;
  assign n1985 = n174 & ~n1984 ;
  assign n1986 = ~x129 & n312 ;
  assign n1987 = ~x129 & n314 ;
  assign n1988 = ~n1986 & ~n1987 ;
  assign n1989 = x129 & n342 ;
  assign n1990 = x129 & n344 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = n1988 & n1991 ;
  assign n1993 = n187 & ~n1992 ;
  assign n1994 = ~n1985 & ~n1993 ;
  assign n1995 = n1977 & n1994 ;
  assign n1996 = n351 & ~n1995 ;
  assign n1997 = ~n1960 & ~n1996 ;
  assign n1998 = n1924 & n1997 ;
  assign n1999 = ~x134 & ~n1998 ;
  assign n2000 = ~x129 & n163 ;
  assign n2001 = ~x129 & n165 ;
  assign n2002 = ~n2000 & ~n2001 ;
  assign n2003 = x129 & n466 ;
  assign n2004 = x129 & n468 ;
  assign n2005 = ~n2003 & ~n2004 ;
  assign n2006 = n2002 & n2005 ;
  assign n2007 = n147 & ~n2006 ;
  assign n2008 = ~x129 & n461 ;
  assign n2009 = ~x129 & n463 ;
  assign n2010 = ~n2008 & ~n2009 ;
  assign n2011 = x129 & n478 ;
  assign n2012 = x129 & n480 ;
  assign n2013 = ~n2011 & ~n2012 ;
  assign n2014 = n2010 & n2013 ;
  assign n2015 = n160 & ~n2014 ;
  assign n2016 = ~n2007 & ~n2015 ;
  assign n2017 = ~x129 & n498 ;
  assign n2018 = ~x129 & n500 ;
  assign n2019 = ~n2017 & ~n2018 ;
  assign n2020 = x129 & n491 ;
  assign n2021 = x129 & n493 ;
  assign n2022 = ~n2020 & ~n2021 ;
  assign n2023 = n2019 & n2022 ;
  assign n2024 = n174 & ~n2023 ;
  assign n2025 = ~x129 & n473 ;
  assign n2026 = ~x129 & n475 ;
  assign n2027 = ~n2025 & ~n2026 ;
  assign n2028 = x129 & n503 ;
  assign n2029 = x129 & n505 ;
  assign n2030 = ~n2028 & ~n2029 ;
  assign n2031 = n2027 & n2030 ;
  assign n2032 = n187 & ~n2031 ;
  assign n2033 = ~n2024 & ~n2032 ;
  assign n2034 = n2016 & n2033 ;
  assign n2035 = n298 & ~n2034 ;
  assign n2036 = ~x129 & n433 ;
  assign n2037 = ~x129 & n435 ;
  assign n2038 = ~n2036 & ~n2037 ;
  assign n2039 = x129 & n361 ;
  assign n2040 = x129 & n363 ;
  assign n2041 = ~n2039 & ~n2040 ;
  assign n2042 = n2038 & n2041 ;
  assign n2043 = n147 & ~n2042 ;
  assign n2044 = ~x129 & n356 ;
  assign n2045 = ~x129 & n358 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = x129 & n373 ;
  assign n2048 = x129 & n375 ;
  assign n2049 = ~n2047 & ~n2048 ;
  assign n2050 = n2046 & n2049 ;
  assign n2051 = n160 & ~n2050 ;
  assign n2052 = ~n2043 & ~n2051 ;
  assign n2053 = ~x129 & n393 ;
  assign n2054 = ~x129 & n395 ;
  assign n2055 = ~n2053 & ~n2054 ;
  assign n2056 = x129 & n386 ;
  assign n2057 = x129 & n388 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2059 = n2055 & n2058 ;
  assign n2060 = n174 & ~n2059 ;
  assign n2061 = ~x129 & n368 ;
  assign n2062 = ~x129 & n370 ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = x129 & n398 ;
  assign n2065 = x129 & n400 ;
  assign n2066 = ~n2064 & ~n2065 ;
  assign n2067 = n2063 & n2066 ;
  assign n2068 = n187 & ~n2067 ;
  assign n2069 = ~n2060 & ~n2068 ;
  assign n2070 = n2052 & n2069 ;
  assign n2071 = n191 & ~n2070 ;
  assign n2072 = ~n2035 & ~n2071 ;
  assign n2073 = ~x129 & n486 ;
  assign n2074 = ~x129 & n488 ;
  assign n2075 = ~n2073 & ~n2074 ;
  assign n2076 = x129 & n518 ;
  assign n2077 = x129 & n520 ;
  assign n2078 = ~n2076 & ~n2077 ;
  assign n2079 = n2075 & n2078 ;
  assign n2080 = n147 & ~n2079 ;
  assign n2081 = x129 & n532 ;
  assign n2082 = x129 & n530 ;
  assign n2083 = ~n2081 & ~n2082 ;
  assign n2084 = ~x129 & n515 ;
  assign n2085 = ~x129 & n513 ;
  assign n2086 = ~n2084 & ~n2085 ;
  assign n2087 = n2083 & n2086 ;
  assign n2088 = n160 & ~n2087 ;
  assign n2089 = ~n2080 & ~n2088 ;
  assign n2090 = ~x129 & n552 ;
  assign n2091 = ~x129 & n557 ;
  assign n2092 = ~n2090 & ~n2091 ;
  assign n2093 = x129 & n543 ;
  assign n2094 = x129 & n545 ;
  assign n2095 = ~n2093 & ~n2094 ;
  assign n2096 = n2092 & n2095 ;
  assign n2097 = n174 & ~n2096 ;
  assign n2098 = ~x129 & n525 ;
  assign n2099 = ~x129 & n527 ;
  assign n2100 = ~n2098 & ~n2099 ;
  assign n2101 = x129 & n555 ;
  assign n2102 = x129 & n550 ;
  assign n2103 = ~n2101 & ~n2102 ;
  assign n2104 = n2100 & n2103 ;
  assign n2105 = n187 & ~n2104 ;
  assign n2106 = ~n2097 & ~n2105 ;
  assign n2107 = n2089 & n2106 ;
  assign n2108 = n351 & ~n2107 ;
  assign n2109 = ~x129 & n538 ;
  assign n2110 = ~x129 & n540 ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = x129 & n413 ;
  assign n2113 = x129 & n415 ;
  assign n2114 = ~n2112 & ~n2113 ;
  assign n2115 = n2111 & n2114 ;
  assign n2116 = n147 & ~n2115 ;
  assign n2117 = ~x129 & n408 ;
  assign n2118 = ~x129 & n410 ;
  assign n2119 = ~n2117 & ~n2118 ;
  assign n2120 = x129 & n425 ;
  assign n2121 = x129 & n427 ;
  assign n2122 = ~n2120 & ~n2121 ;
  assign n2123 = n2119 & n2122 ;
  assign n2124 = n160 & ~n2123 ;
  assign n2125 = ~n2116 & ~n2124 ;
  assign n2126 = ~x129 & n445 ;
  assign n2127 = ~x129 & n447 ;
  assign n2128 = ~n2126 & ~n2127 ;
  assign n2129 = x129 & n438 ;
  assign n2130 = x129 & n440 ;
  assign n2131 = ~n2129 & ~n2130 ;
  assign n2132 = n2128 & n2131 ;
  assign n2133 = n174 & ~n2132 ;
  assign n2134 = ~x129 & n420 ;
  assign n2135 = ~x129 & n422 ;
  assign n2136 = ~n2134 & ~n2135 ;
  assign n2137 = x129 & n450 ;
  assign n2138 = x129 & n452 ;
  assign n2139 = ~n2137 & ~n2138 ;
  assign n2140 = n2136 & n2139 ;
  assign n2141 = n187 & ~n2140 ;
  assign n2142 = ~n2133 & ~n2141 ;
  assign n2143 = n2125 & n2142 ;
  assign n2144 = n244 & ~n2143 ;
  assign n2145 = ~n2108 & ~n2144 ;
  assign n2146 = n2072 & n2145 ;
  assign n2147 = x134 & ~n2146 ;
  assign n2148 = ~n1999 & ~n2147 ;
  assign n2447 = ~n2148 & x137 ;
  assign n2149 = x129 & n646 ;
  assign n2150 = x129 & n648 ;
  assign n2151 = ~n2149 & ~n2150 ;
  assign n2152 = ~x129 & n574 ;
  assign n2153 = ~x129 & n576 ;
  assign n2154 = ~n2152 & ~n2153 ;
  assign n2155 = n2151 & n2154 ;
  assign n2156 = n174 & ~n2155 ;
  assign n2157 = x129 & n569 ;
  assign n2158 = x129 & n571 ;
  assign n2159 = ~n2157 & ~n2158 ;
  assign n2160 = ~x129 & n586 ;
  assign n2161 = ~x129 & n588 ;
  assign n2162 = ~n2160 & ~n2161 ;
  assign n2163 = n2159 & n2162 ;
  assign n2164 = n187 & ~n2163 ;
  assign n2165 = ~n2156 & ~n2164 ;
  assign n2166 = x129 & n606 ;
  assign n2167 = x129 & n608 ;
  assign n2168 = ~n2166 & ~n2167 ;
  assign n2169 = ~x129 & n599 ;
  assign n2170 = ~x129 & n601 ;
  assign n2171 = ~n2169 & ~n2170 ;
  assign n2172 = n2168 & n2171 ;
  assign n2173 = n147 & ~n2172 ;
  assign n2174 = x129 & n581 ;
  assign n2175 = x129 & n583 ;
  assign n2176 = ~n2174 & ~n2175 ;
  assign n2177 = ~x129 & n611 ;
  assign n2178 = ~x129 & n613 ;
  assign n2179 = ~n2177 & ~n2178 ;
  assign n2180 = n2176 & n2179 ;
  assign n2181 = n160 & ~n2180 ;
  assign n2182 = ~n2173 & ~n2181 ;
  assign n2183 = n2165 & n2182 ;
  assign n2184 = n298 & ~n2183 ;
  assign n2185 = x129 & n751 ;
  assign n2186 = x129 & n753 ;
  assign n2187 = ~n2185 & ~n2186 ;
  assign n2188 = ~x129 & n626 ;
  assign n2189 = ~x129 & n628 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2191 = n2187 & n2190 ;
  assign n2192 = n174 & ~n2191 ;
  assign n2193 = x129 & n621 ;
  assign n2194 = x129 & n623 ;
  assign n2195 = ~n2193 & ~n2194 ;
  assign n2196 = ~x129 & n638 ;
  assign n2197 = ~x129 & n640 ;
  assign n2198 = ~n2196 & ~n2197 ;
  assign n2199 = n2195 & n2198 ;
  assign n2200 = n187 & ~n2199 ;
  assign n2201 = ~n2192 & ~n2200 ;
  assign n2202 = x129 & n658 ;
  assign n2203 = x129 & n660 ;
  assign n2204 = ~n2202 & ~n2203 ;
  assign n2205 = ~x129 & n651 ;
  assign n2206 = ~x129 & n653 ;
  assign n2207 = ~n2205 & ~n2206 ;
  assign n2208 = n2204 & n2207 ;
  assign n2209 = n147 & ~n2208 ;
  assign n2210 = x129 & n633 ;
  assign n2211 = x129 & n635 ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2213 = ~x129 & n663 ;
  assign n2214 = ~x129 & n665 ;
  assign n2215 = ~n2213 & ~n2214 ;
  assign n2216 = n2212 & n2215 ;
  assign n2217 = n160 & ~n2216 ;
  assign n2218 = ~n2209 & ~n2217 ;
  assign n2219 = n2201 & n2218 ;
  assign n2220 = n351 & ~n2219 ;
  assign n2221 = ~n2184 & ~n2220 ;
  assign n2222 = x129 & n806 ;
  assign n2223 = x129 & n808 ;
  assign n2224 = ~n2222 & ~n2223 ;
  assign n2225 = ~x129 & n679 ;
  assign n2226 = ~x129 & n681 ;
  assign n2227 = ~n2225 & ~n2226 ;
  assign n2228 = n2224 & n2227 ;
  assign n2229 = n174 & ~n2228 ;
  assign n2230 = x129 & n674 ;
  assign n2231 = x129 & n676 ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = ~x129 & n691 ;
  assign n2234 = ~x129 & n693 ;
  assign n2235 = ~n2233 & ~n2234 ;
  assign n2236 = n2232 & n2235 ;
  assign n2237 = n187 & ~n2236 ;
  assign n2238 = ~n2229 & ~n2237 ;
  assign n2239 = x129 & n711 ;
  assign n2240 = x129 & n713 ;
  assign n2241 = ~n2239 & ~n2240 ;
  assign n2242 = ~x129 & n704 ;
  assign n2243 = ~x129 & n706 ;
  assign n2244 = ~n2242 & ~n2243 ;
  assign n2245 = n2241 & n2244 ;
  assign n2246 = n147 & ~n2245 ;
  assign n2247 = x129 & n686 ;
  assign n2248 = x129 & n688 ;
  assign n2249 = ~n2247 & ~n2248 ;
  assign n2250 = ~x129 & n716 ;
  assign n2251 = ~x129 & n718 ;
  assign n2252 = ~n2250 & ~n2251 ;
  assign n2253 = n2249 & n2252 ;
  assign n2254 = n160 & ~n2253 ;
  assign n2255 = ~n2246 & ~n2254 ;
  assign n2256 = n2238 & n2255 ;
  assign n2257 = n191 & ~n2256 ;
  assign n2258 = x129 & n699 ;
  assign n2259 = x129 & n701 ;
  assign n2260 = ~n2258 & ~n2259 ;
  assign n2261 = ~x129 & n731 ;
  assign n2262 = ~x129 & n733 ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2264 = n2260 & n2263 ;
  assign n2265 = n174 & ~n2264 ;
  assign n2266 = x129 & n726 ;
  assign n2267 = x129 & n728 ;
  assign n2268 = ~n2266 & ~n2267 ;
  assign n2269 = ~x129 & n743 ;
  assign n2270 = ~x129 & n745 ;
  assign n2271 = ~n2269 & ~n2270 ;
  assign n2272 = n2268 & n2271 ;
  assign n2273 = n187 & ~n2272 ;
  assign n2274 = ~n2265 & ~n2273 ;
  assign n2275 = x129 & n763 ;
  assign n2276 = x129 & n765 ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = ~x129 & n756 ;
  assign n2279 = ~x129 & n758 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = n2277 & n2280 ;
  assign n2282 = n147 & ~n2281 ;
  assign n2283 = x129 & n738 ;
  assign n2284 = x129 & n740 ;
  assign n2285 = ~n2283 & ~n2284 ;
  assign n2286 = ~x129 & n768 ;
  assign n2287 = ~x129 & n770 ;
  assign n2288 = ~n2286 & ~n2287 ;
  assign n2289 = n2285 & n2288 ;
  assign n2290 = n160 & ~n2289 ;
  assign n2291 = ~n2282 & ~n2290 ;
  assign n2292 = n2274 & n2291 ;
  assign n2293 = n244 & ~n2292 ;
  assign n2294 = ~n2257 & ~n2293 ;
  assign n2295 = n2221 & n2294 ;
  assign n2296 = x134 & ~n2295 ;
  assign n2297 = x129 & n594 ;
  assign n2298 = x129 & n596 ;
  assign n2299 = ~n2297 & ~n2298 ;
  assign n2300 = ~x129 & n891 ;
  assign n2301 = ~x129 & n893 ;
  assign n2302 = ~n2300 & ~n2301 ;
  assign n2303 = n2299 & n2302 ;
  assign n2304 = n174 & ~n2303 ;
  assign n2305 = x129 & n886 ;
  assign n2306 = x129 & n888 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = ~x129 & n903 ;
  assign n2309 = ~x129 & n905 ;
  assign n2310 = ~n2308 & ~n2309 ;
  assign n2311 = n2307 & n2310 ;
  assign n2312 = n187 & ~n2311 ;
  assign n2313 = ~n2304 & ~n2312 ;
  assign n2314 = x129 & n923 ;
  assign n2315 = x129 & n925 ;
  assign n2316 = ~n2314 & ~n2315 ;
  assign n2317 = ~x129 & n916 ;
  assign n2318 = ~x129 & n918 ;
  assign n2319 = ~n2317 & ~n2318 ;
  assign n2320 = n2316 & n2319 ;
  assign n2321 = n147 & ~n2320 ;
  assign n2322 = x129 & n898 ;
  assign n2323 = x129 & n900 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = ~x129 & n928 ;
  assign n2326 = ~x129 & n930 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = n2324 & n2327 ;
  assign n2329 = n160 & ~n2328 ;
  assign n2330 = ~n2321 & ~n2329 ;
  assign n2331 = n2313 & n2330 ;
  assign n2332 = n191 & ~n2331 ;
  assign n2333 = x129 & n858 ;
  assign n2334 = x129 & n860 ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = ~x129 & n786 ;
  assign n2337 = ~x129 & n788 ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = n2335 & n2338 ;
  assign n2340 = n174 & ~n2339 ;
  assign n2341 = x129 & n781 ;
  assign n2342 = x129 & n783 ;
  assign n2343 = ~n2341 & ~n2342 ;
  assign n2344 = ~x129 & n798 ;
  assign n2345 = ~x129 & n800 ;
  assign n2346 = ~n2344 & ~n2345 ;
  assign n2347 = n2343 & n2346 ;
  assign n2348 = n187 & ~n2347 ;
  assign n2349 = ~n2340 & ~n2348 ;
  assign n2350 = x129 & n818 ;
  assign n2351 = x129 & n820 ;
  assign n2352 = ~n2350 & ~n2351 ;
  assign n2353 = ~x129 & n811 ;
  assign n2354 = ~x129 & n813 ;
  assign n2355 = ~n2353 & ~n2354 ;
  assign n2356 = n2352 & n2355 ;
  assign n2357 = n147 & ~n2356 ;
  assign n2358 = x129 & n793 ;
  assign n2359 = x129 & n795 ;
  assign n2360 = ~n2358 & ~n2359 ;
  assign n2361 = ~x129 & n823 ;
  assign n2362 = ~x129 & n825 ;
  assign n2363 = ~n2361 & ~n2362 ;
  assign n2364 = n2360 & n2363 ;
  assign n2365 = n160 & ~n2364 ;
  assign n2366 = ~n2357 & ~n2365 ;
  assign n2367 = n2349 & n2366 ;
  assign n2368 = n298 & ~n2367 ;
  assign n2369 = ~n2332 & ~n2368 ;
  assign n2370 = x129 & n911 ;
  assign n2371 = x129 & n913 ;
  assign n2372 = ~n2370 & ~n2371 ;
  assign n2373 = ~x129 & n943 ;
  assign n2374 = ~x129 & n945 ;
  assign n2375 = ~n2373 & ~n2374 ;
  assign n2376 = n2372 & n2375 ;
  assign n2377 = n174 & ~n2376 ;
  assign n2378 = ~x129 & n957 ;
  assign n2379 = ~x129 & n955 ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = x129 & n940 ;
  assign n2382 = x129 & n938 ;
  assign n2383 = ~n2381 & ~n2382 ;
  assign n2384 = n2380 & n2383 ;
  assign n2385 = n187 & ~n2384 ;
  assign n2386 = ~n2377 & ~n2385 ;
  assign n2387 = x129 & n977 ;
  assign n2388 = x129 & n982 ;
  assign n2389 = ~n2387 & ~n2388 ;
  assign n2390 = ~x129 & n968 ;
  assign n2391 = ~x129 & n970 ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = n2389 & n2392 ;
  assign n2394 = n147 & ~n2393 ;
  assign n2395 = x129 & n950 ;
  assign n2396 = x129 & n952 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = ~x129 & n980 ;
  assign n2399 = ~x129 & n975 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = n2397 & n2400 ;
  assign n2402 = n160 & ~n2401 ;
  assign n2403 = ~n2394 & ~n2402 ;
  assign n2404 = n2386 & n2403 ;
  assign n2405 = n244 & ~n2404 ;
  assign n2406 = x129 & n963 ;
  assign n2407 = x129 & n965 ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = ~x129 & n838 ;
  assign n2410 = ~x129 & n840 ;
  assign n2411 = ~n2409 & ~n2410 ;
  assign n2412 = n2408 & n2411 ;
  assign n2413 = n174 & ~n2412 ;
  assign n2414 = x129 & n833 ;
  assign n2415 = x129 & n835 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = ~x129 & n850 ;
  assign n2418 = ~x129 & n852 ;
  assign n2419 = ~n2417 & ~n2418 ;
  assign n2420 = n2416 & n2419 ;
  assign n2421 = n187 & ~n2420 ;
  assign n2422 = ~n2413 & ~n2421 ;
  assign n2423 = x129 & n870 ;
  assign n2424 = x129 & n872 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = ~x129 & n863 ;
  assign n2427 = ~x129 & n865 ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign n2429 = n2425 & n2428 ;
  assign n2430 = n147 & ~n2429 ;
  assign n2431 = x129 & n845 ;
  assign n2432 = x129 & n847 ;
  assign n2433 = ~n2431 & ~n2432 ;
  assign n2434 = ~x129 & n875 ;
  assign n2435 = ~x129 & n877 ;
  assign n2436 = ~n2434 & ~n2435 ;
  assign n2437 = n2433 & n2436 ;
  assign n2438 = n160 & ~n2437 ;
  assign n2439 = ~n2430 & ~n2438 ;
  assign n2440 = n2422 & n2439 ;
  assign n2441 = n351 & ~n2440 ;
  assign n2442 = ~n2405 & ~n2441 ;
  assign n2443 = n2369 & n2442 ;
  assign n2444 = ~x134 & ~n2443 ;
  assign n2445 = ~n2296 & ~n2444 ;
  assign n2448 = n2445 & ~x137 ;
  assign n2449 = ~n2447 & ~n2448 ;
  assign n2450 = x129 & n1155 ;
  assign n2451 = ~x129 & n1130 ;
  assign n2452 = ~n2450 & ~n2451 ;
  assign n2453 = x129 & n1160 ;
  assign n2454 = ~x129 & n1135 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2456 = n2452 & n2455 ;
  assign n2457 = n147 & ~n2456 ;
  assign n2458 = x129 & n1167 ;
  assign n2459 = ~x129 & n1157 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = x129 & n1172 ;
  assign n2462 = ~x129 & n1162 ;
  assign n2463 = ~n2461 & ~n2462 ;
  assign n2464 = n2460 & n2463 ;
  assign n2465 = n160 & ~n2464 ;
  assign n2466 = ~n2457 & ~n2465 ;
  assign n2467 = x129 & n1180 ;
  assign n2468 = ~x129 & n1194 ;
  assign n2469 = ~n2467 & ~n2468 ;
  assign n2470 = x129 & n1185 ;
  assign n2471 = ~x129 & n1199 ;
  assign n2472 = ~n2470 & ~n2471 ;
  assign n2473 = n2469 & n2472 ;
  assign n2474 = n174 & ~n2473 ;
  assign n2475 = x129 & n1192 ;
  assign n2476 = ~x129 & n1169 ;
  assign n2477 = ~n2475 & ~n2476 ;
  assign n2478 = x129 & n1197 ;
  assign n2479 = ~x129 & n1174 ;
  assign n2480 = ~n2478 & ~n2479 ;
  assign n2481 = n2477 & n2480 ;
  assign n2482 = n187 & ~n2481 ;
  assign n2483 = ~n2474 & ~n2482 ;
  assign n2484 = n2466 & n2483 ;
  assign n2485 = n351 & ~n2484 ;
  assign n2486 = x129 & n1050 ;
  assign n2487 = ~x129 & n1182 ;
  assign n2488 = ~n2486 & ~n2487 ;
  assign n2489 = x129 & n1055 ;
  assign n2490 = ~x129 & n1187 ;
  assign n2491 = ~n2489 & ~n2490 ;
  assign n2492 = n2488 & n2491 ;
  assign n2493 = n147 & ~n2492 ;
  assign n2494 = x129 & n1062 ;
  assign n2495 = ~x129 & n1052 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = x129 & n1067 ;
  assign n2498 = ~x129 & n1057 ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = n2496 & n2499 ;
  assign n2501 = n160 & ~n2500 ;
  assign n2502 = ~n2493 & ~n2501 ;
  assign n2503 = x129 & n1075 ;
  assign n2504 = ~x129 & n1089 ;
  assign n2505 = ~n2503 & ~n2504 ;
  assign n2506 = x129 & n1080 ;
  assign n2507 = ~x129 & n1094 ;
  assign n2508 = ~n2506 & ~n2507 ;
  assign n2509 = n2505 & n2508 ;
  assign n2510 = n174 & ~n2509 ;
  assign n2511 = x129 & n1087 ;
  assign n2512 = ~x129 & n1064 ;
  assign n2513 = ~n2511 & ~n2512 ;
  assign n2514 = x129 & n1092 ;
  assign n2515 = ~x129 & n1069 ;
  assign n2516 = ~n2514 & ~n2515 ;
  assign n2517 = n2513 & n2516 ;
  assign n2518 = n187 & ~n2517 ;
  assign n2519 = ~n2510 & ~n2518 ;
  assign n2520 = n2502 & n2519 ;
  assign n2521 = n244 & ~n2520 ;
  assign n2522 = ~n2485 & ~n2521 ;
  assign n2523 = x129 & n1103 ;
  assign n2524 = ~x129 & n1289 ;
  assign n2525 = ~n2523 & ~n2524 ;
  assign n2526 = x129 & n1108 ;
  assign n2527 = ~x129 & n1294 ;
  assign n2528 = ~n2526 & ~n2527 ;
  assign n2529 = n2525 & n2528 ;
  assign n2530 = n147 & ~n2529 ;
  assign n2531 = x129 & n1115 ;
  assign n2532 = ~x129 & n1105 ;
  assign n2533 = ~n2531 & ~n2532 ;
  assign n2534 = x129 & n1120 ;
  assign n2535 = ~x129 & n1110 ;
  assign n2536 = ~n2534 & ~n2535 ;
  assign n2537 = n2533 & n2536 ;
  assign n2538 = n160 & ~n2537 ;
  assign n2539 = ~n2530 & ~n2538 ;
  assign n2540 = x129 & n1128 ;
  assign n2541 = ~x129 & n1142 ;
  assign n2542 = ~n2540 & ~n2541 ;
  assign n2543 = x129 & n1133 ;
  assign n2544 = ~x129 & n1147 ;
  assign n2545 = ~n2543 & ~n2544 ;
  assign n2546 = n2542 & n2545 ;
  assign n2547 = n174 & ~n2546 ;
  assign n2548 = x129 & n1140 ;
  assign n2549 = ~x129 & n1117 ;
  assign n2550 = ~n2548 & ~n2549 ;
  assign n2551 = x129 & n1145 ;
  assign n2552 = ~x129 & n1122 ;
  assign n2553 = ~n2551 & ~n2552 ;
  assign n2554 = n2550 & n2553 ;
  assign n2555 = n187 & ~n2554 ;
  assign n2556 = ~n2547 & ~n2555 ;
  assign n2557 = n2539 & n2556 ;
  assign n2558 = n298 & ~n2557 ;
  assign n2559 = x129 & n998 ;
  assign n2560 = ~x129 & n1077 ;
  assign n2561 = ~n2559 & ~n2560 ;
  assign n2562 = x129 & n1003 ;
  assign n2563 = ~x129 & n1082 ;
  assign n2564 = ~n2562 & ~n2563 ;
  assign n2565 = n2561 & n2564 ;
  assign n2566 = n147 & ~n2565 ;
  assign n2567 = x129 & n1010 ;
  assign n2568 = ~x129 & n1000 ;
  assign n2569 = ~n2567 & ~n2568 ;
  assign n2570 = x129 & n1015 ;
  assign n2571 = ~x129 & n1005 ;
  assign n2572 = ~n2570 & ~n2571 ;
  assign n2573 = n2569 & n2572 ;
  assign n2574 = n160 & ~n2573 ;
  assign n2575 = ~n2566 & ~n2574 ;
  assign n2576 = x129 & n1023 ;
  assign n2577 = ~x129 & n1037 ;
  assign n2578 = ~n2576 & ~n2577 ;
  assign n2579 = x129 & n1028 ;
  assign n2580 = ~x129 & n1042 ;
  assign n2581 = ~n2579 & ~n2580 ;
  assign n2582 = n2578 & n2581 ;
  assign n2583 = n174 & ~n2582 ;
  assign n2584 = x129 & n1035 ;
  assign n2585 = ~x129 & n1012 ;
  assign n2586 = ~n2584 & ~n2585 ;
  assign n2587 = x129 & n1040 ;
  assign n2588 = ~x129 & n1017 ;
  assign n2589 = ~n2587 & ~n2588 ;
  assign n2590 = n2586 & n2589 ;
  assign n2591 = n187 & ~n2590 ;
  assign n2592 = ~n2583 & ~n2591 ;
  assign n2593 = n2575 & n2592 ;
  assign n2594 = n191 & ~n2593 ;
  assign n2595 = ~n2558 & ~n2594 ;
  assign n2596 = n2522 & n2595 ;
  assign n2597 = ~x134 & ~n2596 ;
  assign n2598 = x129 & n1210 ;
  assign n2599 = ~x129 & n1025 ;
  assign n2600 = ~n2598 & ~n2599 ;
  assign n2601 = x129 & n1215 ;
  assign n2602 = ~x129 & n1030 ;
  assign n2603 = ~n2601 & ~n2602 ;
  assign n2604 = n2600 & n2603 ;
  assign n2605 = n147 & ~n2604 ;
  assign n2606 = x129 & n1222 ;
  assign n2607 = ~x129 & n1212 ;
  assign n2608 = ~n2606 & ~n2607 ;
  assign n2609 = x129 & n1227 ;
  assign n2610 = ~x129 & n1217 ;
  assign n2611 = ~n2609 & ~n2610 ;
  assign n2612 = n2608 & n2611 ;
  assign n2613 = n160 & ~n2612 ;
  assign n2614 = ~n2605 & ~n2613 ;
  assign n2615 = x129 & n1235 ;
  assign n2616 = ~x129 & n1249 ;
  assign n2617 = ~n2615 & ~n2616 ;
  assign n2618 = x129 & n1240 ;
  assign n2619 = ~x129 & n1254 ;
  assign n2620 = ~n2618 & ~n2619 ;
  assign n2621 = n2617 & n2620 ;
  assign n2622 = n174 & ~n2621 ;
  assign n2623 = x129 & n1247 ;
  assign n2624 = ~x129 & n1224 ;
  assign n2625 = ~n2623 & ~n2624 ;
  assign n2626 = x129 & n1252 ;
  assign n2627 = ~x129 & n1229 ;
  assign n2628 = ~n2626 & ~n2627 ;
  assign n2629 = n2625 & n2628 ;
  assign n2630 = n187 & ~n2629 ;
  assign n2631 = ~n2622 & ~n2630 ;
  assign n2632 = n2614 & n2631 ;
  assign n2633 = n298 & ~n2632 ;
  assign n2634 = x129 & n1315 ;
  assign n2635 = ~x129 & n1237 ;
  assign n2636 = ~n2634 & ~n2635 ;
  assign n2637 = x129 & n1320 ;
  assign n2638 = ~x129 & n1242 ;
  assign n2639 = ~n2637 & ~n2638 ;
  assign n2640 = n2636 & n2639 ;
  assign n2641 = n147 & ~n2640 ;
  assign n2642 = x129 & n1334 ;
  assign n2643 = x129 & n1332 ;
  assign n2644 = ~n2642 & ~n2643 ;
  assign n2645 = ~x129 & n1322 ;
  assign n2646 = ~x129 & n1317 ;
  assign n2647 = ~n2645 & ~n2646 ;
  assign n2648 = n2644 & n2647 ;
  assign n2649 = n160 & ~n2648 ;
  assign n2650 = ~n2641 & ~n2649 ;
  assign n2651 = x129 & n1340 ;
  assign n2652 = ~x129 & n1359 ;
  assign n2653 = ~n2651 & ~n2652 ;
  assign n2654 = x129 & n1345 ;
  assign n2655 = ~x129 & n1357 ;
  assign n2656 = ~n2654 & ~n2655 ;
  assign n2657 = n2653 & n2656 ;
  assign n2658 = n174 & ~n2657 ;
  assign n2659 = x129 & n1352 ;
  assign n2660 = ~x129 & n1327 ;
  assign n2661 = ~n2659 & ~n2660 ;
  assign n2662 = x129 & n1354 ;
  assign n2663 = ~x129 & n1329 ;
  assign n2664 = ~n2662 & ~n2663 ;
  assign n2665 = n2661 & n2664 ;
  assign n2666 = n187 & ~n2665 ;
  assign n2667 = ~n2658 & ~n2666 ;
  assign n2668 = n2650 & n2667 ;
  assign n2669 = n351 & ~n2668 ;
  assign n2670 = ~n2633 & ~n2669 ;
  assign n2671 = x129 & n1262 ;
  assign n2672 = ~x129 & n1394 ;
  assign n2673 = ~n2671 & ~n2672 ;
  assign n2674 = x129 & n1267 ;
  assign n2675 = ~x129 & n1399 ;
  assign n2676 = ~n2674 & ~n2675 ;
  assign n2677 = n2673 & n2676 ;
  assign n2678 = n147 & ~n2677 ;
  assign n2679 = x129 & n1274 ;
  assign n2680 = ~x129 & n1264 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = x129 & n1279 ;
  assign n2683 = ~x129 & n1269 ;
  assign n2684 = ~n2682 & ~n2683 ;
  assign n2685 = n2681 & n2684 ;
  assign n2686 = n160 & ~n2685 ;
  assign n2687 = ~n2678 & ~n2686 ;
  assign n2688 = x129 & n1287 ;
  assign n2689 = ~x129 & n1301 ;
  assign n2690 = ~n2688 & ~n2689 ;
  assign n2691 = x129 & n1292 ;
  assign n2692 = ~x129 & n1306 ;
  assign n2693 = ~n2691 & ~n2692 ;
  assign n2694 = n2690 & n2693 ;
  assign n2695 = n174 & ~n2694 ;
  assign n2696 = x129 & n1299 ;
  assign n2697 = ~x129 & n1276 ;
  assign n2698 = ~n2696 & ~n2697 ;
  assign n2699 = x129 & n1304 ;
  assign n2700 = ~x129 & n1281 ;
  assign n2701 = ~n2699 & ~n2700 ;
  assign n2702 = n2698 & n2701 ;
  assign n2703 = n187 & ~n2702 ;
  assign n2704 = ~n2695 & ~n2703 ;
  assign n2705 = n2687 & n2704 ;
  assign n2706 = n191 & ~n2705 ;
  assign n2707 = x129 & n1367 ;
  assign n2708 = ~x129 & n1342 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = x129 & n1372 ;
  assign n2711 = ~x129 & n1347 ;
  assign n2712 = ~n2710 & ~n2711 ;
  assign n2713 = n2709 & n2712 ;
  assign n2714 = n147 & ~n2713 ;
  assign n2715 = x129 & n1379 ;
  assign n2716 = ~x129 & n1369 ;
  assign n2717 = ~n2715 & ~n2716 ;
  assign n2718 = x129 & n1384 ;
  assign n2719 = ~x129 & n1374 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2721 = n2717 & n2720 ;
  assign n2722 = n160 & ~n2721 ;
  assign n2723 = ~n2714 & ~n2722 ;
  assign n2724 = x129 & n1392 ;
  assign n2725 = ~x129 & n1406 ;
  assign n2726 = ~n2724 & ~n2725 ;
  assign n2727 = x129 & n1397 ;
  assign n2728 = ~x129 & n1411 ;
  assign n2729 = ~n2727 & ~n2728 ;
  assign n2730 = n2726 & n2729 ;
  assign n2731 = n174 & ~n2730 ;
  assign n2732 = x129 & n1404 ;
  assign n2733 = ~x129 & n1381 ;
  assign n2734 = ~n2732 & ~n2733 ;
  assign n2735 = x129 & n1409 ;
  assign n2736 = ~x129 & n1386 ;
  assign n2737 = ~n2735 & ~n2736 ;
  assign n2738 = n2734 & n2737 ;
  assign n2739 = n187 & ~n2738 ;
  assign n2740 = ~n2731 & ~n2739 ;
  assign n2741 = n2723 & n2740 ;
  assign n2742 = n244 & ~n2741 ;
  assign n2743 = ~n2706 & ~n2742 ;
  assign n2744 = n2670 & n2743 ;
  assign n2745 = x134 & ~n2744 ;
  assign n2746 = ~n2597 & ~n2745 ;
  assign n3045 = ~n2746 & x138 ;
  assign n2747 = ~x129 & n1580 ;
  assign n2748 = x129 & n1555 ;
  assign n2749 = ~n2747 & ~n2748 ;
  assign n2750 = ~x129 & n1585 ;
  assign n2751 = x129 & n1560 ;
  assign n2752 = ~n2750 & ~n2751 ;
  assign n2753 = n2749 & n2752 ;
  assign n2754 = n174 & ~n2753 ;
  assign n2755 = ~x129 & n1592 ;
  assign n2756 = x129 & n1582 ;
  assign n2757 = ~n2755 & ~n2756 ;
  assign n2758 = ~x129 & n1597 ;
  assign n2759 = x129 & n1587 ;
  assign n2760 = ~n2758 & ~n2759 ;
  assign n2761 = n2757 & n2760 ;
  assign n2762 = n187 & ~n2761 ;
  assign n2763 = ~n2754 & ~n2762 ;
  assign n2764 = ~x129 & n1605 ;
  assign n2765 = x129 & n1619 ;
  assign n2766 = ~n2764 & ~n2765 ;
  assign n2767 = ~x129 & n1610 ;
  assign n2768 = x129 & n1624 ;
  assign n2769 = ~n2767 & ~n2768 ;
  assign n2770 = n2766 & n2769 ;
  assign n2771 = n147 & ~n2770 ;
  assign n2772 = ~x129 & n1617 ;
  assign n2773 = x129 & n1594 ;
  assign n2774 = ~n2772 & ~n2773 ;
  assign n2775 = ~x129 & n1622 ;
  assign n2776 = x129 & n1599 ;
  assign n2777 = ~n2775 & ~n2776 ;
  assign n2778 = n2774 & n2777 ;
  assign n2779 = n160 & ~n2778 ;
  assign n2780 = ~n2771 & ~n2779 ;
  assign n2781 = n2763 & n2780 ;
  assign n2782 = n244 & ~n2781 ;
  assign n2783 = ~x129 & n1475 ;
  assign n2784 = x129 & n1607 ;
  assign n2785 = ~n2783 & ~n2784 ;
  assign n2786 = ~x129 & n1480 ;
  assign n2787 = x129 & n1612 ;
  assign n2788 = ~n2786 & ~n2787 ;
  assign n2789 = n2785 & n2788 ;
  assign n2790 = n174 & ~n2789 ;
  assign n2791 = ~x129 & n1487 ;
  assign n2792 = x129 & n1477 ;
  assign n2793 = ~n2791 & ~n2792 ;
  assign n2794 = ~x129 & n1492 ;
  assign n2795 = x129 & n1482 ;
  assign n2796 = ~n2794 & ~n2795 ;
  assign n2797 = n2793 & n2796 ;
  assign n2798 = n187 & ~n2797 ;
  assign n2799 = ~n2790 & ~n2798 ;
  assign n2800 = ~x129 & n1500 ;
  assign n2801 = x129 & n1514 ;
  assign n2802 = ~n2800 & ~n2801 ;
  assign n2803 = ~x129 & n1505 ;
  assign n2804 = x129 & n1519 ;
  assign n2805 = ~n2803 & ~n2804 ;
  assign n2806 = n2802 & n2805 ;
  assign n2807 = n147 & ~n2806 ;
  assign n2808 = ~x129 & n1512 ;
  assign n2809 = x129 & n1489 ;
  assign n2810 = ~n2808 & ~n2809 ;
  assign n2811 = ~x129 & n1517 ;
  assign n2812 = x129 & n1494 ;
  assign n2813 = ~n2811 & ~n2812 ;
  assign n2814 = n2810 & n2813 ;
  assign n2815 = n160 & ~n2814 ;
  assign n2816 = ~n2807 & ~n2815 ;
  assign n2817 = n2799 & n2816 ;
  assign n2818 = n351 & ~n2817 ;
  assign n2819 = ~n2782 & ~n2818 ;
  assign n2820 = ~x129 & n1528 ;
  assign n2821 = x129 & n1714 ;
  assign n2822 = ~n2820 & ~n2821 ;
  assign n2823 = ~x129 & n1533 ;
  assign n2824 = x129 & n1719 ;
  assign n2825 = ~n2823 & ~n2824 ;
  assign n2826 = n2822 & n2825 ;
  assign n2827 = n174 & ~n2826 ;
  assign n2828 = ~x129 & n1540 ;
  assign n2829 = x129 & n1530 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = ~x129 & n1545 ;
  assign n2832 = x129 & n1535 ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2834 = n2830 & n2833 ;
  assign n2835 = n187 & ~n2834 ;
  assign n2836 = ~n2827 & ~n2835 ;
  assign n2837 = ~x129 & n1553 ;
  assign n2838 = x129 & n1567 ;
  assign n2839 = ~n2837 & ~n2838 ;
  assign n2840 = ~x129 & n1558 ;
  assign n2841 = x129 & n1572 ;
  assign n2842 = ~n2840 & ~n2841 ;
  assign n2843 = n2839 & n2842 ;
  assign n2844 = n147 & ~n2843 ;
  assign n2845 = ~x129 & n1565 ;
  assign n2846 = x129 & n1542 ;
  assign n2847 = ~n2845 & ~n2846 ;
  assign n2848 = ~x129 & n1570 ;
  assign n2849 = x129 & n1547 ;
  assign n2850 = ~n2848 & ~n2849 ;
  assign n2851 = n2847 & n2850 ;
  assign n2852 = n160 & ~n2851 ;
  assign n2853 = ~n2844 & ~n2852 ;
  assign n2854 = n2836 & n2853 ;
  assign n2855 = n191 & ~n2854 ;
  assign n2856 = ~x129 & n1423 ;
  assign n2857 = x129 & n1502 ;
  assign n2858 = ~n2856 & ~n2857 ;
  assign n2859 = ~x129 & n1428 ;
  assign n2860 = x129 & n1507 ;
  assign n2861 = ~n2859 & ~n2860 ;
  assign n2862 = n2858 & n2861 ;
  assign n2863 = n174 & ~n2862 ;
  assign n2864 = ~x129 & n1435 ;
  assign n2865 = x129 & n1425 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = ~x129 & n1440 ;
  assign n2868 = x129 & n1430 ;
  assign n2869 = ~n2867 & ~n2868 ;
  assign n2870 = n2866 & n2869 ;
  assign n2871 = n187 & ~n2870 ;
  assign n2872 = ~n2863 & ~n2871 ;
  assign n2873 = ~x129 & n1448 ;
  assign n2874 = x129 & n1462 ;
  assign n2875 = ~n2873 & ~n2874 ;
  assign n2876 = ~x129 & n1453 ;
  assign n2877 = x129 & n1467 ;
  assign n2878 = ~n2876 & ~n2877 ;
  assign n2879 = n2875 & n2878 ;
  assign n2880 = n147 & ~n2879 ;
  assign n2881 = ~x129 & n1460 ;
  assign n2882 = x129 & n1437 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = ~x129 & n1465 ;
  assign n2885 = x129 & n1442 ;
  assign n2886 = ~n2884 & ~n2885 ;
  assign n2887 = n2883 & n2886 ;
  assign n2888 = n160 & ~n2887 ;
  assign n2889 = ~n2880 & ~n2888 ;
  assign n2890 = n2872 & n2889 ;
  assign n2891 = n298 & ~n2890 ;
  assign n2892 = ~n2855 & ~n2891 ;
  assign n2893 = n2819 & n2892 ;
  assign n2894 = x134 & ~n2893 ;
  assign n2895 = ~x129 & n1635 ;
  assign n2896 = x129 & n1450 ;
  assign n2897 = ~n2895 & ~n2896 ;
  assign n2898 = ~x129 & n1640 ;
  assign n2899 = x129 & n1455 ;
  assign n2900 = ~n2898 & ~n2899 ;
  assign n2901 = n2897 & n2900 ;
  assign n2902 = n174 & ~n2901 ;
  assign n2903 = ~x129 & n1647 ;
  assign n2904 = x129 & n1637 ;
  assign n2905 = ~n2903 & ~n2904 ;
  assign n2906 = ~x129 & n1652 ;
  assign n2907 = x129 & n1642 ;
  assign n2908 = ~n2906 & ~n2907 ;
  assign n2909 = n2905 & n2908 ;
  assign n2910 = n187 & ~n2909 ;
  assign n2911 = ~n2902 & ~n2910 ;
  assign n2912 = ~x129 & n1660 ;
  assign n2913 = x129 & n1674 ;
  assign n2914 = ~n2912 & ~n2913 ;
  assign n2915 = ~x129 & n1665 ;
  assign n2916 = x129 & n1679 ;
  assign n2917 = ~n2915 & ~n2916 ;
  assign n2918 = n2914 & n2917 ;
  assign n2919 = n147 & ~n2918 ;
  assign n2920 = ~x129 & n1672 ;
  assign n2921 = x129 & n1649 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~x129 & n1677 ;
  assign n2924 = x129 & n1654 ;
  assign n2925 = ~n2923 & ~n2924 ;
  assign n2926 = n2922 & n2925 ;
  assign n2927 = n160 & ~n2926 ;
  assign n2928 = ~n2919 & ~n2927 ;
  assign n2929 = n2911 & n2928 ;
  assign n2930 = n191 & ~n2929 ;
  assign n2931 = ~x129 & n1740 ;
  assign n2932 = x129 & n1662 ;
  assign n2933 = ~n2931 & ~n2932 ;
  assign n2934 = ~x129 & n1745 ;
  assign n2935 = x129 & n1667 ;
  assign n2936 = ~n2934 & ~n2935 ;
  assign n2937 = n2933 & n2936 ;
  assign n2938 = n174 & ~n2937 ;
  assign n2939 = ~x129 & n1759 ;
  assign n2940 = ~x129 & n1757 ;
  assign n2941 = ~n2939 & ~n2940 ;
  assign n2942 = x129 & n1747 ;
  assign n2943 = x129 & n1742 ;
  assign n2944 = ~n2942 & ~n2943 ;
  assign n2945 = n2941 & n2944 ;
  assign n2946 = n187 & ~n2945 ;
  assign n2947 = ~n2938 & ~n2946 ;
  assign n2948 = ~x129 & n1765 ;
  assign n2949 = x129 & n1784 ;
  assign n2950 = ~n2948 & ~n2949 ;
  assign n2951 = ~x129 & n1770 ;
  assign n2952 = x129 & n1782 ;
  assign n2953 = ~n2951 & ~n2952 ;
  assign n2954 = n2950 & n2953 ;
  assign n2955 = n147 & ~n2954 ;
  assign n2956 = ~x129 & n1777 ;
  assign n2957 = x129 & n1752 ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = ~x129 & n1779 ;
  assign n2960 = x129 & n1754 ;
  assign n2961 = ~n2959 & ~n2960 ;
  assign n2962 = n2958 & n2961 ;
  assign n2963 = n160 & ~n2962 ;
  assign n2964 = ~n2955 & ~n2963 ;
  assign n2965 = n2947 & n2964 ;
  assign n2966 = n244 & ~n2965 ;
  assign n2967 = ~n2930 & ~n2966 ;
  assign n2968 = ~x129 & n1687 ;
  assign n2969 = x129 & n1819 ;
  assign n2970 = ~n2968 & ~n2969 ;
  assign n2971 = ~x129 & n1692 ;
  assign n2972 = x129 & n1824 ;
  assign n2973 = ~n2971 & ~n2972 ;
  assign n2974 = n2970 & n2973 ;
  assign n2975 = n174 & ~n2974 ;
  assign n2976 = ~x129 & n1699 ;
  assign n2977 = x129 & n1689 ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = ~x129 & n1704 ;
  assign n2980 = x129 & n1694 ;
  assign n2981 = ~n2979 & ~n2980 ;
  assign n2982 = n2978 & n2981 ;
  assign n2983 = n187 & ~n2982 ;
  assign n2984 = ~n2975 & ~n2983 ;
  assign n2985 = ~x129 & n1712 ;
  assign n2986 = x129 & n1726 ;
  assign n2987 = ~n2985 & ~n2986 ;
  assign n2988 = ~x129 & n1717 ;
  assign n2989 = x129 & n1731 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = n2987 & n2990 ;
  assign n2992 = n147 & ~n2991 ;
  assign n2993 = ~x129 & n1724 ;
  assign n2994 = x129 & n1701 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = ~x129 & n1729 ;
  assign n2997 = x129 & n1706 ;
  assign n2998 = ~n2996 & ~n2997 ;
  assign n2999 = n2995 & n2998 ;
  assign n3000 = n160 & ~n2999 ;
  assign n3001 = ~n2992 & ~n3000 ;
  assign n3002 = n2984 & n3001 ;
  assign n3003 = n298 & ~n3002 ;
  assign n3004 = ~x129 & n1792 ;
  assign n3005 = x129 & n1767 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = ~x129 & n1797 ;
  assign n3008 = x129 & n1772 ;
  assign n3009 = ~n3007 & ~n3008 ;
  assign n3010 = n3006 & n3009 ;
  assign n3011 = n174 & ~n3010 ;
  assign n3012 = ~x129 & n1804 ;
  assign n3013 = x129 & n1794 ;
  assign n3014 = ~n3012 & ~n3013 ;
  assign n3015 = ~x129 & n1809 ;
  assign n3016 = x129 & n1799 ;
  assign n3017 = ~n3015 & ~n3016 ;
  assign n3018 = n3014 & n3017 ;
  assign n3019 = n187 & ~n3018 ;
  assign n3020 = ~n3011 & ~n3019 ;
  assign n3021 = ~x129 & n1817 ;
  assign n3022 = x129 & n1831 ;
  assign n3023 = ~n3021 & ~n3022 ;
  assign n3024 = ~x129 & n1822 ;
  assign n3025 = x129 & n1836 ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = n3023 & n3026 ;
  assign n3028 = n147 & ~n3027 ;
  assign n3029 = ~x129 & n1829 ;
  assign n3030 = x129 & n1806 ;
  assign n3031 = ~n3029 & ~n3030 ;
  assign n3032 = ~x129 & n1834 ;
  assign n3033 = x129 & n1811 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = n3031 & n3034 ;
  assign n3036 = n160 & ~n3035 ;
  assign n3037 = ~n3028 & ~n3036 ;
  assign n3038 = n3020 & n3037 ;
  assign n3039 = n351 & ~n3038 ;
  assign n3040 = ~n3003 & ~n3039 ;
  assign n3041 = n2967 & n3040 ;
  assign n3042 = ~x134 & ~n3041 ;
  assign n3043 = ~n2894 & ~n3042 ;
  assign n3046 = n3043 & ~x138 ;
  assign n3047 = ~n3045 & ~n3046 ;
  assign n3048 = n147 & ~n228 ;
  assign n3049 = ~n146 & n160 ;
  assign n3050 = ~n3048 & ~n3049 ;
  assign n3051 = n174 & ~n186 ;
  assign n3052 = ~n159 & n187 ;
  assign n3053 = ~n3051 & ~n3052 ;
  assign n3054 = n3050 & n3053 ;
  assign n3055 = n191 & ~n3054 ;
  assign n3056 = n147 & ~n335 ;
  assign n3057 = n160 & ~n203 ;
  assign n3058 = ~n3056 & ~n3057 ;
  assign n3059 = n174 & ~n240 ;
  assign n3060 = n187 & ~n215 ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3062 = n3058 & n3061 ;
  assign n3063 = n244 & ~n3062 ;
  assign n3064 = ~n3055 & ~n3063 ;
  assign n3065 = n147 & ~n391 ;
  assign n3066 = n160 & ~n257 ;
  assign n3067 = ~n3065 & ~n3066 ;
  assign n3068 = n174 & ~n294 ;
  assign n3069 = n187 & ~n269 ;
  assign n3070 = ~n3068 & ~n3069 ;
  assign n3071 = n3067 & n3070 ;
  assign n3072 = n298 & ~n3071 ;
  assign n3073 = n147 & ~n282 ;
  assign n3074 = n160 & ~n310 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = n174 & ~n347 ;
  assign n3077 = n187 & ~n322 ;
  assign n3078 = ~n3076 & ~n3077 ;
  assign n3079 = n3075 & n3078 ;
  assign n3080 = n351 & ~n3079 ;
  assign n3081 = ~n3072 & ~n3080 ;
  assign n3082 = n3064 & n3081 ;
  assign n3083 = ~x134 & ~n3082 ;
  assign n3084 = n147 & ~n496 ;
  assign n3085 = n160 & ~n523 ;
  assign n3086 = ~n3084 & ~n3085 ;
  assign n3087 = n174 & ~n560 ;
  assign n3088 = n187 & ~n535 ;
  assign n3089 = ~n3087 & ~n3088 ;
  assign n3090 = n3086 & n3089 ;
  assign n3091 = n351 & ~n3090 ;
  assign n3092 = n147 & ~n173 ;
  assign n3093 = n160 & ~n471 ;
  assign n3094 = ~n3092 & ~n3093 ;
  assign n3095 = n174 & ~n508 ;
  assign n3096 = n187 & ~n483 ;
  assign n3097 = ~n3095 & ~n3096 ;
  assign n3098 = n3094 & n3097 ;
  assign n3099 = n298 & ~n3098 ;
  assign n3100 = ~n3091 & ~n3099 ;
  assign n3101 = n147 & ~n548 ;
  assign n3102 = n160 & ~n418 ;
  assign n3103 = ~n3101 & ~n3102 ;
  assign n3104 = n174 & ~n455 ;
  assign n3105 = n187 & ~n430 ;
  assign n3106 = ~n3104 & ~n3105 ;
  assign n3107 = n3103 & n3106 ;
  assign n3108 = n244 & ~n3107 ;
  assign n3109 = n147 & ~n443 ;
  assign n3110 = n160 & ~n366 ;
  assign n3111 = ~n3109 & ~n3110 ;
  assign n3112 = n174 & ~n403 ;
  assign n3113 = n187 & ~n378 ;
  assign n3114 = ~n3112 & ~n3113 ;
  assign n3115 = n3111 & n3114 ;
  assign n3116 = n191 & ~n3115 ;
  assign n3117 = ~n3108 & ~n3116 ;
  assign n3118 = n3100 & n3117 ;
  assign n3119 = x134 & ~n3118 ;
  assign n3120 = ~n3083 & ~n3119 ;
  assign n3195 = ~n3120 & x139 ;
  assign n3121 = n174 & ~n656 ;
  assign n3122 = n187 & ~n579 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = n147 & ~n616 ;
  assign n3125 = n160 & ~n591 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = n3123 & n3126 ;
  assign n3128 = n298 & ~n3127 ;
  assign n3129 = n174 & ~n761 ;
  assign n3130 = n187 & ~n631 ;
  assign n3131 = ~n3129 & ~n3130 ;
  assign n3132 = n147 & ~n668 ;
  assign n3133 = n160 & ~n643 ;
  assign n3134 = ~n3132 & ~n3133 ;
  assign n3135 = n3131 & n3134 ;
  assign n3136 = n351 & ~n3135 ;
  assign n3137 = ~n3128 & ~n3136 ;
  assign n3138 = n174 & ~n816 ;
  assign n3139 = n187 & ~n684 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3141 = n147 & ~n721 ;
  assign n3142 = n160 & ~n696 ;
  assign n3143 = ~n3141 & ~n3142 ;
  assign n3144 = n3140 & n3143 ;
  assign n3145 = n191 & ~n3144 ;
  assign n3146 = n174 & ~n709 ;
  assign n3147 = n187 & ~n736 ;
  assign n3148 = ~n3146 & ~n3147 ;
  assign n3149 = n147 & ~n773 ;
  assign n3150 = n160 & ~n748 ;
  assign n3151 = ~n3149 & ~n3150 ;
  assign n3152 = n3148 & n3151 ;
  assign n3153 = n244 & ~n3152 ;
  assign n3154 = ~n3145 & ~n3153 ;
  assign n3155 = n3137 & n3154 ;
  assign n3156 = x134 & ~n3155 ;
  assign n3157 = n174 & ~n921 ;
  assign n3158 = n187 & ~n948 ;
  assign n3159 = ~n3157 & ~n3158 ;
  assign n3160 = n147 & ~n985 ;
  assign n3161 = n160 & ~n960 ;
  assign n3162 = ~n3160 & ~n3161 ;
  assign n3163 = n3159 & n3162 ;
  assign n3164 = n244 & ~n3163 ;
  assign n3165 = n174 & ~n604 ;
  assign n3166 = n187 & ~n896 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = n147 & ~n933 ;
  assign n3169 = n160 & ~n908 ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = n3167 & n3170 ;
  assign n3172 = n191 & ~n3171 ;
  assign n3173 = ~n3164 & ~n3172 ;
  assign n3174 = n174 & ~n973 ;
  assign n3175 = n187 & ~n843 ;
  assign n3176 = ~n3174 & ~n3175 ;
  assign n3177 = n147 & ~n880 ;
  assign n3178 = n160 & ~n855 ;
  assign n3179 = ~n3177 & ~n3178 ;
  assign n3180 = n3176 & n3179 ;
  assign n3181 = n351 & ~n3180 ;
  assign n3182 = n174 & ~n868 ;
  assign n3183 = n187 & ~n791 ;
  assign n3184 = ~n3182 & ~n3183 ;
  assign n3185 = n147 & ~n828 ;
  assign n3186 = n160 & ~n803 ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = n3184 & n3187 ;
  assign n3189 = n298 & ~n3188 ;
  assign n3190 = ~n3181 & ~n3189 ;
  assign n3191 = n3173 & n3190 ;
  assign n3192 = ~x134 & ~n3191 ;
  assign n3193 = ~n3156 & ~n3192 ;
  assign n3196 = n3193 & ~x139 ;
  assign n3197 = ~n3195 & ~n3196 ;
  assign n3198 = n147 & ~n1085 ;
  assign n3199 = n160 & ~n1008 ;
  assign n3200 = ~n3198 & ~n3199 ;
  assign n3201 = n174 & ~n1045 ;
  assign n3202 = n187 & ~n1020 ;
  assign n3203 = ~n3201 & ~n3202 ;
  assign n3204 = n3200 & n3203 ;
  assign n3205 = n191 & ~n3204 ;
  assign n3206 = n147 & ~n1190 ;
  assign n3207 = n160 & ~n1060 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = n174 & ~n1097 ;
  assign n3210 = n187 & ~n1072 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = n3208 & n3211 ;
  assign n3213 = n244 & ~n3212 ;
  assign n3214 = ~n3205 & ~n3213 ;
  assign n3215 = n147 & ~n1297 ;
  assign n3216 = n160 & ~n1113 ;
  assign n3217 = ~n3215 & ~n3216 ;
  assign n3218 = n174 & ~n1150 ;
  assign n3219 = n187 & ~n1125 ;
  assign n3220 = ~n3218 & ~n3219 ;
  assign n3221 = n3217 & n3220 ;
  assign n3222 = n298 & ~n3221 ;
  assign n3223 = n147 & ~n1138 ;
  assign n3224 = n160 & ~n1165 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = n174 & ~n1202 ;
  assign n3227 = n187 & ~n1177 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = n3225 & n3228 ;
  assign n3230 = n351 & ~n3229 ;
  assign n3231 = ~n3222 & ~n3230 ;
  assign n3232 = n3214 & n3231 ;
  assign n3233 = ~x134 & ~n3232 ;
  assign n3234 = n147 & ~n1245 ;
  assign n3235 = n160 & ~n1325 ;
  assign n3236 = ~n3234 & ~n3235 ;
  assign n3237 = n174 & ~n1362 ;
  assign n3238 = n187 & ~n1337 ;
  assign n3239 = ~n3237 & ~n3238 ;
  assign n3240 = n3236 & n3239 ;
  assign n3241 = n351 & ~n3240 ;
  assign n3242 = n147 & ~n1033 ;
  assign n3243 = n160 & ~n1220 ;
  assign n3244 = ~n3242 & ~n3243 ;
  assign n3245 = n174 & ~n1257 ;
  assign n3246 = n187 & ~n1232 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = n3244 & n3247 ;
  assign n3249 = n298 & ~n3248 ;
  assign n3250 = ~n3241 & ~n3249 ;
  assign n3251 = n147 & ~n1350 ;
  assign n3252 = n160 & ~n1377 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = n174 & ~n1414 ;
  assign n3255 = n187 & ~n1389 ;
  assign n3256 = ~n3254 & ~n3255 ;
  assign n3257 = n3253 & n3256 ;
  assign n3258 = n244 & ~n3257 ;
  assign n3259 = n147 & ~n1402 ;
  assign n3260 = n160 & ~n1272 ;
  assign n3261 = ~n3259 & ~n3260 ;
  assign n3262 = n174 & ~n1309 ;
  assign n3263 = n187 & ~n1284 ;
  assign n3264 = ~n3262 & ~n3263 ;
  assign n3265 = n3261 & n3264 ;
  assign n3266 = n191 & ~n3265 ;
  assign n3267 = ~n3258 & ~n3266 ;
  assign n3268 = n3250 & n3267 ;
  assign n3269 = x134 & ~n3268 ;
  assign n3270 = ~n3233 & ~n3269 ;
  assign n3345 = ~n3270 & x140 ;
  assign n3271 = n174 & ~n1510 ;
  assign n3272 = n187 & ~n1433 ;
  assign n3273 = ~n3271 & ~n3272 ;
  assign n3274 = n147 & ~n1470 ;
  assign n3275 = n160 & ~n1445 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign n3277 = n3273 & n3276 ;
  assign n3278 = n298 & ~n3277 ;
  assign n3279 = n174 & ~n1615 ;
  assign n3280 = n187 & ~n1485 ;
  assign n3281 = ~n3279 & ~n3280 ;
  assign n3282 = n147 & ~n1522 ;
  assign n3283 = n160 & ~n1497 ;
  assign n3284 = ~n3282 & ~n3283 ;
  assign n3285 = n3281 & n3284 ;
  assign n3286 = n351 & ~n3285 ;
  assign n3287 = ~n3278 & ~n3286 ;
  assign n3288 = n174 & ~n1722 ;
  assign n3289 = n187 & ~n1538 ;
  assign n3290 = ~n3288 & ~n3289 ;
  assign n3291 = n147 & ~n1575 ;
  assign n3292 = n160 & ~n1550 ;
  assign n3293 = ~n3291 & ~n3292 ;
  assign n3294 = n3290 & n3293 ;
  assign n3295 = n191 & ~n3294 ;
  assign n3296 = n174 & ~n1563 ;
  assign n3297 = n187 & ~n1590 ;
  assign n3298 = ~n3296 & ~n3297 ;
  assign n3299 = n147 & ~n1627 ;
  assign n3300 = n160 & ~n1602 ;
  assign n3301 = ~n3299 & ~n3300 ;
  assign n3302 = n3298 & n3301 ;
  assign n3303 = n244 & ~n3302 ;
  assign n3304 = ~n3295 & ~n3303 ;
  assign n3305 = n3287 & n3304 ;
  assign n3306 = x134 & ~n3305 ;
  assign n3307 = n174 & ~n1670 ;
  assign n3308 = n187 & ~n1750 ;
  assign n3309 = ~n3307 & ~n3308 ;
  assign n3310 = n147 & ~n1787 ;
  assign n3311 = n160 & ~n1762 ;
  assign n3312 = ~n3310 & ~n3311 ;
  assign n3313 = n3309 & n3312 ;
  assign n3314 = n244 & ~n3313 ;
  assign n3315 = n174 & ~n1458 ;
  assign n3316 = n187 & ~n1645 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = n147 & ~n1682 ;
  assign n3319 = n160 & ~n1657 ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = n3317 & n3320 ;
  assign n3322 = n191 & ~n3321 ;
  assign n3323 = ~n3314 & ~n3322 ;
  assign n3324 = n174 & ~n1775 ;
  assign n3325 = n187 & ~n1802 ;
  assign n3326 = ~n3324 & ~n3325 ;
  assign n3327 = n147 & ~n1839 ;
  assign n3328 = n160 & ~n1814 ;
  assign n3329 = ~n3327 & ~n3328 ;
  assign n3330 = n3326 & n3329 ;
  assign n3331 = n351 & ~n3330 ;
  assign n3332 = n174 & ~n1827 ;
  assign n3333 = n187 & ~n1697 ;
  assign n3334 = ~n3332 & ~n3333 ;
  assign n3335 = n147 & ~n1734 ;
  assign n3336 = n160 & ~n1709 ;
  assign n3337 = ~n3335 & ~n3336 ;
  assign n3338 = n3334 & n3337 ;
  assign n3339 = n298 & ~n3338 ;
  assign n3340 = ~n3331 & ~n3339 ;
  assign n3341 = n3323 & n3340 ;
  assign n3342 = ~x134 & ~n3341 ;
  assign n3343 = ~n3306 & ~n3342 ;
  assign n3346 = n3343 & ~x140 ;
  assign n3347 = ~n3345 & ~n3346 ;
  assign n3348 = n147 & ~n1911 ;
  assign n3349 = n160 & ~n1858 ;
  assign n3350 = ~n3348 & ~n3349 ;
  assign n3351 = n174 & ~n1883 ;
  assign n3352 = n187 & ~n1866 ;
  assign n3353 = ~n3351 & ~n3352 ;
  assign n3354 = n3350 & n3353 ;
  assign n3355 = n191 & ~n3354 ;
  assign n3356 = n147 & ~n1984 ;
  assign n3357 = n160 & ~n1894 ;
  assign n3358 = ~n3356 & ~n3357 ;
  assign n3359 = n174 & ~n1919 ;
  assign n3360 = n187 & ~n1902 ;
  assign n3361 = ~n3359 & ~n3360 ;
  assign n3362 = n3358 & n3361 ;
  assign n3363 = n244 & ~n3362 ;
  assign n3364 = ~n3355 & ~n3363 ;
  assign n3365 = n147 & ~n2059 ;
  assign n3366 = n160 & ~n1931 ;
  assign n3367 = ~n3365 & ~n3366 ;
  assign n3368 = n174 & ~n1956 ;
  assign n3369 = n187 & ~n1939 ;
  assign n3370 = ~n3368 & ~n3369 ;
  assign n3371 = n3367 & n3370 ;
  assign n3372 = n298 & ~n3371 ;
  assign n3373 = n147 & ~n1948 ;
  assign n3374 = n160 & ~n1967 ;
  assign n3375 = ~n3373 & ~n3374 ;
  assign n3376 = n174 & ~n1992 ;
  assign n3377 = n187 & ~n1975 ;
  assign n3378 = ~n3376 & ~n3377 ;
  assign n3379 = n3375 & n3378 ;
  assign n3380 = n351 & ~n3379 ;
  assign n3381 = ~n3372 & ~n3380 ;
  assign n3382 = n3364 & n3381 ;
  assign n3383 = ~x134 & ~n3382 ;
  assign n3384 = n147 & ~n2023 ;
  assign n3385 = n160 & ~n2079 ;
  assign n3386 = ~n3384 & ~n3385 ;
  assign n3387 = n174 & ~n2104 ;
  assign n3388 = n187 & ~n2087 ;
  assign n3389 = ~n3387 & ~n3388 ;
  assign n3390 = n3386 & n3389 ;
  assign n3391 = n351 & ~n3390 ;
  assign n3392 = n147 & ~n1875 ;
  assign n3393 = n160 & ~n2006 ;
  assign n3394 = ~n3392 & ~n3393 ;
  assign n3395 = n174 & ~n2031 ;
  assign n3396 = n187 & ~n2014 ;
  assign n3397 = ~n3395 & ~n3396 ;
  assign n3398 = n3394 & n3397 ;
  assign n3399 = n298 & ~n3398 ;
  assign n3400 = ~n3391 & ~n3399 ;
  assign n3401 = n147 & ~n2096 ;
  assign n3402 = n160 & ~n2115 ;
  assign n3403 = ~n3401 & ~n3402 ;
  assign n3404 = n174 & ~n2140 ;
  assign n3405 = n187 & ~n2123 ;
  assign n3406 = ~n3404 & ~n3405 ;
  assign n3407 = n3403 & n3406 ;
  assign n3408 = n244 & ~n3407 ;
  assign n3409 = n147 & ~n2132 ;
  assign n3410 = n160 & ~n2042 ;
  assign n3411 = ~n3409 & ~n3410 ;
  assign n3412 = n174 & ~n2067 ;
  assign n3413 = n187 & ~n2050 ;
  assign n3414 = ~n3412 & ~n3413 ;
  assign n3415 = n3411 & n3414 ;
  assign n3416 = n191 & ~n3415 ;
  assign n3417 = ~n3408 & ~n3416 ;
  assign n3418 = n3400 & n3417 ;
  assign n3419 = x134 & ~n3418 ;
  assign n3420 = ~n3383 & ~n3419 ;
  assign n3495 = ~n3420 & x141 ;
  assign n3421 = n174 & ~n2208 ;
  assign n3422 = n187 & ~n2155 ;
  assign n3423 = ~n3421 & ~n3422 ;
  assign n3424 = n147 & ~n2180 ;
  assign n3425 = n160 & ~n2163 ;
  assign n3426 = ~n3424 & ~n3425 ;
  assign n3427 = n3423 & n3426 ;
  assign n3428 = n298 & ~n3427 ;
  assign n3429 = n174 & ~n2281 ;
  assign n3430 = n187 & ~n2191 ;
  assign n3431 = ~n3429 & ~n3430 ;
  assign n3432 = n147 & ~n2216 ;
  assign n3433 = n160 & ~n2199 ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3435 = n3431 & n3434 ;
  assign n3436 = n351 & ~n3435 ;
  assign n3437 = ~n3428 & ~n3436 ;
  assign n3438 = n174 & ~n2356 ;
  assign n3439 = n187 & ~n2228 ;
  assign n3440 = ~n3438 & ~n3439 ;
  assign n3441 = n147 & ~n2253 ;
  assign n3442 = n160 & ~n2236 ;
  assign n3443 = ~n3441 & ~n3442 ;
  assign n3444 = n3440 & n3443 ;
  assign n3445 = n191 & ~n3444 ;
  assign n3446 = n174 & ~n2245 ;
  assign n3447 = n187 & ~n2264 ;
  assign n3448 = ~n3446 & ~n3447 ;
  assign n3449 = n147 & ~n2289 ;
  assign n3450 = n160 & ~n2272 ;
  assign n3451 = ~n3449 & ~n3450 ;
  assign n3452 = n3448 & n3451 ;
  assign n3453 = n244 & ~n3452 ;
  assign n3454 = ~n3445 & ~n3453 ;
  assign n3455 = n3437 & n3454 ;
  assign n3456 = x134 & ~n3455 ;
  assign n3457 = n174 & ~n2320 ;
  assign n3458 = n187 & ~n2376 ;
  assign n3459 = ~n3457 & ~n3458 ;
  assign n3460 = n147 & ~n2401 ;
  assign n3461 = n160 & ~n2384 ;
  assign n3462 = ~n3460 & ~n3461 ;
  assign n3463 = n3459 & n3462 ;
  assign n3464 = n244 & ~n3463 ;
  assign n3465 = n174 & ~n2172 ;
  assign n3466 = n187 & ~n2303 ;
  assign n3467 = ~n3465 & ~n3466 ;
  assign n3468 = n147 & ~n2328 ;
  assign n3469 = n160 & ~n2311 ;
  assign n3470 = ~n3468 & ~n3469 ;
  assign n3471 = n3467 & n3470 ;
  assign n3472 = n191 & ~n3471 ;
  assign n3473 = ~n3464 & ~n3472 ;
  assign n3474 = n174 & ~n2393 ;
  assign n3475 = n187 & ~n2412 ;
  assign n3476 = ~n3474 & ~n3475 ;
  assign n3477 = n147 & ~n2437 ;
  assign n3478 = n160 & ~n2420 ;
  assign n3479 = ~n3477 & ~n3478 ;
  assign n3480 = n3476 & n3479 ;
  assign n3481 = n351 & ~n3480 ;
  assign n3482 = n174 & ~n2429 ;
  assign n3483 = n187 & ~n2339 ;
  assign n3484 = ~n3482 & ~n3483 ;
  assign n3485 = n147 & ~n2364 ;
  assign n3486 = n160 & ~n2347 ;
  assign n3487 = ~n3485 & ~n3486 ;
  assign n3488 = n3484 & n3487 ;
  assign n3489 = n298 & ~n3488 ;
  assign n3490 = ~n3481 & ~n3489 ;
  assign n3491 = n3473 & n3490 ;
  assign n3492 = ~x134 & ~n3491 ;
  assign n3493 = ~n3456 & ~n3492 ;
  assign n3496 = n3493 & ~x141 ;
  assign n3497 = ~n3495 & ~n3496 ;
  assign n3498 = n147 & ~n2509 ;
  assign n3499 = n160 & ~n2565 ;
  assign n3500 = ~n3498 & ~n3499 ;
  assign n3501 = n174 & ~n2590 ;
  assign n3502 = n187 & ~n2573 ;
  assign n3503 = ~n3501 & ~n3502 ;
  assign n3504 = n3500 & n3503 ;
  assign n3505 = n191 & ~n3504 ;
  assign n3506 = n147 & ~n2473 ;
  assign n3507 = n160 & ~n2492 ;
  assign n3508 = ~n3506 & ~n3507 ;
  assign n3509 = n174 & ~n2517 ;
  assign n3510 = n187 & ~n2500 ;
  assign n3511 = ~n3509 & ~n3510 ;
  assign n3512 = n3508 & n3511 ;
  assign n3513 = n244 & ~n3512 ;
  assign n3514 = ~n3505 & ~n3513 ;
  assign n3515 = n147 & ~n2694 ;
  assign n3516 = n160 & ~n2529 ;
  assign n3517 = ~n3515 & ~n3516 ;
  assign n3518 = n174 & ~n2554 ;
  assign n3519 = n187 & ~n2537 ;
  assign n3520 = ~n3518 & ~n3519 ;
  assign n3521 = n3517 & n3520 ;
  assign n3522 = n298 & ~n3521 ;
  assign n3523 = n147 & ~n2546 ;
  assign n3524 = n160 & ~n2456 ;
  assign n3525 = ~n3523 & ~n3524 ;
  assign n3526 = n174 & ~n2481 ;
  assign n3527 = n187 & ~n2464 ;
  assign n3528 = ~n3526 & ~n3527 ;
  assign n3529 = n3525 & n3528 ;
  assign n3530 = n351 & ~n3529 ;
  assign n3531 = ~n3522 & ~n3530 ;
  assign n3532 = n3514 & n3531 ;
  assign n3533 = ~x134 & ~n3532 ;
  assign n3534 = n160 & ~n2640 ;
  assign n3535 = n187 & ~n2648 ;
  assign n3536 = ~n3534 & ~n3535 ;
  assign n3537 = n174 & ~n2665 ;
  assign n3538 = n147 & ~n2621 ;
  assign n3539 = ~n3537 & ~n3538 ;
  assign n3540 = n3536 & n3539 ;
  assign n3541 = n351 & ~n3540 ;
  assign n3542 = n147 & ~n2582 ;
  assign n3543 = n160 & ~n2604 ;
  assign n3544 = ~n3542 & ~n3543 ;
  assign n3545 = n174 & ~n2629 ;
  assign n3546 = n187 & ~n2612 ;
  assign n3547 = ~n3545 & ~n3546 ;
  assign n3548 = n3544 & n3547 ;
  assign n3549 = n298 & ~n3548 ;
  assign n3550 = ~n3541 & ~n3549 ;
  assign n3551 = n147 & ~n2657 ;
  assign n3552 = n160 & ~n2713 ;
  assign n3553 = ~n3551 & ~n3552 ;
  assign n3554 = n174 & ~n2738 ;
  assign n3555 = n187 & ~n2721 ;
  assign n3556 = ~n3554 & ~n3555 ;
  assign n3557 = n3553 & n3556 ;
  assign n3558 = n244 & ~n3557 ;
  assign n3559 = n147 & ~n2730 ;
  assign n3560 = n160 & ~n2677 ;
  assign n3561 = ~n3559 & ~n3560 ;
  assign n3562 = n174 & ~n2702 ;
  assign n3563 = n187 & ~n2685 ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = n3561 & n3564 ;
  assign n3566 = n191 & ~n3565 ;
  assign n3567 = ~n3558 & ~n3566 ;
  assign n3568 = n3550 & n3567 ;
  assign n3569 = x134 & ~n3568 ;
  assign n3570 = ~n3533 & ~n3569 ;
  assign n3645 = ~n3570 & x142 ;
  assign n3571 = n174 & ~n2806 ;
  assign n3572 = n187 & ~n2862 ;
  assign n3573 = ~n3571 & ~n3572 ;
  assign n3574 = n147 & ~n2887 ;
  assign n3575 = n160 & ~n2870 ;
  assign n3576 = ~n3574 & ~n3575 ;
  assign n3577 = n3573 & n3576 ;
  assign n3578 = n298 & ~n3577 ;
  assign n3579 = n174 & ~n2770 ;
  assign n3580 = n187 & ~n2789 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = n147 & ~n2814 ;
  assign n3583 = n160 & ~n2797 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = n3581 & n3584 ;
  assign n3586 = n351 & ~n3585 ;
  assign n3587 = ~n3578 & ~n3586 ;
  assign n3588 = n174 & ~n2991 ;
  assign n3589 = n187 & ~n2826 ;
  assign n3590 = ~n3588 & ~n3589 ;
  assign n3591 = n147 & ~n2851 ;
  assign n3592 = n160 & ~n2834 ;
  assign n3593 = ~n3591 & ~n3592 ;
  assign n3594 = n3590 & n3593 ;
  assign n3595 = n191 & ~n3594 ;
  assign n3596 = n174 & ~n2843 ;
  assign n3597 = n187 & ~n2753 ;
  assign n3598 = ~n3596 & ~n3597 ;
  assign n3599 = n147 & ~n2778 ;
  assign n3600 = n160 & ~n2761 ;
  assign n3601 = ~n3599 & ~n3600 ;
  assign n3602 = n3598 & n3601 ;
  assign n3603 = n244 & ~n3602 ;
  assign n3604 = ~n3595 & ~n3603 ;
  assign n3605 = n3587 & n3604 ;
  assign n3606 = x134 & ~n3605 ;
  assign n3607 = n187 & ~n2937 ;
  assign n3608 = n160 & ~n2945 ;
  assign n3609 = ~n3607 & ~n3608 ;
  assign n3610 = n147 & ~n2962 ;
  assign n3611 = n174 & ~n2918 ;
  assign n3612 = ~n3610 & ~n3611 ;
  assign n3613 = n3609 & n3612 ;
  assign n3614 = n244 & ~n3613 ;
  assign n3615 = n174 & ~n2879 ;
  assign n3616 = n187 & ~n2901 ;
  assign n3617 = ~n3615 & ~n3616 ;
  assign n3618 = n147 & ~n2926 ;
  assign n3619 = n160 & ~n2909 ;
  assign n3620 = ~n3618 & ~n3619 ;
  assign n3621 = n3617 & n3620 ;
  assign n3622 = n191 & ~n3621 ;
  assign n3623 = ~n3614 & ~n3622 ;
  assign n3624 = n174 & ~n2954 ;
  assign n3625 = n187 & ~n3010 ;
  assign n3626 = ~n3624 & ~n3625 ;
  assign n3627 = n147 & ~n3035 ;
  assign n3628 = n160 & ~n3018 ;
  assign n3629 = ~n3627 & ~n3628 ;
  assign n3630 = n3626 & n3629 ;
  assign n3631 = n351 & ~n3630 ;
  assign n3632 = n174 & ~n3027 ;
  assign n3633 = n187 & ~n2974 ;
  assign n3634 = ~n3632 & ~n3633 ;
  assign n3635 = n147 & ~n2999 ;
  assign n3636 = n160 & ~n2982 ;
  assign n3637 = ~n3635 & ~n3636 ;
  assign n3638 = n3634 & n3637 ;
  assign n3639 = n298 & ~n3638 ;
  assign n3640 = ~n3631 & ~n3639 ;
  assign n3641 = n3623 & n3640 ;
  assign n3642 = ~x134 & ~n3641 ;
  assign n3643 = ~n3606 & ~n3642 ;
  assign n3646 = n3643 & ~x142 ;
  assign n3647 = ~n3645 & ~n3646 ;
  assign n3648 = n147 & ~n240 ;
  assign n3649 = n160 & ~n228 ;
  assign n3650 = ~n3648 & ~n3649 ;
  assign n3651 = ~n159 & n174 ;
  assign n3652 = ~n146 & n187 ;
  assign n3653 = ~n3651 & ~n3652 ;
  assign n3654 = n3650 & n3653 ;
  assign n3655 = n191 & ~n3654 ;
  assign n3656 = n147 & ~n347 ;
  assign n3657 = n160 & ~n335 ;
  assign n3658 = ~n3656 & ~n3657 ;
  assign n3659 = n174 & ~n215 ;
  assign n3660 = n187 & ~n203 ;
  assign n3661 = ~n3659 & ~n3660 ;
  assign n3662 = n3658 & n3661 ;
  assign n3663 = n244 & ~n3662 ;
  assign n3664 = ~n3655 & ~n3663 ;
  assign n3665 = n147 & ~n403 ;
  assign n3666 = n160 & ~n391 ;
  assign n3667 = ~n3665 & ~n3666 ;
  assign n3668 = n174 & ~n269 ;
  assign n3669 = n187 & ~n257 ;
  assign n3670 = ~n3668 & ~n3669 ;
  assign n3671 = n3667 & n3670 ;
  assign n3672 = n298 & ~n3671 ;
  assign n3673 = n147 & ~n294 ;
  assign n3674 = n160 & ~n282 ;
  assign n3675 = ~n3673 & ~n3674 ;
  assign n3676 = n174 & ~n322 ;
  assign n3677 = n187 & ~n310 ;
  assign n3678 = ~n3676 & ~n3677 ;
  assign n3679 = n3675 & n3678 ;
  assign n3680 = n351 & ~n3679 ;
  assign n3681 = ~n3672 & ~n3680 ;
  assign n3682 = n3664 & n3681 ;
  assign n3683 = ~x134 & ~n3682 ;
  assign n3684 = n147 & ~n508 ;
  assign n3685 = n160 & ~n496 ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = n174 & ~n535 ;
  assign n3688 = n187 & ~n523 ;
  assign n3689 = ~n3687 & ~n3688 ;
  assign n3690 = n3686 & n3689 ;
  assign n3691 = n351 & ~n3690 ;
  assign n3692 = n147 & ~n186 ;
  assign n3693 = n160 & ~n173 ;
  assign n3694 = ~n3692 & ~n3693 ;
  assign n3695 = n174 & ~n483 ;
  assign n3696 = n187 & ~n471 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3698 = n3694 & n3697 ;
  assign n3699 = n298 & ~n3698 ;
  assign n3700 = ~n3691 & ~n3699 ;
  assign n3701 = n147 & ~n560 ;
  assign n3702 = n160 & ~n548 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = n174 & ~n430 ;
  assign n3705 = n187 & ~n418 ;
  assign n3706 = ~n3704 & ~n3705 ;
  assign n3707 = n3703 & n3706 ;
  assign n3708 = n244 & ~n3707 ;
  assign n3709 = n147 & ~n455 ;
  assign n3710 = n160 & ~n443 ;
  assign n3711 = ~n3709 & ~n3710 ;
  assign n3712 = n174 & ~n378 ;
  assign n3713 = n187 & ~n366 ;
  assign n3714 = ~n3712 & ~n3713 ;
  assign n3715 = n3711 & n3714 ;
  assign n3716 = n191 & ~n3715 ;
  assign n3717 = ~n3708 & ~n3716 ;
  assign n3718 = n3700 & n3717 ;
  assign n3719 = x134 & ~n3718 ;
  assign n3720 = ~n3683 & ~n3719 ;
  assign n3795 = ~n3720 & x143 ;
  assign n3721 = n174 & ~n668 ;
  assign n3722 = n187 & ~n656 ;
  assign n3723 = ~n3721 & ~n3722 ;
  assign n3724 = n147 & ~n591 ;
  assign n3725 = n160 & ~n579 ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3727 = n3723 & n3726 ;
  assign n3728 = n298 & ~n3727 ;
  assign n3729 = n174 & ~n773 ;
  assign n3730 = n187 & ~n761 ;
  assign n3731 = ~n3729 & ~n3730 ;
  assign n3732 = n147 & ~n643 ;
  assign n3733 = n160 & ~n631 ;
  assign n3734 = ~n3732 & ~n3733 ;
  assign n3735 = n3731 & n3734 ;
  assign n3736 = n351 & ~n3735 ;
  assign n3737 = ~n3728 & ~n3736 ;
  assign n3738 = n174 & ~n828 ;
  assign n3739 = n187 & ~n816 ;
  assign n3740 = ~n3738 & ~n3739 ;
  assign n3741 = n147 & ~n696 ;
  assign n3742 = n160 & ~n684 ;
  assign n3743 = ~n3741 & ~n3742 ;
  assign n3744 = n3740 & n3743 ;
  assign n3745 = n191 & ~n3744 ;
  assign n3746 = n174 & ~n721 ;
  assign n3747 = n187 & ~n709 ;
  assign n3748 = ~n3746 & ~n3747 ;
  assign n3749 = n147 & ~n748 ;
  assign n3750 = n160 & ~n736 ;
  assign n3751 = ~n3749 & ~n3750 ;
  assign n3752 = n3748 & n3751 ;
  assign n3753 = n244 & ~n3752 ;
  assign n3754 = ~n3745 & ~n3753 ;
  assign n3755 = n3737 & n3754 ;
  assign n3756 = x134 & ~n3755 ;
  assign n3757 = n174 & ~n933 ;
  assign n3758 = n187 & ~n921 ;
  assign n3759 = ~n3757 & ~n3758 ;
  assign n3760 = n147 & ~n960 ;
  assign n3761 = n160 & ~n948 ;
  assign n3762 = ~n3760 & ~n3761 ;
  assign n3763 = n3759 & n3762 ;
  assign n3764 = n244 & ~n3763 ;
  assign n3765 = n174 & ~n616 ;
  assign n3766 = n187 & ~n604 ;
  assign n3767 = ~n3765 & ~n3766 ;
  assign n3768 = n147 & ~n908 ;
  assign n3769 = n160 & ~n896 ;
  assign n3770 = ~n3768 & ~n3769 ;
  assign n3771 = n3767 & n3770 ;
  assign n3772 = n191 & ~n3771 ;
  assign n3773 = ~n3764 & ~n3772 ;
  assign n3774 = n174 & ~n985 ;
  assign n3775 = n187 & ~n973 ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3777 = n147 & ~n855 ;
  assign n3778 = n160 & ~n843 ;
  assign n3779 = ~n3777 & ~n3778 ;
  assign n3780 = n3776 & n3779 ;
  assign n3781 = n351 & ~n3780 ;
  assign n3782 = n174 & ~n880 ;
  assign n3783 = n187 & ~n868 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = n147 & ~n803 ;
  assign n3786 = n160 & ~n791 ;
  assign n3787 = ~n3785 & ~n3786 ;
  assign n3788 = n3784 & n3787 ;
  assign n3789 = n298 & ~n3788 ;
  assign n3790 = ~n3781 & ~n3789 ;
  assign n3791 = n3773 & n3790 ;
  assign n3792 = ~x134 & ~n3791 ;
  assign n3793 = ~n3756 & ~n3792 ;
  assign n3796 = n3793 & ~x143 ;
  assign n3797 = ~n3795 & ~n3796 ;
  assign n3798 = n147 & ~n1097 ;
  assign n3799 = n160 & ~n1085 ;
  assign n3800 = ~n3798 & ~n3799 ;
  assign n3801 = n174 & ~n1020 ;
  assign n3802 = n187 & ~n1008 ;
  assign n3803 = ~n3801 & ~n3802 ;
  assign n3804 = n3800 & n3803 ;
  assign n3805 = n191 & ~n3804 ;
  assign n3806 = n147 & ~n1202 ;
  assign n3807 = n160 & ~n1190 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = n174 & ~n1072 ;
  assign n3810 = n187 & ~n1060 ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = n3808 & n3811 ;
  assign n3813 = n244 & ~n3812 ;
  assign n3814 = ~n3805 & ~n3813 ;
  assign n3815 = n147 & ~n1309 ;
  assign n3816 = n160 & ~n1297 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = n174 & ~n1125 ;
  assign n3819 = n187 & ~n1113 ;
  assign n3820 = ~n3818 & ~n3819 ;
  assign n3821 = n3817 & n3820 ;
  assign n3822 = n298 & ~n3821 ;
  assign n3823 = n147 & ~n1150 ;
  assign n3824 = n160 & ~n1138 ;
  assign n3825 = ~n3823 & ~n3824 ;
  assign n3826 = n174 & ~n1177 ;
  assign n3827 = n187 & ~n1165 ;
  assign n3828 = ~n3826 & ~n3827 ;
  assign n3829 = n3825 & n3828 ;
  assign n3830 = n351 & ~n3829 ;
  assign n3831 = ~n3822 & ~n3830 ;
  assign n3832 = n3814 & n3831 ;
  assign n3833 = ~x134 & ~n3832 ;
  assign n3834 = n147 & ~n1257 ;
  assign n3835 = n160 & ~n1245 ;
  assign n3836 = ~n3834 & ~n3835 ;
  assign n3837 = n174 & ~n1337 ;
  assign n3838 = n187 & ~n1325 ;
  assign n3839 = ~n3837 & ~n3838 ;
  assign n3840 = n3836 & n3839 ;
  assign n3841 = n351 & ~n3840 ;
  assign n3842 = n147 & ~n1045 ;
  assign n3843 = n160 & ~n1033 ;
  assign n3844 = ~n3842 & ~n3843 ;
  assign n3845 = n174 & ~n1232 ;
  assign n3846 = n187 & ~n1220 ;
  assign n3847 = ~n3845 & ~n3846 ;
  assign n3848 = n3844 & n3847 ;
  assign n3849 = n298 & ~n3848 ;
  assign n3850 = ~n3841 & ~n3849 ;
  assign n3851 = n147 & ~n1362 ;
  assign n3852 = n160 & ~n1350 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = n174 & ~n1389 ;
  assign n3855 = n187 & ~n1377 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = n3853 & n3856 ;
  assign n3858 = n244 & ~n3857 ;
  assign n3859 = n147 & ~n1414 ;
  assign n3860 = n160 & ~n1402 ;
  assign n3861 = ~n3859 & ~n3860 ;
  assign n3862 = n174 & ~n1284 ;
  assign n3863 = n187 & ~n1272 ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = n3861 & n3864 ;
  assign n3866 = n191 & ~n3865 ;
  assign n3867 = ~n3858 & ~n3866 ;
  assign n3868 = n3850 & n3867 ;
  assign n3869 = x134 & ~n3868 ;
  assign n3870 = ~n3833 & ~n3869 ;
  assign n3945 = ~n3870 & x144 ;
  assign n3871 = n174 & ~n1522 ;
  assign n3872 = n187 & ~n1510 ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = n147 & ~n1445 ;
  assign n3875 = n160 & ~n1433 ;
  assign n3876 = ~n3874 & ~n3875 ;
  assign n3877 = n3873 & n3876 ;
  assign n3878 = n298 & ~n3877 ;
  assign n3879 = n174 & ~n1627 ;
  assign n3880 = n187 & ~n1615 ;
  assign n3881 = ~n3879 & ~n3880 ;
  assign n3882 = n147 & ~n1497 ;
  assign n3883 = n160 & ~n1485 ;
  assign n3884 = ~n3882 & ~n3883 ;
  assign n3885 = n3881 & n3884 ;
  assign n3886 = n351 & ~n3885 ;
  assign n3887 = ~n3878 & ~n3886 ;
  assign n3888 = n174 & ~n1734 ;
  assign n3889 = n187 & ~n1722 ;
  assign n3890 = ~n3888 & ~n3889 ;
  assign n3891 = n147 & ~n1550 ;
  assign n3892 = n160 & ~n1538 ;
  assign n3893 = ~n3891 & ~n3892 ;
  assign n3894 = n3890 & n3893 ;
  assign n3895 = n191 & ~n3894 ;
  assign n3896 = n174 & ~n1575 ;
  assign n3897 = n187 & ~n1563 ;
  assign n3898 = ~n3896 & ~n3897 ;
  assign n3899 = n147 & ~n1602 ;
  assign n3900 = n160 & ~n1590 ;
  assign n3901 = ~n3899 & ~n3900 ;
  assign n3902 = n3898 & n3901 ;
  assign n3903 = n244 & ~n3902 ;
  assign n3904 = ~n3895 & ~n3903 ;
  assign n3905 = n3887 & n3904 ;
  assign n3906 = x134 & ~n3905 ;
  assign n3907 = n174 & ~n1682 ;
  assign n3908 = n187 & ~n1670 ;
  assign n3909 = ~n3907 & ~n3908 ;
  assign n3910 = n147 & ~n1762 ;
  assign n3911 = n160 & ~n1750 ;
  assign n3912 = ~n3910 & ~n3911 ;
  assign n3913 = n3909 & n3912 ;
  assign n3914 = n244 & ~n3913 ;
  assign n3915 = n174 & ~n1470 ;
  assign n3916 = n187 & ~n1458 ;
  assign n3917 = ~n3915 & ~n3916 ;
  assign n3918 = n147 & ~n1657 ;
  assign n3919 = n160 & ~n1645 ;
  assign n3920 = ~n3918 & ~n3919 ;
  assign n3921 = n3917 & n3920 ;
  assign n3922 = n191 & ~n3921 ;
  assign n3923 = ~n3914 & ~n3922 ;
  assign n3924 = n174 & ~n1787 ;
  assign n3925 = n187 & ~n1775 ;
  assign n3926 = ~n3924 & ~n3925 ;
  assign n3927 = n147 & ~n1814 ;
  assign n3928 = n160 & ~n1802 ;
  assign n3929 = ~n3927 & ~n3928 ;
  assign n3930 = n3926 & n3929 ;
  assign n3931 = n351 & ~n3930 ;
  assign n3932 = n174 & ~n1839 ;
  assign n3933 = n187 & ~n1827 ;
  assign n3934 = ~n3932 & ~n3933 ;
  assign n3935 = n147 & ~n1709 ;
  assign n3936 = n160 & ~n1697 ;
  assign n3937 = ~n3935 & ~n3936 ;
  assign n3938 = n3934 & n3937 ;
  assign n3939 = n298 & ~n3938 ;
  assign n3940 = ~n3931 & ~n3939 ;
  assign n3941 = n3923 & n3940 ;
  assign n3942 = ~x134 & ~n3941 ;
  assign n3943 = ~n3906 & ~n3942 ;
  assign n3946 = n3943 & ~x144 ;
  assign n3947 = ~n3945 & ~n3946 ;
  assign n3948 = n147 & ~n1919 ;
  assign n3949 = n160 & ~n1911 ;
  assign n3950 = ~n3948 & ~n3949 ;
  assign n3951 = n174 & ~n1866 ;
  assign n3952 = n187 & ~n1858 ;
  assign n3953 = ~n3951 & ~n3952 ;
  assign n3954 = n3950 & n3953 ;
  assign n3955 = n191 & ~n3954 ;
  assign n3956 = n147 & ~n1992 ;
  assign n3957 = n160 & ~n1984 ;
  assign n3958 = ~n3956 & ~n3957 ;
  assign n3959 = n174 & ~n1902 ;
  assign n3960 = n187 & ~n1894 ;
  assign n3961 = ~n3959 & ~n3960 ;
  assign n3962 = n3958 & n3961 ;
  assign n3963 = n244 & ~n3962 ;
  assign n3964 = ~n3955 & ~n3963 ;
  assign n3965 = n147 & ~n2067 ;
  assign n3966 = n160 & ~n2059 ;
  assign n3967 = ~n3965 & ~n3966 ;
  assign n3968 = n174 & ~n1939 ;
  assign n3969 = n187 & ~n1931 ;
  assign n3970 = ~n3968 & ~n3969 ;
  assign n3971 = n3967 & n3970 ;
  assign n3972 = n298 & ~n3971 ;
  assign n3973 = n147 & ~n1956 ;
  assign n3974 = n160 & ~n1948 ;
  assign n3975 = ~n3973 & ~n3974 ;
  assign n3976 = n174 & ~n1975 ;
  assign n3977 = n187 & ~n1967 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = n3975 & n3978 ;
  assign n3980 = n351 & ~n3979 ;
  assign n3981 = ~n3972 & ~n3980 ;
  assign n3982 = n3964 & n3981 ;
  assign n3983 = ~x134 & ~n3982 ;
  assign n3984 = n147 & ~n2031 ;
  assign n3985 = n160 & ~n2023 ;
  assign n3986 = ~n3984 & ~n3985 ;
  assign n3987 = n174 & ~n2087 ;
  assign n3988 = n187 & ~n2079 ;
  assign n3989 = ~n3987 & ~n3988 ;
  assign n3990 = n3986 & n3989 ;
  assign n3991 = n351 & ~n3990 ;
  assign n3992 = n147 & ~n1883 ;
  assign n3993 = n160 & ~n1875 ;
  assign n3994 = ~n3992 & ~n3993 ;
  assign n3995 = n174 & ~n2014 ;
  assign n3996 = n187 & ~n2006 ;
  assign n3997 = ~n3995 & ~n3996 ;
  assign n3998 = n3994 & n3997 ;
  assign n3999 = n298 & ~n3998 ;
  assign n4000 = ~n3991 & ~n3999 ;
  assign n4001 = n147 & ~n2104 ;
  assign n4002 = n160 & ~n2096 ;
  assign n4003 = ~n4001 & ~n4002 ;
  assign n4004 = n174 & ~n2123 ;
  assign n4005 = n187 & ~n2115 ;
  assign n4006 = ~n4004 & ~n4005 ;
  assign n4007 = n4003 & n4006 ;
  assign n4008 = n244 & ~n4007 ;
  assign n4009 = n147 & ~n2140 ;
  assign n4010 = n160 & ~n2132 ;
  assign n4011 = ~n4009 & ~n4010 ;
  assign n4012 = n174 & ~n2050 ;
  assign n4013 = n187 & ~n2042 ;
  assign n4014 = ~n4012 & ~n4013 ;
  assign n4015 = n4011 & n4014 ;
  assign n4016 = n191 & ~n4015 ;
  assign n4017 = ~n4008 & ~n4016 ;
  assign n4018 = n4000 & n4017 ;
  assign n4019 = x134 & ~n4018 ;
  assign n4020 = ~n3983 & ~n4019 ;
  assign n4095 = ~n4020 & x145 ;
  assign n4021 = n174 & ~n2216 ;
  assign n4022 = n187 & ~n2208 ;
  assign n4023 = ~n4021 & ~n4022 ;
  assign n4024 = n147 & ~n2163 ;
  assign n4025 = n160 & ~n2155 ;
  assign n4026 = ~n4024 & ~n4025 ;
  assign n4027 = n4023 & n4026 ;
  assign n4028 = n298 & ~n4027 ;
  assign n4029 = n174 & ~n2289 ;
  assign n4030 = n187 & ~n2281 ;
  assign n4031 = ~n4029 & ~n4030 ;
  assign n4032 = n147 & ~n2199 ;
  assign n4033 = n160 & ~n2191 ;
  assign n4034 = ~n4032 & ~n4033 ;
  assign n4035 = n4031 & n4034 ;
  assign n4036 = n351 & ~n4035 ;
  assign n4037 = ~n4028 & ~n4036 ;
  assign n4038 = n174 & ~n2364 ;
  assign n4039 = n187 & ~n2356 ;
  assign n4040 = ~n4038 & ~n4039 ;
  assign n4041 = n147 & ~n2236 ;
  assign n4042 = n160 & ~n2228 ;
  assign n4043 = ~n4041 & ~n4042 ;
  assign n4044 = n4040 & n4043 ;
  assign n4045 = n191 & ~n4044 ;
  assign n4046 = n174 & ~n2253 ;
  assign n4047 = n187 & ~n2245 ;
  assign n4048 = ~n4046 & ~n4047 ;
  assign n4049 = n147 & ~n2272 ;
  assign n4050 = n160 & ~n2264 ;
  assign n4051 = ~n4049 & ~n4050 ;
  assign n4052 = n4048 & n4051 ;
  assign n4053 = n244 & ~n4052 ;
  assign n4054 = ~n4045 & ~n4053 ;
  assign n4055 = n4037 & n4054 ;
  assign n4056 = x134 & ~n4055 ;
  assign n4057 = n174 & ~n2328 ;
  assign n4058 = n187 & ~n2320 ;
  assign n4059 = ~n4057 & ~n4058 ;
  assign n4060 = n147 & ~n2384 ;
  assign n4061 = n160 & ~n2376 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = n4059 & n4062 ;
  assign n4064 = n244 & ~n4063 ;
  assign n4065 = n174 & ~n2180 ;
  assign n4066 = n187 & ~n2172 ;
  assign n4067 = ~n4065 & ~n4066 ;
  assign n4068 = n147 & ~n2311 ;
  assign n4069 = n160 & ~n2303 ;
  assign n4070 = ~n4068 & ~n4069 ;
  assign n4071 = n4067 & n4070 ;
  assign n4072 = n191 & ~n4071 ;
  assign n4073 = ~n4064 & ~n4072 ;
  assign n4074 = n174 & ~n2401 ;
  assign n4075 = n187 & ~n2393 ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = n147 & ~n2420 ;
  assign n4078 = n160 & ~n2412 ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = n4076 & n4079 ;
  assign n4081 = n351 & ~n4080 ;
  assign n4082 = n174 & ~n2437 ;
  assign n4083 = n187 & ~n2429 ;
  assign n4084 = ~n4082 & ~n4083 ;
  assign n4085 = n147 & ~n2347 ;
  assign n4086 = n160 & ~n2339 ;
  assign n4087 = ~n4085 & ~n4086 ;
  assign n4088 = n4084 & n4087 ;
  assign n4089 = n298 & ~n4088 ;
  assign n4090 = ~n4081 & ~n4089 ;
  assign n4091 = n4073 & n4090 ;
  assign n4092 = ~x134 & ~n4091 ;
  assign n4093 = ~n4056 & ~n4092 ;
  assign n4096 = n4093 & ~x145 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = n147 & ~n2517 ;
  assign n4099 = n160 & ~n2509 ;
  assign n4100 = ~n4098 & ~n4099 ;
  assign n4101 = n174 & ~n2573 ;
  assign n4102 = n187 & ~n2565 ;
  assign n4103 = ~n4101 & ~n4102 ;
  assign n4104 = n4100 & n4103 ;
  assign n4105 = n191 & ~n4104 ;
  assign n4106 = n147 & ~n2481 ;
  assign n4107 = n160 & ~n2473 ;
  assign n4108 = ~n4106 & ~n4107 ;
  assign n4109 = n174 & ~n2500 ;
  assign n4110 = n187 & ~n2492 ;
  assign n4111 = ~n4109 & ~n4110 ;
  assign n4112 = n4108 & n4111 ;
  assign n4113 = n244 & ~n4112 ;
  assign n4114 = ~n4105 & ~n4113 ;
  assign n4115 = n147 & ~n2702 ;
  assign n4116 = n160 & ~n2694 ;
  assign n4117 = ~n4115 & ~n4116 ;
  assign n4118 = n174 & ~n2537 ;
  assign n4119 = n187 & ~n2529 ;
  assign n4120 = ~n4118 & ~n4119 ;
  assign n4121 = n4117 & n4120 ;
  assign n4122 = n298 & ~n4121 ;
  assign n4123 = n147 & ~n2554 ;
  assign n4124 = n160 & ~n2546 ;
  assign n4125 = ~n4123 & ~n4124 ;
  assign n4126 = n174 & ~n2464 ;
  assign n4127 = n187 & ~n2456 ;
  assign n4128 = ~n4126 & ~n4127 ;
  assign n4129 = n4125 & n4128 ;
  assign n4130 = n351 & ~n4129 ;
  assign n4131 = ~n4122 & ~n4130 ;
  assign n4132 = n4114 & n4131 ;
  assign n4133 = ~x134 & ~n4132 ;
  assign n4134 = n147 & ~n2629 ;
  assign n4135 = n187 & ~n2640 ;
  assign n4136 = ~n4134 & ~n4135 ;
  assign n4137 = n174 & ~n2648 ;
  assign n4138 = n160 & ~n2621 ;
  assign n4139 = ~n4137 & ~n4138 ;
  assign n4140 = n4136 & n4139 ;
  assign n4141 = n351 & ~n4140 ;
  assign n4142 = n147 & ~n2590 ;
  assign n4143 = n160 & ~n2582 ;
  assign n4144 = ~n4142 & ~n4143 ;
  assign n4145 = n174 & ~n2612 ;
  assign n4146 = n187 & ~n2604 ;
  assign n4147 = ~n4145 & ~n4146 ;
  assign n4148 = n4144 & n4147 ;
  assign n4149 = n298 & ~n4148 ;
  assign n4150 = ~n4141 & ~n4149 ;
  assign n4151 = n147 & ~n2665 ;
  assign n4152 = n160 & ~n2657 ;
  assign n4153 = ~n4151 & ~n4152 ;
  assign n4154 = n174 & ~n2721 ;
  assign n4155 = n187 & ~n2713 ;
  assign n4156 = ~n4154 & ~n4155 ;
  assign n4157 = n4153 & n4156 ;
  assign n4158 = n244 & ~n4157 ;
  assign n4159 = n147 & ~n2738 ;
  assign n4160 = n160 & ~n2730 ;
  assign n4161 = ~n4159 & ~n4160 ;
  assign n4162 = n174 & ~n2685 ;
  assign n4163 = n187 & ~n2677 ;
  assign n4164 = ~n4162 & ~n4163 ;
  assign n4165 = n4161 & n4164 ;
  assign n4166 = n191 & ~n4165 ;
  assign n4167 = ~n4158 & ~n4166 ;
  assign n4168 = n4150 & n4167 ;
  assign n4169 = x134 & ~n4168 ;
  assign n4170 = ~n4133 & ~n4169 ;
  assign n4245 = ~n4170 & x146 ;
  assign n4171 = n174 & ~n2814 ;
  assign n4172 = n187 & ~n2806 ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4174 = n147 & ~n2870 ;
  assign n4175 = n160 & ~n2862 ;
  assign n4176 = ~n4174 & ~n4175 ;
  assign n4177 = n4173 & n4176 ;
  assign n4178 = n298 & ~n4177 ;
  assign n4179 = n174 & ~n2778 ;
  assign n4180 = n187 & ~n2770 ;
  assign n4181 = ~n4179 & ~n4180 ;
  assign n4182 = n147 & ~n2797 ;
  assign n4183 = n160 & ~n2789 ;
  assign n4184 = ~n4182 & ~n4183 ;
  assign n4185 = n4181 & n4184 ;
  assign n4186 = n351 & ~n4185 ;
  assign n4187 = ~n4178 & ~n4186 ;
  assign n4188 = n174 & ~n2999 ;
  assign n4189 = n187 & ~n2991 ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = n147 & ~n2834 ;
  assign n4192 = n160 & ~n2826 ;
  assign n4193 = ~n4191 & ~n4192 ;
  assign n4194 = n4190 & n4193 ;
  assign n4195 = n191 & ~n4194 ;
  assign n4196 = n174 & ~n2851 ;
  assign n4197 = n187 & ~n2843 ;
  assign n4198 = ~n4196 & ~n4197 ;
  assign n4199 = n147 & ~n2761 ;
  assign n4200 = n160 & ~n2753 ;
  assign n4201 = ~n4199 & ~n4200 ;
  assign n4202 = n4198 & n4201 ;
  assign n4203 = n244 & ~n4202 ;
  assign n4204 = ~n4195 & ~n4203 ;
  assign n4205 = n4187 & n4204 ;
  assign n4206 = x134 & ~n4205 ;
  assign n4207 = n174 & ~n2926 ;
  assign n4208 = n160 & ~n2937 ;
  assign n4209 = ~n4207 & ~n4208 ;
  assign n4210 = n147 & ~n2945 ;
  assign n4211 = n187 & ~n2918 ;
  assign n4212 = ~n4210 & ~n4211 ;
  assign n4213 = n4209 & n4212 ;
  assign n4214 = n244 & ~n4213 ;
  assign n4215 = n174 & ~n2887 ;
  assign n4216 = n187 & ~n2879 ;
  assign n4217 = ~n4215 & ~n4216 ;
  assign n4218 = n147 & ~n2909 ;
  assign n4219 = n160 & ~n2901 ;
  assign n4220 = ~n4218 & ~n4219 ;
  assign n4221 = n4217 & n4220 ;
  assign n4222 = n191 & ~n4221 ;
  assign n4223 = ~n4214 & ~n4222 ;
  assign n4224 = n174 & ~n2962 ;
  assign n4225 = n187 & ~n2954 ;
  assign n4226 = ~n4224 & ~n4225 ;
  assign n4227 = n147 & ~n3018 ;
  assign n4228 = n160 & ~n3010 ;
  assign n4229 = ~n4227 & ~n4228 ;
  assign n4230 = n4226 & n4229 ;
  assign n4231 = n351 & ~n4230 ;
  assign n4232 = n174 & ~n3035 ;
  assign n4233 = n187 & ~n3027 ;
  assign n4234 = ~n4232 & ~n4233 ;
  assign n4235 = n147 & ~n2982 ;
  assign n4236 = n160 & ~n2974 ;
  assign n4237 = ~n4235 & ~n4236 ;
  assign n4238 = n4234 & n4237 ;
  assign n4239 = n298 & ~n4238 ;
  assign n4240 = ~n4231 & ~n4239 ;
  assign n4241 = n4223 & n4240 ;
  assign n4242 = ~x134 & ~n4241 ;
  assign n4243 = ~n4206 & ~n4242 ;
  assign n4246 = n4243 & ~x146 ;
  assign n4247 = ~n4245 & ~n4246 ;
  assign n4248 = n147 & ~n215 ;
  assign n4249 = n160 & ~n240 ;
  assign n4250 = ~n4248 & ~n4249 ;
  assign n4251 = ~n146 & n174 ;
  assign n4252 = n187 & ~n228 ;
  assign n4253 = ~n4251 & ~n4252 ;
  assign n4254 = n4250 & n4253 ;
  assign n4255 = n191 & ~n4254 ;
  assign n4256 = n147 & ~n322 ;
  assign n4257 = n160 & ~n347 ;
  assign n4258 = ~n4256 & ~n4257 ;
  assign n4259 = n174 & ~n203 ;
  assign n4260 = n187 & ~n335 ;
  assign n4261 = ~n4259 & ~n4260 ;
  assign n4262 = n4258 & n4261 ;
  assign n4263 = n244 & ~n4262 ;
  assign n4264 = ~n4255 & ~n4263 ;
  assign n4265 = n147 & ~n378 ;
  assign n4266 = n160 & ~n403 ;
  assign n4267 = ~n4265 & ~n4266 ;
  assign n4268 = n174 & ~n257 ;
  assign n4269 = n187 & ~n391 ;
  assign n4270 = ~n4268 & ~n4269 ;
  assign n4271 = n4267 & n4270 ;
  assign n4272 = n298 & ~n4271 ;
  assign n4273 = n147 & ~n269 ;
  assign n4274 = n160 & ~n294 ;
  assign n4275 = ~n4273 & ~n4274 ;
  assign n4276 = n174 & ~n310 ;
  assign n4277 = n187 & ~n282 ;
  assign n4278 = ~n4276 & ~n4277 ;
  assign n4279 = n4275 & n4278 ;
  assign n4280 = n351 & ~n4279 ;
  assign n4281 = ~n4272 & ~n4280 ;
  assign n4282 = n4264 & n4281 ;
  assign n4283 = ~x134 & ~n4282 ;
  assign n4284 = n147 & ~n483 ;
  assign n4285 = n160 & ~n508 ;
  assign n4286 = ~n4284 & ~n4285 ;
  assign n4287 = n174 & ~n523 ;
  assign n4288 = n187 & ~n496 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = n4286 & n4289 ;
  assign n4291 = n351 & ~n4290 ;
  assign n4292 = n147 & ~n159 ;
  assign n4293 = n160 & ~n186 ;
  assign n4294 = ~n4292 & ~n4293 ;
  assign n4295 = n174 & ~n471 ;
  assign n4296 = ~n173 & n187 ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4298 = n4294 & n4297 ;
  assign n4299 = n298 & ~n4298 ;
  assign n4300 = ~n4291 & ~n4299 ;
  assign n4301 = n147 & ~n535 ;
  assign n4302 = n160 & ~n560 ;
  assign n4303 = ~n4301 & ~n4302 ;
  assign n4304 = n174 & ~n418 ;
  assign n4305 = n187 & ~n548 ;
  assign n4306 = ~n4304 & ~n4305 ;
  assign n4307 = n4303 & n4306 ;
  assign n4308 = n244 & ~n4307 ;
  assign n4309 = n147 & ~n430 ;
  assign n4310 = n160 & ~n455 ;
  assign n4311 = ~n4309 & ~n4310 ;
  assign n4312 = n174 & ~n366 ;
  assign n4313 = n187 & ~n443 ;
  assign n4314 = ~n4312 & ~n4313 ;
  assign n4315 = n4311 & n4314 ;
  assign n4316 = n191 & ~n4315 ;
  assign n4317 = ~n4308 & ~n4316 ;
  assign n4318 = n4300 & n4317 ;
  assign n4319 = x134 & ~n4318 ;
  assign n4320 = ~n4283 & ~n4319 ;
  assign n4395 = ~n4320 & x147 ;
  assign n4321 = n174 & ~n643 ;
  assign n4322 = n187 & ~n668 ;
  assign n4323 = ~n4321 & ~n4322 ;
  assign n4324 = n147 & ~n579 ;
  assign n4325 = n160 & ~n656 ;
  assign n4326 = ~n4324 & ~n4325 ;
  assign n4327 = n4323 & n4326 ;
  assign n4328 = n298 & ~n4327 ;
  assign n4329 = n174 & ~n748 ;
  assign n4330 = n187 & ~n773 ;
  assign n4331 = ~n4329 & ~n4330 ;
  assign n4332 = n147 & ~n631 ;
  assign n4333 = n160 & ~n761 ;
  assign n4334 = ~n4332 & ~n4333 ;
  assign n4335 = n4331 & n4334 ;
  assign n4336 = n351 & ~n4335 ;
  assign n4337 = ~n4328 & ~n4336 ;
  assign n4338 = n174 & ~n803 ;
  assign n4339 = n187 & ~n828 ;
  assign n4340 = ~n4338 & ~n4339 ;
  assign n4341 = n147 & ~n684 ;
  assign n4342 = n160 & ~n816 ;
  assign n4343 = ~n4341 & ~n4342 ;
  assign n4344 = n4340 & n4343 ;
  assign n4345 = n191 & ~n4344 ;
  assign n4346 = n174 & ~n696 ;
  assign n4347 = n187 & ~n721 ;
  assign n4348 = ~n4346 & ~n4347 ;
  assign n4349 = n147 & ~n736 ;
  assign n4350 = n160 & ~n709 ;
  assign n4351 = ~n4349 & ~n4350 ;
  assign n4352 = n4348 & n4351 ;
  assign n4353 = n244 & ~n4352 ;
  assign n4354 = ~n4345 & ~n4353 ;
  assign n4355 = n4337 & n4354 ;
  assign n4356 = x134 & ~n4355 ;
  assign n4357 = n174 & ~n908 ;
  assign n4358 = n187 & ~n933 ;
  assign n4359 = ~n4357 & ~n4358 ;
  assign n4360 = n147 & ~n948 ;
  assign n4361 = n160 & ~n921 ;
  assign n4362 = ~n4360 & ~n4361 ;
  assign n4363 = n4359 & n4362 ;
  assign n4364 = n244 & ~n4363 ;
  assign n4365 = n174 & ~n591 ;
  assign n4366 = n187 & ~n616 ;
  assign n4367 = ~n4365 & ~n4366 ;
  assign n4368 = n147 & ~n896 ;
  assign n4369 = n160 & ~n604 ;
  assign n4370 = ~n4368 & ~n4369 ;
  assign n4371 = n4367 & n4370 ;
  assign n4372 = n191 & ~n4371 ;
  assign n4373 = ~n4364 & ~n4372 ;
  assign n4374 = n174 & ~n960 ;
  assign n4375 = n187 & ~n985 ;
  assign n4376 = ~n4374 & ~n4375 ;
  assign n4377 = n147 & ~n843 ;
  assign n4378 = n160 & ~n973 ;
  assign n4379 = ~n4377 & ~n4378 ;
  assign n4380 = n4376 & n4379 ;
  assign n4381 = n351 & ~n4380 ;
  assign n4382 = n174 & ~n855 ;
  assign n4383 = n187 & ~n880 ;
  assign n4384 = ~n4382 & ~n4383 ;
  assign n4385 = n147 & ~n791 ;
  assign n4386 = n160 & ~n868 ;
  assign n4387 = ~n4385 & ~n4386 ;
  assign n4388 = n4384 & n4387 ;
  assign n4389 = n298 & ~n4388 ;
  assign n4390 = ~n4381 & ~n4389 ;
  assign n4391 = n4373 & n4390 ;
  assign n4392 = ~x134 & ~n4391 ;
  assign n4393 = ~n4356 & ~n4392 ;
  assign n4396 = n4393 & ~x147 ;
  assign n4397 = ~n4395 & ~n4396 ;
  assign n4398 = n147 & ~n1072 ;
  assign n4399 = n160 & ~n1097 ;
  assign n4400 = ~n4398 & ~n4399 ;
  assign n4401 = n174 & ~n1008 ;
  assign n4402 = n187 & ~n1085 ;
  assign n4403 = ~n4401 & ~n4402 ;
  assign n4404 = n4400 & n4403 ;
  assign n4405 = n191 & ~n4404 ;
  assign n4406 = n147 & ~n1177 ;
  assign n4407 = n160 & ~n1202 ;
  assign n4408 = ~n4406 & ~n4407 ;
  assign n4409 = n174 & ~n1060 ;
  assign n4410 = n187 & ~n1190 ;
  assign n4411 = ~n4409 & ~n4410 ;
  assign n4412 = n4408 & n4411 ;
  assign n4413 = n244 & ~n4412 ;
  assign n4414 = ~n4405 & ~n4413 ;
  assign n4415 = n147 & ~n1284 ;
  assign n4416 = n160 & ~n1309 ;
  assign n4417 = ~n4415 & ~n4416 ;
  assign n4418 = n174 & ~n1113 ;
  assign n4419 = n187 & ~n1297 ;
  assign n4420 = ~n4418 & ~n4419 ;
  assign n4421 = n4417 & n4420 ;
  assign n4422 = n298 & ~n4421 ;
  assign n4423 = n147 & ~n1125 ;
  assign n4424 = n160 & ~n1150 ;
  assign n4425 = ~n4423 & ~n4424 ;
  assign n4426 = n174 & ~n1165 ;
  assign n4427 = n187 & ~n1138 ;
  assign n4428 = ~n4426 & ~n4427 ;
  assign n4429 = n4425 & n4428 ;
  assign n4430 = n351 & ~n4429 ;
  assign n4431 = ~n4422 & ~n4430 ;
  assign n4432 = n4414 & n4431 ;
  assign n4433 = ~x134 & ~n4432 ;
  assign n4434 = n147 & ~n1232 ;
  assign n4435 = n160 & ~n1257 ;
  assign n4436 = ~n4434 & ~n4435 ;
  assign n4437 = n174 & ~n1325 ;
  assign n4438 = n187 & ~n1245 ;
  assign n4439 = ~n4437 & ~n4438 ;
  assign n4440 = n4436 & n4439 ;
  assign n4441 = n351 & ~n4440 ;
  assign n4442 = n147 & ~n1020 ;
  assign n4443 = n160 & ~n1045 ;
  assign n4444 = ~n4442 & ~n4443 ;
  assign n4445 = n174 & ~n1220 ;
  assign n4446 = n187 & ~n1033 ;
  assign n4447 = ~n4445 & ~n4446 ;
  assign n4448 = n4444 & n4447 ;
  assign n4449 = n298 & ~n4448 ;
  assign n4450 = ~n4441 & ~n4449 ;
  assign n4451 = n147 & ~n1337 ;
  assign n4452 = n160 & ~n1362 ;
  assign n4453 = ~n4451 & ~n4452 ;
  assign n4454 = n174 & ~n1377 ;
  assign n4455 = n187 & ~n1350 ;
  assign n4456 = ~n4454 & ~n4455 ;
  assign n4457 = n4453 & n4456 ;
  assign n4458 = n244 & ~n4457 ;
  assign n4459 = n147 & ~n1389 ;
  assign n4460 = n160 & ~n1414 ;
  assign n4461 = ~n4459 & ~n4460 ;
  assign n4462 = n174 & ~n1272 ;
  assign n4463 = n187 & ~n1402 ;
  assign n4464 = ~n4462 & ~n4463 ;
  assign n4465 = n4461 & n4464 ;
  assign n4466 = n191 & ~n4465 ;
  assign n4467 = ~n4458 & ~n4466 ;
  assign n4468 = n4450 & n4467 ;
  assign n4469 = x134 & ~n4468 ;
  assign n4470 = ~n4433 & ~n4469 ;
  assign n4545 = ~n4470 & x148 ;
  assign n4471 = n174 & ~n1497 ;
  assign n4472 = n187 & ~n1522 ;
  assign n4473 = ~n4471 & ~n4472 ;
  assign n4474 = n147 & ~n1433 ;
  assign n4475 = n160 & ~n1510 ;
  assign n4476 = ~n4474 & ~n4475 ;
  assign n4477 = n4473 & n4476 ;
  assign n4478 = n298 & ~n4477 ;
  assign n4479 = n174 & ~n1602 ;
  assign n4480 = n187 & ~n1627 ;
  assign n4481 = ~n4479 & ~n4480 ;
  assign n4482 = n147 & ~n1485 ;
  assign n4483 = n160 & ~n1615 ;
  assign n4484 = ~n4482 & ~n4483 ;
  assign n4485 = n4481 & n4484 ;
  assign n4486 = n351 & ~n4485 ;
  assign n4487 = ~n4478 & ~n4486 ;
  assign n4488 = n174 & ~n1709 ;
  assign n4489 = n187 & ~n1734 ;
  assign n4490 = ~n4488 & ~n4489 ;
  assign n4491 = n147 & ~n1538 ;
  assign n4492 = n160 & ~n1722 ;
  assign n4493 = ~n4491 & ~n4492 ;
  assign n4494 = n4490 & n4493 ;
  assign n4495 = n191 & ~n4494 ;
  assign n4496 = n174 & ~n1550 ;
  assign n4497 = n187 & ~n1575 ;
  assign n4498 = ~n4496 & ~n4497 ;
  assign n4499 = n147 & ~n1590 ;
  assign n4500 = n160 & ~n1563 ;
  assign n4501 = ~n4499 & ~n4500 ;
  assign n4502 = n4498 & n4501 ;
  assign n4503 = n244 & ~n4502 ;
  assign n4504 = ~n4495 & ~n4503 ;
  assign n4505 = n4487 & n4504 ;
  assign n4506 = x134 & ~n4505 ;
  assign n4507 = n174 & ~n1657 ;
  assign n4508 = n187 & ~n1682 ;
  assign n4509 = ~n4507 & ~n4508 ;
  assign n4510 = n147 & ~n1750 ;
  assign n4511 = n160 & ~n1670 ;
  assign n4512 = ~n4510 & ~n4511 ;
  assign n4513 = n4509 & n4512 ;
  assign n4514 = n244 & ~n4513 ;
  assign n4515 = n174 & ~n1445 ;
  assign n4516 = n187 & ~n1470 ;
  assign n4517 = ~n4515 & ~n4516 ;
  assign n4518 = n147 & ~n1645 ;
  assign n4519 = n160 & ~n1458 ;
  assign n4520 = ~n4518 & ~n4519 ;
  assign n4521 = n4517 & n4520 ;
  assign n4522 = n191 & ~n4521 ;
  assign n4523 = ~n4514 & ~n4522 ;
  assign n4524 = n174 & ~n1762 ;
  assign n4525 = n187 & ~n1787 ;
  assign n4526 = ~n4524 & ~n4525 ;
  assign n4527 = n147 & ~n1802 ;
  assign n4528 = n160 & ~n1775 ;
  assign n4529 = ~n4527 & ~n4528 ;
  assign n4530 = n4526 & n4529 ;
  assign n4531 = n351 & ~n4530 ;
  assign n4532 = n174 & ~n1814 ;
  assign n4533 = n187 & ~n1839 ;
  assign n4534 = ~n4532 & ~n4533 ;
  assign n4535 = n147 & ~n1697 ;
  assign n4536 = n160 & ~n1827 ;
  assign n4537 = ~n4535 & ~n4536 ;
  assign n4538 = n4534 & n4537 ;
  assign n4539 = n298 & ~n4538 ;
  assign n4540 = ~n4531 & ~n4539 ;
  assign n4541 = n4523 & n4540 ;
  assign n4542 = ~x134 & ~n4541 ;
  assign n4543 = ~n4506 & ~n4542 ;
  assign n4546 = n4543 & ~x148 ;
  assign n4547 = ~n4545 & ~n4546 ;
  assign n4548 = n147 & ~n1902 ;
  assign n4549 = n160 & ~n1919 ;
  assign n4550 = ~n4548 & ~n4549 ;
  assign n4551 = n174 & ~n1858 ;
  assign n4552 = n187 & ~n1911 ;
  assign n4553 = ~n4551 & ~n4552 ;
  assign n4554 = n4550 & n4553 ;
  assign n4555 = n191 & ~n4554 ;
  assign n4556 = n147 & ~n1975 ;
  assign n4557 = n160 & ~n1992 ;
  assign n4558 = ~n4556 & ~n4557 ;
  assign n4559 = n174 & ~n1894 ;
  assign n4560 = n187 & ~n1984 ;
  assign n4561 = ~n4559 & ~n4560 ;
  assign n4562 = n4558 & n4561 ;
  assign n4563 = n244 & ~n4562 ;
  assign n4564 = ~n4555 & ~n4563 ;
  assign n4565 = n147 & ~n2050 ;
  assign n4566 = n160 & ~n2067 ;
  assign n4567 = ~n4565 & ~n4566 ;
  assign n4568 = n174 & ~n1931 ;
  assign n4569 = n187 & ~n2059 ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = n4567 & n4570 ;
  assign n4572 = n298 & ~n4571 ;
  assign n4573 = n147 & ~n1939 ;
  assign n4574 = n160 & ~n1956 ;
  assign n4575 = ~n4573 & ~n4574 ;
  assign n4576 = n174 & ~n1967 ;
  assign n4577 = n187 & ~n1948 ;
  assign n4578 = ~n4576 & ~n4577 ;
  assign n4579 = n4575 & n4578 ;
  assign n4580 = n351 & ~n4579 ;
  assign n4581 = ~n4572 & ~n4580 ;
  assign n4582 = n4564 & n4581 ;
  assign n4583 = ~x134 & ~n4582 ;
  assign n4584 = n147 & ~n2014 ;
  assign n4585 = n160 & ~n2031 ;
  assign n4586 = ~n4584 & ~n4585 ;
  assign n4587 = n174 & ~n2079 ;
  assign n4588 = n187 & ~n2023 ;
  assign n4589 = ~n4587 & ~n4588 ;
  assign n4590 = n4586 & n4589 ;
  assign n4591 = n351 & ~n4590 ;
  assign n4592 = n147 & ~n1866 ;
  assign n4593 = n160 & ~n1883 ;
  assign n4594 = ~n4592 & ~n4593 ;
  assign n4595 = n174 & ~n2006 ;
  assign n4596 = n187 & ~n1875 ;
  assign n4597 = ~n4595 & ~n4596 ;
  assign n4598 = n4594 & n4597 ;
  assign n4599 = n298 & ~n4598 ;
  assign n4600 = ~n4591 & ~n4599 ;
  assign n4601 = n147 & ~n2087 ;
  assign n4602 = n160 & ~n2104 ;
  assign n4603 = ~n4601 & ~n4602 ;
  assign n4604 = n174 & ~n2115 ;
  assign n4605 = n187 & ~n2096 ;
  assign n4606 = ~n4604 & ~n4605 ;
  assign n4607 = n4603 & n4606 ;
  assign n4608 = n244 & ~n4607 ;
  assign n4609 = n147 & ~n2123 ;
  assign n4610 = n160 & ~n2140 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = n174 & ~n2042 ;
  assign n4613 = n187 & ~n2132 ;
  assign n4614 = ~n4612 & ~n4613 ;
  assign n4615 = n4611 & n4614 ;
  assign n4616 = n191 & ~n4615 ;
  assign n4617 = ~n4608 & ~n4616 ;
  assign n4618 = n4600 & n4617 ;
  assign n4619 = x134 & ~n4618 ;
  assign n4620 = ~n4583 & ~n4619 ;
  assign n4695 = ~n4620 & x149 ;
  assign n4621 = n174 & ~n2199 ;
  assign n4622 = n187 & ~n2216 ;
  assign n4623 = ~n4621 & ~n4622 ;
  assign n4624 = n147 & ~n2155 ;
  assign n4625 = n160 & ~n2208 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = n4623 & n4626 ;
  assign n4628 = n298 & ~n4627 ;
  assign n4629 = n174 & ~n2272 ;
  assign n4630 = n187 & ~n2289 ;
  assign n4631 = ~n4629 & ~n4630 ;
  assign n4632 = n147 & ~n2191 ;
  assign n4633 = n160 & ~n2281 ;
  assign n4634 = ~n4632 & ~n4633 ;
  assign n4635 = n4631 & n4634 ;
  assign n4636 = n351 & ~n4635 ;
  assign n4637 = ~n4628 & ~n4636 ;
  assign n4638 = n174 & ~n2347 ;
  assign n4639 = n187 & ~n2364 ;
  assign n4640 = ~n4638 & ~n4639 ;
  assign n4641 = n147 & ~n2228 ;
  assign n4642 = n160 & ~n2356 ;
  assign n4643 = ~n4641 & ~n4642 ;
  assign n4644 = n4640 & n4643 ;
  assign n4645 = n191 & ~n4644 ;
  assign n4646 = n174 & ~n2236 ;
  assign n4647 = n187 & ~n2253 ;
  assign n4648 = ~n4646 & ~n4647 ;
  assign n4649 = n147 & ~n2264 ;
  assign n4650 = n160 & ~n2245 ;
  assign n4651 = ~n4649 & ~n4650 ;
  assign n4652 = n4648 & n4651 ;
  assign n4653 = n244 & ~n4652 ;
  assign n4654 = ~n4645 & ~n4653 ;
  assign n4655 = n4637 & n4654 ;
  assign n4656 = x134 & ~n4655 ;
  assign n4657 = n174 & ~n2311 ;
  assign n4658 = n187 & ~n2328 ;
  assign n4659 = ~n4657 & ~n4658 ;
  assign n4660 = n147 & ~n2376 ;
  assign n4661 = n160 & ~n2320 ;
  assign n4662 = ~n4660 & ~n4661 ;
  assign n4663 = n4659 & n4662 ;
  assign n4664 = n244 & ~n4663 ;
  assign n4665 = n174 & ~n2163 ;
  assign n4666 = n187 & ~n2180 ;
  assign n4667 = ~n4665 & ~n4666 ;
  assign n4668 = n147 & ~n2303 ;
  assign n4669 = n160 & ~n2172 ;
  assign n4670 = ~n4668 & ~n4669 ;
  assign n4671 = n4667 & n4670 ;
  assign n4672 = n191 & ~n4671 ;
  assign n4673 = ~n4664 & ~n4672 ;
  assign n4674 = n174 & ~n2384 ;
  assign n4675 = n187 & ~n2401 ;
  assign n4676 = ~n4674 & ~n4675 ;
  assign n4677 = n147 & ~n2412 ;
  assign n4678 = n160 & ~n2393 ;
  assign n4679 = ~n4677 & ~n4678 ;
  assign n4680 = n4676 & n4679 ;
  assign n4681 = n351 & ~n4680 ;
  assign n4682 = n174 & ~n2420 ;
  assign n4683 = n187 & ~n2437 ;
  assign n4684 = ~n4682 & ~n4683 ;
  assign n4685 = n147 & ~n2339 ;
  assign n4686 = n160 & ~n2429 ;
  assign n4687 = ~n4685 & ~n4686 ;
  assign n4688 = n4684 & n4687 ;
  assign n4689 = n298 & ~n4688 ;
  assign n4690 = ~n4681 & ~n4689 ;
  assign n4691 = n4673 & n4690 ;
  assign n4692 = ~x134 & ~n4691 ;
  assign n4693 = ~n4656 & ~n4692 ;
  assign n4696 = n4693 & ~x149 ;
  assign n4697 = ~n4695 & ~n4696 ;
  assign n4698 = n147 & ~n2500 ;
  assign n4699 = n160 & ~n2517 ;
  assign n4700 = ~n4698 & ~n4699 ;
  assign n4701 = n174 & ~n2565 ;
  assign n4702 = n187 & ~n2509 ;
  assign n4703 = ~n4701 & ~n4702 ;
  assign n4704 = n4700 & n4703 ;
  assign n4705 = n191 & ~n4704 ;
  assign n4706 = n147 & ~n2464 ;
  assign n4707 = n160 & ~n2481 ;
  assign n4708 = ~n4706 & ~n4707 ;
  assign n4709 = n174 & ~n2492 ;
  assign n4710 = n187 & ~n2473 ;
  assign n4711 = ~n4709 & ~n4710 ;
  assign n4712 = n4708 & n4711 ;
  assign n4713 = n244 & ~n4712 ;
  assign n4714 = ~n4705 & ~n4713 ;
  assign n4715 = n147 & ~n2685 ;
  assign n4716 = n160 & ~n2702 ;
  assign n4717 = ~n4715 & ~n4716 ;
  assign n4718 = n174 & ~n2529 ;
  assign n4719 = n187 & ~n2694 ;
  assign n4720 = ~n4718 & ~n4719 ;
  assign n4721 = n4717 & n4720 ;
  assign n4722 = n298 & ~n4721 ;
  assign n4723 = n147 & ~n2537 ;
  assign n4724 = n160 & ~n2554 ;
  assign n4725 = ~n4723 & ~n4724 ;
  assign n4726 = n174 & ~n2456 ;
  assign n4727 = n187 & ~n2546 ;
  assign n4728 = ~n4726 & ~n4727 ;
  assign n4729 = n4725 & n4728 ;
  assign n4730 = n351 & ~n4729 ;
  assign n4731 = ~n4722 & ~n4730 ;
  assign n4732 = n4714 & n4731 ;
  assign n4733 = ~x134 & ~n4732 ;
  assign n4734 = n147 & ~n2612 ;
  assign n4735 = n160 & ~n2629 ;
  assign n4736 = ~n4734 & ~n4735 ;
  assign n4737 = n174 & ~n2640 ;
  assign n4738 = n187 & ~n2621 ;
  assign n4739 = ~n4737 & ~n4738 ;
  assign n4740 = n4736 & n4739 ;
  assign n4741 = n351 & ~n4740 ;
  assign n4742 = n147 & ~n2573 ;
  assign n4743 = n160 & ~n2590 ;
  assign n4744 = ~n4742 & ~n4743 ;
  assign n4745 = n174 & ~n2604 ;
  assign n4746 = n187 & ~n2582 ;
  assign n4747 = ~n4745 & ~n4746 ;
  assign n4748 = n4744 & n4747 ;
  assign n4749 = n298 & ~n4748 ;
  assign n4750 = ~n4741 & ~n4749 ;
  assign n4751 = n147 & ~n2648 ;
  assign n4752 = n160 & ~n2665 ;
  assign n4753 = ~n4751 & ~n4752 ;
  assign n4754 = n174 & ~n2713 ;
  assign n4755 = n187 & ~n2657 ;
  assign n4756 = ~n4754 & ~n4755 ;
  assign n4757 = n4753 & n4756 ;
  assign n4758 = n244 & ~n4757 ;
  assign n4759 = n147 & ~n2721 ;
  assign n4760 = n160 & ~n2738 ;
  assign n4761 = ~n4759 & ~n4760 ;
  assign n4762 = n174 & ~n2677 ;
  assign n4763 = n187 & ~n2730 ;
  assign n4764 = ~n4762 & ~n4763 ;
  assign n4765 = n4761 & n4764 ;
  assign n4766 = n191 & ~n4765 ;
  assign n4767 = ~n4758 & ~n4766 ;
  assign n4768 = n4750 & n4767 ;
  assign n4769 = x134 & ~n4768 ;
  assign n4770 = ~n4733 & ~n4769 ;
  assign n4845 = ~n4770 & x150 ;
  assign n4771 = n174 & ~n2797 ;
  assign n4772 = n187 & ~n2814 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = n147 & ~n2862 ;
  assign n4775 = n160 & ~n2806 ;
  assign n4776 = ~n4774 & ~n4775 ;
  assign n4777 = n4773 & n4776 ;
  assign n4778 = n298 & ~n4777 ;
  assign n4779 = n174 & ~n2761 ;
  assign n4780 = n187 & ~n2778 ;
  assign n4781 = ~n4779 & ~n4780 ;
  assign n4782 = n147 & ~n2789 ;
  assign n4783 = n160 & ~n2770 ;
  assign n4784 = ~n4782 & ~n4783 ;
  assign n4785 = n4781 & n4784 ;
  assign n4786 = n351 & ~n4785 ;
  assign n4787 = ~n4778 & ~n4786 ;
  assign n4788 = n174 & ~n2982 ;
  assign n4789 = n187 & ~n2999 ;
  assign n4790 = ~n4788 & ~n4789 ;
  assign n4791 = n147 & ~n2826 ;
  assign n4792 = n160 & ~n2991 ;
  assign n4793 = ~n4791 & ~n4792 ;
  assign n4794 = n4790 & n4793 ;
  assign n4795 = n191 & ~n4794 ;
  assign n4796 = n174 & ~n2834 ;
  assign n4797 = n187 & ~n2851 ;
  assign n4798 = ~n4796 & ~n4797 ;
  assign n4799 = n147 & ~n2753 ;
  assign n4800 = n160 & ~n2843 ;
  assign n4801 = ~n4799 & ~n4800 ;
  assign n4802 = n4798 & n4801 ;
  assign n4803 = n244 & ~n4802 ;
  assign n4804 = ~n4795 & ~n4803 ;
  assign n4805 = n4787 & n4804 ;
  assign n4806 = x134 & ~n4805 ;
  assign n4807 = n174 & ~n2909 ;
  assign n4808 = n187 & ~n2926 ;
  assign n4809 = ~n4807 & ~n4808 ;
  assign n4810 = n147 & ~n2937 ;
  assign n4811 = n160 & ~n2918 ;
  assign n4812 = ~n4810 & ~n4811 ;
  assign n4813 = n4809 & n4812 ;
  assign n4814 = n244 & ~n4813 ;
  assign n4815 = n174 & ~n2870 ;
  assign n4816 = n187 & ~n2887 ;
  assign n4817 = ~n4815 & ~n4816 ;
  assign n4818 = n147 & ~n2901 ;
  assign n4819 = n160 & ~n2879 ;
  assign n4820 = ~n4818 & ~n4819 ;
  assign n4821 = n4817 & n4820 ;
  assign n4822 = n191 & ~n4821 ;
  assign n4823 = ~n4814 & ~n4822 ;
  assign n4824 = n174 & ~n2945 ;
  assign n4825 = n187 & ~n2962 ;
  assign n4826 = ~n4824 & ~n4825 ;
  assign n4827 = n147 & ~n3010 ;
  assign n4828 = n160 & ~n2954 ;
  assign n4829 = ~n4827 & ~n4828 ;
  assign n4830 = n4826 & n4829 ;
  assign n4831 = n351 & ~n4830 ;
  assign n4832 = n174 & ~n3018 ;
  assign n4833 = n187 & ~n3035 ;
  assign n4834 = ~n4832 & ~n4833 ;
  assign n4835 = n147 & ~n2974 ;
  assign n4836 = n160 & ~n3027 ;
  assign n4837 = ~n4835 & ~n4836 ;
  assign n4838 = n4834 & n4837 ;
  assign n4839 = n298 & ~n4838 ;
  assign n4840 = ~n4831 & ~n4839 ;
  assign n4841 = n4823 & n4840 ;
  assign n4842 = ~x134 & ~n4841 ;
  assign n4843 = ~n4806 & ~n4842 ;
  assign n4846 = n4843 & ~x150 ;
  assign n4847 = ~n4845 & ~n4846 ;
  assign n4848 = n191 & ~n243 ;
  assign n4849 = n244 & ~n350 ;
  assign n4850 = ~n4848 & ~n4849 ;
  assign n4851 = n298 & ~n406 ;
  assign n4852 = ~n297 & n351 ;
  assign n4853 = ~n4851 & ~n4852 ;
  assign n4854 = n4850 & n4853 ;
  assign n4855 = ~x134 & ~n4854 ;
  assign n4856 = ~n190 & n298 ;
  assign n4857 = n191 & ~n458 ;
  assign n4858 = ~n4856 & ~n4857 ;
  assign n4859 = n351 & ~n511 ;
  assign n4860 = n244 & ~n563 ;
  assign n4861 = ~n4859 & ~n4860 ;
  assign n4862 = n4858 & n4861 ;
  assign n4863 = x134 & ~n4862 ;
  assign n4864 = ~n4855 & ~n4863 ;
  assign n4883 = ~n4864 & x151 ;
  assign n4865 = n298 & ~n671 ;
  assign n4866 = n351 & ~n776 ;
  assign n4867 = ~n4865 & ~n4866 ;
  assign n4868 = n191 & ~n831 ;
  assign n4869 = n244 & ~n724 ;
  assign n4870 = ~n4868 & ~n4869 ;
  assign n4871 = n4867 & n4870 ;
  assign n4872 = x134 & ~n4871 ;
  assign n4873 = n191 & ~n619 ;
  assign n4874 = n298 & ~n883 ;
  assign n4875 = ~n4873 & ~n4874 ;
  assign n4876 = n244 & ~n936 ;
  assign n4877 = n351 & ~n988 ;
  assign n4878 = ~n4876 & ~n4877 ;
  assign n4879 = n4875 & n4878 ;
  assign n4880 = ~x134 & ~n4879 ;
  assign n4881 = ~n4872 & ~n4880 ;
  assign n4884 = n4881 & ~x151 ;
  assign n4885 = ~n4883 & ~n4884 ;
  assign n4886 = n191 & ~n1100 ;
  assign n4887 = n244 & ~n1205 ;
  assign n4888 = ~n4886 & ~n4887 ;
  assign n4889 = n298 & ~n1312 ;
  assign n4890 = n351 & ~n1153 ;
  assign n4891 = ~n4889 & ~n4890 ;
  assign n4892 = n4888 & n4891 ;
  assign n4893 = ~x134 & ~n4892 ;
  assign n4894 = n351 & ~n1260 ;
  assign n4895 = n298 & ~n1048 ;
  assign n4896 = ~n4894 & ~n4895 ;
  assign n4897 = n244 & ~n1365 ;
  assign n4898 = n191 & ~n1417 ;
  assign n4899 = ~n4897 & ~n4898 ;
  assign n4900 = n4896 & n4899 ;
  assign n4901 = x134 & ~n4900 ;
  assign n4902 = ~n4893 & ~n4901 ;
  assign n4921 = ~n4902 & x152 ;
  assign n4903 = n298 & ~n1525 ;
  assign n4904 = n351 & ~n1630 ;
  assign n4905 = ~n4903 & ~n4904 ;
  assign n4906 = n191 & ~n1737 ;
  assign n4907 = n244 & ~n1578 ;
  assign n4908 = ~n4906 & ~n4907 ;
  assign n4909 = n4905 & n4908 ;
  assign n4910 = x134 & ~n4909 ;
  assign n4911 = n244 & ~n1685 ;
  assign n4912 = n191 & ~n1473 ;
  assign n4913 = ~n4911 & ~n4912 ;
  assign n4914 = n351 & ~n1790 ;
  assign n4915 = n298 & ~n1842 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4917 = n4913 & n4916 ;
  assign n4918 = ~x134 & ~n4917 ;
  assign n4919 = ~n4910 & ~n4918 ;
  assign n4922 = n4919 & ~x152 ;
  assign n4923 = ~n4921 & ~n4922 ;
  assign n4924 = n191 & ~n1922 ;
  assign n4925 = n244 & ~n1995 ;
  assign n4926 = ~n4924 & ~n4925 ;
  assign n4927 = n298 & ~n2070 ;
  assign n4928 = n351 & ~n1959 ;
  assign n4929 = ~n4927 & ~n4928 ;
  assign n4930 = n4926 & n4929 ;
  assign n4931 = ~x134 & ~n4930 ;
  assign n4932 = n351 & ~n2034 ;
  assign n4933 = n298 & ~n1886 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = n244 & ~n2107 ;
  assign n4936 = n191 & ~n2143 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = n4934 & n4937 ;
  assign n4939 = x134 & ~n4938 ;
  assign n4940 = ~n4931 & ~n4939 ;
  assign n4959 = ~n4940 & x153 ;
  assign n4941 = n298 & ~n2219 ;
  assign n4942 = n351 & ~n2292 ;
  assign n4943 = ~n4941 & ~n4942 ;
  assign n4944 = n191 & ~n2367 ;
  assign n4945 = n244 & ~n2256 ;
  assign n4946 = ~n4944 & ~n4945 ;
  assign n4947 = n4943 & n4946 ;
  assign n4948 = x134 & ~n4947 ;
  assign n4949 = n244 & ~n2331 ;
  assign n4950 = n191 & ~n2183 ;
  assign n4951 = ~n4949 & ~n4950 ;
  assign n4952 = n351 & ~n2404 ;
  assign n4953 = n298 & ~n2440 ;
  assign n4954 = ~n4952 & ~n4953 ;
  assign n4955 = n4951 & n4954 ;
  assign n4956 = ~x134 & ~n4955 ;
  assign n4957 = ~n4948 & ~n4956 ;
  assign n4960 = n4957 & ~x153 ;
  assign n4961 = ~n4959 & ~n4960 ;
  assign n4962 = n244 & ~n2484 ;
  assign n4963 = n191 & ~n2520 ;
  assign n4964 = ~n4962 & ~n4963 ;
  assign n4965 = n351 & ~n2557 ;
  assign n4966 = n298 & ~n2705 ;
  assign n4967 = ~n4965 & ~n4966 ;
  assign n4968 = n4964 & n4967 ;
  assign n4969 = ~x134 & ~n4968 ;
  assign n4970 = n351 & ~n2632 ;
  assign n4971 = n298 & ~n2593 ;
  assign n4972 = ~n4970 & ~n4971 ;
  assign n4973 = n191 & ~n2741 ;
  assign n4974 = n244 & ~n2668 ;
  assign n4975 = ~n4973 & ~n4974 ;
  assign n4976 = n4972 & n4975 ;
  assign n4977 = x134 & ~n4976 ;
  assign n4978 = ~n4969 & ~n4977 ;
  assign n4997 = ~n4978 & x154 ;
  assign n4979 = n351 & ~n2781 ;
  assign n4980 = n298 & ~n2817 ;
  assign n4981 = ~n4979 & ~n4980 ;
  assign n4982 = n244 & ~n2854 ;
  assign n4983 = n191 & ~n3002 ;
  assign n4984 = ~n4982 & ~n4983 ;
  assign n4985 = n4981 & n4984 ;
  assign n4986 = x134 & ~n4985 ;
  assign n4987 = n244 & ~n2929 ;
  assign n4988 = n191 & ~n2890 ;
  assign n4989 = ~n4987 & ~n4988 ;
  assign n4990 = n298 & ~n3038 ;
  assign n4991 = n351 & ~n2965 ;
  assign n4992 = ~n4990 & ~n4991 ;
  assign n4993 = n4989 & n4992 ;
  assign n4994 = ~x134 & ~n4993 ;
  assign n4995 = ~n4986 & ~n4994 ;
  assign n4998 = n4995 & ~x154 ;
  assign n4999 = ~n4997 & ~n4998 ;
  assign n5000 = n191 & ~n3062 ;
  assign n5001 = n244 & ~n3079 ;
  assign n5002 = ~n5000 & ~n5001 ;
  assign n5003 = n298 & ~n3115 ;
  assign n5004 = n351 & ~n3071 ;
  assign n5005 = ~n5003 & ~n5004 ;
  assign n5006 = n5002 & n5005 ;
  assign n5007 = ~x134 & ~n5006 ;
  assign n5008 = n298 & ~n3054 ;
  assign n5009 = n244 & ~n3090 ;
  assign n5010 = ~n5008 & ~n5009 ;
  assign n5011 = n191 & ~n3107 ;
  assign n5012 = n351 & ~n3098 ;
  assign n5013 = ~n5011 & ~n5012 ;
  assign n5014 = n5010 & n5013 ;
  assign n5015 = x134 & ~n5014 ;
  assign n5016 = ~n5007 & ~n5015 ;
  assign n5035 = ~n5016 & x155 ;
  assign n5017 = n298 & ~n3135 ;
  assign n5018 = n351 & ~n3152 ;
  assign n5019 = ~n5017 & ~n5018 ;
  assign n5020 = n191 & ~n3188 ;
  assign n5021 = n244 & ~n3144 ;
  assign n5022 = ~n5020 & ~n5021 ;
  assign n5023 = n5019 & n5022 ;
  assign n5024 = x134 & ~n5023 ;
  assign n5025 = n191 & ~n3127 ;
  assign n5026 = n351 & ~n3163 ;
  assign n5027 = ~n5025 & ~n5026 ;
  assign n5028 = n298 & ~n3180 ;
  assign n5029 = n244 & ~n3171 ;
  assign n5030 = ~n5028 & ~n5029 ;
  assign n5031 = n5027 & n5030 ;
  assign n5032 = ~x134 & ~n5031 ;
  assign n5033 = ~n5024 & ~n5032 ;
  assign n5036 = n5033 & ~x155 ;
  assign n5037 = ~n5035 & ~n5036 ;
  assign n5038 = n191 & ~n3212 ;
  assign n5039 = n244 & ~n3229 ;
  assign n5040 = ~n5038 & ~n5039 ;
  assign n5041 = n298 & ~n3265 ;
  assign n5042 = n351 & ~n3221 ;
  assign n5043 = ~n5041 & ~n5042 ;
  assign n5044 = n5040 & n5043 ;
  assign n5045 = ~x134 & ~n5044 ;
  assign n5046 = n298 & ~n3204 ;
  assign n5047 = n244 & ~n3240 ;
  assign n5048 = ~n5046 & ~n5047 ;
  assign n5049 = n191 & ~n3257 ;
  assign n5050 = n351 & ~n3248 ;
  assign n5051 = ~n5049 & ~n5050 ;
  assign n5052 = n5048 & n5051 ;
  assign n5053 = x134 & ~n5052 ;
  assign n5054 = ~n5045 & ~n5053 ;
  assign n5073 = ~n5054 & x156 ;
  assign n5055 = n298 & ~n3285 ;
  assign n5056 = n351 & ~n3302 ;
  assign n5057 = ~n5055 & ~n5056 ;
  assign n5058 = n191 & ~n3338 ;
  assign n5059 = n244 & ~n3294 ;
  assign n5060 = ~n5058 & ~n5059 ;
  assign n5061 = n5057 & n5060 ;
  assign n5062 = x134 & ~n5061 ;
  assign n5063 = n191 & ~n3277 ;
  assign n5064 = n351 & ~n3313 ;
  assign n5065 = ~n5063 & ~n5064 ;
  assign n5066 = n298 & ~n3330 ;
  assign n5067 = n244 & ~n3321 ;
  assign n5068 = ~n5066 & ~n5067 ;
  assign n5069 = n5065 & n5068 ;
  assign n5070 = ~x134 & ~n5069 ;
  assign n5071 = ~n5062 & ~n5070 ;
  assign n5074 = n5071 & ~x156 ;
  assign n5075 = ~n5073 & ~n5074 ;
  assign n5076 = n191 & ~n3362 ;
  assign n5077 = n244 & ~n3379 ;
  assign n5078 = ~n5076 & ~n5077 ;
  assign n5079 = n298 & ~n3415 ;
  assign n5080 = n351 & ~n3371 ;
  assign n5081 = ~n5079 & ~n5080 ;
  assign n5082 = n5078 & n5081 ;
  assign n5083 = ~x134 & ~n5082 ;
  assign n5084 = n298 & ~n3354 ;
  assign n5085 = n244 & ~n3390 ;
  assign n5086 = ~n5084 & ~n5085 ;
  assign n5087 = n191 & ~n3407 ;
  assign n5088 = n351 & ~n3398 ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5090 = n5086 & n5089 ;
  assign n5091 = x134 & ~n5090 ;
  assign n5092 = ~n5083 & ~n5091 ;
  assign n5111 = ~n5092 & x157 ;
  assign n5093 = n298 & ~n3435 ;
  assign n5094 = n351 & ~n3452 ;
  assign n5095 = ~n5093 & ~n5094 ;
  assign n5096 = n191 & ~n3488 ;
  assign n5097 = n244 & ~n3444 ;
  assign n5098 = ~n5096 & ~n5097 ;
  assign n5099 = n5095 & n5098 ;
  assign n5100 = x134 & ~n5099 ;
  assign n5101 = n191 & ~n3427 ;
  assign n5102 = n351 & ~n3463 ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = n298 & ~n3480 ;
  assign n5105 = n244 & ~n3471 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = n5103 & n5106 ;
  assign n5108 = ~x134 & ~n5107 ;
  assign n5109 = ~n5100 & ~n5108 ;
  assign n5112 = n5109 & ~x157 ;
  assign n5113 = ~n5111 & ~n5112 ;
  assign n5114 = n191 & ~n3512 ;
  assign n5115 = n298 & ~n3565 ;
  assign n5116 = ~n5114 & ~n5115 ;
  assign n5117 = n351 & ~n3521 ;
  assign n5118 = n244 & ~n3529 ;
  assign n5119 = ~n5117 & ~n5118 ;
  assign n5120 = n5116 & n5119 ;
  assign n5121 = ~x134 & ~n5120 ;
  assign n5122 = n244 & ~n3540 ;
  assign n5123 = n351 & ~n3548 ;
  assign n5124 = ~n5122 & ~n5123 ;
  assign n5125 = n191 & ~n3557 ;
  assign n5126 = n298 & ~n3504 ;
  assign n5127 = ~n5125 & ~n5126 ;
  assign n5128 = n5124 & n5127 ;
  assign n5129 = x134 & ~n5128 ;
  assign n5130 = ~n5121 & ~n5129 ;
  assign n5149 = ~n5130 & x158 ;
  assign n5131 = n298 & ~n3585 ;
  assign n5132 = n191 & ~n3638 ;
  assign n5133 = ~n5131 & ~n5132 ;
  assign n5134 = n244 & ~n3594 ;
  assign n5135 = n351 & ~n3602 ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = n5133 & n5136 ;
  assign n5138 = x134 & ~n5137 ;
  assign n5139 = n351 & ~n3613 ;
  assign n5140 = n244 & ~n3621 ;
  assign n5141 = ~n5139 & ~n5140 ;
  assign n5142 = n298 & ~n3630 ;
  assign n5143 = n191 & ~n3577 ;
  assign n5144 = ~n5142 & ~n5143 ;
  assign n5145 = n5141 & n5144 ;
  assign n5146 = ~x134 & ~n5145 ;
  assign n5147 = ~n5138 & ~n5146 ;
  assign n5150 = n5147 & ~x158 ;
  assign n5151 = ~n5149 & ~n5150 ;
  assign n5152 = n191 & ~n3662 ;
  assign n5153 = n298 & ~n3715 ;
  assign n5154 = ~n5152 & ~n5153 ;
  assign n5155 = n351 & ~n3671 ;
  assign n5156 = n244 & ~n3679 ;
  assign n5157 = ~n5155 & ~n5156 ;
  assign n5158 = n5154 & n5157 ;
  assign n5159 = ~x134 & ~n5158 ;
  assign n5160 = n244 & ~n3690 ;
  assign n5161 = n351 & ~n3698 ;
  assign n5162 = ~n5160 & ~n5161 ;
  assign n5163 = n191 & ~n3707 ;
  assign n5164 = n298 & ~n3654 ;
  assign n5165 = ~n5163 & ~n5164 ;
  assign n5166 = n5162 & n5165 ;
  assign n5167 = x134 & ~n5166 ;
  assign n5168 = ~n5159 & ~n5167 ;
  assign n5187 = ~n5168 & x159 ;
  assign n5169 = n298 & ~n3735 ;
  assign n5170 = n191 & ~n3788 ;
  assign n5171 = ~n5169 & ~n5170 ;
  assign n5172 = n244 & ~n3744 ;
  assign n5173 = n351 & ~n3752 ;
  assign n5174 = ~n5172 & ~n5173 ;
  assign n5175 = n5171 & n5174 ;
  assign n5176 = x134 & ~n5175 ;
  assign n5177 = n351 & ~n3763 ;
  assign n5178 = n244 & ~n3771 ;
  assign n5179 = ~n5177 & ~n5178 ;
  assign n5180 = n298 & ~n3780 ;
  assign n5181 = n191 & ~n3727 ;
  assign n5182 = ~n5180 & ~n5181 ;
  assign n5183 = n5179 & n5182 ;
  assign n5184 = ~x134 & ~n5183 ;
  assign n5185 = ~n5176 & ~n5184 ;
  assign n5188 = n5185 & ~x159 ;
  assign n5189 = ~n5187 & ~n5188 ;
  assign n5190 = n191 & ~n3812 ;
  assign n5191 = n298 & ~n3865 ;
  assign n5192 = ~n5190 & ~n5191 ;
  assign n5193 = n351 & ~n3821 ;
  assign n5194 = n244 & ~n3829 ;
  assign n5195 = ~n5193 & ~n5194 ;
  assign n5196 = n5192 & n5195 ;
  assign n5197 = ~x134 & ~n5196 ;
  assign n5198 = n244 & ~n3840 ;
  assign n5199 = n351 & ~n3848 ;
  assign n5200 = ~n5198 & ~n5199 ;
  assign n5201 = n191 & ~n3857 ;
  assign n5202 = n298 & ~n3804 ;
  assign n5203 = ~n5201 & ~n5202 ;
  assign n5204 = n5200 & n5203 ;
  assign n5205 = x134 & ~n5204 ;
  assign n5206 = ~n5197 & ~n5205 ;
  assign n5225 = ~n5206 & x160 ;
  assign n5207 = n298 & ~n3885 ;
  assign n5208 = n191 & ~n3938 ;
  assign n5209 = ~n5207 & ~n5208 ;
  assign n5210 = n244 & ~n3894 ;
  assign n5211 = n351 & ~n3902 ;
  assign n5212 = ~n5210 & ~n5211 ;
  assign n5213 = n5209 & n5212 ;
  assign n5214 = x134 & ~n5213 ;
  assign n5215 = n351 & ~n3913 ;
  assign n5216 = n244 & ~n3921 ;
  assign n5217 = ~n5215 & ~n5216 ;
  assign n5218 = n298 & ~n3930 ;
  assign n5219 = n191 & ~n3877 ;
  assign n5220 = ~n5218 & ~n5219 ;
  assign n5221 = n5217 & n5220 ;
  assign n5222 = ~x134 & ~n5221 ;
  assign n5223 = ~n5214 & ~n5222 ;
  assign n5226 = n5223 & ~x160 ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5228 = n191 & ~n3962 ;
  assign n5229 = n244 & ~n3979 ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5231 = n298 & ~n4015 ;
  assign n5232 = n351 & ~n3971 ;
  assign n5233 = ~n5231 & ~n5232 ;
  assign n5234 = n5230 & n5233 ;
  assign n5235 = ~x134 & ~n5234 ;
  assign n5236 = n244 & ~n3990 ;
  assign n5237 = n351 & ~n3998 ;
  assign n5238 = ~n5236 & ~n5237 ;
  assign n5239 = n191 & ~n4007 ;
  assign n5240 = n298 & ~n3954 ;
  assign n5241 = ~n5239 & ~n5240 ;
  assign n5242 = n5238 & n5241 ;
  assign n5243 = x134 & ~n5242 ;
  assign n5244 = ~n5235 & ~n5243 ;
  assign n5263 = ~n5244 & x161 ;
  assign n5245 = n298 & ~n4035 ;
  assign n5246 = n351 & ~n4052 ;
  assign n5247 = ~n5245 & ~n5246 ;
  assign n5248 = n191 & ~n4088 ;
  assign n5249 = n244 & ~n4044 ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = n5247 & n5250 ;
  assign n5252 = x134 & ~n5251 ;
  assign n5253 = n351 & ~n4063 ;
  assign n5254 = n244 & ~n4071 ;
  assign n5255 = ~n5253 & ~n5254 ;
  assign n5256 = n298 & ~n4080 ;
  assign n5257 = n191 & ~n4027 ;
  assign n5258 = ~n5256 & ~n5257 ;
  assign n5259 = n5255 & n5258 ;
  assign n5260 = ~x134 & ~n5259 ;
  assign n5261 = ~n5252 & ~n5260 ;
  assign n5264 = n5261 & ~x161 ;
  assign n5265 = ~n5263 & ~n5264 ;
  assign n5266 = n191 & ~n4112 ;
  assign n5267 = n244 & ~n4129 ;
  assign n5268 = ~n5266 & ~n5267 ;
  assign n5269 = n298 & ~n4165 ;
  assign n5270 = n351 & ~n4121 ;
  assign n5271 = ~n5269 & ~n5270 ;
  assign n5272 = n5268 & n5271 ;
  assign n5273 = ~x134 & ~n5272 ;
  assign n5274 = n244 & ~n4140 ;
  assign n5275 = n351 & ~n4148 ;
  assign n5276 = ~n5274 & ~n5275 ;
  assign n5277 = n191 & ~n4157 ;
  assign n5278 = n298 & ~n4104 ;
  assign n5279 = ~n5277 & ~n5278 ;
  assign n5280 = n5276 & n5279 ;
  assign n5281 = x134 & ~n5280 ;
  assign n5282 = ~n5273 & ~n5281 ;
  assign n5301 = ~n5282 & x162 ;
  assign n5283 = n298 & ~n4185 ;
  assign n5284 = n351 & ~n4202 ;
  assign n5285 = ~n5283 & ~n5284 ;
  assign n5286 = n191 & ~n4238 ;
  assign n5287 = n244 & ~n4194 ;
  assign n5288 = ~n5286 & ~n5287 ;
  assign n5289 = n5285 & n5288 ;
  assign n5290 = x134 & ~n5289 ;
  assign n5291 = n351 & ~n4213 ;
  assign n5292 = n244 & ~n4221 ;
  assign n5293 = ~n5291 & ~n5292 ;
  assign n5294 = n298 & ~n4230 ;
  assign n5295 = n191 & ~n4177 ;
  assign n5296 = ~n5294 & ~n5295 ;
  assign n5297 = n5293 & n5296 ;
  assign n5298 = ~x134 & ~n5297 ;
  assign n5299 = ~n5290 & ~n5298 ;
  assign n5302 = n5299 & ~x162 ;
  assign n5303 = ~n5301 & ~n5302 ;
  assign n5304 = n191 & ~n4262 ;
  assign n5305 = n244 & ~n4279 ;
  assign n5306 = ~n5304 & ~n5305 ;
  assign n5307 = n298 & ~n4315 ;
  assign n5308 = n351 & ~n4271 ;
  assign n5309 = ~n5307 & ~n5308 ;
  assign n5310 = n5306 & n5309 ;
  assign n5311 = ~x134 & ~n5310 ;
  assign n5312 = n244 & ~n4290 ;
  assign n5313 = n351 & ~n4298 ;
  assign n5314 = ~n5312 & ~n5313 ;
  assign n5315 = n191 & ~n4307 ;
  assign n5316 = n298 & ~n4254 ;
  assign n5317 = ~n5315 & ~n5316 ;
  assign n5318 = n5314 & n5317 ;
  assign n5319 = x134 & ~n5318 ;
  assign n5320 = ~n5311 & ~n5319 ;
  assign n5339 = ~n5320 & x163 ;
  assign n5321 = n298 & ~n4335 ;
  assign n5322 = n351 & ~n4352 ;
  assign n5323 = ~n5321 & ~n5322 ;
  assign n5324 = n191 & ~n4388 ;
  assign n5325 = n244 & ~n4344 ;
  assign n5326 = ~n5324 & ~n5325 ;
  assign n5327 = n5323 & n5326 ;
  assign n5328 = x134 & ~n5327 ;
  assign n5329 = n351 & ~n4363 ;
  assign n5330 = n244 & ~n4371 ;
  assign n5331 = ~n5329 & ~n5330 ;
  assign n5332 = n298 & ~n4380 ;
  assign n5333 = n191 & ~n4327 ;
  assign n5334 = ~n5332 & ~n5333 ;
  assign n5335 = n5331 & n5334 ;
  assign n5336 = ~x134 & ~n5335 ;
  assign n5337 = ~n5328 & ~n5336 ;
  assign n5340 = n5337 & ~x163 ;
  assign n5341 = ~n5339 & ~n5340 ;
  assign n5342 = n191 & ~n4412 ;
  assign n5343 = n244 & ~n4429 ;
  assign n5344 = ~n5342 & ~n5343 ;
  assign n5345 = n298 & ~n4465 ;
  assign n5346 = n351 & ~n4421 ;
  assign n5347 = ~n5345 & ~n5346 ;
  assign n5348 = n5344 & n5347 ;
  assign n5349 = ~x134 & ~n5348 ;
  assign n5350 = n244 & ~n4440 ;
  assign n5351 = n351 & ~n4448 ;
  assign n5352 = ~n5350 & ~n5351 ;
  assign n5353 = n191 & ~n4457 ;
  assign n5354 = n298 & ~n4404 ;
  assign n5355 = ~n5353 & ~n5354 ;
  assign n5356 = n5352 & n5355 ;
  assign n5357 = x134 & ~n5356 ;
  assign n5358 = ~n5349 & ~n5357 ;
  assign n5377 = ~n5358 & x164 ;
  assign n5359 = n298 & ~n4485 ;
  assign n5360 = n351 & ~n4502 ;
  assign n5361 = ~n5359 & ~n5360 ;
  assign n5362 = n191 & ~n4538 ;
  assign n5363 = n244 & ~n4494 ;
  assign n5364 = ~n5362 & ~n5363 ;
  assign n5365 = n5361 & n5364 ;
  assign n5366 = x134 & ~n5365 ;
  assign n5367 = n351 & ~n4513 ;
  assign n5368 = n244 & ~n4521 ;
  assign n5369 = ~n5367 & ~n5368 ;
  assign n5370 = n298 & ~n4530 ;
  assign n5371 = n191 & ~n4477 ;
  assign n5372 = ~n5370 & ~n5371 ;
  assign n5373 = n5369 & n5372 ;
  assign n5374 = ~x134 & ~n5373 ;
  assign n5375 = ~n5366 & ~n5374 ;
  assign n5378 = n5375 & ~x164 ;
  assign n5379 = ~n5377 & ~n5378 ;
  assign n5380 = n191 & ~n4562 ;
  assign n5381 = n244 & ~n4579 ;
  assign n5382 = ~n5380 & ~n5381 ;
  assign n5383 = n298 & ~n4615 ;
  assign n5384 = n351 & ~n4571 ;
  assign n5385 = ~n5383 & ~n5384 ;
  assign n5386 = n5382 & n5385 ;
  assign n5387 = ~x134 & ~n5386 ;
  assign n5388 = n244 & ~n4590 ;
  assign n5389 = n351 & ~n4598 ;
  assign n5390 = ~n5388 & ~n5389 ;
  assign n5391 = n191 & ~n4607 ;
  assign n5392 = n298 & ~n4554 ;
  assign n5393 = ~n5391 & ~n5392 ;
  assign n5394 = n5390 & n5393 ;
  assign n5395 = x134 & ~n5394 ;
  assign n5396 = ~n5387 & ~n5395 ;
  assign n5415 = ~n5396 & x165 ;
  assign n5397 = n298 & ~n4635 ;
  assign n5398 = n351 & ~n4652 ;
  assign n5399 = ~n5397 & ~n5398 ;
  assign n5400 = n191 & ~n4688 ;
  assign n5401 = n244 & ~n4644 ;
  assign n5402 = ~n5400 & ~n5401 ;
  assign n5403 = n5399 & n5402 ;
  assign n5404 = x134 & ~n5403 ;
  assign n5405 = n351 & ~n4663 ;
  assign n5406 = n244 & ~n4671 ;
  assign n5407 = ~n5405 & ~n5406 ;
  assign n5408 = n298 & ~n4680 ;
  assign n5409 = n191 & ~n4627 ;
  assign n5410 = ~n5408 & ~n5409 ;
  assign n5411 = n5407 & n5410 ;
  assign n5412 = ~x134 & ~n5411 ;
  assign n5413 = ~n5404 & ~n5412 ;
  assign n5416 = n5413 & ~x165 ;
  assign n5417 = ~n5415 & ~n5416 ;
  assign n5418 = n191 & ~n4712 ;
  assign n5419 = n244 & ~n4729 ;
  assign n5420 = ~n5418 & ~n5419 ;
  assign n5421 = n298 & ~n4765 ;
  assign n5422 = n351 & ~n4721 ;
  assign n5423 = ~n5421 & ~n5422 ;
  assign n5424 = n5420 & n5423 ;
  assign n5425 = ~x134 & ~n5424 ;
  assign n5426 = n244 & ~n4740 ;
  assign n5427 = n351 & ~n4748 ;
  assign n5428 = ~n5426 & ~n5427 ;
  assign n5429 = n191 & ~n4757 ;
  assign n5430 = n298 & ~n4704 ;
  assign n5431 = ~n5429 & ~n5430 ;
  assign n5432 = n5428 & n5431 ;
  assign n5433 = x134 & ~n5432 ;
  assign n5434 = ~n5425 & ~n5433 ;
  assign n5453 = ~n5434 & x166 ;
  assign n5435 = n298 & ~n4785 ;
  assign n5436 = n351 & ~n4802 ;
  assign n5437 = ~n5435 & ~n5436 ;
  assign n5438 = n191 & ~n4838 ;
  assign n5439 = n244 & ~n4794 ;
  assign n5440 = ~n5438 & ~n5439 ;
  assign n5441 = n5437 & n5440 ;
  assign n5442 = x134 & ~n5441 ;
  assign n5443 = n351 & ~n4813 ;
  assign n5444 = n244 & ~n4821 ;
  assign n5445 = ~n5443 & ~n5444 ;
  assign n5446 = n298 & ~n4830 ;
  assign n5447 = n191 & ~n4777 ;
  assign n5448 = ~n5446 & ~n5447 ;
  assign n5449 = n5445 & n5448 ;
  assign n5450 = ~x134 & ~n5449 ;
  assign n5451 = ~n5442 & ~n5450 ;
  assign n5454 = n5451 & ~x166 ;
  assign n5455 = ~n5453 & ~n5454 ;
  assign n5456 = n191 & ~n350 ;
  assign n5457 = n244 & ~n297 ;
  assign n5458 = ~n5456 & ~n5457 ;
  assign n5459 = n298 & ~n458 ;
  assign n5460 = n351 & ~n406 ;
  assign n5461 = ~n5459 & ~n5460 ;
  assign n5462 = n5458 & n5461 ;
  assign n5463 = ~x134 & ~n5462 ;
  assign n5464 = ~n190 & n351 ;
  assign n5465 = ~n243 & n298 ;
  assign n5466 = ~n5464 & ~n5465 ;
  assign n5467 = n244 & ~n511 ;
  assign n5468 = n191 & ~n563 ;
  assign n5469 = ~n5467 & ~n5468 ;
  assign n5470 = n5466 & n5469 ;
  assign n5471 = x134 & ~n5470 ;
  assign n5472 = ~n5463 & ~n5471 ;
  assign n5491 = ~n5472 & x167 ;
  assign n5473 = n298 & ~n776 ;
  assign n5474 = n351 & ~n724 ;
  assign n5475 = ~n5473 & ~n5474 ;
  assign n5476 = n191 & ~n883 ;
  assign n5477 = n244 & ~n831 ;
  assign n5478 = ~n5476 & ~n5477 ;
  assign n5479 = n5475 & n5478 ;
  assign n5480 = x134 & ~n5479 ;
  assign n5481 = n244 & ~n619 ;
  assign n5482 = n191 & ~n671 ;
  assign n5483 = ~n5481 & ~n5482 ;
  assign n5484 = n351 & ~n936 ;
  assign n5485 = n298 & ~n988 ;
  assign n5486 = ~n5484 & ~n5485 ;
  assign n5487 = n5483 & n5486 ;
  assign n5488 = ~x134 & ~n5487 ;
  assign n5489 = ~n5480 & ~n5488 ;
  assign n5492 = n5489 & ~x167 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = n191 & ~n1205 ;
  assign n5495 = n244 & ~n1153 ;
  assign n5496 = ~n5494 & ~n5495 ;
  assign n5497 = n298 & ~n1417 ;
  assign n5498 = n351 & ~n1312 ;
  assign n5499 = ~n5497 & ~n5498 ;
  assign n5500 = n5496 & n5499 ;
  assign n5501 = ~x134 & ~n5500 ;
  assign n5502 = n244 & ~n1260 ;
  assign n5503 = n351 & ~n1048 ;
  assign n5504 = ~n5502 & ~n5503 ;
  assign n5505 = n191 & ~n1365 ;
  assign n5506 = n298 & ~n1100 ;
  assign n5507 = ~n5505 & ~n5506 ;
  assign n5508 = n5504 & n5507 ;
  assign n5509 = x134 & ~n5508 ;
  assign n5510 = ~n5501 & ~n5509 ;
  assign n5529 = ~n5510 & x168 ;
  assign n5511 = n298 & ~n1630 ;
  assign n5512 = n351 & ~n1578 ;
  assign n5513 = ~n5511 & ~n5512 ;
  assign n5514 = n191 & ~n1842 ;
  assign n5515 = n244 & ~n1737 ;
  assign n5516 = ~n5514 & ~n5515 ;
  assign n5517 = n5513 & n5516 ;
  assign n5518 = x134 & ~n5517 ;
  assign n5519 = n351 & ~n1685 ;
  assign n5520 = n244 & ~n1473 ;
  assign n5521 = ~n5519 & ~n5520 ;
  assign n5522 = n298 & ~n1790 ;
  assign n5523 = n191 & ~n1525 ;
  assign n5524 = ~n5522 & ~n5523 ;
  assign n5525 = n5521 & n5524 ;
  assign n5526 = ~x134 & ~n5525 ;
  assign n5527 = ~n5518 & ~n5526 ;
  assign n5530 = n5527 & ~x168 ;
  assign n5531 = ~n5529 & ~n5530 ;
  assign n5532 = n191 & ~n1995 ;
  assign n5533 = n244 & ~n1959 ;
  assign n5534 = ~n5532 & ~n5533 ;
  assign n5535 = n298 & ~n2143 ;
  assign n5536 = n351 & ~n2070 ;
  assign n5537 = ~n5535 & ~n5536 ;
  assign n5538 = n5534 & n5537 ;
  assign n5539 = ~x134 & ~n5538 ;
  assign n5540 = n244 & ~n2034 ;
  assign n5541 = n351 & ~n1886 ;
  assign n5542 = ~n5540 & ~n5541 ;
  assign n5543 = n191 & ~n2107 ;
  assign n5544 = n298 & ~n1922 ;
  assign n5545 = ~n5543 & ~n5544 ;
  assign n5546 = n5542 & n5545 ;
  assign n5547 = x134 & ~n5546 ;
  assign n5548 = ~n5539 & ~n5547 ;
  assign n5567 = ~n5548 & x169 ;
  assign n5549 = n298 & ~n2292 ;
  assign n5550 = n351 & ~n2256 ;
  assign n5551 = ~n5549 & ~n5550 ;
  assign n5552 = n191 & ~n2440 ;
  assign n5553 = n244 & ~n2367 ;
  assign n5554 = ~n5552 & ~n5553 ;
  assign n5555 = n5551 & n5554 ;
  assign n5556 = x134 & ~n5555 ;
  assign n5557 = n351 & ~n2331 ;
  assign n5558 = n244 & ~n2183 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5560 = n298 & ~n2404 ;
  assign n5561 = n191 & ~n2219 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5563 = n5559 & n5562 ;
  assign n5564 = ~x134 & ~n5563 ;
  assign n5565 = ~n5556 & ~n5564 ;
  assign n5568 = n5565 & ~x169 ;
  assign n5569 = ~n5567 & ~n5568 ;
  assign n5570 = n191 & ~n2484 ;
  assign n5571 = n298 & ~n2741 ;
  assign n5572 = ~n5570 & ~n5571 ;
  assign n5573 = n244 & ~n2557 ;
  assign n5574 = n351 & ~n2705 ;
  assign n5575 = ~n5573 & ~n5574 ;
  assign n5576 = n5572 & n5575 ;
  assign n5577 = ~x134 & ~n5576 ;
  assign n5578 = n244 & ~n2632 ;
  assign n5579 = n298 & ~n2520 ;
  assign n5580 = ~n5578 & ~n5579 ;
  assign n5581 = n191 & ~n2668 ;
  assign n5582 = n351 & ~n2593 ;
  assign n5583 = ~n5581 & ~n5582 ;
  assign n5584 = n5580 & n5583 ;
  assign n5585 = x134 & ~n5584 ;
  assign n5586 = ~n5577 & ~n5585 ;
  assign n5605 = ~n5586 & x170 ;
  assign n5587 = n298 & ~n2781 ;
  assign n5588 = n191 & ~n3038 ;
  assign n5589 = ~n5587 & ~n5588 ;
  assign n5590 = n351 & ~n2854 ;
  assign n5591 = n244 & ~n3002 ;
  assign n5592 = ~n5590 & ~n5591 ;
  assign n5593 = n5589 & n5592 ;
  assign n5594 = x134 & ~n5593 ;
  assign n5595 = n351 & ~n2929 ;
  assign n5596 = n191 & ~n2817 ;
  assign n5597 = ~n5595 & ~n5596 ;
  assign n5598 = n298 & ~n2965 ;
  assign n5599 = n244 & ~n2890 ;
  assign n5600 = ~n5598 & ~n5599 ;
  assign n5601 = n5597 & n5600 ;
  assign n5602 = ~x134 & ~n5601 ;
  assign n5603 = ~n5594 & ~n5602 ;
  assign n5606 = n5603 & ~x170 ;
  assign n5607 = ~n5605 & ~n5606 ;
  assign n5608 = n191 & ~n3079 ;
  assign n5609 = n244 & ~n3071 ;
  assign n5610 = ~n5608 & ~n5609 ;
  assign n5611 = n298 & ~n3107 ;
  assign n5612 = n351 & ~n3115 ;
  assign n5613 = ~n5611 & ~n5612 ;
  assign n5614 = n5610 & n5613 ;
  assign n5615 = ~x134 & ~n5614 ;
  assign n5616 = n351 & ~n3054 ;
  assign n5617 = n298 & ~n3062 ;
  assign n5618 = ~n5616 & ~n5617 ;
  assign n5619 = n244 & ~n3098 ;
  assign n5620 = n191 & ~n3090 ;
  assign n5621 = ~n5619 & ~n5620 ;
  assign n5622 = n5618 & n5621 ;
  assign n5623 = x134 & ~n5622 ;
  assign n5624 = ~n5615 & ~n5623 ;
  assign n5643 = ~n5624 & x171 ;
  assign n5625 = n298 & ~n3152 ;
  assign n5626 = n351 & ~n3144 ;
  assign n5627 = ~n5625 & ~n5626 ;
  assign n5628 = n191 & ~n3180 ;
  assign n5629 = n244 & ~n3188 ;
  assign n5630 = ~n5628 & ~n5629 ;
  assign n5631 = n5627 & n5630 ;
  assign n5632 = x134 & ~n5631 ;
  assign n5633 = n244 & ~n3127 ;
  assign n5634 = n191 & ~n3135 ;
  assign n5635 = ~n5633 & ~n5634 ;
  assign n5636 = n351 & ~n3171 ;
  assign n5637 = n298 & ~n3163 ;
  assign n5638 = ~n5636 & ~n5637 ;
  assign n5639 = n5635 & n5638 ;
  assign n5640 = ~x134 & ~n5639 ;
  assign n5641 = ~n5632 & ~n5640 ;
  assign n5644 = n5641 & ~x171 ;
  assign n5645 = ~n5643 & ~n5644 ;
  assign n5646 = n191 & ~n3229 ;
  assign n5647 = n244 & ~n3221 ;
  assign n5648 = ~n5646 & ~n5647 ;
  assign n5649 = n298 & ~n3257 ;
  assign n5650 = n351 & ~n3265 ;
  assign n5651 = ~n5649 & ~n5650 ;
  assign n5652 = n5648 & n5651 ;
  assign n5653 = ~x134 & ~n5652 ;
  assign n5654 = n351 & ~n3204 ;
  assign n5655 = n298 & ~n3212 ;
  assign n5656 = ~n5654 & ~n5655 ;
  assign n5657 = n244 & ~n3248 ;
  assign n5658 = n191 & ~n3240 ;
  assign n5659 = ~n5657 & ~n5658 ;
  assign n5660 = n5656 & n5659 ;
  assign n5661 = x134 & ~n5660 ;
  assign n5662 = ~n5653 & ~n5661 ;
  assign n5681 = ~n5662 & x172 ;
  assign n5663 = n298 & ~n3302 ;
  assign n5664 = n351 & ~n3294 ;
  assign n5665 = ~n5663 & ~n5664 ;
  assign n5666 = n191 & ~n3330 ;
  assign n5667 = n244 & ~n3338 ;
  assign n5668 = ~n5666 & ~n5667 ;
  assign n5669 = n5665 & n5668 ;
  assign n5670 = x134 & ~n5669 ;
  assign n5671 = n244 & ~n3277 ;
  assign n5672 = n191 & ~n3285 ;
  assign n5673 = ~n5671 & ~n5672 ;
  assign n5674 = n351 & ~n3321 ;
  assign n5675 = n298 & ~n3313 ;
  assign n5676 = ~n5674 & ~n5675 ;
  assign n5677 = n5673 & n5676 ;
  assign n5678 = ~x134 & ~n5677 ;
  assign n5679 = ~n5670 & ~n5678 ;
  assign n5682 = n5679 & ~x172 ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5684 = n191 & ~n3379 ;
  assign n5685 = n244 & ~n3371 ;
  assign n5686 = ~n5684 & ~n5685 ;
  assign n5687 = n298 & ~n3407 ;
  assign n5688 = n351 & ~n3415 ;
  assign n5689 = ~n5687 & ~n5688 ;
  assign n5690 = n5686 & n5689 ;
  assign n5691 = ~x134 & ~n5690 ;
  assign n5692 = n351 & ~n3354 ;
  assign n5693 = n298 & ~n3362 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = n244 & ~n3398 ;
  assign n5696 = n191 & ~n3390 ;
  assign n5697 = ~n5695 & ~n5696 ;
  assign n5698 = n5694 & n5697 ;
  assign n5699 = x134 & ~n5698 ;
  assign n5700 = ~n5691 & ~n5699 ;
  assign n5719 = ~n5700 & x173 ;
  assign n5701 = n298 & ~n3452 ;
  assign n5702 = n351 & ~n3444 ;
  assign n5703 = ~n5701 & ~n5702 ;
  assign n5704 = n191 & ~n3480 ;
  assign n5705 = n244 & ~n3488 ;
  assign n5706 = ~n5704 & ~n5705 ;
  assign n5707 = n5703 & n5706 ;
  assign n5708 = x134 & ~n5707 ;
  assign n5709 = n244 & ~n3427 ;
  assign n5710 = n191 & ~n3435 ;
  assign n5711 = ~n5709 & ~n5710 ;
  assign n5712 = n351 & ~n3471 ;
  assign n5713 = n298 & ~n3463 ;
  assign n5714 = ~n5712 & ~n5713 ;
  assign n5715 = n5711 & n5714 ;
  assign n5716 = ~x134 & ~n5715 ;
  assign n5717 = ~n5708 & ~n5716 ;
  assign n5720 = n5717 & ~x173 ;
  assign n5721 = ~n5719 & ~n5720 ;
  assign n5722 = n351 & ~n3565 ;
  assign n5723 = n298 & ~n3557 ;
  assign n5724 = ~n5722 & ~n5723 ;
  assign n5725 = n244 & ~n3521 ;
  assign n5726 = n191 & ~n3529 ;
  assign n5727 = ~n5725 & ~n5726 ;
  assign n5728 = n5724 & n5727 ;
  assign n5729 = ~x134 & ~n5728 ;
  assign n5730 = n191 & ~n3540 ;
  assign n5731 = n244 & ~n3548 ;
  assign n5732 = ~n5730 & ~n5731 ;
  assign n5733 = n298 & ~n3512 ;
  assign n5734 = n351 & ~n3504 ;
  assign n5735 = ~n5733 & ~n5734 ;
  assign n5736 = n5732 & n5735 ;
  assign n5737 = x134 & ~n5736 ;
  assign n5738 = ~n5729 & ~n5737 ;
  assign n5757 = ~n5738 & x174 ;
  assign n5739 = n244 & ~n3638 ;
  assign n5740 = n191 & ~n3630 ;
  assign n5741 = ~n5739 & ~n5740 ;
  assign n5742 = n351 & ~n3594 ;
  assign n5743 = n298 & ~n3602 ;
  assign n5744 = ~n5742 & ~n5743 ;
  assign n5745 = n5741 & n5744 ;
  assign n5746 = x134 & ~n5745 ;
  assign n5747 = n298 & ~n3613 ;
  assign n5748 = n351 & ~n3621 ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5750 = n191 & ~n3585 ;
  assign n5751 = n244 & ~n3577 ;
  assign n5752 = ~n5750 & ~n5751 ;
  assign n5753 = n5749 & n5752 ;
  assign n5754 = ~x134 & ~n5753 ;
  assign n5755 = ~n5746 & ~n5754 ;
  assign n5758 = n5755 & ~x174 ;
  assign n5759 = ~n5757 & ~n5758 ;
  assign n5760 = n351 & ~n3715 ;
  assign n5761 = n298 & ~n3707 ;
  assign n5762 = ~n5760 & ~n5761 ;
  assign n5763 = n244 & ~n3671 ;
  assign n5764 = n191 & ~n3679 ;
  assign n5765 = ~n5763 & ~n5764 ;
  assign n5766 = n5762 & n5765 ;
  assign n5767 = ~x134 & ~n5766 ;
  assign n5768 = n191 & ~n3690 ;
  assign n5769 = n244 & ~n3698 ;
  assign n5770 = ~n5768 & ~n5769 ;
  assign n5771 = n298 & ~n3662 ;
  assign n5772 = n351 & ~n3654 ;
  assign n5773 = ~n5771 & ~n5772 ;
  assign n5774 = n5770 & n5773 ;
  assign n5775 = x134 & ~n5774 ;
  assign n5776 = ~n5767 & ~n5775 ;
  assign n5795 = ~n5776 & x175 ;
  assign n5777 = n244 & ~n3788 ;
  assign n5778 = n191 & ~n3780 ;
  assign n5779 = ~n5777 & ~n5778 ;
  assign n5780 = n351 & ~n3744 ;
  assign n5781 = n298 & ~n3752 ;
  assign n5782 = ~n5780 & ~n5781 ;
  assign n5783 = n5779 & n5782 ;
  assign n5784 = x134 & ~n5783 ;
  assign n5785 = n298 & ~n3763 ;
  assign n5786 = n351 & ~n3771 ;
  assign n5787 = ~n5785 & ~n5786 ;
  assign n5788 = n191 & ~n3735 ;
  assign n5789 = n244 & ~n3727 ;
  assign n5790 = ~n5788 & ~n5789 ;
  assign n5791 = n5787 & n5790 ;
  assign n5792 = ~x134 & ~n5791 ;
  assign n5793 = ~n5784 & ~n5792 ;
  assign n5796 = n5793 & ~x175 ;
  assign n5797 = ~n5795 & ~n5796 ;
  assign n5798 = n351 & ~n3865 ;
  assign n5799 = n298 & ~n3857 ;
  assign n5800 = ~n5798 & ~n5799 ;
  assign n5801 = n244 & ~n3821 ;
  assign n5802 = n191 & ~n3829 ;
  assign n5803 = ~n5801 & ~n5802 ;
  assign n5804 = n5800 & n5803 ;
  assign n5805 = ~x134 & ~n5804 ;
  assign n5806 = n191 & ~n3840 ;
  assign n5807 = n244 & ~n3848 ;
  assign n5808 = ~n5806 & ~n5807 ;
  assign n5809 = n298 & ~n3812 ;
  assign n5810 = n351 & ~n3804 ;
  assign n5811 = ~n5809 & ~n5810 ;
  assign n5812 = n5808 & n5811 ;
  assign n5813 = x134 & ~n5812 ;
  assign n5814 = ~n5805 & ~n5813 ;
  assign n5833 = ~n5814 & x176 ;
  assign n5815 = n244 & ~n3938 ;
  assign n5816 = n191 & ~n3930 ;
  assign n5817 = ~n5815 & ~n5816 ;
  assign n5818 = n351 & ~n3894 ;
  assign n5819 = n298 & ~n3902 ;
  assign n5820 = ~n5818 & ~n5819 ;
  assign n5821 = n5817 & n5820 ;
  assign n5822 = x134 & ~n5821 ;
  assign n5823 = n298 & ~n3913 ;
  assign n5824 = n351 & ~n3921 ;
  assign n5825 = ~n5823 & ~n5824 ;
  assign n5826 = n191 & ~n3885 ;
  assign n5827 = n244 & ~n3877 ;
  assign n5828 = ~n5826 & ~n5827 ;
  assign n5829 = n5825 & n5828 ;
  assign n5830 = ~x134 & ~n5829 ;
  assign n5831 = ~n5822 & ~n5830 ;
  assign n5834 = n5831 & ~x176 ;
  assign n5835 = ~n5833 & ~n5834 ;
  assign n5836 = n191 & ~n3979 ;
  assign n5837 = n244 & ~n3971 ;
  assign n5838 = ~n5836 & ~n5837 ;
  assign n5839 = n298 & ~n4007 ;
  assign n5840 = n351 & ~n4015 ;
  assign n5841 = ~n5839 & ~n5840 ;
  assign n5842 = n5838 & n5841 ;
  assign n5843 = ~x134 & ~n5842 ;
  assign n5844 = n191 & ~n3990 ;
  assign n5845 = n244 & ~n3998 ;
  assign n5846 = ~n5844 & ~n5845 ;
  assign n5847 = n298 & ~n3962 ;
  assign n5848 = n351 & ~n3954 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = n5846 & n5849 ;
  assign n5851 = x134 & ~n5850 ;
  assign n5852 = ~n5843 & ~n5851 ;
  assign n5871 = ~n5852 & x177 ;
  assign n5853 = n298 & ~n4052 ;
  assign n5854 = n351 & ~n4044 ;
  assign n5855 = ~n5853 & ~n5854 ;
  assign n5856 = n191 & ~n4080 ;
  assign n5857 = n244 & ~n4088 ;
  assign n5858 = ~n5856 & ~n5857 ;
  assign n5859 = n5855 & n5858 ;
  assign n5860 = x134 & ~n5859 ;
  assign n5861 = n298 & ~n4063 ;
  assign n5862 = n351 & ~n4071 ;
  assign n5863 = ~n5861 & ~n5862 ;
  assign n5864 = n191 & ~n4035 ;
  assign n5865 = n244 & ~n4027 ;
  assign n5866 = ~n5864 & ~n5865 ;
  assign n5867 = n5863 & n5866 ;
  assign n5868 = ~x134 & ~n5867 ;
  assign n5869 = ~n5860 & ~n5868 ;
  assign n5872 = n5869 & ~x177 ;
  assign n5873 = ~n5871 & ~n5872 ;
  assign n5874 = n191 & ~n4129 ;
  assign n5875 = n244 & ~n4121 ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = n298 & ~n4157 ;
  assign n5878 = n351 & ~n4165 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = n5876 & n5879 ;
  assign n5881 = ~x134 & ~n5880 ;
  assign n5882 = n191 & ~n4140 ;
  assign n5883 = n244 & ~n4148 ;
  assign n5884 = ~n5882 & ~n5883 ;
  assign n5885 = n298 & ~n4112 ;
  assign n5886 = n351 & ~n4104 ;
  assign n5887 = ~n5885 & ~n5886 ;
  assign n5888 = n5884 & n5887 ;
  assign n5889 = x134 & ~n5888 ;
  assign n5890 = ~n5881 & ~n5889 ;
  assign n5909 = ~n5890 & x178 ;
  assign n5891 = n298 & ~n4202 ;
  assign n5892 = n351 & ~n4194 ;
  assign n5893 = ~n5891 & ~n5892 ;
  assign n5894 = n191 & ~n4230 ;
  assign n5895 = n244 & ~n4238 ;
  assign n5896 = ~n5894 & ~n5895 ;
  assign n5897 = n5893 & n5896 ;
  assign n5898 = x134 & ~n5897 ;
  assign n5899 = n298 & ~n4213 ;
  assign n5900 = n351 & ~n4221 ;
  assign n5901 = ~n5899 & ~n5900 ;
  assign n5902 = n191 & ~n4185 ;
  assign n5903 = n244 & ~n4177 ;
  assign n5904 = ~n5902 & ~n5903 ;
  assign n5905 = n5901 & n5904 ;
  assign n5906 = ~x134 & ~n5905 ;
  assign n5907 = ~n5898 & ~n5906 ;
  assign n5910 = n5907 & ~x178 ;
  assign n5911 = ~n5909 & ~n5910 ;
  assign n5912 = n191 & ~n4279 ;
  assign n5913 = n244 & ~n4271 ;
  assign n5914 = ~n5912 & ~n5913 ;
  assign n5915 = n298 & ~n4307 ;
  assign n5916 = n351 & ~n4315 ;
  assign n5917 = ~n5915 & ~n5916 ;
  assign n5918 = n5914 & n5917 ;
  assign n5919 = ~x134 & ~n5918 ;
  assign n5920 = n191 & ~n4290 ;
  assign n5921 = n244 & ~n4298 ;
  assign n5922 = ~n5920 & ~n5921 ;
  assign n5923 = n298 & ~n4262 ;
  assign n5924 = n351 & ~n4254 ;
  assign n5925 = ~n5923 & ~n5924 ;
  assign n5926 = n5922 & n5925 ;
  assign n5927 = x134 & ~n5926 ;
  assign n5928 = ~n5919 & ~n5927 ;
  assign n5947 = ~n5928 & x179 ;
  assign n5929 = n298 & ~n4352 ;
  assign n5930 = n351 & ~n4344 ;
  assign n5931 = ~n5929 & ~n5930 ;
  assign n5932 = n191 & ~n4380 ;
  assign n5933 = n244 & ~n4388 ;
  assign n5934 = ~n5932 & ~n5933 ;
  assign n5935 = n5931 & n5934 ;
  assign n5936 = x134 & ~n5935 ;
  assign n5937 = n298 & ~n4363 ;
  assign n5938 = n351 & ~n4371 ;
  assign n5939 = ~n5937 & ~n5938 ;
  assign n5940 = n191 & ~n4335 ;
  assign n5941 = n244 & ~n4327 ;
  assign n5942 = ~n5940 & ~n5941 ;
  assign n5943 = n5939 & n5942 ;
  assign n5944 = ~x134 & ~n5943 ;
  assign n5945 = ~n5936 & ~n5944 ;
  assign n5948 = n5945 & ~x179 ;
  assign n5949 = ~n5947 & ~n5948 ;
  assign n5950 = n191 & ~n4429 ;
  assign n5951 = n244 & ~n4421 ;
  assign n5952 = ~n5950 & ~n5951 ;
  assign n5953 = n298 & ~n4457 ;
  assign n5954 = n351 & ~n4465 ;
  assign n5955 = ~n5953 & ~n5954 ;
  assign n5956 = n5952 & n5955 ;
  assign n5957 = ~x134 & ~n5956 ;
  assign n5958 = n191 & ~n4440 ;
  assign n5959 = n244 & ~n4448 ;
  assign n5960 = ~n5958 & ~n5959 ;
  assign n5961 = n298 & ~n4412 ;
  assign n5962 = n351 & ~n4404 ;
  assign n5963 = ~n5961 & ~n5962 ;
  assign n5964 = n5960 & n5963 ;
  assign n5965 = x134 & ~n5964 ;
  assign n5966 = ~n5957 & ~n5965 ;
  assign n5985 = ~n5966 & x180 ;
  assign n5967 = n298 & ~n4502 ;
  assign n5968 = n351 & ~n4494 ;
  assign n5969 = ~n5967 & ~n5968 ;
  assign n5970 = n191 & ~n4530 ;
  assign n5971 = n244 & ~n4538 ;
  assign n5972 = ~n5970 & ~n5971 ;
  assign n5973 = n5969 & n5972 ;
  assign n5974 = x134 & ~n5973 ;
  assign n5975 = n298 & ~n4513 ;
  assign n5976 = n351 & ~n4521 ;
  assign n5977 = ~n5975 & ~n5976 ;
  assign n5978 = n191 & ~n4485 ;
  assign n5979 = n244 & ~n4477 ;
  assign n5980 = ~n5978 & ~n5979 ;
  assign n5981 = n5977 & n5980 ;
  assign n5982 = ~x134 & ~n5981 ;
  assign n5983 = ~n5974 & ~n5982 ;
  assign n5986 = n5983 & ~x180 ;
  assign n5987 = ~n5985 & ~n5986 ;
  assign n5988 = n191 & ~n4579 ;
  assign n5989 = n244 & ~n4571 ;
  assign n5990 = ~n5988 & ~n5989 ;
  assign n5991 = n298 & ~n4607 ;
  assign n5992 = n351 & ~n4615 ;
  assign n5993 = ~n5991 & ~n5992 ;
  assign n5994 = n5990 & n5993 ;
  assign n5995 = ~x134 & ~n5994 ;
  assign n5996 = n191 & ~n4590 ;
  assign n5997 = n244 & ~n4598 ;
  assign n5998 = ~n5996 & ~n5997 ;
  assign n5999 = n298 & ~n4562 ;
  assign n6000 = n351 & ~n4554 ;
  assign n6001 = ~n5999 & ~n6000 ;
  assign n6002 = n5998 & n6001 ;
  assign n6003 = x134 & ~n6002 ;
  assign n6004 = ~n5995 & ~n6003 ;
  assign n6023 = ~n6004 & x181 ;
  assign n6005 = n298 & ~n4652 ;
  assign n6006 = n351 & ~n4644 ;
  assign n6007 = ~n6005 & ~n6006 ;
  assign n6008 = n191 & ~n4680 ;
  assign n6009 = n244 & ~n4688 ;
  assign n6010 = ~n6008 & ~n6009 ;
  assign n6011 = n6007 & n6010 ;
  assign n6012 = x134 & ~n6011 ;
  assign n6013 = n298 & ~n4663 ;
  assign n6014 = n351 & ~n4671 ;
  assign n6015 = ~n6013 & ~n6014 ;
  assign n6016 = n191 & ~n4635 ;
  assign n6017 = n244 & ~n4627 ;
  assign n6018 = ~n6016 & ~n6017 ;
  assign n6019 = n6015 & n6018 ;
  assign n6020 = ~x134 & ~n6019 ;
  assign n6021 = ~n6012 & ~n6020 ;
  assign n6024 = n6021 & ~x181 ;
  assign n6025 = ~n6023 & ~n6024 ;
  assign n6026 = n191 & ~n4729 ;
  assign n6027 = n244 & ~n4721 ;
  assign n6028 = ~n6026 & ~n6027 ;
  assign n6029 = n298 & ~n4757 ;
  assign n6030 = n351 & ~n4765 ;
  assign n6031 = ~n6029 & ~n6030 ;
  assign n6032 = n6028 & n6031 ;
  assign n6033 = ~x134 & ~n6032 ;
  assign n6034 = n191 & ~n4740 ;
  assign n6035 = n244 & ~n4748 ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = n298 & ~n4712 ;
  assign n6038 = n351 & ~n4704 ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6040 = n6036 & n6039 ;
  assign n6041 = x134 & ~n6040 ;
  assign n6042 = ~n6033 & ~n6041 ;
  assign n6061 = ~n6042 & x182 ;
  assign n6043 = n298 & ~n4802 ;
  assign n6044 = n351 & ~n4794 ;
  assign n6045 = ~n6043 & ~n6044 ;
  assign n6046 = n191 & ~n4830 ;
  assign n6047 = n244 & ~n4838 ;
  assign n6048 = ~n6046 & ~n6047 ;
  assign n6049 = n6045 & n6048 ;
  assign n6050 = x134 & ~n6049 ;
  assign n6051 = n298 & ~n4813 ;
  assign n6052 = n351 & ~n4821 ;
  assign n6053 = ~n6051 & ~n6052 ;
  assign n6054 = n191 & ~n4785 ;
  assign n6055 = n244 & ~n4777 ;
  assign n6056 = ~n6054 & ~n6055 ;
  assign n6057 = n6053 & n6056 ;
  assign n6058 = ~x134 & ~n6057 ;
  assign n6059 = ~n6050 & ~n6058 ;
  assign n6062 = n6059 & ~x182 ;
  assign n6063 = ~n6061 & ~n6062 ;
  assign n6064 = n191 & ~n297 ;
  assign n6065 = n244 & ~n406 ;
  assign n6066 = ~n6064 & ~n6065 ;
  assign n6067 = n298 & ~n563 ;
  assign n6068 = n351 & ~n458 ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6070 = n6066 & n6069 ;
  assign n6071 = ~x134 & ~n6070 ;
  assign n6072 = ~n190 & n244 ;
  assign n6073 = ~n243 & n351 ;
  assign n6074 = ~n6072 & ~n6073 ;
  assign n6075 = n191 & ~n511 ;
  assign n6076 = n298 & ~n350 ;
  assign n6077 = ~n6075 & ~n6076 ;
  assign n6078 = n6074 & n6077 ;
  assign n6079 = x134 & ~n6078 ;
  assign n6080 = ~n6071 & ~n6079 ;
  assign n6099 = ~n6080 & x183 ;
  assign n6081 = n298 & ~n724 ;
  assign n6082 = n351 & ~n831 ;
  assign n6083 = ~n6081 & ~n6082 ;
  assign n6084 = n191 & ~n988 ;
  assign n6085 = n244 & ~n883 ;
  assign n6086 = ~n6084 & ~n6085 ;
  assign n6087 = n6083 & n6086 ;
  assign n6088 = x134 & ~n6087 ;
  assign n6089 = n351 & ~n619 ;
  assign n6090 = n244 & ~n671 ;
  assign n6091 = ~n6089 & ~n6090 ;
  assign n6092 = n298 & ~n936 ;
  assign n6093 = n191 & ~n776 ;
  assign n6094 = ~n6092 & ~n6093 ;
  assign n6095 = n6091 & n6094 ;
  assign n6096 = ~x134 & ~n6095 ;
  assign n6097 = ~n6088 & ~n6096 ;
  assign n6100 = n6097 & ~x183 ;
  assign n6101 = ~n6099 & ~n6100 ;
  assign n6102 = n191 & ~n1153 ;
  assign n6103 = n244 & ~n1312 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6105 = n298 & ~n1365 ;
  assign n6106 = n351 & ~n1417 ;
  assign n6107 = ~n6105 & ~n6106 ;
  assign n6108 = n6104 & n6107 ;
  assign n6109 = ~x134 & ~n6108 ;
  assign n6110 = n191 & ~n1260 ;
  assign n6111 = n244 & ~n1048 ;
  assign n6112 = ~n6110 & ~n6111 ;
  assign n6113 = n298 & ~n1205 ;
  assign n6114 = n351 & ~n1100 ;
  assign n6115 = ~n6113 & ~n6114 ;
  assign n6116 = n6112 & n6115 ;
  assign n6117 = x134 & ~n6116 ;
  assign n6118 = ~n6109 & ~n6117 ;
  assign n6137 = ~n6118 & x184 ;
  assign n6119 = n298 & ~n1578 ;
  assign n6120 = n351 & ~n1737 ;
  assign n6121 = ~n6119 & ~n6120 ;
  assign n6122 = n191 & ~n1790 ;
  assign n6123 = n244 & ~n1842 ;
  assign n6124 = ~n6122 & ~n6123 ;
  assign n6125 = n6121 & n6124 ;
  assign n6126 = x134 & ~n6125 ;
  assign n6127 = n298 & ~n1685 ;
  assign n6128 = n351 & ~n1473 ;
  assign n6129 = ~n6127 & ~n6128 ;
  assign n6130 = n191 & ~n1630 ;
  assign n6131 = n244 & ~n1525 ;
  assign n6132 = ~n6130 & ~n6131 ;
  assign n6133 = n6129 & n6132 ;
  assign n6134 = ~x134 & ~n6133 ;
  assign n6135 = ~n6126 & ~n6134 ;
  assign n6138 = n6135 & ~x184 ;
  assign n6139 = ~n6137 & ~n6138 ;
  assign n6140 = n191 & ~n1959 ;
  assign n6141 = n244 & ~n2070 ;
  assign n6142 = ~n6140 & ~n6141 ;
  assign n6143 = n298 & ~n2107 ;
  assign n6144 = n351 & ~n2143 ;
  assign n6145 = ~n6143 & ~n6144 ;
  assign n6146 = n6142 & n6145 ;
  assign n6147 = ~x134 & ~n6146 ;
  assign n6148 = n191 & ~n2034 ;
  assign n6149 = n244 & ~n1886 ;
  assign n6150 = ~n6148 & ~n6149 ;
  assign n6151 = n298 & ~n1995 ;
  assign n6152 = n351 & ~n1922 ;
  assign n6153 = ~n6151 & ~n6152 ;
  assign n6154 = n6150 & n6153 ;
  assign n6155 = x134 & ~n6154 ;
  assign n6156 = ~n6147 & ~n6155 ;
  assign n6175 = ~n6156 & x185 ;
  assign n6157 = n298 & ~n2256 ;
  assign n6158 = n351 & ~n2367 ;
  assign n6159 = ~n6157 & ~n6158 ;
  assign n6160 = n191 & ~n2404 ;
  assign n6161 = n244 & ~n2440 ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6163 = n6159 & n6162 ;
  assign n6164 = x134 & ~n6163 ;
  assign n6165 = n298 & ~n2331 ;
  assign n6166 = n351 & ~n2183 ;
  assign n6167 = ~n6165 & ~n6166 ;
  assign n6168 = n191 & ~n2292 ;
  assign n6169 = n244 & ~n2219 ;
  assign n6170 = ~n6168 & ~n6169 ;
  assign n6171 = n6167 & n6170 ;
  assign n6172 = ~x134 & ~n6171 ;
  assign n6173 = ~n6164 & ~n6172 ;
  assign n6176 = n6173 & ~x185 ;
  assign n6177 = ~n6175 & ~n6176 ;
  assign n6178 = n298 & ~n2668 ;
  assign n6179 = n351 & ~n2741 ;
  assign n6180 = ~n6178 & ~n6179 ;
  assign n6181 = n191 & ~n2557 ;
  assign n6182 = n244 & ~n2705 ;
  assign n6183 = ~n6181 & ~n6182 ;
  assign n6184 = n6180 & n6183 ;
  assign n6185 = ~x134 & ~n6184 ;
  assign n6186 = n191 & ~n2632 ;
  assign n6187 = n298 & ~n2484 ;
  assign n6188 = ~n6186 & ~n6187 ;
  assign n6189 = n244 & ~n2593 ;
  assign n6190 = n351 & ~n2520 ;
  assign n6191 = ~n6189 & ~n6190 ;
  assign n6192 = n6188 & n6191 ;
  assign n6193 = x134 & ~n6192 ;
  assign n6194 = ~n6185 & ~n6193 ;
  assign n6213 = ~n6194 & x186 ;
  assign n6195 = n191 & ~n2965 ;
  assign n6196 = n244 & ~n3038 ;
  assign n6197 = ~n6195 & ~n6196 ;
  assign n6198 = n298 & ~n2854 ;
  assign n6199 = n351 & ~n3002 ;
  assign n6200 = ~n6198 & ~n6199 ;
  assign n6201 = n6197 & n6200 ;
  assign n6202 = x134 & ~n6201 ;
  assign n6203 = n298 & ~n2929 ;
  assign n6204 = n191 & ~n2781 ;
  assign n6205 = ~n6203 & ~n6204 ;
  assign n6206 = n351 & ~n2890 ;
  assign n6207 = n244 & ~n2817 ;
  assign n6208 = ~n6206 & ~n6207 ;
  assign n6209 = n6205 & n6208 ;
  assign n6210 = ~x134 & ~n6209 ;
  assign n6211 = ~n6202 & ~n6210 ;
  assign n6214 = n6211 & ~x186 ;
  assign n6215 = ~n6213 & ~n6214 ;
  assign n6216 = n298 & ~n3090 ;
  assign n6217 = n191 & ~n3071 ;
  assign n6218 = ~n6216 & ~n6217 ;
  assign n6219 = n351 & ~n3107 ;
  assign n6220 = n244 & ~n3115 ;
  assign n6221 = ~n6219 & ~n6220 ;
  assign n6222 = n6218 & n6221 ;
  assign n6223 = ~x134 & ~n6222 ;
  assign n6224 = n244 & ~n3054 ;
  assign n6225 = n351 & ~n3062 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = n298 & ~n3079 ;
  assign n6228 = n191 & ~n3098 ;
  assign n6229 = ~n6227 & ~n6228 ;
  assign n6230 = n6226 & n6229 ;
  assign n6231 = x134 & ~n6230 ;
  assign n6232 = ~n6223 & ~n6231 ;
  assign n6251 = ~n6232 & x187 ;
  assign n6233 = n191 & ~n3163 ;
  assign n6234 = n298 & ~n3144 ;
  assign n6235 = ~n6233 & ~n6234 ;
  assign n6236 = n244 & ~n3180 ;
  assign n6237 = n351 & ~n3188 ;
  assign n6238 = ~n6236 & ~n6237 ;
  assign n6239 = n6235 & n6238 ;
  assign n6240 = x134 & ~n6239 ;
  assign n6241 = n351 & ~n3127 ;
  assign n6242 = n244 & ~n3135 ;
  assign n6243 = ~n6241 & ~n6242 ;
  assign n6244 = n191 & ~n3152 ;
  assign n6245 = n298 & ~n3171 ;
  assign n6246 = ~n6244 & ~n6245 ;
  assign n6247 = n6243 & n6246 ;
  assign n6248 = ~x134 & ~n6247 ;
  assign n6249 = ~n6240 & ~n6248 ;
  assign n6252 = n6249 & ~x187 ;
  assign n6253 = ~n6251 & ~n6252 ;
  assign n6254 = n298 & ~n3240 ;
  assign n6255 = n191 & ~n3221 ;
  assign n6256 = ~n6254 & ~n6255 ;
  assign n6257 = n351 & ~n3257 ;
  assign n6258 = n244 & ~n3265 ;
  assign n6259 = ~n6257 & ~n6258 ;
  assign n6260 = n6256 & n6259 ;
  assign n6261 = ~x134 & ~n6260 ;
  assign n6262 = n244 & ~n3204 ;
  assign n6263 = n351 & ~n3212 ;
  assign n6264 = ~n6262 & ~n6263 ;
  assign n6265 = n298 & ~n3229 ;
  assign n6266 = n191 & ~n3248 ;
  assign n6267 = ~n6265 & ~n6266 ;
  assign n6268 = n6264 & n6267 ;
  assign n6269 = x134 & ~n6268 ;
  assign n6270 = ~n6261 & ~n6269 ;
  assign n6289 = ~n6270 & x188 ;
  assign n6271 = n191 & ~n3313 ;
  assign n6272 = n298 & ~n3294 ;
  assign n6273 = ~n6271 & ~n6272 ;
  assign n6274 = n244 & ~n3330 ;
  assign n6275 = n351 & ~n3338 ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6277 = n6273 & n6276 ;
  assign n6278 = x134 & ~n6277 ;
  assign n6279 = n351 & ~n3277 ;
  assign n6280 = n244 & ~n3285 ;
  assign n6281 = ~n6279 & ~n6280 ;
  assign n6282 = n191 & ~n3302 ;
  assign n6283 = n298 & ~n3321 ;
  assign n6284 = ~n6282 & ~n6283 ;
  assign n6285 = n6281 & n6284 ;
  assign n6286 = ~x134 & ~n6285 ;
  assign n6287 = ~n6278 & ~n6286 ;
  assign n6290 = n6287 & ~x188 ;
  assign n6291 = ~n6289 & ~n6290 ;
  assign n6292 = n298 & ~n3390 ;
  assign n6293 = n191 & ~n3371 ;
  assign n6294 = ~n6292 & ~n6293 ;
  assign n6295 = n351 & ~n3407 ;
  assign n6296 = n244 & ~n3415 ;
  assign n6297 = ~n6295 & ~n6296 ;
  assign n6298 = n6294 & n6297 ;
  assign n6299 = ~x134 & ~n6298 ;
  assign n6300 = n244 & ~n3354 ;
  assign n6301 = n351 & ~n3362 ;
  assign n6302 = ~n6300 & ~n6301 ;
  assign n6303 = n298 & ~n3379 ;
  assign n6304 = n191 & ~n3398 ;
  assign n6305 = ~n6303 & ~n6304 ;
  assign n6306 = n6302 & n6305 ;
  assign n6307 = x134 & ~n6306 ;
  assign n6308 = ~n6299 & ~n6307 ;
  assign n6327 = ~n6308 & x189 ;
  assign n6309 = n191 & ~n3463 ;
  assign n6310 = n298 & ~n3444 ;
  assign n6311 = ~n6309 & ~n6310 ;
  assign n6312 = n244 & ~n3480 ;
  assign n6313 = n351 & ~n3488 ;
  assign n6314 = ~n6312 & ~n6313 ;
  assign n6315 = n6311 & n6314 ;
  assign n6316 = x134 & ~n6315 ;
  assign n6317 = n351 & ~n3427 ;
  assign n6318 = n244 & ~n3435 ;
  assign n6319 = ~n6317 & ~n6318 ;
  assign n6320 = n191 & ~n3452 ;
  assign n6321 = n298 & ~n3471 ;
  assign n6322 = ~n6320 & ~n6321 ;
  assign n6323 = n6319 & n6322 ;
  assign n6324 = ~x134 & ~n6323 ;
  assign n6325 = ~n6316 & ~n6324 ;
  assign n6328 = n6325 & ~x189 ;
  assign n6329 = ~n6327 & ~n6328 ;
  assign n6330 = n298 & ~n3540 ;
  assign n6331 = n244 & ~n3565 ;
  assign n6332 = ~n6330 & ~n6331 ;
  assign n6333 = n191 & ~n3521 ;
  assign n6334 = n351 & ~n3557 ;
  assign n6335 = ~n6333 & ~n6334 ;
  assign n6336 = n6332 & n6335 ;
  assign n6337 = ~x134 & ~n6336 ;
  assign n6338 = n191 & ~n3548 ;
  assign n6339 = n244 & ~n3504 ;
  assign n6340 = ~n6338 & ~n6339 ;
  assign n6341 = n298 & ~n3529 ;
  assign n6342 = n351 & ~n3512 ;
  assign n6343 = ~n6341 & ~n6342 ;
  assign n6344 = n6340 & n6343 ;
  assign n6345 = x134 & ~n6344 ;
  assign n6346 = ~n6337 & ~n6345 ;
  assign n6365 = ~n6346 & x190 ;
  assign n6347 = n191 & ~n3613 ;
  assign n6348 = n351 & ~n3638 ;
  assign n6349 = ~n6347 & ~n6348 ;
  assign n6350 = n298 & ~n3594 ;
  assign n6351 = n244 & ~n3630 ;
  assign n6352 = ~n6350 & ~n6351 ;
  assign n6353 = n6349 & n6352 ;
  assign n6354 = x134 & ~n6353 ;
  assign n6355 = n298 & ~n3621 ;
  assign n6356 = n351 & ~n3577 ;
  assign n6357 = ~n6355 & ~n6356 ;
  assign n6358 = n191 & ~n3602 ;
  assign n6359 = n244 & ~n3585 ;
  assign n6360 = ~n6358 & ~n6359 ;
  assign n6361 = n6357 & n6360 ;
  assign n6362 = ~x134 & ~n6361 ;
  assign n6363 = ~n6354 & ~n6362 ;
  assign n6366 = n6363 & ~x190 ;
  assign n6367 = ~n6365 & ~n6366 ;
  assign n6368 = n298 & ~n3690 ;
  assign n6369 = n244 & ~n3715 ;
  assign n6370 = ~n6368 & ~n6369 ;
  assign n6371 = n191 & ~n3671 ;
  assign n6372 = n351 & ~n3707 ;
  assign n6373 = ~n6371 & ~n6372 ;
  assign n6374 = n6370 & n6373 ;
  assign n6375 = ~x134 & ~n6374 ;
  assign n6376 = n191 & ~n3698 ;
  assign n6377 = n244 & ~n3654 ;
  assign n6378 = ~n6376 & ~n6377 ;
  assign n6379 = n298 & ~n3679 ;
  assign n6380 = n351 & ~n3662 ;
  assign n6381 = ~n6379 & ~n6380 ;
  assign n6382 = n6378 & n6381 ;
  assign n6383 = x134 & ~n6382 ;
  assign n6384 = ~n6375 & ~n6383 ;
  assign n6403 = ~n6384 & x191 ;
  assign n6385 = n191 & ~n3763 ;
  assign n6386 = n351 & ~n3788 ;
  assign n6387 = ~n6385 & ~n6386 ;
  assign n6388 = n298 & ~n3744 ;
  assign n6389 = n244 & ~n3780 ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = n6387 & n6390 ;
  assign n6392 = x134 & ~n6391 ;
  assign n6393 = n298 & ~n3771 ;
  assign n6394 = n351 & ~n3727 ;
  assign n6395 = ~n6393 & ~n6394 ;
  assign n6396 = n191 & ~n3752 ;
  assign n6397 = n244 & ~n3735 ;
  assign n6398 = ~n6396 & ~n6397 ;
  assign n6399 = n6395 & n6398 ;
  assign n6400 = ~x134 & ~n6399 ;
  assign n6401 = ~n6392 & ~n6400 ;
  assign n6404 = n6401 & ~x191 ;
  assign n6405 = ~n6403 & ~n6404 ;
  assign n6406 = n298 & ~n3840 ;
  assign n6407 = n244 & ~n3865 ;
  assign n6408 = ~n6406 & ~n6407 ;
  assign n6409 = n191 & ~n3821 ;
  assign n6410 = n351 & ~n3857 ;
  assign n6411 = ~n6409 & ~n6410 ;
  assign n6412 = n6408 & n6411 ;
  assign n6413 = ~x134 & ~n6412 ;
  assign n6414 = n191 & ~n3848 ;
  assign n6415 = n244 & ~n3804 ;
  assign n6416 = ~n6414 & ~n6415 ;
  assign n6417 = n298 & ~n3829 ;
  assign n6418 = n351 & ~n3812 ;
  assign n6419 = ~n6417 & ~n6418 ;
  assign n6420 = n6416 & n6419 ;
  assign n6421 = x134 & ~n6420 ;
  assign n6422 = ~n6413 & ~n6421 ;
  assign n6441 = ~n6422 & x192 ;
  assign n6423 = n191 & ~n3913 ;
  assign n6424 = n351 & ~n3938 ;
  assign n6425 = ~n6423 & ~n6424 ;
  assign n6426 = n298 & ~n3894 ;
  assign n6427 = n244 & ~n3930 ;
  assign n6428 = ~n6426 & ~n6427 ;
  assign n6429 = n6425 & n6428 ;
  assign n6430 = x134 & ~n6429 ;
  assign n6431 = n298 & ~n3921 ;
  assign n6432 = n351 & ~n3877 ;
  assign n6433 = ~n6431 & ~n6432 ;
  assign n6434 = n191 & ~n3902 ;
  assign n6435 = n244 & ~n3885 ;
  assign n6436 = ~n6434 & ~n6435 ;
  assign n6437 = n6433 & n6436 ;
  assign n6438 = ~x134 & ~n6437 ;
  assign n6439 = ~n6430 & ~n6438 ;
  assign n6442 = n6439 & ~x192 ;
  assign n6443 = ~n6441 & ~n6442 ;
  assign n6444 = n298 & ~n3990 ;
  assign n6445 = n191 & ~n3971 ;
  assign n6446 = ~n6444 & ~n6445 ;
  assign n6447 = n351 & ~n4007 ;
  assign n6448 = n244 & ~n4015 ;
  assign n6449 = ~n6447 & ~n6448 ;
  assign n6450 = n6446 & n6449 ;
  assign n6451 = ~x134 & ~n6450 ;
  assign n6452 = n191 & ~n3998 ;
  assign n6453 = n244 & ~n3954 ;
  assign n6454 = ~n6452 & ~n6453 ;
  assign n6455 = n298 & ~n3979 ;
  assign n6456 = n351 & ~n3962 ;
  assign n6457 = ~n6455 & ~n6456 ;
  assign n6458 = n6454 & n6457 ;
  assign n6459 = x134 & ~n6458 ;
  assign n6460 = ~n6451 & ~n6459 ;
  assign n6479 = ~n6460 & x193 ;
  assign n6461 = n191 & ~n4063 ;
  assign n6462 = n298 & ~n4044 ;
  assign n6463 = ~n6461 & ~n6462 ;
  assign n6464 = n244 & ~n4080 ;
  assign n6465 = n351 & ~n4088 ;
  assign n6466 = ~n6464 & ~n6465 ;
  assign n6467 = n6463 & n6466 ;
  assign n6468 = x134 & ~n6467 ;
  assign n6469 = n298 & ~n4071 ;
  assign n6470 = n351 & ~n4027 ;
  assign n6471 = ~n6469 & ~n6470 ;
  assign n6472 = n191 & ~n4052 ;
  assign n6473 = n244 & ~n4035 ;
  assign n6474 = ~n6472 & ~n6473 ;
  assign n6475 = n6471 & n6474 ;
  assign n6476 = ~x134 & ~n6475 ;
  assign n6477 = ~n6468 & ~n6476 ;
  assign n6480 = n6477 & ~x193 ;
  assign n6481 = ~n6479 & ~n6480 ;
  assign n6482 = n298 & ~n4140 ;
  assign n6483 = n191 & ~n4121 ;
  assign n6484 = ~n6482 & ~n6483 ;
  assign n6485 = n351 & ~n4157 ;
  assign n6486 = n244 & ~n4165 ;
  assign n6487 = ~n6485 & ~n6486 ;
  assign n6488 = n6484 & n6487 ;
  assign n6489 = ~x134 & ~n6488 ;
  assign n6490 = n191 & ~n4148 ;
  assign n6491 = n244 & ~n4104 ;
  assign n6492 = ~n6490 & ~n6491 ;
  assign n6493 = n298 & ~n4129 ;
  assign n6494 = n351 & ~n4112 ;
  assign n6495 = ~n6493 & ~n6494 ;
  assign n6496 = n6492 & n6495 ;
  assign n6497 = x134 & ~n6496 ;
  assign n6498 = ~n6489 & ~n6497 ;
  assign n6517 = ~n6498 & x194 ;
  assign n6499 = n191 & ~n4213 ;
  assign n6500 = n298 & ~n4194 ;
  assign n6501 = ~n6499 & ~n6500 ;
  assign n6502 = n244 & ~n4230 ;
  assign n6503 = n351 & ~n4238 ;
  assign n6504 = ~n6502 & ~n6503 ;
  assign n6505 = n6501 & n6504 ;
  assign n6506 = x134 & ~n6505 ;
  assign n6507 = n298 & ~n4221 ;
  assign n6508 = n351 & ~n4177 ;
  assign n6509 = ~n6507 & ~n6508 ;
  assign n6510 = n191 & ~n4202 ;
  assign n6511 = n244 & ~n4185 ;
  assign n6512 = ~n6510 & ~n6511 ;
  assign n6513 = n6509 & n6512 ;
  assign n6514 = ~x134 & ~n6513 ;
  assign n6515 = ~n6506 & ~n6514 ;
  assign n6518 = n6515 & ~x194 ;
  assign n6519 = ~n6517 & ~n6518 ;
  assign n6520 = n298 & ~n4290 ;
  assign n6521 = n191 & ~n4271 ;
  assign n6522 = ~n6520 & ~n6521 ;
  assign n6523 = n351 & ~n4307 ;
  assign n6524 = n244 & ~n4315 ;
  assign n6525 = ~n6523 & ~n6524 ;
  assign n6526 = n6522 & n6525 ;
  assign n6527 = ~x134 & ~n6526 ;
  assign n6528 = n191 & ~n4298 ;
  assign n6529 = n244 & ~n4254 ;
  assign n6530 = ~n6528 & ~n6529 ;
  assign n6531 = n298 & ~n4279 ;
  assign n6532 = n351 & ~n4262 ;
  assign n6533 = ~n6531 & ~n6532 ;
  assign n6534 = n6530 & n6533 ;
  assign n6535 = x134 & ~n6534 ;
  assign n6536 = ~n6527 & ~n6535 ;
  assign n6555 = ~n6536 & x195 ;
  assign n6537 = n191 & ~n4363 ;
  assign n6538 = n298 & ~n4344 ;
  assign n6539 = ~n6537 & ~n6538 ;
  assign n6540 = n244 & ~n4380 ;
  assign n6541 = n351 & ~n4388 ;
  assign n6542 = ~n6540 & ~n6541 ;
  assign n6543 = n6539 & n6542 ;
  assign n6544 = x134 & ~n6543 ;
  assign n6545 = n298 & ~n4371 ;
  assign n6546 = n351 & ~n4327 ;
  assign n6547 = ~n6545 & ~n6546 ;
  assign n6548 = n191 & ~n4352 ;
  assign n6549 = n244 & ~n4335 ;
  assign n6550 = ~n6548 & ~n6549 ;
  assign n6551 = n6547 & n6550 ;
  assign n6552 = ~x134 & ~n6551 ;
  assign n6553 = ~n6544 & ~n6552 ;
  assign n6556 = n6553 & ~x195 ;
  assign n6557 = ~n6555 & ~n6556 ;
  assign n6558 = n298 & ~n4440 ;
  assign n6559 = n191 & ~n4421 ;
  assign n6560 = ~n6558 & ~n6559 ;
  assign n6561 = n351 & ~n4457 ;
  assign n6562 = n244 & ~n4465 ;
  assign n6563 = ~n6561 & ~n6562 ;
  assign n6564 = n6560 & n6563 ;
  assign n6565 = ~x134 & ~n6564 ;
  assign n6566 = n191 & ~n4448 ;
  assign n6567 = n244 & ~n4404 ;
  assign n6568 = ~n6566 & ~n6567 ;
  assign n6569 = n298 & ~n4429 ;
  assign n6570 = n351 & ~n4412 ;
  assign n6571 = ~n6569 & ~n6570 ;
  assign n6572 = n6568 & n6571 ;
  assign n6573 = x134 & ~n6572 ;
  assign n6574 = ~n6565 & ~n6573 ;
  assign n6593 = ~n6574 & x196 ;
  assign n6575 = n191 & ~n4513 ;
  assign n6576 = n298 & ~n4494 ;
  assign n6577 = ~n6575 & ~n6576 ;
  assign n6578 = n244 & ~n4530 ;
  assign n6579 = n351 & ~n4538 ;
  assign n6580 = ~n6578 & ~n6579 ;
  assign n6581 = n6577 & n6580 ;
  assign n6582 = x134 & ~n6581 ;
  assign n6583 = n298 & ~n4521 ;
  assign n6584 = n351 & ~n4477 ;
  assign n6585 = ~n6583 & ~n6584 ;
  assign n6586 = n191 & ~n4502 ;
  assign n6587 = n244 & ~n4485 ;
  assign n6588 = ~n6586 & ~n6587 ;
  assign n6589 = n6585 & n6588 ;
  assign n6590 = ~x134 & ~n6589 ;
  assign n6591 = ~n6582 & ~n6590 ;
  assign n6594 = n6591 & ~x196 ;
  assign n6595 = ~n6593 & ~n6594 ;
  assign n6596 = n298 & ~n4590 ;
  assign n6597 = n191 & ~n4571 ;
  assign n6598 = ~n6596 & ~n6597 ;
  assign n6599 = n351 & ~n4607 ;
  assign n6600 = n244 & ~n4615 ;
  assign n6601 = ~n6599 & ~n6600 ;
  assign n6602 = n6598 & n6601 ;
  assign n6603 = ~x134 & ~n6602 ;
  assign n6604 = n191 & ~n4598 ;
  assign n6605 = n244 & ~n4554 ;
  assign n6606 = ~n6604 & ~n6605 ;
  assign n6607 = n298 & ~n4579 ;
  assign n6608 = n351 & ~n4562 ;
  assign n6609 = ~n6607 & ~n6608 ;
  assign n6610 = n6606 & n6609 ;
  assign n6611 = x134 & ~n6610 ;
  assign n6612 = ~n6603 & ~n6611 ;
  assign n6631 = ~n6612 & x197 ;
  assign n6613 = n191 & ~n4663 ;
  assign n6614 = n298 & ~n4644 ;
  assign n6615 = ~n6613 & ~n6614 ;
  assign n6616 = n244 & ~n4680 ;
  assign n6617 = n351 & ~n4688 ;
  assign n6618 = ~n6616 & ~n6617 ;
  assign n6619 = n6615 & n6618 ;
  assign n6620 = x134 & ~n6619 ;
  assign n6621 = n298 & ~n4671 ;
  assign n6622 = n351 & ~n4627 ;
  assign n6623 = ~n6621 & ~n6622 ;
  assign n6624 = n191 & ~n4652 ;
  assign n6625 = n244 & ~n4635 ;
  assign n6626 = ~n6624 & ~n6625 ;
  assign n6627 = n6623 & n6626 ;
  assign n6628 = ~x134 & ~n6627 ;
  assign n6629 = ~n6620 & ~n6628 ;
  assign n6632 = n6629 & ~x197 ;
  assign n6633 = ~n6631 & ~n6632 ;
  assign n6634 = n298 & ~n4740 ;
  assign n6635 = n191 & ~n4721 ;
  assign n6636 = ~n6634 & ~n6635 ;
  assign n6637 = n351 & ~n4757 ;
  assign n6638 = n244 & ~n4765 ;
  assign n6639 = ~n6637 & ~n6638 ;
  assign n6640 = n6636 & n6639 ;
  assign n6641 = ~x134 & ~n6640 ;
  assign n6642 = n191 & ~n4748 ;
  assign n6643 = n244 & ~n4704 ;
  assign n6644 = ~n6642 & ~n6643 ;
  assign n6645 = n298 & ~n4729 ;
  assign n6646 = n351 & ~n4712 ;
  assign n6647 = ~n6645 & ~n6646 ;
  assign n6648 = n6644 & n6647 ;
  assign n6649 = x134 & ~n6648 ;
  assign n6650 = ~n6641 & ~n6649 ;
  assign n6669 = ~n6650 & x198 ;
  assign n6651 = n191 & ~n4813 ;
  assign n6652 = n298 & ~n4794 ;
  assign n6653 = ~n6651 & ~n6652 ;
  assign n6654 = n244 & ~n4830 ;
  assign n6655 = n351 & ~n4838 ;
  assign n6656 = ~n6654 & ~n6655 ;
  assign n6657 = n6653 & n6656 ;
  assign n6658 = x134 & ~n6657 ;
  assign n6659 = n298 & ~n4821 ;
  assign n6660 = n351 & ~n4777 ;
  assign n6661 = ~n6659 & ~n6660 ;
  assign n6662 = n191 & ~n4802 ;
  assign n6663 = n244 & ~n4785 ;
  assign n6664 = ~n6662 & ~n6663 ;
  assign n6665 = n6661 & n6664 ;
  assign n6666 = ~x134 & ~n6665 ;
  assign n6667 = ~n6658 & ~n6666 ;
  assign n6670 = n6667 & ~x198 ;
  assign n6671 = ~n6669 & ~n6670 ;
  assign n6672 = ~x134 & ~n566 ;
  assign n6673 = x134 & ~n354 ;
  assign n6674 = ~n6672 & ~n6673 ;
  assign n6679 = ~n6674 & x199 ;
  assign n6675 = x134 & ~n991 ;
  assign n6676 = ~x134 & ~n779 ;
  assign n6677 = ~n6675 & ~n6676 ;
  assign n6680 = n6677 & ~x199 ;
  assign n6681 = ~n6679 & ~n6680 ;
  assign n6682 = ~x134 & ~n1420 ;
  assign n6683 = x134 & ~n1208 ;
  assign n6684 = ~n6682 & ~n6683 ;
  assign n6689 = ~n6684 & x200 ;
  assign n6685 = x134 & ~n1845 ;
  assign n6686 = ~x134 & ~n1633 ;
  assign n6687 = ~n6685 & ~n6686 ;
  assign n6690 = n6687 & ~x200 ;
  assign n6691 = ~n6689 & ~n6690 ;
  assign n6692 = ~x134 & ~n2146 ;
  assign n6693 = x134 & ~n1998 ;
  assign n6694 = ~n6692 & ~n6693 ;
  assign n6699 = ~n6694 & x201 ;
  assign n6695 = x134 & ~n2443 ;
  assign n6696 = ~x134 & ~n2295 ;
  assign n6697 = ~n6695 & ~n6696 ;
  assign n6700 = n6697 & ~x201 ;
  assign n6701 = ~n6699 & ~n6700 ;
  assign n6702 = ~x134 & ~n2744 ;
  assign n6703 = x134 & ~n2596 ;
  assign n6704 = ~n6702 & ~n6703 ;
  assign n6709 = ~n6704 & x202 ;
  assign n6705 = x134 & ~n3041 ;
  assign n6706 = ~x134 & ~n2893 ;
  assign n6707 = ~n6705 & ~n6706 ;
  assign n6710 = n6707 & ~x202 ;
  assign n6711 = ~n6709 & ~n6710 ;
  assign n6712 = ~x134 & ~n3118 ;
  assign n6713 = x134 & ~n3082 ;
  assign n6714 = ~n6712 & ~n6713 ;
  assign n6719 = ~n6714 & x203 ;
  assign n6715 = x134 & ~n3191 ;
  assign n6716 = ~x134 & ~n3155 ;
  assign n6717 = ~n6715 & ~n6716 ;
  assign n6720 = n6717 & ~x203 ;
  assign n6721 = ~n6719 & ~n6720 ;
  assign n6722 = ~x134 & ~n3268 ;
  assign n6723 = x134 & ~n3232 ;
  assign n6724 = ~n6722 & ~n6723 ;
  assign n6729 = ~n6724 & x204 ;
  assign n6725 = x134 & ~n3341 ;
  assign n6726 = ~x134 & ~n3305 ;
  assign n6727 = ~n6725 & ~n6726 ;
  assign n6730 = n6727 & ~x204 ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6732 = ~x134 & ~n3418 ;
  assign n6733 = x134 & ~n3382 ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6739 = ~n6734 & x205 ;
  assign n6735 = x134 & ~n3491 ;
  assign n6736 = ~x134 & ~n3455 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6740 = n6737 & ~x205 ;
  assign n6741 = ~n6739 & ~n6740 ;
  assign n6742 = ~x134 & ~n3568 ;
  assign n6743 = x134 & ~n3532 ;
  assign n6744 = ~n6742 & ~n6743 ;
  assign n6749 = ~n6744 & x206 ;
  assign n6745 = x134 & ~n3641 ;
  assign n6746 = ~x134 & ~n3605 ;
  assign n6747 = ~n6745 & ~n6746 ;
  assign n6750 = n6747 & ~x206 ;
  assign n6751 = ~n6749 & ~n6750 ;
  assign n6752 = ~x134 & ~n3718 ;
  assign n6753 = x134 & ~n3682 ;
  assign n6754 = ~n6752 & ~n6753 ;
  assign n6759 = ~n6754 & x207 ;
  assign n6755 = x134 & ~n3791 ;
  assign n6756 = ~x134 & ~n3755 ;
  assign n6757 = ~n6755 & ~n6756 ;
  assign n6760 = n6757 & ~x207 ;
  assign n6761 = ~n6759 & ~n6760 ;
  assign n6762 = ~x134 & ~n3868 ;
  assign n6763 = x134 & ~n3832 ;
  assign n6764 = ~n6762 & ~n6763 ;
  assign n6769 = ~n6764 & x208 ;
  assign n6765 = x134 & ~n3941 ;
  assign n6766 = ~x134 & ~n3905 ;
  assign n6767 = ~n6765 & ~n6766 ;
  assign n6770 = n6767 & ~x208 ;
  assign n6771 = ~n6769 & ~n6770 ;
  assign n6772 = ~x134 & ~n4018 ;
  assign n6773 = x134 & ~n3982 ;
  assign n6774 = ~n6772 & ~n6773 ;
  assign n6779 = ~n6774 & x209 ;
  assign n6775 = x134 & ~n4091 ;
  assign n6776 = ~x134 & ~n4055 ;
  assign n6777 = ~n6775 & ~n6776 ;
  assign n6780 = n6777 & ~x209 ;
  assign n6781 = ~n6779 & ~n6780 ;
  assign n6782 = ~x134 & ~n4168 ;
  assign n6783 = x134 & ~n4132 ;
  assign n6784 = ~n6782 & ~n6783 ;
  assign n6789 = ~n6784 & x210 ;
  assign n6785 = x134 & ~n4241 ;
  assign n6786 = ~x134 & ~n4205 ;
  assign n6787 = ~n6785 & ~n6786 ;
  assign n6790 = n6787 & ~x210 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = ~x134 & ~n4318 ;
  assign n6793 = x134 & ~n4282 ;
  assign n6794 = ~n6792 & ~n6793 ;
  assign n6799 = ~n6794 & x211 ;
  assign n6795 = x134 & ~n4391 ;
  assign n6796 = ~x134 & ~n4355 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6800 = n6797 & ~x211 ;
  assign n6801 = ~n6799 & ~n6800 ;
  assign n6802 = ~x134 & ~n4468 ;
  assign n6803 = x134 & ~n4432 ;
  assign n6804 = ~n6802 & ~n6803 ;
  assign n6809 = ~n6804 & x212 ;
  assign n6805 = x134 & ~n4541 ;
  assign n6806 = ~x134 & ~n4505 ;
  assign n6807 = ~n6805 & ~n6806 ;
  assign n6810 = n6807 & ~x212 ;
  assign n6811 = ~n6809 & ~n6810 ;
  assign n6812 = ~x134 & ~n4618 ;
  assign n6813 = x134 & ~n4582 ;
  assign n6814 = ~n6812 & ~n6813 ;
  assign n6819 = ~n6814 & x213 ;
  assign n6815 = x134 & ~n4691 ;
  assign n6816 = ~x134 & ~n4655 ;
  assign n6817 = ~n6815 & ~n6816 ;
  assign n6820 = n6817 & ~x213 ;
  assign n6821 = ~n6819 & ~n6820 ;
  assign n6822 = ~x134 & ~n4768 ;
  assign n6823 = x134 & ~n4732 ;
  assign n6824 = ~n6822 & ~n6823 ;
  assign n6829 = ~n6824 & x214 ;
  assign n6825 = x134 & ~n4841 ;
  assign n6826 = ~x134 & ~n4805 ;
  assign n6827 = ~n6825 & ~n6826 ;
  assign n6830 = n6827 & ~x214 ;
  assign n6831 = ~n6829 & ~n6830 ;
  assign n6832 = ~x134 & ~n4862 ;
  assign n6833 = x134 & ~n4854 ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6839 = ~n6834 & x215 ;
  assign n6835 = x134 & ~n4879 ;
  assign n6836 = ~x134 & ~n4871 ;
  assign n6837 = ~n6835 & ~n6836 ;
  assign n6840 = n6837 & ~x215 ;
  assign n6841 = ~n6839 & ~n6840 ;
  assign n6842 = ~x134 & ~n4900 ;
  assign n6843 = x134 & ~n4892 ;
  assign n6844 = ~n6842 & ~n6843 ;
  assign n6849 = ~n6844 & x216 ;
  assign n6845 = x134 & ~n4917 ;
  assign n6846 = ~x134 & ~n4909 ;
  assign n6847 = ~n6845 & ~n6846 ;
  assign n6850 = n6847 & ~x216 ;
  assign n6851 = ~n6849 & ~n6850 ;
  assign n6852 = ~x134 & ~n4938 ;
  assign n6853 = x134 & ~n4930 ;
  assign n6854 = ~n6852 & ~n6853 ;
  assign n6859 = ~n6854 & x217 ;
  assign n6855 = x134 & ~n4955 ;
  assign n6856 = ~x134 & ~n4947 ;
  assign n6857 = ~n6855 & ~n6856 ;
  assign n6860 = n6857 & ~x217 ;
  assign n6861 = ~n6859 & ~n6860 ;
  assign n6862 = ~x134 & ~n4976 ;
  assign n6863 = x134 & ~n4968 ;
  assign n6864 = ~n6862 & ~n6863 ;
  assign n6869 = ~n6864 & x218 ;
  assign n6865 = x134 & ~n4993 ;
  assign n6866 = ~x134 & ~n4985 ;
  assign n6867 = ~n6865 & ~n6866 ;
  assign n6870 = n6867 & ~x218 ;
  assign n6871 = ~n6869 & ~n6870 ;
  assign n6872 = ~x134 & ~n5014 ;
  assign n6873 = x134 & ~n5006 ;
  assign n6874 = ~n6872 & ~n6873 ;
  assign n6879 = ~n6874 & x219 ;
  assign n6875 = x134 & ~n5031 ;
  assign n6876 = ~x134 & ~n5023 ;
  assign n6877 = ~n6875 & ~n6876 ;
  assign n6880 = n6877 & ~x219 ;
  assign n6881 = ~n6879 & ~n6880 ;
  assign n6882 = ~x134 & ~n5052 ;
  assign n6883 = x134 & ~n5044 ;
  assign n6884 = ~n6882 & ~n6883 ;
  assign n6889 = ~n6884 & x220 ;
  assign n6885 = x134 & ~n5069 ;
  assign n6886 = ~x134 & ~n5061 ;
  assign n6887 = ~n6885 & ~n6886 ;
  assign n6890 = n6887 & ~x220 ;
  assign n6891 = ~n6889 & ~n6890 ;
  assign n6892 = ~x134 & ~n5090 ;
  assign n6893 = x134 & ~n5082 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6899 = ~n6894 & x221 ;
  assign n6895 = x134 & ~n5107 ;
  assign n6896 = ~x134 & ~n5099 ;
  assign n6897 = ~n6895 & ~n6896 ;
  assign n6900 = n6897 & ~x221 ;
  assign n6901 = ~n6899 & ~n6900 ;
  assign n6902 = ~x134 & ~n5128 ;
  assign n6903 = x134 & ~n5120 ;
  assign n6904 = ~n6902 & ~n6903 ;
  assign n6909 = ~n6904 & x222 ;
  assign n6905 = x134 & ~n5145 ;
  assign n6906 = ~x134 & ~n5137 ;
  assign n6907 = ~n6905 & ~n6906 ;
  assign n6910 = n6907 & ~x222 ;
  assign n6911 = ~n6909 & ~n6910 ;
  assign n6912 = ~x134 & ~n5166 ;
  assign n6913 = x134 & ~n5158 ;
  assign n6914 = ~n6912 & ~n6913 ;
  assign n6919 = ~n6914 & x223 ;
  assign n6915 = x134 & ~n5183 ;
  assign n6916 = ~x134 & ~n5175 ;
  assign n6917 = ~n6915 & ~n6916 ;
  assign n6920 = n6917 & ~x223 ;
  assign n6921 = ~n6919 & ~n6920 ;
  assign n6922 = ~x134 & ~n5204 ;
  assign n6923 = x134 & ~n5196 ;
  assign n6924 = ~n6922 & ~n6923 ;
  assign n6929 = ~n6924 & x224 ;
  assign n6925 = x134 & ~n5221 ;
  assign n6926 = ~x134 & ~n5213 ;
  assign n6927 = ~n6925 & ~n6926 ;
  assign n6930 = n6927 & ~x224 ;
  assign n6931 = ~n6929 & ~n6930 ;
  assign n6932 = ~x134 & ~n5242 ;
  assign n6933 = x134 & ~n5234 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6939 = ~n6934 & x225 ;
  assign n6935 = x134 & ~n5259 ;
  assign n6936 = ~x134 & ~n5251 ;
  assign n6937 = ~n6935 & ~n6936 ;
  assign n6940 = n6937 & ~x225 ;
  assign n6941 = ~n6939 & ~n6940 ;
  assign n6942 = ~x134 & ~n5280 ;
  assign n6943 = x134 & ~n5272 ;
  assign n6944 = ~n6942 & ~n6943 ;
  assign n6949 = ~n6944 & x226 ;
  assign n6945 = x134 & ~n5297 ;
  assign n6946 = ~x134 & ~n5289 ;
  assign n6947 = ~n6945 & ~n6946 ;
  assign n6950 = n6947 & ~x226 ;
  assign n6951 = ~n6949 & ~n6950 ;
  assign n6952 = ~x134 & ~n5318 ;
  assign n6953 = x134 & ~n5310 ;
  assign n6954 = ~n6952 & ~n6953 ;
  assign n6959 = ~n6954 & x227 ;
  assign n6955 = x134 & ~n5335 ;
  assign n6956 = ~x134 & ~n5327 ;
  assign n6957 = ~n6955 & ~n6956 ;
  assign n6960 = n6957 & ~x227 ;
  assign n6961 = ~n6959 & ~n6960 ;
  assign n6962 = ~x134 & ~n5356 ;
  assign n6963 = x134 & ~n5348 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6969 = ~n6964 & x228 ;
  assign n6965 = x134 & ~n5373 ;
  assign n6966 = ~x134 & ~n5365 ;
  assign n6967 = ~n6965 & ~n6966 ;
  assign n6970 = n6967 & ~x228 ;
  assign n6971 = ~n6969 & ~n6970 ;
  assign n6972 = ~x134 & ~n5394 ;
  assign n6973 = x134 & ~n5386 ;
  assign n6974 = ~n6972 & ~n6973 ;
  assign n6979 = ~n6974 & x229 ;
  assign n6975 = x134 & ~n5411 ;
  assign n6976 = ~x134 & ~n5403 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6980 = n6977 & ~x229 ;
  assign n6981 = ~n6979 & ~n6980 ;
  assign n6982 = ~x134 & ~n5432 ;
  assign n6983 = x134 & ~n5424 ;
  assign n6984 = ~n6982 & ~n6983 ;
  assign n6989 = ~n6984 & x230 ;
  assign n6985 = x134 & ~n5449 ;
  assign n6986 = ~x134 & ~n5441 ;
  assign n6987 = ~n6985 & ~n6986 ;
  assign n6990 = n6987 & ~x230 ;
  assign n6991 = ~n6989 & ~n6990 ;
  assign n6992 = ~x134 & ~n5470 ;
  assign n6993 = x134 & ~n5462 ;
  assign n6994 = ~n6992 & ~n6993 ;
  assign n6999 = ~n6994 & x231 ;
  assign n6995 = x134 & ~n5487 ;
  assign n6996 = ~x134 & ~n5479 ;
  assign n6997 = ~n6995 & ~n6996 ;
  assign n7000 = n6997 & ~x231 ;
  assign n7001 = ~n6999 & ~n7000 ;
  assign n7002 = ~x134 & ~n5508 ;
  assign n7003 = x134 & ~n5500 ;
  assign n7004 = ~n7002 & ~n7003 ;
  assign n7009 = ~n7004 & x232 ;
  assign n7005 = x134 & ~n5525 ;
  assign n7006 = ~x134 & ~n5517 ;
  assign n7007 = ~n7005 & ~n7006 ;
  assign n7010 = n7007 & ~x232 ;
  assign n7011 = ~n7009 & ~n7010 ;
  assign n7012 = ~x134 & ~n5546 ;
  assign n7013 = x134 & ~n5538 ;
  assign n7014 = ~n7012 & ~n7013 ;
  assign n7019 = ~n7014 & x233 ;
  assign n7015 = x134 & ~n5563 ;
  assign n7016 = ~x134 & ~n5555 ;
  assign n7017 = ~n7015 & ~n7016 ;
  assign n7020 = n7017 & ~x233 ;
  assign n7021 = ~n7019 & ~n7020 ;
  assign n7022 = ~x134 & ~n5584 ;
  assign n7023 = x134 & ~n5576 ;
  assign n7024 = ~n7022 & ~n7023 ;
  assign n7029 = ~n7024 & x234 ;
  assign n7025 = x134 & ~n5601 ;
  assign n7026 = ~x134 & ~n5593 ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7030 = n7027 & ~x234 ;
  assign n7031 = ~n7029 & ~n7030 ;
  assign n7032 = ~x134 & ~n5622 ;
  assign n7033 = x134 & ~n5614 ;
  assign n7034 = ~n7032 & ~n7033 ;
  assign n7039 = ~n7034 & x235 ;
  assign n7035 = x134 & ~n5639 ;
  assign n7036 = ~x134 & ~n5631 ;
  assign n7037 = ~n7035 & ~n7036 ;
  assign n7040 = n7037 & ~x235 ;
  assign n7041 = ~n7039 & ~n7040 ;
  assign n7042 = ~x134 & ~n5660 ;
  assign n7043 = x134 & ~n5652 ;
  assign n7044 = ~n7042 & ~n7043 ;
  assign n7049 = ~n7044 & x236 ;
  assign n7045 = x134 & ~n5677 ;
  assign n7046 = ~x134 & ~n5669 ;
  assign n7047 = ~n7045 & ~n7046 ;
  assign n7050 = n7047 & ~x236 ;
  assign n7051 = ~n7049 & ~n7050 ;
  assign n7052 = ~x134 & ~n5698 ;
  assign n7053 = x134 & ~n5690 ;
  assign n7054 = ~n7052 & ~n7053 ;
  assign n7059 = ~n7054 & x237 ;
  assign n7055 = x134 & ~n5715 ;
  assign n7056 = ~x134 & ~n5707 ;
  assign n7057 = ~n7055 & ~n7056 ;
  assign n7060 = n7057 & ~x237 ;
  assign n7061 = ~n7059 & ~n7060 ;
  assign n7062 = ~x134 & ~n5736 ;
  assign n7063 = x134 & ~n5728 ;
  assign n7064 = ~n7062 & ~n7063 ;
  assign n7069 = ~n7064 & x238 ;
  assign n7065 = x134 & ~n5753 ;
  assign n7066 = ~x134 & ~n5745 ;
  assign n7067 = ~n7065 & ~n7066 ;
  assign n7070 = n7067 & ~x238 ;
  assign n7071 = ~n7069 & ~n7070 ;
  assign n7072 = ~x134 & ~n5774 ;
  assign n7073 = x134 & ~n5766 ;
  assign n7074 = ~n7072 & ~n7073 ;
  assign n7079 = ~n7074 & x239 ;
  assign n7075 = x134 & ~n5791 ;
  assign n7076 = ~x134 & ~n5783 ;
  assign n7077 = ~n7075 & ~n7076 ;
  assign n7080 = n7077 & ~x239 ;
  assign n7081 = ~n7079 & ~n7080 ;
  assign n7082 = ~x134 & ~n5812 ;
  assign n7083 = x134 & ~n5804 ;
  assign n7084 = ~n7082 & ~n7083 ;
  assign n7089 = ~n7084 & x240 ;
  assign n7085 = x134 & ~n5829 ;
  assign n7086 = ~x134 & ~n5821 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7090 = n7087 & ~x240 ;
  assign n7091 = ~n7089 & ~n7090 ;
  assign n7092 = ~x134 & ~n5850 ;
  assign n7093 = x134 & ~n5842 ;
  assign n7094 = ~n7092 & ~n7093 ;
  assign n7099 = ~n7094 & x241 ;
  assign n7095 = x134 & ~n5867 ;
  assign n7096 = ~x134 & ~n5859 ;
  assign n7097 = ~n7095 & ~n7096 ;
  assign n7100 = n7097 & ~x241 ;
  assign n7101 = ~n7099 & ~n7100 ;
  assign n7102 = ~x134 & ~n5888 ;
  assign n7103 = x134 & ~n5880 ;
  assign n7104 = ~n7102 & ~n7103 ;
  assign n7109 = ~n7104 & x242 ;
  assign n7105 = x134 & ~n5905 ;
  assign n7106 = ~x134 & ~n5897 ;
  assign n7107 = ~n7105 & ~n7106 ;
  assign n7110 = n7107 & ~x242 ;
  assign n7111 = ~n7109 & ~n7110 ;
  assign n7112 = ~x134 & ~n5926 ;
  assign n7113 = x134 & ~n5918 ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7119 = ~n7114 & x243 ;
  assign n7115 = x134 & ~n5943 ;
  assign n7116 = ~x134 & ~n5935 ;
  assign n7117 = ~n7115 & ~n7116 ;
  assign n7120 = n7117 & ~x243 ;
  assign n7121 = ~n7119 & ~n7120 ;
  assign n7122 = ~x134 & ~n5964 ;
  assign n7123 = x134 & ~n5956 ;
  assign n7124 = ~n7122 & ~n7123 ;
  assign n7129 = ~n7124 & x244 ;
  assign n7125 = x134 & ~n5981 ;
  assign n7126 = ~x134 & ~n5973 ;
  assign n7127 = ~n7125 & ~n7126 ;
  assign n7130 = n7127 & ~x244 ;
  assign n7131 = ~n7129 & ~n7130 ;
  assign n7132 = ~x134 & ~n6002 ;
  assign n7133 = x134 & ~n5994 ;
  assign n7134 = ~n7132 & ~n7133 ;
  assign n7139 = ~n7134 & x245 ;
  assign n7135 = x134 & ~n6019 ;
  assign n7136 = ~x134 & ~n6011 ;
  assign n7137 = ~n7135 & ~n7136 ;
  assign n7140 = n7137 & ~x245 ;
  assign n7141 = ~n7139 & ~n7140 ;
  assign n7142 = ~x134 & ~n6040 ;
  assign n7143 = x134 & ~n6032 ;
  assign n7144 = ~n7142 & ~n7143 ;
  assign n7149 = ~n7144 & x246 ;
  assign n7145 = x134 & ~n6057 ;
  assign n7146 = ~x134 & ~n6049 ;
  assign n7147 = ~n7145 & ~n7146 ;
  assign n7150 = n7147 & ~x246 ;
  assign n7151 = ~n7149 & ~n7150 ;
  assign n7152 = ~x134 & ~n6078 ;
  assign n7153 = x134 & ~n6070 ;
  assign n7154 = ~n7152 & ~n7153 ;
  assign n7159 = ~n7154 & x247 ;
  assign n7155 = x134 & ~n6095 ;
  assign n7156 = ~x134 & ~n6087 ;
  assign n7157 = ~n7155 & ~n7156 ;
  assign n7160 = n7157 & ~x247 ;
  assign n7161 = ~n7159 & ~n7160 ;
  assign n7162 = ~x134 & ~n6116 ;
  assign n7163 = x134 & ~n6108 ;
  assign n7164 = ~n7162 & ~n7163 ;
  assign n7169 = ~n7164 & x248 ;
  assign n7165 = x134 & ~n6133 ;
  assign n7166 = ~x134 & ~n6125 ;
  assign n7167 = ~n7165 & ~n7166 ;
  assign n7170 = n7167 & ~x248 ;
  assign n7171 = ~n7169 & ~n7170 ;
  assign n7172 = ~x134 & ~n6154 ;
  assign n7173 = x134 & ~n6146 ;
  assign n7174 = ~n7172 & ~n7173 ;
  assign n7179 = ~n7174 & x249 ;
  assign n7175 = x134 & ~n6171 ;
  assign n7176 = ~x134 & ~n6163 ;
  assign n7177 = ~n7175 & ~n7176 ;
  assign n7180 = n7177 & ~x249 ;
  assign n7181 = ~n7179 & ~n7180 ;
  assign n7182 = ~x134 & ~n6192 ;
  assign n7183 = x134 & ~n6184 ;
  assign n7184 = ~n7182 & ~n7183 ;
  assign n7189 = ~n7184 & x250 ;
  assign n7185 = x134 & ~n6209 ;
  assign n7186 = ~x134 & ~n6201 ;
  assign n7187 = ~n7185 & ~n7186 ;
  assign n7190 = n7187 & ~x250 ;
  assign n7191 = ~n7189 & ~n7190 ;
  assign n7192 = ~x134 & ~n6230 ;
  assign n7193 = x134 & ~n6222 ;
  assign n7194 = ~n7192 & ~n7193 ;
  assign n7199 = ~n7194 & x251 ;
  assign n7195 = x134 & ~n6247 ;
  assign n7196 = ~x134 & ~n6239 ;
  assign n7197 = ~n7195 & ~n7196 ;
  assign n7200 = n7197 & ~x251 ;
  assign n7201 = ~n7199 & ~n7200 ;
  assign n7202 = ~x134 & ~n6268 ;
  assign n7203 = x134 & ~n6260 ;
  assign n7204 = ~n7202 & ~n7203 ;
  assign n7209 = ~n7204 & x252 ;
  assign n7205 = x134 & ~n6285 ;
  assign n7206 = ~x134 & ~n6277 ;
  assign n7207 = ~n7205 & ~n7206 ;
  assign n7210 = n7207 & ~x252 ;
  assign n7211 = ~n7209 & ~n7210 ;
  assign n7212 = ~x134 & ~n6306 ;
  assign n7213 = x134 & ~n6298 ;
  assign n7214 = ~n7212 & ~n7213 ;
  assign n7219 = ~n7214 & x253 ;
  assign n7215 = x134 & ~n6323 ;
  assign n7216 = ~x134 & ~n6315 ;
  assign n7217 = ~n7215 & ~n7216 ;
  assign n7220 = n7217 & ~x253 ;
  assign n7221 = ~n7219 & ~n7220 ;
  assign n7222 = ~x134 & ~n6344 ;
  assign n7223 = x134 & ~n6336 ;
  assign n7224 = ~n7222 & ~n7223 ;
  assign n7229 = ~n7224 & x254 ;
  assign n7225 = x134 & ~n6361 ;
  assign n7226 = ~x134 & ~n6353 ;
  assign n7227 = ~n7225 & ~n7226 ;
  assign n7230 = n7227 & ~x254 ;
  assign n7231 = ~n7229 & ~n7230 ;
  assign n7232 = ~x134 & ~n6382 ;
  assign n7233 = x134 & ~n6374 ;
  assign n7234 = ~n7232 & ~n7233 ;
  assign n7239 = ~n7234 & x255 ;
  assign n7235 = x134 & ~n6399 ;
  assign n7236 = ~x134 & ~n6391 ;
  assign n7237 = ~n7235 & ~n7236 ;
  assign n7240 = n7237 & ~x255 ;
  assign n7241 = ~n7239 & ~n7240 ;
  assign n7242 = ~x134 & ~n6420 ;
  assign n7243 = x134 & ~n6412 ;
  assign n7244 = ~n7242 & ~n7243 ;
  assign n7249 = ~n7244 & x256 ;
  assign n7245 = x134 & ~n6437 ;
  assign n7246 = ~x134 & ~n6429 ;
  assign n7247 = ~n7245 & ~n7246 ;
  assign n7250 = n7247 & ~x256 ;
  assign n7251 = ~n7249 & ~n7250 ;
  assign n7252 = ~x134 & ~n6458 ;
  assign n7253 = x134 & ~n6450 ;
  assign n7254 = ~n7252 & ~n7253 ;
  assign n7259 = ~n7254 & x257 ;
  assign n7255 = x134 & ~n6475 ;
  assign n7256 = ~x134 & ~n6467 ;
  assign n7257 = ~n7255 & ~n7256 ;
  assign n7260 = n7257 & ~x257 ;
  assign n7261 = ~n7259 & ~n7260 ;
  assign n7262 = ~x134 & ~n6496 ;
  assign n7263 = x134 & ~n6488 ;
  assign n7264 = ~n7262 & ~n7263 ;
  assign n7269 = ~n7264 & x258 ;
  assign n7265 = x134 & ~n6513 ;
  assign n7266 = ~x134 & ~n6505 ;
  assign n7267 = ~n7265 & ~n7266 ;
  assign n7270 = n7267 & ~x258 ;
  assign n7271 = ~n7269 & ~n7270 ;
  assign n7272 = ~x134 & ~n6534 ;
  assign n7273 = x134 & ~n6526 ;
  assign n7274 = ~n7272 & ~n7273 ;
  assign n7279 = ~n7274 & x259 ;
  assign n7275 = x134 & ~n6551 ;
  assign n7276 = ~x134 & ~n6543 ;
  assign n7277 = ~n7275 & ~n7276 ;
  assign n7280 = n7277 & ~x259 ;
  assign n7281 = ~n7279 & ~n7280 ;
  assign n7282 = ~x134 & ~n6572 ;
  assign n7283 = x134 & ~n6564 ;
  assign n7284 = ~n7282 & ~n7283 ;
  assign n7289 = ~n7284 & x260 ;
  assign n7285 = x134 & ~n6589 ;
  assign n7286 = ~x134 & ~n6581 ;
  assign n7287 = ~n7285 & ~n7286 ;
  assign n7290 = n7287 & ~x260 ;
  assign n7291 = ~n7289 & ~n7290 ;
  assign n7292 = ~x134 & ~n6610 ;
  assign n7293 = x134 & ~n6602 ;
  assign n7294 = ~n7292 & ~n7293 ;
  assign n7299 = ~n7294 & x261 ;
  assign n7295 = x134 & ~n6627 ;
  assign n7296 = ~x134 & ~n6619 ;
  assign n7297 = ~n7295 & ~n7296 ;
  assign n7300 = n7297 & ~x261 ;
  assign n7301 = ~n7299 & ~n7300 ;
  assign n7302 = ~x134 & ~n6648 ;
  assign n7303 = x134 & ~n6640 ;
  assign n7304 = ~n7302 & ~n7303 ;
  assign n7309 = ~n7304 & x262 ;
  assign n7305 = x134 & ~n6665 ;
  assign n7306 = ~x134 & ~n6657 ;
  assign n7307 = ~n7305 & ~n7306 ;
  assign n7310 = n7307 & ~x262 ;
  assign n7311 = ~n7309 & ~n7310 ;
  assign y0 = ~n997 ;
  assign y1 = ~n1851 ;
  assign y2 = ~n2449 ;
  assign y3 = ~n3047 ;
  assign y4 = ~n3197 ;
  assign y5 = ~n3347 ;
  assign y6 = ~n3497 ;
  assign y7 = ~n3647 ;
  assign y8 = ~n3797 ;
  assign y9 = ~n3947 ;
  assign y10 = ~n4097 ;
  assign y11 = ~n4247 ;
  assign y12 = ~n4397 ;
  assign y13 = ~n4547 ;
  assign y14 = ~n4697 ;
  assign y15 = ~n4847 ;
  assign y16 = ~n4885 ;
  assign y17 = ~n4923 ;
  assign y18 = ~n4961 ;
  assign y19 = ~n4999 ;
  assign y20 = ~n5037 ;
  assign y21 = ~n5075 ;
  assign y22 = ~n5113 ;
  assign y23 = ~n5151 ;
  assign y24 = ~n5189 ;
  assign y25 = ~n5227 ;
  assign y26 = ~n5265 ;
  assign y27 = ~n5303 ;
  assign y28 = ~n5341 ;
  assign y29 = ~n5379 ;
  assign y30 = ~n5417 ;
  assign y31 = ~n5455 ;
  assign y32 = ~n5493 ;
  assign y33 = ~n5531 ;
  assign y34 = ~n5569 ;
  assign y35 = ~n5607 ;
  assign y36 = ~n5645 ;
  assign y37 = ~n5683 ;
  assign y38 = ~n5721 ;
  assign y39 = ~n5759 ;
  assign y40 = ~n5797 ;
  assign y41 = ~n5835 ;
  assign y42 = ~n5873 ;
  assign y43 = ~n5911 ;
  assign y44 = ~n5949 ;
  assign y45 = ~n5987 ;
  assign y46 = ~n6025 ;
  assign y47 = ~n6063 ;
  assign y48 = ~n6101 ;
  assign y49 = ~n6139 ;
  assign y50 = ~n6177 ;
  assign y51 = ~n6215 ;
  assign y52 = ~n6253 ;
  assign y53 = ~n6291 ;
  assign y54 = ~n6329 ;
  assign y55 = ~n6367 ;
  assign y56 = ~n6405 ;
  assign y57 = ~n6443 ;
  assign y58 = ~n6481 ;
  assign y59 = ~n6519 ;
  assign y60 = ~n6557 ;
  assign y61 = ~n6595 ;
  assign y62 = ~n6633 ;
  assign y63 = ~n6671 ;
  assign y64 = ~n6681 ;
  assign y65 = ~n6691 ;
  assign y66 = ~n6701 ;
  assign y67 = ~n6711 ;
  assign y68 = ~n6721 ;
  assign y69 = ~n6731 ;
  assign y70 = ~n6741 ;
  assign y71 = ~n6751 ;
  assign y72 = ~n6761 ;
  assign y73 = ~n6771 ;
  assign y74 = ~n6781 ;
  assign y75 = ~n6791 ;
  assign y76 = ~n6801 ;
  assign y77 = ~n6811 ;
  assign y78 = ~n6821 ;
  assign y79 = ~n6831 ;
  assign y80 = ~n6841 ;
  assign y81 = ~n6851 ;
  assign y82 = ~n6861 ;
  assign y83 = ~n6871 ;
  assign y84 = ~n6881 ;
  assign y85 = ~n6891 ;
  assign y86 = ~n6901 ;
  assign y87 = ~n6911 ;
  assign y88 = ~n6921 ;
  assign y89 = ~n6931 ;
  assign y90 = ~n6941 ;
  assign y91 = ~n6951 ;
  assign y92 = ~n6961 ;
  assign y93 = ~n6971 ;
  assign y94 = ~n6981 ;
  assign y95 = ~n6991 ;
  assign y96 = ~n7001 ;
  assign y97 = ~n7011 ;
  assign y98 = ~n7021 ;
  assign y99 = ~n7031 ;
  assign y100 = ~n7041 ;
  assign y101 = ~n7051 ;
  assign y102 = ~n7061 ;
  assign y103 = ~n7071 ;
  assign y104 = ~n7081 ;
  assign y105 = ~n7091 ;
  assign y106 = ~n7101 ;
  assign y107 = ~n7111 ;
  assign y108 = ~n7121 ;
  assign y109 = ~n7131 ;
  assign y110 = ~n7141 ;
  assign y111 = ~n7151 ;
  assign y112 = ~n7161 ;
  assign y113 = ~n7171 ;
  assign y114 = ~n7181 ;
  assign y115 = ~n7191 ;
  assign y116 = ~n7201 ;
  assign y117 = ~n7211 ;
  assign y118 = ~n7221 ;
  assign y119 = ~n7231 ;
  assign y120 = ~n7241 ;
  assign y121 = ~n7251 ;
  assign y122 = ~n7261 ;
  assign y123 = ~n7271 ;
  assign y124 = ~n7281 ;
  assign y125 = ~n7291 ;
  assign y126 = ~n7301 ;
  assign y127 = ~n7311 ;
endmodule
