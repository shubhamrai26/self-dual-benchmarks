module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 ;
  assign n256 = x233 ^ x103 ^ x6 ;
  assign n257 = x77 & x159 ;
  assign n258 = n257 ^ x238 ^ 1'b0 ;
  assign n259 = n258 ^ x135 ^ x99 ;
  assign n260 = x30 ^ x26 ^ x23 ;
  assign n261 = x240 ^ x127 ^ 1'b0 ;
  assign n262 = ~n260 & n261 ;
  assign n263 = n262 ^ x231 ^ x177 ;
  assign n264 = n263 ^ x191 ^ x32 ;
  assign n265 = ( ~x98 & x143 ) | ( ~x98 & x233 ) | ( x143 & x233 ) ;
  assign n266 = x207 ^ x2 ^ 1'b0 ;
  assign n267 = x211 & n266 ;
  assign n268 = n267 ^ x67 ^ 1'b0 ;
  assign n269 = x58 & n268 ;
  assign n270 = ( x33 & x117 ) | ( x33 & ~x215 ) | ( x117 & ~x215 ) ;
  assign n271 = ( x25 & x222 ) | ( x25 & ~n270 ) | ( x222 & ~n270 ) ;
  assign n272 = ( x25 & x88 ) | ( x25 & ~x134 ) | ( x88 & ~x134 ) ;
  assign n273 = n272 ^ x243 ^ x95 ;
  assign n274 = x29 & x219 ;
  assign n275 = ~x180 & n274 ;
  assign n276 = x118 ^ x89 ^ 1'b0 ;
  assign n277 = ( x29 & ~x211 ) | ( x29 & n276 ) | ( ~x211 & n276 ) ;
  assign n278 = x237 ^ x115 ^ x70 ;
  assign n279 = ( ~x49 & x159 ) | ( ~x49 & n269 ) | ( x159 & n269 ) ;
  assign n280 = x234 ^ x226 ^ x13 ;
  assign n281 = n280 ^ x247 ^ x112 ;
  assign n282 = n281 ^ x254 ^ x25 ;
  assign n283 = ( x44 & ~x132 ) | ( x44 & x238 ) | ( ~x132 & x238 ) ;
  assign n284 = ( ~x73 & x244 ) | ( ~x73 & n283 ) | ( x244 & n283 ) ;
  assign n285 = x92 ^ x13 ^ 1'b0 ;
  assign n286 = x50 & n285 ;
  assign n287 = ( ~x80 & x221 ) | ( ~x80 & n286 ) | ( x221 & n286 ) ;
  assign n288 = x231 ^ x135 ^ x85 ;
  assign n289 = x99 & x247 ;
  assign n290 = n289 ^ x97 ^ 1'b0 ;
  assign n291 = x62 ^ x53 ^ 1'b0 ;
  assign n292 = x11 & n291 ;
  assign n293 = ( ~x108 & x138 ) | ( ~x108 & n292 ) | ( x138 & n292 ) ;
  assign n294 = n293 ^ x104 ^ x79 ;
  assign n295 = ( ~x7 & x13 ) | ( ~x7 & x104 ) | ( x13 & x104 ) ;
  assign n296 = ( x61 & x140 ) | ( x61 & ~n295 ) | ( x140 & ~n295 ) ;
  assign n297 = ( ~x191 & x197 ) | ( ~x191 & n296 ) | ( x197 & n296 ) ;
  assign n298 = x44 & x254 ;
  assign n299 = ~x235 & n298 ;
  assign n300 = x195 & x234 ;
  assign n301 = n288 & n300 ;
  assign n302 = n301 ^ x136 ^ x131 ;
  assign n303 = ( x96 & ~x101 ) | ( x96 & x184 ) | ( ~x101 & x184 ) ;
  assign n304 = ( x203 & ~x216 ) | ( x203 & n303 ) | ( ~x216 & n303 ) ;
  assign n305 = x125 ^ x84 ^ x68 ;
  assign n306 = n305 ^ n258 ^ x112 ;
  assign n307 = n306 ^ x194 ^ x135 ;
  assign n308 = x213 ^ x165 ^ 1'b0 ;
  assign n309 = x10 & n308 ;
  assign n310 = n309 ^ x110 ^ 1'b0 ;
  assign n311 = ( x3 & ~n256 ) | ( x3 & n310 ) | ( ~n256 & n310 ) ;
  assign n312 = n260 ^ x139 ^ x93 ;
  assign n313 = ( x7 & ~x120 ) | ( x7 & n312 ) | ( ~x120 & n312 ) ;
  assign n314 = x191 & x220 ;
  assign n315 = n314 ^ x145 ^ 1'b0 ;
  assign n316 = ( ~x34 & x143 ) | ( ~x34 & n315 ) | ( x143 & n315 ) ;
  assign n317 = x63 ^ x58 ^ x1 ;
  assign n318 = n317 ^ n316 ^ x240 ;
  assign n320 = n258 ^ x118 ^ x95 ;
  assign n319 = ( x162 & ~x179 ) | ( x162 & n303 ) | ( ~x179 & n303 ) ;
  assign n321 = n320 ^ n319 ^ x156 ;
  assign n322 = x202 & x247 ;
  assign n323 = n322 ^ x38 ^ 1'b0 ;
  assign n324 = ( ~x43 & x88 ) | ( ~x43 & x196 ) | ( x88 & x196 ) ;
  assign n325 = x217 ^ x122 ^ 1'b0 ;
  assign n326 = x232 & n325 ;
  assign n327 = ( x48 & ~n324 ) | ( x48 & n326 ) | ( ~n324 & n326 ) ;
  assign n328 = ( ~x107 & x229 ) | ( ~x107 & n308 ) | ( x229 & n308 ) ;
  assign n329 = x143 ^ x141 ^ 1'b0 ;
  assign n330 = x118 & n329 ;
  assign n331 = ( x33 & x122 ) | ( x33 & ~n330 ) | ( x122 & ~n330 ) ;
  assign n332 = ( x82 & ~x148 ) | ( x82 & n331 ) | ( ~x148 & n331 ) ;
  assign n333 = ( x159 & x176 ) | ( x159 & ~n332 ) | ( x176 & ~n332 ) ;
  assign n334 = x91 ^ x82 ^ x35 ;
  assign n335 = n334 ^ x205 ^ x24 ;
  assign n339 = ( x18 & x171 ) | ( x18 & ~x195 ) | ( x171 & ~x195 ) ;
  assign n340 = n339 ^ x205 ^ x150 ;
  assign n341 = n340 ^ n258 ^ x94 ;
  assign n337 = ( x24 & x38 ) | ( x24 & ~x145 ) | ( x38 & ~x145 ) ;
  assign n336 = x204 ^ x127 ^ 1'b0 ;
  assign n338 = n337 ^ n336 ^ x84 ;
  assign n342 = n341 ^ n338 ^ x172 ;
  assign n346 = ( x124 & ~x138 ) | ( x124 & n324 ) | ( ~x138 & n324 ) ;
  assign n348 = ( ~x120 & x198 ) | ( ~x120 & x234 ) | ( x198 & x234 ) ;
  assign n347 = x104 ^ x31 ^ x5 ;
  assign n349 = n348 ^ n347 ^ 1'b0 ;
  assign n350 = x109 & ~n349 ;
  assign n351 = x171 & n350 ;
  assign n352 = n351 ^ x130 ^ 1'b0 ;
  assign n353 = ( x9 & n346 ) | ( x9 & n352 ) | ( n346 & n352 ) ;
  assign n344 = x58 ^ x45 ^ 1'b0 ;
  assign n345 = x172 & n344 ;
  assign n343 = x208 ^ x153 ^ x13 ;
  assign n354 = n353 ^ n345 ^ n343 ;
  assign n358 = n297 ^ x79 ^ 1'b0 ;
  assign n359 = ~n305 & n358 ;
  assign n355 = ( x82 & x235 ) | ( x82 & ~x241 ) | ( x235 & ~x241 ) ;
  assign n356 = ( x130 & ~n293 ) | ( x130 & n355 ) | ( ~n293 & n355 ) ;
  assign n357 = n356 ^ n324 ^ x154 ;
  assign n360 = n359 ^ n357 ^ 1'b0 ;
  assign n361 = n276 & ~n360 ;
  assign n362 = ( ~x109 & x129 ) | ( ~x109 & x165 ) | ( x129 & x165 ) ;
  assign n363 = ( x39 & ~x204 ) | ( x39 & n362 ) | ( ~x204 & n362 ) ;
  assign n364 = ( ~x142 & x173 ) | ( ~x142 & n363 ) | ( x173 & n363 ) ;
  assign n365 = x186 & ~n354 ;
  assign n370 = x163 ^ x154 ^ x22 ;
  assign n368 = ( ~x13 & x224 ) | ( ~x13 & n283 ) | ( x224 & n283 ) ;
  assign n366 = ( x18 & ~x249 ) | ( x18 & x254 ) | ( ~x249 & x254 ) ;
  assign n367 = n366 ^ x225 ^ x93 ;
  assign n369 = n368 ^ n367 ^ x232 ;
  assign n371 = n370 ^ n369 ^ n366 ;
  assign n372 = x206 ^ x114 ^ x107 ;
  assign n373 = ( ~x14 & x157 ) | ( ~x14 & x209 ) | ( x157 & x209 ) ;
  assign n374 = ( n333 & n372 ) | ( n333 & n373 ) | ( n372 & n373 ) ;
  assign n375 = ( x31 & x226 ) | ( x31 & ~x227 ) | ( x226 & ~x227 ) ;
  assign n378 = n263 ^ x109 ^ x17 ;
  assign n376 = x216 & ~n273 ;
  assign n377 = ~x81 & n376 ;
  assign n379 = n378 ^ n377 ^ x112 ;
  assign n380 = n370 ^ n333 ^ 1'b0 ;
  assign n381 = x111 & x126 ;
  assign n382 = ~x31 & n381 ;
  assign n383 = ( n282 & ~n320 ) | ( n282 & n366 ) | ( ~n320 & n366 ) ;
  assign n384 = ( x115 & n382 ) | ( x115 & ~n383 ) | ( n382 & ~n383 ) ;
  assign n391 = n317 ^ x90 ^ x18 ;
  assign n392 = ( ~x78 & n296 ) | ( ~x78 & n391 ) | ( n296 & n391 ) ;
  assign n388 = ( x115 & ~x167 ) | ( x115 & n259 ) | ( ~x167 & n259 ) ;
  assign n389 = n388 ^ n271 ^ x5 ;
  assign n385 = ~x106 & x254 ;
  assign n386 = x61 & x203 ;
  assign n387 = n385 & n386 ;
  assign n390 = n389 ^ n387 ^ x241 ;
  assign n393 = n392 ^ n390 ^ x80 ;
  assign n394 = ( ~x208 & x215 ) | ( ~x208 & n292 ) | ( x215 & n292 ) ;
  assign n395 = ( x91 & ~x201 ) | ( x91 & x237 ) | ( ~x201 & x237 ) ;
  assign n396 = x105 ^ x103 ^ x53 ;
  assign n397 = x203 | n396 ;
  assign n398 = n395 & n397 ;
  assign n399 = n398 ^ x8 ^ 1'b0 ;
  assign n400 = ( x15 & ~x231 ) | ( x15 & n399 ) | ( ~x231 & n399 ) ;
  assign n401 = x202 ^ x65 ^ x2 ;
  assign n402 = ( x95 & n369 ) | ( x95 & n401 ) | ( n369 & n401 ) ;
  assign n403 = n336 ^ x44 ^ 1'b0 ;
  assign n404 = x13 & x80 ;
  assign n405 = n404 ^ n321 ^ 1'b0 ;
  assign n406 = x89 ^ x66 ^ x25 ;
  assign n407 = ( x12 & x141 ) | ( x12 & n406 ) | ( x141 & n406 ) ;
  assign n408 = n306 | n407 ;
  assign n409 = n299 ^ x26 ^ 1'b0 ;
  assign n410 = ( ~x53 & x152 ) | ( ~x53 & n409 ) | ( x152 & n409 ) ;
  assign n414 = ( x68 & x175 ) | ( x68 & ~x218 ) | ( x175 & ~x218 ) ;
  assign n412 = n312 ^ x97 ^ x52 ;
  assign n411 = n366 ^ x166 ^ x96 ;
  assign n413 = n412 ^ n411 ^ x169 ;
  assign n415 = n414 ^ n413 ^ x200 ;
  assign n416 = n415 ^ n272 ^ x30 ;
  assign n417 = ( x233 & n364 ) | ( x233 & n416 ) | ( n364 & n416 ) ;
  assign n418 = ( x171 & ~n391 ) | ( x171 & n417 ) | ( ~n391 & n417 ) ;
  assign n419 = n418 ^ x86 ^ 1'b0 ;
  assign n420 = ~n410 & n419 ;
  assign n423 = x240 ^ x209 ^ x54 ;
  assign n424 = x227 | n423 ;
  assign n425 = ( ~x34 & x203 ) | ( ~x34 & x223 ) | ( x203 & x223 ) ;
  assign n426 = ( ~x113 & n312 ) | ( ~x113 & n425 ) | ( n312 & n425 ) ;
  assign n427 = ( ~x215 & n424 ) | ( ~x215 & n426 ) | ( n424 & n426 ) ;
  assign n421 = n414 ^ x156 ^ 1'b0 ;
  assign n422 = x25 & n421 ;
  assign n428 = n427 ^ n422 ^ 1'b0 ;
  assign n435 = x12 & x151 ;
  assign n436 = ~x252 & n435 ;
  assign n429 = x59 & x200 ;
  assign n430 = n429 ^ x216 ^ 1'b0 ;
  assign n431 = ( x82 & x164 ) | ( x82 & n430 ) | ( x164 & n430 ) ;
  assign n432 = x252 ^ x109 ^ 1'b0 ;
  assign n433 = x242 & n432 ;
  assign n434 = ~n431 & n433 ;
  assign n437 = n436 ^ n434 ^ n341 ;
  assign n438 = x152 ^ x25 ^ 1'b0 ;
  assign n439 = n437 & n438 ;
  assign n440 = ( x130 & ~x235 ) | ( x130 & x252 ) | ( ~x235 & x252 ) ;
  assign n444 = x240 & ~n315 ;
  assign n445 = n444 ^ x81 ^ 1'b0 ;
  assign n442 = ( x8 & ~n271 ) | ( x8 & n302 ) | ( ~n271 & n302 ) ;
  assign n441 = x210 ^ x7 ^ x6 ;
  assign n443 = n442 ^ n441 ^ x192 ;
  assign n446 = n445 ^ n443 ^ 1'b0 ;
  assign n447 = ( x5 & n440 ) | ( x5 & n446 ) | ( n440 & n446 ) ;
  assign n450 = x9 & n267 ;
  assign n451 = ~x246 & n450 ;
  assign n448 = ( ~x28 & x215 ) | ( ~x28 & x242 ) | ( x215 & x242 ) ;
  assign n449 = ~n370 & n448 ;
  assign n452 = n451 ^ n449 ^ 1'b0 ;
  assign n453 = ( n272 & n383 ) | ( n272 & n452 ) | ( n383 & n452 ) ;
  assign n454 = x70 & n345 ;
  assign n455 = ~x250 & n454 ;
  assign n456 = x187 ^ x20 ^ 1'b0 ;
  assign n457 = x185 & n456 ;
  assign n458 = ~n315 & n457 ;
  assign n459 = n423 & n458 ;
  assign n460 = n459 ^ n301 ^ x175 ;
  assign n461 = ( ~x39 & x130 ) | ( ~x39 & x203 ) | ( x130 & x203 ) ;
  assign n462 = ( ~x108 & n307 ) | ( ~x108 & n461 ) | ( n307 & n461 ) ;
  assign n464 = ( x72 & ~x172 ) | ( x72 & x177 ) | ( ~x172 & x177 ) ;
  assign n465 = ( x44 & ~x63 ) | ( x44 & n464 ) | ( ~x63 & n464 ) ;
  assign n463 = n336 ^ x150 ^ x67 ;
  assign n466 = n465 ^ n463 ^ x92 ;
  assign n467 = x80 & ~n323 ;
  assign n468 = ~n308 & n467 ;
  assign n469 = ( x5 & x59 ) | ( x5 & ~x97 ) | ( x59 & ~x97 ) ;
  assign n470 = x171 ^ x122 ^ 1'b0 ;
  assign n471 = x132 & n470 ;
  assign n472 = ( x144 & n370 ) | ( x144 & n471 ) | ( n370 & n471 ) ;
  assign n473 = n414 ^ x215 ^ x85 ;
  assign n474 = ( x127 & x243 ) | ( x127 & n473 ) | ( x243 & n473 ) ;
  assign n475 = x247 ^ x172 ^ x82 ;
  assign n476 = ( x19 & x222 ) | ( x19 & n475 ) | ( x222 & n475 ) ;
  assign n477 = ( x237 & n474 ) | ( x237 & ~n476 ) | ( n474 & ~n476 ) ;
  assign n478 = ( n395 & n472 ) | ( n395 & ~n477 ) | ( n472 & ~n477 ) ;
  assign n479 = x11 & ~n478 ;
  assign n480 = ~x134 & x138 ;
  assign n481 = x149 & x219 ;
  assign n482 = ~x61 & n481 ;
  assign n483 = x192 & n313 ;
  assign n484 = ~x97 & n483 ;
  assign n485 = n484 ^ n355 ^ x176 ;
  assign n486 = ( x80 & n482 ) | ( x80 & n485 ) | ( n482 & n485 ) ;
  assign n487 = n486 ^ n468 ^ x118 ;
  assign n488 = ( ~x26 & n480 ) | ( ~x26 & n487 ) | ( n480 & n487 ) ;
  assign n489 = x101 & n457 ;
  assign n490 = ~x102 & n489 ;
  assign n491 = ( ~x109 & n337 ) | ( ~x109 & n490 ) | ( n337 & n490 ) ;
  assign n492 = ( x179 & ~n350 ) | ( x179 & n491 ) | ( ~n350 & n491 ) ;
  assign n493 = x219 & ~n327 ;
  assign n494 = ( ~n294 & n492 ) | ( ~n294 & n493 ) | ( n492 & n493 ) ;
  assign n495 = ( ~x246 & n312 ) | ( ~x246 & n494 ) | ( n312 & n494 ) ;
  assign n496 = x237 ^ x234 ^ x171 ;
  assign n497 = n496 ^ n409 ^ 1'b0 ;
  assign n498 = n393 & n497 ;
  assign n499 = x115 & ~n263 ;
  assign n500 = n499 ^ x134 ^ 1'b0 ;
  assign n501 = n500 ^ n432 ^ x115 ;
  assign n502 = x237 ^ x217 ^ x155 ;
  assign n503 = ( x43 & n501 ) | ( x43 & n502 ) | ( n501 & n502 ) ;
  assign n504 = ( x181 & ~n498 ) | ( x181 & n503 ) | ( ~n498 & n503 ) ;
  assign n505 = ( x27 & x99 ) | ( x27 & ~x238 ) | ( x99 & ~x238 ) ;
  assign n506 = n505 ^ n354 ^ x215 ;
  assign n507 = n506 ^ x156 ^ 1'b0 ;
  assign n508 = n504 & ~n507 ;
  assign n509 = x167 & n476 ;
  assign n510 = x166 & x204 ;
  assign n511 = ~x240 & n510 ;
  assign n512 = ( n492 & n509 ) | ( n492 & ~n511 ) | ( n509 & ~n511 ) ;
  assign n513 = n312 ^ x167 ^ 1'b0 ;
  assign n514 = ~n389 & n513 ;
  assign n515 = x27 & x86 ;
  assign n516 = ~x166 & n515 ;
  assign n517 = n516 ^ x170 ^ x83 ;
  assign n518 = ( x209 & x232 ) | ( x209 & ~x252 ) | ( x232 & ~x252 ) ;
  assign n519 = n518 ^ x98 ^ x13 ;
  assign n520 = x136 & ~n389 ;
  assign n521 = ~x70 & n520 ;
  assign n522 = ( ~n484 & n519 ) | ( ~n484 & n521 ) | ( n519 & n521 ) ;
  assign n523 = ( n514 & n517 ) | ( n514 & n522 ) | ( n517 & n522 ) ;
  assign n524 = n276 & ~n315 ;
  assign n525 = ~x24 & n524 ;
  assign n526 = n525 ^ n493 ^ 1'b0 ;
  assign n527 = x224 ^ x163 ^ 1'b0 ;
  assign n528 = x106 & n527 ;
  assign n529 = n312 ^ n258 ^ n256 ;
  assign n530 = ( x168 & ~x201 ) | ( x168 & x232 ) | ( ~x201 & x232 ) ;
  assign n531 = ( ~x130 & n529 ) | ( ~x130 & n530 ) | ( n529 & n530 ) ;
  assign n532 = ( x27 & ~n528 ) | ( x27 & n531 ) | ( ~n528 & n531 ) ;
  assign n533 = x165 & ~n318 ;
  assign n534 = n533 ^ x79 ^ 1'b0 ;
  assign n535 = n388 & n534 ;
  assign n536 = ( x151 & ~x201 ) | ( x151 & n482 ) | ( ~x201 & n482 ) ;
  assign n537 = n536 ^ x205 ^ x72 ;
  assign n538 = ( x171 & n535 ) | ( x171 & ~n537 ) | ( n535 & ~n537 ) ;
  assign n539 = ( x142 & n281 ) | ( x142 & ~n327 ) | ( n281 & ~n327 ) ;
  assign n546 = n530 ^ n283 ^ x129 ;
  assign n540 = ( x8 & ~x119 ) | ( x8 & x173 ) | ( ~x119 & x173 ) ;
  assign n542 = ( ~x0 & x62 ) | ( ~x0 & x97 ) | ( x62 & x97 ) ;
  assign n541 = x222 ^ x73 ^ x53 ;
  assign n543 = n542 ^ n541 ^ n490 ;
  assign n544 = n540 & n543 ;
  assign n545 = n544 ^ n490 ^ x82 ;
  assign n547 = n546 ^ n545 ^ n382 ;
  assign n548 = ( x156 & n539 ) | ( x156 & ~n547 ) | ( n539 & ~n547 ) ;
  assign n549 = ( ~n286 & n315 ) | ( ~n286 & n384 ) | ( n315 & n384 ) ;
  assign n550 = n335 & ~n549 ;
  assign n551 = n550 ^ x99 ^ 1'b0 ;
  assign n552 = ( ~x140 & x212 ) | ( ~x140 & n348 ) | ( x212 & n348 ) ;
  assign n553 = n346 ^ n328 ^ 1'b0 ;
  assign n554 = x36 | n273 ;
  assign n555 = n554 ^ x236 ^ x28 ;
  assign n556 = ( n552 & n553 ) | ( n552 & n555 ) | ( n553 & n555 ) ;
  assign n557 = ( x122 & n267 ) | ( x122 & ~n556 ) | ( n267 & ~n556 ) ;
  assign n560 = x63 & x206 ;
  assign n561 = n560 ^ n465 ^ 1'b0 ;
  assign n562 = ( x168 & n414 ) | ( x168 & n561 ) | ( n414 & n561 ) ;
  assign n563 = x67 & n562 ;
  assign n564 = ~x114 & n563 ;
  assign n558 = ( x101 & n345 ) | ( x101 & n475 ) | ( n345 & n475 ) ;
  assign n559 = x96 & n558 ;
  assign n565 = n564 ^ n559 ^ x87 ;
  assign n566 = ( ~x25 & n372 ) | ( ~x25 & n565 ) | ( n372 & n565 ) ;
  assign n567 = n281 ^ x134 ^ x68 ;
  assign n568 = n269 ^ x248 ^ x134 ;
  assign n569 = ( x6 & n567 ) | ( x6 & n568 ) | ( n567 & n568 ) ;
  assign n570 = x187 & ~n569 ;
  assign n571 = n570 ^ n308 ^ 1'b0 ;
  assign n572 = n418 & n571 ;
  assign n584 = x15 & x16 ;
  assign n585 = n584 ^ x219 ^ 1'b0 ;
  assign n586 = n585 ^ n348 ^ 1'b0 ;
  assign n587 = n352 | n586 ;
  assign n588 = n587 ^ n413 ^ x89 ;
  assign n573 = x75 & x139 ;
  assign n574 = n573 ^ x134 ^ 1'b0 ;
  assign n575 = n574 ^ n301 ^ x120 ;
  assign n576 = n575 ^ n272 ^ x214 ;
  assign n577 = n576 ^ x7 ^ 1'b0 ;
  assign n578 = n577 ^ x122 ^ x70 ;
  assign n579 = x189 ^ x34 ^ x33 ;
  assign n580 = n579 ^ n330 ^ x241 ;
  assign n581 = ( x227 & n308 ) | ( x227 & ~n580 ) | ( n308 & ~n580 ) ;
  assign n582 = ( n272 & ~n284 ) | ( n272 & n581 ) | ( ~n284 & n581 ) ;
  assign n583 = ( ~n328 & n578 ) | ( ~n328 & n582 ) | ( n578 & n582 ) ;
  assign n589 = n588 ^ n583 ^ 1'b0 ;
  assign n596 = ( ~x39 & x76 ) | ( ~x39 & n492 ) | ( x76 & n492 ) ;
  assign n594 = x230 ^ x198 ^ x14 ;
  assign n595 = n594 ^ x158 ^ 1'b0 ;
  assign n590 = ( x125 & n299 ) | ( x125 & n471 ) | ( n299 & n471 ) ;
  assign n591 = ~n506 & n590 ;
  assign n592 = ~n503 & n591 ;
  assign n593 = ( ~x34 & x100 ) | ( ~x34 & n592 ) | ( x100 & n592 ) ;
  assign n597 = n596 ^ n595 ^ n593 ;
  assign n598 = n597 ^ n492 ^ 1'b0 ;
  assign n599 = n589 & ~n598 ;
  assign n601 = ( ~x184 & n260 ) | ( ~x184 & n461 ) | ( n260 & n461 ) ;
  assign n600 = x128 ^ x32 ^ 1'b0 ;
  assign n602 = n601 ^ n600 ^ n554 ;
  assign n603 = x106 & ~n317 ;
  assign n604 = ~x121 & n603 ;
  assign n605 = n406 ^ x52 ^ 1'b0 ;
  assign n606 = n604 | n605 ;
  assign n611 = n367 ^ x172 ^ x162 ;
  assign n607 = n368 ^ x187 ^ 1'b0 ;
  assign n608 = n607 ^ n540 ^ n332 ;
  assign n609 = n283 ^ x249 ^ 1'b0 ;
  assign n610 = ~n608 & n609 ;
  assign n612 = n611 ^ n610 ^ x80 ;
  assign n613 = ( ~x42 & x57 ) | ( ~x42 & n331 ) | ( x57 & n331 ) ;
  assign n614 = ( x3 & ~x43 ) | ( x3 & n422 ) | ( ~x43 & n422 ) ;
  assign n615 = n614 ^ n611 ^ 1'b0 ;
  assign n616 = x81 & x92 ;
  assign n617 = ~x43 & n616 ;
  assign n618 = x27 & n464 ;
  assign n619 = n618 ^ x10 ^ 1'b0 ;
  assign n620 = ( n525 & n617 ) | ( n525 & ~n619 ) | ( n617 & ~n619 ) ;
  assign n625 = x184 ^ x43 ^ 1'b0 ;
  assign n626 = n519 & n625 ;
  assign n623 = n271 ^ x149 ^ x48 ;
  assign n621 = n440 ^ n346 ^ x254 ;
  assign n622 = ( x234 & n455 ) | ( x234 & ~n621 ) | ( n455 & ~n621 ) ;
  assign n624 = n623 ^ n622 ^ 1'b0 ;
  assign n627 = n626 ^ n624 ^ 1'b0 ;
  assign n628 = n324 & ~n627 ;
  assign n631 = x217 ^ x54 ^ 1'b0 ;
  assign n629 = x193 ^ x42 ^ 1'b0 ;
  assign n630 = n596 | n629 ;
  assign n632 = n631 ^ n630 ^ x167 ;
  assign n634 = n579 ^ x143 ^ x16 ;
  assign n633 = n292 ^ x236 ^ x60 ;
  assign n635 = n634 ^ n633 ^ n601 ;
  assign n636 = ( ~x30 & x145 ) | ( ~x30 & n319 ) | ( x145 & n319 ) ;
  assign n637 = n636 ^ x191 ^ x163 ;
  assign n638 = n331 & ~n637 ;
  assign n639 = n638 ^ n286 ^ 1'b0 ;
  assign n640 = ( x180 & n635 ) | ( x180 & n639 ) | ( n635 & n639 ) ;
  assign n641 = ( x72 & ~x176 ) | ( x72 & n640 ) | ( ~x176 & n640 ) ;
  assign n643 = ( ~x123 & n281 ) | ( ~x123 & n370 ) | ( n281 & n370 ) ;
  assign n644 = n643 ^ n490 ^ x197 ;
  assign n642 = n364 ^ x49 ^ x0 ;
  assign n645 = n644 ^ n642 ^ 1'b0 ;
  assign n646 = x241 ^ x35 ^ x19 ;
  assign n647 = ( n279 & ~n532 ) | ( n279 & n646 ) | ( ~n532 & n646 ) ;
  assign n660 = x203 ^ x158 ^ x156 ;
  assign n661 = ( x1 & n273 ) | ( x1 & ~n660 ) | ( n273 & ~n660 ) ;
  assign n655 = x81 ^ x31 ^ x26 ;
  assign n656 = ( x205 & ~x227 ) | ( x205 & n279 ) | ( ~x227 & n279 ) ;
  assign n657 = ~n315 & n656 ;
  assign n658 = n655 & n657 ;
  assign n654 = ( x29 & x88 ) | ( x29 & ~x178 ) | ( x88 & ~x178 ) ;
  assign n652 = ( x68 & ~x141 ) | ( x68 & x153 ) | ( ~x141 & x153 ) ;
  assign n653 = ( n346 & n354 ) | ( n346 & ~n652 ) | ( n354 & ~n652 ) ;
  assign n659 = n658 ^ n654 ^ n653 ;
  assign n648 = ( n332 & n410 ) | ( n332 & n634 ) | ( n410 & n634 ) ;
  assign n649 = ( x209 & n334 ) | ( x209 & n648 ) | ( n334 & n648 ) ;
  assign n650 = n292 & n649 ;
  assign n651 = ~x3 & n650 ;
  assign n662 = n661 ^ n659 ^ n651 ;
  assign n663 = n662 ^ x239 ^ x90 ;
  assign n664 = x135 & n297 ;
  assign n665 = n664 ^ x192 ^ 1'b0 ;
  assign n666 = n665 ^ x173 ^ x165 ;
  assign n667 = n666 ^ x153 ^ x141 ;
  assign n668 = x121 ^ x55 ^ 1'b0 ;
  assign n669 = x127 & n668 ;
  assign n670 = ( x83 & n464 ) | ( x83 & ~n669 ) | ( n464 & ~n669 ) ;
  assign n671 = n333 ^ n304 ^ x70 ;
  assign n672 = ( ~x57 & x103 ) | ( ~x57 & n258 ) | ( x103 & n258 ) ;
  assign n673 = n672 ^ n265 ^ x153 ;
  assign n674 = x74 & n673 ;
  assign n675 = n674 ^ n316 ^ 1'b0 ;
  assign n676 = ( n277 & n671 ) | ( n277 & n675 ) | ( n671 & n675 ) ;
  assign n677 = x6 & x181 ;
  assign n678 = n677 ^ n308 ^ 1'b0 ;
  assign n684 = x47 & ~n561 ;
  assign n685 = n484 & n684 ;
  assign n686 = ( x248 & n387 ) | ( x248 & ~n685 ) | ( n387 & ~n685 ) ;
  assign n687 = n686 ^ n434 ^ x154 ;
  assign n681 = n339 ^ x249 ^ x168 ;
  assign n679 = n375 & ~n491 ;
  assign n680 = n679 ^ x108 ^ 1'b0 ;
  assign n682 = n681 ^ n680 ^ n293 ;
  assign n683 = x194 | n682 ;
  assign n688 = n687 ^ n683 ^ n477 ;
  assign n690 = ( ~x32 & x66 ) | ( ~x32 & x220 ) | ( x66 & x220 ) ;
  assign n689 = ~x86 & x234 ;
  assign n691 = n690 ^ n689 ^ n317 ;
  assign n692 = n691 ^ n269 ^ 1'b0 ;
  assign n693 = n581 ^ x39 ^ 1'b0 ;
  assign n694 = n330 ^ x246 ^ x115 ;
  assign n695 = n694 ^ n437 ^ x228 ;
  assign n696 = n568 ^ x88 ^ x41 ;
  assign n697 = ( x3 & n516 ) | ( x3 & ~n690 ) | ( n516 & ~n690 ) ;
  assign n699 = ( ~x40 & x106 ) | ( ~x40 & x250 ) | ( x106 & x250 ) ;
  assign n700 = ( ~x83 & n472 ) | ( ~x83 & n699 ) | ( n472 & n699 ) ;
  assign n698 = x123 & n424 ;
  assign n701 = n700 ^ n698 ^ x236 ;
  assign n702 = ( x249 & n697 ) | ( x249 & ~n701 ) | ( n697 & ~n701 ) ;
  assign n703 = ( n307 & n387 ) | ( n307 & n541 ) | ( n387 & n541 ) ;
  assign n707 = ~x85 & x178 ;
  assign n704 = x192 ^ x191 ^ x132 ;
  assign n705 = ( x68 & ~x166 ) | ( x68 & n704 ) | ( ~x166 & n704 ) ;
  assign n706 = n705 ^ n482 ^ x169 ;
  assign n708 = n707 ^ n706 ^ n361 ;
  assign n709 = ( n354 & ~n445 ) | ( n354 & n708 ) | ( ~n445 & n708 ) ;
  assign n710 = n443 | n492 ;
  assign n711 = ( n317 & n565 ) | ( n317 & n710 ) | ( n565 & n710 ) ;
  assign n712 = n711 ^ x174 ^ 1'b0 ;
  assign n713 = x220 & n712 ;
  assign n714 = ( x172 & n306 ) | ( x172 & n713 ) | ( n306 & n713 ) ;
  assign n715 = ( ~x150 & x253 ) | ( ~x150 & n501 ) | ( x253 & n501 ) ;
  assign n716 = n715 ^ x162 ^ 1'b0 ;
  assign n717 = ~n382 & n716 ;
  assign n718 = ~x8 & n717 ;
  assign n719 = ( x35 & ~n707 ) | ( x35 & n718 ) | ( ~n707 & n718 ) ;
  assign n720 = ( n317 & n417 ) | ( n317 & n671 ) | ( n417 & n671 ) ;
  assign n721 = n719 | n720 ;
  assign n722 = x128 ^ x4 ^ 1'b0 ;
  assign n729 = n275 ^ x185 ^ 1'b0 ;
  assign n723 = n656 ^ x251 ^ 1'b0 ;
  assign n724 = x7 & n723 ;
  assign n725 = ( ~x97 & x233 ) | ( ~x97 & n724 ) | ( x233 & n724 ) ;
  assign n726 = n304 ^ x224 ^ 1'b0 ;
  assign n727 = n725 & n726 ;
  assign n728 = ( ~x97 & n472 ) | ( ~x97 & n727 ) | ( n472 & n727 ) ;
  assign n730 = n729 ^ n728 ^ x202 ;
  assign n731 = x125 & n730 ;
  assign n732 = n722 & n731 ;
  assign n733 = n559 ^ n286 ^ x63 ;
  assign n734 = ( x224 & n262 ) | ( x224 & n733 ) | ( n262 & n733 ) ;
  assign n735 = x182 ^ x181 ^ x6 ;
  assign n736 = n735 ^ n411 ^ n353 ;
  assign n737 = ( ~x34 & x160 ) | ( ~x34 & n736 ) | ( x160 & n736 ) ;
  assign n738 = x221 & ~n737 ;
  assign n739 = n519 & n738 ;
  assign n740 = n729 ^ n633 ^ x145 ;
  assign n741 = n740 ^ n377 ^ 1'b0 ;
  assign n742 = ~n739 & n741 ;
  assign n743 = x118 & x187 ;
  assign n744 = n743 ^ n514 ^ x227 ;
  assign n745 = n744 ^ x57 ^ 1'b0 ;
  assign n756 = ( ~x100 & x156 ) | ( ~x100 & n544 ) | ( x156 & n544 ) ;
  assign n748 = x171 ^ x30 ^ x9 ;
  assign n749 = n748 ^ n652 ^ x166 ;
  assign n750 = x99 & x101 ;
  assign n751 = n750 ^ x88 ^ 1'b0 ;
  assign n752 = n751 ^ n293 ^ x137 ;
  assign n753 = ( n644 & n749 ) | ( n644 & n752 ) | ( n749 & n752 ) ;
  assign n746 = n310 ^ x49 ^ 1'b0 ;
  assign n747 = n746 ^ n479 ^ 1'b0 ;
  assign n754 = n753 ^ n747 ^ 1'b0 ;
  assign n755 = n464 & n754 ;
  assign n757 = n756 ^ n755 ^ x175 ;
  assign n759 = x227 & ~n519 ;
  assign n760 = ~x242 & n759 ;
  assign n758 = x66 & n293 ;
  assign n761 = n760 ^ n758 ^ 1'b0 ;
  assign n762 = n525 ^ x212 ^ 1'b0 ;
  assign n763 = n561 | n762 ;
  assign n764 = ( ~x118 & n761 ) | ( ~x118 & n763 ) | ( n761 & n763 ) ;
  assign n765 = x175 & n331 ;
  assign n766 = ~x127 & n765 ;
  assign n767 = n528 ^ n459 ^ n279 ;
  assign n768 = ( n643 & ~n766 ) | ( n643 & n767 ) | ( ~n766 & n767 ) ;
  assign n769 = ( x35 & n280 ) | ( x35 & ~n585 ) | ( n280 & ~n585 ) ;
  assign n770 = n769 ^ n287 ^ x166 ;
  assign n771 = ( ~x25 & x127 ) | ( ~x25 & n770 ) | ( x127 & n770 ) ;
  assign n772 = ( x186 & ~n768 ) | ( x186 & n771 ) | ( ~n768 & n771 ) ;
  assign n773 = n464 & n772 ;
  assign n774 = n553 ^ n267 ^ x178 ;
  assign n775 = n506 | n546 ;
  assign n776 = ( ~n323 & n446 ) | ( ~n323 & n581 ) | ( n446 & n581 ) ;
  assign n777 = ( x225 & ~n265 ) | ( x225 & n720 ) | ( ~n265 & n720 ) ;
  assign n778 = n777 ^ n292 ^ x142 ;
  assign n779 = ( n775 & n776 ) | ( n775 & ~n778 ) | ( n776 & ~n778 ) ;
  assign n780 = x140 & x244 ;
  assign n781 = n780 ^ n747 ^ 1'b0 ;
  assign n784 = n504 ^ n442 ^ n409 ;
  assign n782 = ( x28 & n511 ) | ( x28 & ~n528 ) | ( n511 & ~n528 ) ;
  assign n783 = ( x136 & n533 ) | ( x136 & n782 ) | ( n533 & n782 ) ;
  assign n785 = n784 ^ n783 ^ n282 ;
  assign n786 = n659 ^ n402 ^ 1'b0 ;
  assign n787 = x29 & n786 ;
  assign n788 = n714 ^ n424 ^ x114 ;
  assign n789 = ( x13 & n787 ) | ( x13 & n788 ) | ( n787 & n788 ) ;
  assign n797 = ( x146 & x181 ) | ( x146 & n347 ) | ( x181 & n347 ) ;
  assign n798 = ( x44 & ~x211 ) | ( x44 & n797 ) | ( ~x211 & n797 ) ;
  assign n793 = n281 ^ x150 ^ x49 ;
  assign n794 = n793 ^ n270 ^ 1'b0 ;
  assign n795 = n619 ^ n544 ^ 1'b0 ;
  assign n796 = ( x80 & n794 ) | ( x80 & n795 ) | ( n794 & n795 ) ;
  assign n790 = ( ~x59 & x237 ) | ( ~x59 & n396 ) | ( x237 & n396 ) ;
  assign n791 = n568 | n790 ;
  assign n792 = n678 & ~n791 ;
  assign n799 = n798 ^ n796 ^ n792 ;
  assign n800 = ( x50 & n482 ) | ( x50 & n567 ) | ( n482 & n567 ) ;
  assign n801 = ~x56 & x187 ;
  assign n802 = x181 & ~n801 ;
  assign n803 = n802 ^ n343 ^ 1'b0 ;
  assign n804 = ( n282 & n440 ) | ( n282 & ~n803 ) | ( n440 & ~n803 ) ;
  assign n808 = n363 ^ x82 ^ 1'b0 ;
  assign n809 = n324 & n808 ;
  assign n810 = n809 ^ n607 ^ x174 ;
  assign n806 = x108 & n280 ;
  assign n805 = ( x121 & n279 ) | ( x121 & ~n437 ) | ( n279 & ~n437 ) ;
  assign n807 = n806 ^ n805 ^ n735 ;
  assign n811 = n810 ^ n807 ^ n453 ;
  assign n812 = n811 ^ n720 ^ x42 ;
  assign n813 = ( n392 & n804 ) | ( n392 & n812 ) | ( n804 & n812 ) ;
  assign n814 = ( n367 & n800 ) | ( n367 & ~n813 ) | ( n800 & ~n813 ) ;
  assign n818 = n451 ^ n279 ^ x121 ;
  assign n819 = n818 ^ n373 ^ 1'b0 ;
  assign n820 = x188 & n819 ;
  assign n821 = ( x15 & n267 ) | ( x15 & n490 ) | ( n267 & n490 ) ;
  assign n822 = n821 ^ x131 ^ x84 ;
  assign n823 = n822 ^ n416 ^ x31 ;
  assign n824 = ( x93 & x209 ) | ( x93 & n823 ) | ( x209 & n823 ) ;
  assign n825 = ~n604 & n824 ;
  assign n826 = ~n820 & n825 ;
  assign n815 = n748 ^ n697 ^ n315 ;
  assign n816 = n706 ^ n568 ^ 1'b0 ;
  assign n817 = n815 & n816 ;
  assign n827 = n826 ^ n817 ^ x177 ;
  assign n831 = ( ~n366 & n413 ) | ( ~n366 & n432 ) | ( n413 & n432 ) ;
  assign n832 = ( x156 & ~n357 ) | ( x156 & n831 ) | ( ~n357 & n831 ) ;
  assign n828 = ( x148 & ~x213 ) | ( x148 & n623 ) | ( ~x213 & n623 ) ;
  assign n829 = n828 ^ n514 ^ x106 ;
  assign n830 = n829 ^ n743 ^ n552 ;
  assign n833 = n832 ^ n830 ^ x144 ;
  assign n834 = n415 ^ x5 ^ 1'b0 ;
  assign n835 = n539 & n834 ;
  assign n836 = n835 ^ n420 ^ n399 ;
  assign n837 = x201 ^ x0 ^ 1'b0 ;
  assign n838 = ~n306 & n837 ;
  assign n839 = n838 ^ n465 ^ n443 ;
  assign n840 = ( x155 & x169 ) | ( x155 & n484 ) | ( x169 & n484 ) ;
  assign n841 = n714 ^ n665 ^ n342 ;
  assign n842 = ( n839 & n840 ) | ( n839 & n841 ) | ( n840 & n841 ) ;
  assign n843 = x80 & x224 ;
  assign n844 = ~x90 & n843 ;
  assign n847 = n818 ^ n412 ^ n380 ;
  assign n848 = n847 ^ n529 ^ n295 ;
  assign n845 = ( x43 & ~n465 ) | ( x43 & n541 ) | ( ~n465 & n541 ) ;
  assign n846 = ( ~x214 & n556 ) | ( ~x214 & n845 ) | ( n556 & n845 ) ;
  assign n849 = n848 ^ n846 ^ n295 ;
  assign n850 = n632 | n849 ;
  assign n851 = x202 & n402 ;
  assign n852 = n655 ^ n346 ^ n265 ;
  assign n853 = n852 ^ x3 ^ 1'b0 ;
  assign n854 = ( ~n645 & n851 ) | ( ~n645 & n853 ) | ( n851 & n853 ) ;
  assign n855 = ( n844 & n850 ) | ( n844 & n854 ) | ( n850 & n854 ) ;
  assign n856 = x140 ^ x131 ^ x31 ;
  assign n857 = n856 ^ x188 ^ x48 ;
  assign n858 = n857 ^ x127 ^ 1'b0 ;
  assign n859 = n354 ^ n292 ^ 1'b0 ;
  assign n860 = n859 ^ n782 ^ 1'b0 ;
  assign n861 = n634 ^ x112 ^ 1'b0 ;
  assign n862 = ( n623 & ~n860 ) | ( n623 & n861 ) | ( ~n860 & n861 ) ;
  assign n866 = ( x50 & x57 ) | ( x50 & ~x162 ) | ( x57 & ~x162 ) ;
  assign n865 = n281 & n832 ;
  assign n867 = n866 ^ n865 ^ 1'b0 ;
  assign n868 = n867 ^ n551 ^ x242 ;
  assign n864 = ( x58 & x137 ) | ( x58 & n646 ) | ( x137 & n646 ) ;
  assign n863 = ( x168 & ~n600 ) | ( x168 & n656 ) | ( ~n600 & n656 ) ;
  assign n869 = n868 ^ n864 ^ n863 ;
  assign n870 = n595 ^ n459 ^ n333 ;
  assign n871 = ( n512 & ~n686 ) | ( n512 & n870 ) | ( ~n686 & n870 ) ;
  assign n872 = n871 ^ n855 ^ n590 ;
  assign n883 = ( x111 & ~n405 ) | ( x111 & n719 ) | ( ~n405 & n719 ) ;
  assign n884 = ( ~x100 & x198 ) | ( ~x100 & x204 ) | ( x198 & x204 ) ;
  assign n885 = ( n399 & n407 ) | ( n399 & n884 ) | ( n407 & n884 ) ;
  assign n886 = n885 ^ n509 ^ 1'b0 ;
  assign n887 = n883 & n886 ;
  assign n873 = ( n484 & n548 ) | ( n484 & ~n571 ) | ( n548 & ~n571 ) ;
  assign n874 = n831 ^ x254 ^ x175 ;
  assign n875 = ( ~x181 & x193 ) | ( ~x181 & n874 ) | ( x193 & n874 ) ;
  assign n877 = n431 ^ x178 ^ 1'b0 ;
  assign n876 = n365 ^ x241 ^ x11 ;
  assign n878 = n877 ^ n876 ^ 1'b0 ;
  assign n879 = ~n377 & n878 ;
  assign n880 = ( n743 & n875 ) | ( n743 & ~n879 ) | ( n875 & ~n879 ) ;
  assign n881 = ( x51 & x94 ) | ( x51 & ~n880 ) | ( x94 & ~n880 ) ;
  assign n882 = ( n672 & ~n873 ) | ( n672 & n881 ) | ( ~n873 & n881 ) ;
  assign n888 = n887 ^ n882 ^ n651 ;
  assign n889 = ( x242 & n357 ) | ( x242 & n814 ) | ( n357 & n814 ) ;
  assign n890 = n396 ^ n345 ^ x158 ;
  assign n891 = n432 ^ n394 ^ x223 ;
  assign n892 = ( n739 & n797 ) | ( n739 & n891 ) | ( n797 & n891 ) ;
  assign n893 = ( n297 & n807 ) | ( n297 & ~n892 ) | ( n807 & ~n892 ) ;
  assign n894 = ( x131 & x180 ) | ( x131 & ~x235 ) | ( x180 & ~x235 ) ;
  assign n895 = n502 ^ n383 ^ n307 ;
  assign n896 = n531 | n895 ;
  assign n897 = x107 | n896 ;
  assign n898 = ( x6 & x19 ) | ( x6 & ~n394 ) | ( x19 & ~n394 ) ;
  assign n899 = n898 ^ n310 ^ x60 ;
  assign n900 = ( ~x11 & n856 ) | ( ~x11 & n899 ) | ( n856 & n899 ) ;
  assign n901 = ( n894 & ~n897 ) | ( n894 & n900 ) | ( ~n897 & n900 ) ;
  assign n902 = n893 & ~n901 ;
  assign n903 = ~n890 & n902 ;
  assign n904 = ( x138 & n368 ) | ( x138 & ~n414 ) | ( n368 & ~n414 ) ;
  assign n905 = ( x1 & x83 ) | ( x1 & ~n904 ) | ( x83 & ~n904 ) ;
  assign n906 = ( ~x38 & x108 ) | ( ~x38 & n265 ) | ( x108 & n265 ) ;
  assign n907 = ( x36 & ~x114 ) | ( x36 & n906 ) | ( ~x114 & n906 ) ;
  assign n908 = n905 & n907 ;
  assign n909 = n832 ^ n400 ^ 1'b0 ;
  assign n910 = n909 ^ n620 ^ n337 ;
  assign n911 = ( ~x132 & x173 ) | ( ~x132 & n402 ) | ( x173 & n402 ) ;
  assign n912 = n348 ^ x204 ^ x108 ;
  assign n913 = n506 | n912 ;
  assign n914 = n911 | n913 ;
  assign n915 = ( x132 & ~n375 ) | ( x132 & n914 ) | ( ~n375 & n914 ) ;
  assign n916 = n426 ^ x222 ^ x107 ;
  assign n917 = n916 ^ n492 ^ 1'b0 ;
  assign n918 = x7 & n917 ;
  assign n919 = n918 ^ x4 ^ 1'b0 ;
  assign n920 = x84 & n919 ;
  assign n921 = x215 & n330 ;
  assign n922 = n347 & n921 ;
  assign n923 = ( ~n296 & n388 ) | ( ~n296 & n922 ) | ( n388 & n922 ) ;
  assign n924 = ( n424 & n920 ) | ( n424 & n923 ) | ( n920 & n923 ) ;
  assign n930 = n394 & ~n847 ;
  assign n931 = ~n304 & n930 ;
  assign n925 = x18 & x212 ;
  assign n926 = n925 ^ n328 ^ 1'b0 ;
  assign n927 = x219 ^ x131 ^ x57 ;
  assign n928 = n927 ^ n656 ^ x205 ;
  assign n929 = ( n884 & n926 ) | ( n884 & ~n928 ) | ( n926 & ~n928 ) ;
  assign n932 = n931 ^ n929 ^ n659 ;
  assign n933 = x220 & n932 ;
  assign n934 = ( x100 & x254 ) | ( x100 & ~n907 ) | ( x254 & ~n907 ) ;
  assign n935 = n451 | n822 ;
  assign n936 = x59 | n935 ;
  assign n937 = ( ~x32 & n680 ) | ( ~x32 & n715 ) | ( n680 & n715 ) ;
  assign n939 = n672 ^ x195 ^ x2 ;
  assign n938 = ( ~x89 & x142 ) | ( ~x89 & n409 ) | ( x142 & n409 ) ;
  assign n940 = n939 ^ n938 ^ n639 ;
  assign n941 = ( x37 & ~n937 ) | ( x37 & n940 ) | ( ~n937 & n940 ) ;
  assign n942 = n936 & n941 ;
  assign n943 = n942 ^ x25 ^ 1'b0 ;
  assign n944 = ( ~x46 & x143 ) | ( ~x46 & n943 ) | ( x143 & n943 ) ;
  assign n947 = ( x70 & x155 ) | ( x70 & ~n514 ) | ( x155 & ~n514 ) ;
  assign n945 = x136 & x184 ;
  assign n946 = n945 ^ n373 ^ 1'b0 ;
  assign n948 = n947 ^ n946 ^ x53 ;
  assign n949 = n948 ^ n867 ^ n832 ;
  assign n950 = n949 ^ n718 ^ n446 ;
  assign n951 = x200 & n592 ;
  assign n952 = ( n369 & n950 ) | ( n369 & n951 ) | ( n950 & n951 ) ;
  assign n953 = n260 ^ x55 ^ 1'b0 ;
  assign n954 = n953 ^ n845 ^ n385 ;
  assign n955 = x117 & n356 ;
  assign n956 = n954 & n955 ;
  assign n960 = n832 ^ n394 ^ n363 ;
  assign n957 = ( ~x150 & x226 ) | ( ~x150 & n423 ) | ( x226 & n423 ) ;
  assign n958 = n957 ^ x219 ^ x64 ;
  assign n959 = n958 ^ n847 ^ x103 ;
  assign n961 = n960 ^ n959 ^ n339 ;
  assign n962 = ( ~n952 & n956 ) | ( ~n952 & n961 ) | ( n956 & n961 ) ;
  assign n964 = n673 ^ n318 ^ n263 ;
  assign n965 = n540 ^ x159 ^ x130 ;
  assign n966 = n315 & ~n965 ;
  assign n967 = n966 ^ n637 ^ 1'b0 ;
  assign n968 = ~n964 & n967 ;
  assign n963 = ( ~n707 & n743 ) | ( ~n707 & n790 ) | ( n743 & n790 ) ;
  assign n969 = n968 ^ n963 ^ n393 ;
  assign n970 = ( ~x6 & x28 ) | ( ~x6 & n568 ) | ( x28 & n568 ) ;
  assign n971 = n957 ^ n805 ^ n517 ;
  assign n972 = ( n374 & n970 ) | ( n374 & ~n971 ) | ( n970 & ~n971 ) ;
  assign n973 = ( x92 & n318 ) | ( x92 & n972 ) | ( n318 & n972 ) ;
  assign n974 = n287 ^ x155 ^ x82 ;
  assign n975 = n486 & n974 ;
  assign n976 = ( x139 & n370 ) | ( x139 & n975 ) | ( n370 & n975 ) ;
  assign n977 = n976 ^ n768 ^ n659 ;
  assign n980 = ( x31 & x87 ) | ( x31 & ~x235 ) | ( x87 & ~x235 ) ;
  assign n978 = x170 ^ x10 ^ 1'b0 ;
  assign n979 = n713 & n978 ;
  assign n981 = n980 ^ n979 ^ x88 ;
  assign n982 = ( ~n488 & n491 ) | ( ~n488 & n981 ) | ( n491 & n981 ) ;
  assign n988 = ( x43 & ~x148 ) | ( x43 & x203 ) | ( ~x148 & x203 ) ;
  assign n986 = ( x99 & n369 ) | ( x99 & ~n518 ) | ( n369 & ~n518 ) ;
  assign n984 = x251 & ~n655 ;
  assign n985 = n984 ^ n283 ^ 1'b0 ;
  assign n983 = ( x135 & ~x161 ) | ( x135 & n479 ) | ( ~x161 & n479 ) ;
  assign n987 = n986 ^ n985 ^ n983 ;
  assign n989 = n988 ^ n987 ^ n659 ;
  assign n990 = ( n888 & ~n982 ) | ( n888 & n989 ) | ( ~n982 & n989 ) ;
  assign n991 = n264 & n767 ;
  assign n992 = n991 ^ x197 ^ 1'b0 ;
  assign n993 = n992 ^ n821 ^ n651 ;
  assign n994 = n503 & n845 ;
  assign n995 = x37 | n585 ;
  assign n996 = ( x12 & ~n561 ) | ( x12 & n579 ) | ( ~n561 & n579 ) ;
  assign n997 = ( ~x43 & x113 ) | ( ~x43 & n996 ) | ( x113 & n996 ) ;
  assign n998 = n997 ^ x250 ^ x218 ;
  assign n999 = n998 ^ n502 ^ x246 ;
  assign n1000 = n453 & n535 ;
  assign n1001 = ~n918 & n1000 ;
  assign n1002 = ( n317 & n542 ) | ( n317 & ~n614 ) | ( n542 & ~n614 ) ;
  assign n1003 = n607 & ~n1002 ;
  assign n1004 = n1001 & n1003 ;
  assign n1005 = ( n995 & n999 ) | ( n995 & ~n1004 ) | ( n999 & ~n1004 ) ;
  assign n1006 = ( x189 & ~x236 ) | ( x189 & x238 ) | ( ~x236 & x238 ) ;
  assign n1007 = ( x123 & ~n273 ) | ( x123 & n278 ) | ( ~n273 & n278 ) ;
  assign n1008 = ( x23 & ~n1006 ) | ( x23 & n1007 ) | ( ~n1006 & n1007 ) ;
  assign n1009 = ( n531 & n646 ) | ( n531 & ~n790 ) | ( n646 & ~n790 ) ;
  assign n1010 = n400 & n590 ;
  assign n1011 = n929 | n1010 ;
  assign n1012 = n1009 & ~n1011 ;
  assign n1013 = ( n846 & n1008 ) | ( n846 & n1012 ) | ( n1008 & n1012 ) ;
  assign n1015 = n346 ^ x234 ^ x102 ;
  assign n1014 = x8 & ~n566 ;
  assign n1016 = n1015 ^ n1014 ^ 1'b0 ;
  assign n1017 = n1016 ^ n810 ^ 1'b0 ;
  assign n1018 = ( x51 & ~n682 ) | ( x51 & n1017 ) | ( ~n682 & n1017 ) ;
  assign n1020 = ( ~x102 & x116 ) | ( ~x102 & n818 ) | ( x116 & n818 ) ;
  assign n1019 = n414 ^ x216 ^ 1'b0 ;
  assign n1021 = n1020 ^ n1019 ^ n338 ;
  assign n1022 = ( n511 & ~n536 ) | ( n511 & n1021 ) | ( ~n536 & n1021 ) ;
  assign n1024 = ( n671 & ~n705 ) | ( n671 & n832 ) | ( ~n705 & n832 ) ;
  assign n1025 = n1024 ^ x61 ^ 1'b0 ;
  assign n1023 = x15 & ~n860 ;
  assign n1026 = n1025 ^ n1023 ^ x80 ;
  assign n1043 = ( x72 & x223 ) | ( x72 & n436 ) | ( x223 & n436 ) ;
  assign n1044 = ( n473 & n818 ) | ( n473 & ~n1043 ) | ( n818 & ~n1043 ) ;
  assign n1033 = ( n267 & n482 ) | ( n267 & ~n790 ) | ( n482 & ~n790 ) ;
  assign n1034 = x77 & ~n1033 ;
  assign n1035 = n694 | n1034 ;
  assign n1036 = n549 & ~n1035 ;
  assign n1037 = x206 & x220 ;
  assign n1038 = n1036 & n1037 ;
  assign n1039 = ( n392 & n760 ) | ( n392 & n1038 ) | ( n760 & n1038 ) ;
  assign n1040 = ( n521 & ~n940 ) | ( n521 & n1039 ) | ( ~n940 & n1039 ) ;
  assign n1030 = x239 ^ x187 ^ x148 ;
  assign n1028 = ( x81 & n352 ) | ( x81 & ~n411 ) | ( n352 & ~n411 ) ;
  assign n1029 = n1028 ^ n350 ^ x81 ;
  assign n1027 = ( x124 & x169 ) | ( x124 & ~n724 ) | ( x169 & ~n724 ) ;
  assign n1031 = n1030 ^ n1029 ^ n1027 ;
  assign n1032 = n1031 ^ n710 ^ n480 ;
  assign n1041 = n1040 ^ n1032 ^ x23 ;
  assign n1042 = n1041 ^ n472 ^ n399 ;
  assign n1045 = n1044 ^ n1042 ^ x41 ;
  assign n1046 = ( n423 & ~n545 ) | ( n423 & n557 ) | ( ~n545 & n557 ) ;
  assign n1047 = ( ~x249 & n313 ) | ( ~x249 & n1046 ) | ( n313 & n1046 ) ;
  assign n1048 = ( n730 & ~n915 ) | ( n730 & n1047 ) | ( ~n915 & n1047 ) ;
  assign n1049 = ( x72 & ~x242 ) | ( x72 & n662 ) | ( ~x242 & n662 ) ;
  assign n1050 = n334 ^ x152 ^ 1'b0 ;
  assign n1051 = n789 ^ x152 ^ 1'b0 ;
  assign n1052 = ~n1040 & n1051 ;
  assign n1053 = n502 ^ n480 ^ n423 ;
  assign n1054 = n749 & n1053 ;
  assign n1055 = n1054 ^ n649 ^ 1'b0 ;
  assign n1056 = n526 ^ x89 ^ 1'b0 ;
  assign n1057 = ( ~x201 & n557 ) | ( ~x201 & n950 ) | ( n557 & n950 ) ;
  assign n1058 = n1056 & ~n1057 ;
  assign n1059 = ( n463 & ~n697 ) | ( n463 & n821 ) | ( ~n697 & n821 ) ;
  assign n1060 = n1059 ^ n640 ^ n378 ;
  assign n1061 = ( n1055 & n1058 ) | ( n1055 & ~n1060 ) | ( n1058 & ~n1060 ) ;
  assign n1062 = ( n829 & ~n986 ) | ( n829 & n1061 ) | ( ~n986 & n1061 ) ;
  assign n1063 = ~n388 & n695 ;
  assign n1064 = n259 ^ x67 ^ x9 ;
  assign n1065 = ( x62 & ~x72 ) | ( x62 & x176 ) | ( ~x72 & x176 ) ;
  assign n1066 = n1065 ^ n678 ^ n617 ;
  assign n1067 = ( x33 & n1064 ) | ( x33 & n1066 ) | ( n1064 & n1066 ) ;
  assign n1070 = n445 ^ n277 ^ 1'b0 ;
  assign n1071 = n318 | n1070 ;
  assign n1069 = n564 ^ x242 ^ x89 ;
  assign n1068 = ( x196 & ~n442 ) | ( x196 & n979 ) | ( ~n442 & n979 ) ;
  assign n1072 = n1071 ^ n1069 ^ n1068 ;
  assign n1073 = ( x18 & x218 ) | ( x18 & ~n533 ) | ( x218 & ~n533 ) ;
  assign n1074 = n1073 ^ n659 ^ x100 ;
  assign n1075 = ( ~n504 & n753 ) | ( ~n504 & n1074 ) | ( n753 & n1074 ) ;
  assign n1076 = x252 & n297 ;
  assign n1077 = n455 & n1076 ;
  assign n1078 = n1077 ^ x29 ^ 1'b0 ;
  assign n1079 = n1009 ^ x132 ^ x127 ;
  assign n1080 = n1079 ^ n961 ^ n350 ;
  assign n1081 = n849 ^ n463 ^ 1'b0 ;
  assign n1082 = n957 ^ n920 ^ n321 ;
  assign n1083 = ( x189 & ~x215 ) | ( x189 & n838 ) | ( ~x215 & n838 ) ;
  assign n1084 = ( x74 & n1082 ) | ( x74 & n1083 ) | ( n1082 & n1083 ) ;
  assign n1092 = x57 & ~n1025 ;
  assign n1085 = n308 & ~n388 ;
  assign n1086 = x114 & ~n658 ;
  assign n1087 = n1086 ^ n346 ^ 1'b0 ;
  assign n1088 = ( n408 & n715 ) | ( n408 & ~n1087 ) | ( n715 & ~n1087 ) ;
  assign n1089 = ~n621 & n1088 ;
  assign n1090 = ~x179 & n1089 ;
  assign n1091 = ( n521 & ~n1085 ) | ( n521 & n1090 ) | ( ~n1085 & n1090 ) ;
  assign n1093 = n1092 ^ n1091 ^ 1'b0 ;
  assign n1094 = n468 ^ n288 ^ x176 ;
  assign n1095 = ( n414 & n531 ) | ( n414 & n918 ) | ( n531 & n918 ) ;
  assign n1096 = n600 & n1095 ;
  assign n1097 = n1094 & n1096 ;
  assign n1098 = ( n776 & n875 ) | ( n776 & n1097 ) | ( n875 & n1097 ) ;
  assign n1099 = n1098 ^ x75 ^ 1'b0 ;
  assign n1105 = ( x59 & ~x117 ) | ( x59 & n307 ) | ( ~x117 & n307 ) ;
  assign n1104 = ( n405 & n653 ) | ( n405 & ~n1043 ) | ( n653 & ~n1043 ) ;
  assign n1102 = n531 ^ n505 ^ n406 ;
  assign n1101 = n455 ^ x232 ^ x215 ;
  assign n1103 = n1102 ^ n1101 ^ 1'b0 ;
  assign n1106 = n1105 ^ n1104 ^ n1103 ;
  assign n1100 = x252 & ~n745 ;
  assign n1107 = n1106 ^ n1100 ^ 1'b0 ;
  assign n1108 = n1107 ^ x126 ^ 1'b0 ;
  assign n1109 = n735 ^ x1 ^ 1'b0 ;
  assign n1110 = n262 & ~n1109 ;
  assign n1111 = n1110 ^ n634 ^ n262 ;
  assign n1115 = n297 & ~n315 ;
  assign n1116 = n1115 ^ x212 ^ 1'b0 ;
  assign n1112 = x226 & n361 ;
  assign n1113 = ( n287 & n522 ) | ( n287 & ~n1112 ) | ( n522 & ~n1112 ) ;
  assign n1114 = n1113 ^ n751 ^ n466 ;
  assign n1117 = n1116 ^ n1114 ^ n304 ;
  assign n1118 = n447 & n1117 ;
  assign n1119 = n1118 ^ n926 ^ 1'b0 ;
  assign n1120 = n1008 & ~n1119 ;
  assign n1121 = n383 ^ x1 ^ 1'b0 ;
  assign n1122 = n540 & ~n1121 ;
  assign n1123 = ( ~n572 & n870 ) | ( ~n572 & n1122 ) | ( n870 & n1122 ) ;
  assign n1124 = x214 ^ x48 ^ 1'b0 ;
  assign n1125 = n1123 & n1124 ;
  assign n1126 = ( n718 & ~n908 ) | ( n718 & n1125 ) | ( ~n908 & n1125 ) ;
  assign n1127 = n296 ^ x76 ^ x61 ;
  assign n1128 = n1127 ^ n287 ^ x166 ;
  assign n1129 = ( ~x18 & x195 ) | ( ~x18 & n341 ) | ( x195 & n341 ) ;
  assign n1130 = ( ~x72 & n359 ) | ( ~x72 & n1129 ) | ( n359 & n1129 ) ;
  assign n1131 = n1130 ^ x222 ^ x181 ;
  assign n1132 = ( n769 & n1128 ) | ( n769 & ~n1131 ) | ( n1128 & ~n1131 ) ;
  assign n1133 = ( ~n399 & n1126 ) | ( ~n399 & n1132 ) | ( n1126 & n1132 ) ;
  assign n1134 = n333 & ~n1016 ;
  assign n1135 = n1134 ^ n540 ^ n369 ;
  assign n1141 = n634 ^ n457 ^ 1'b0 ;
  assign n1139 = n771 ^ x96 ^ 1'b0 ;
  assign n1140 = n1139 ^ x185 ^ x181 ;
  assign n1136 = ( n728 & ~n875 ) | ( n728 & n1094 ) | ( ~n875 & n1094 ) ;
  assign n1137 = ( x72 & ~n641 ) | ( x72 & n1136 ) | ( ~n641 & n1136 ) ;
  assign n1138 = n1137 ^ n343 ^ x12 ;
  assign n1142 = n1141 ^ n1140 ^ n1138 ;
  assign n1143 = n1142 ^ n283 ^ x43 ;
  assign n1144 = ( x86 & n502 ) | ( x86 & ~n585 ) | ( n502 & ~n585 ) ;
  assign n1145 = n277 ^ x117 ^ x102 ;
  assign n1146 = ( x59 & ~x120 ) | ( x59 & n374 ) | ( ~x120 & n374 ) ;
  assign n1147 = ( n1144 & n1145 ) | ( n1144 & ~n1146 ) | ( n1145 & ~n1146 ) ;
  assign n1148 = n1147 ^ n1084 ^ n815 ;
  assign n1149 = n916 ^ n498 ^ n337 ;
  assign n1150 = ( x151 & x247 ) | ( x151 & ~n1149 ) | ( x247 & ~n1149 ) ;
  assign n1151 = n1150 ^ n592 ^ 1'b0 ;
  assign n1152 = x185 & ~n1151 ;
  assign n1153 = x82 & n544 ;
  assign n1154 = x12 & ~n1153 ;
  assign n1155 = n1154 ^ n1127 ^ 1'b0 ;
  assign n1157 = n427 ^ n267 ^ x242 ;
  assign n1156 = n998 ^ n607 ^ x90 ;
  assign n1158 = n1157 ^ n1156 ^ 1'b0 ;
  assign n1159 = n1155 & ~n1158 ;
  assign n1160 = ( n389 & n1084 ) | ( n389 & n1159 ) | ( n1084 & n1159 ) ;
  assign n1161 = ( ~x140 & x232 ) | ( ~x140 & n313 ) | ( x232 & n313 ) ;
  assign n1163 = n333 ^ x180 ^ 1'b0 ;
  assign n1162 = x128 & ~n363 ;
  assign n1164 = n1163 ^ n1162 ^ n637 ;
  assign n1165 = ( x144 & ~n1161 ) | ( x144 & n1164 ) | ( ~n1161 & n1164 ) ;
  assign n1166 = n1113 ^ n748 ^ x21 ;
  assign n1167 = n1166 ^ n685 ^ 1'b0 ;
  assign n1168 = n508 & n1167 ;
  assign n1169 = ( ~x87 & n1015 ) | ( ~x87 & n1168 ) | ( n1015 & n1168 ) ;
  assign n1170 = n1169 ^ n1161 ^ n1006 ;
  assign n1171 = n801 ^ x126 ^ 1'b0 ;
  assign n1172 = n1170 & ~n1171 ;
  assign n1175 = ( ~x58 & x122 ) | ( ~x58 & n596 ) | ( x122 & n596 ) ;
  assign n1173 = ( ~x34 & n558 ) | ( ~x34 & n874 ) | ( n558 & n874 ) ;
  assign n1174 = ( ~n265 & n761 ) | ( ~n265 & n1173 ) | ( n761 & n1173 ) ;
  assign n1176 = n1175 ^ n1174 ^ 1'b0 ;
  assign n1177 = n1172 & n1176 ;
  assign n1178 = n1177 ^ n305 ^ 1'b0 ;
  assign n1179 = ( x55 & x205 ) | ( x55 & n1178 ) | ( x205 & n1178 ) ;
  assign n1180 = n328 ^ x190 ^ x64 ;
  assign n1181 = ( x57 & x58 ) | ( x57 & ~x112 ) | ( x58 & ~x112 ) ;
  assign n1182 = n1181 ^ n316 ^ x191 ;
  assign n1183 = ( x142 & x199 ) | ( x142 & ~n1182 ) | ( x199 & ~n1182 ) ;
  assign n1184 = ( x51 & n1180 ) | ( x51 & ~n1183 ) | ( n1180 & ~n1183 ) ;
  assign n1185 = ( ~n522 & n857 ) | ( ~n522 & n1184 ) | ( n857 & n1184 ) ;
  assign n1186 = n1185 ^ n417 ^ n390 ;
  assign n1187 = n1186 ^ n692 ^ 1'b0 ;
  assign n1188 = x49 & n733 ;
  assign n1189 = x169 & ~n409 ;
  assign n1190 = ( n400 & ~n947 ) | ( n400 & n1046 ) | ( ~n947 & n1046 ) ;
  assign n1197 = ( n561 & ~n881 ) | ( n561 & n1182 ) | ( ~n881 & n1182 ) ;
  assign n1192 = x137 & n465 ;
  assign n1193 = ~x123 & n1192 ;
  assign n1194 = n1193 ^ x114 ^ x3 ;
  assign n1195 = n1194 ^ n728 ^ x44 ;
  assign n1191 = n1144 ^ n578 ^ x116 ;
  assign n1196 = n1195 ^ n1191 ^ n1088 ;
  assign n1198 = n1197 ^ n1196 ^ n621 ;
  assign n1199 = n997 ^ x21 ^ 1'b0 ;
  assign n1200 = n1199 ^ n380 ^ 1'b0 ;
  assign n1201 = x77 & ~n502 ;
  assign n1202 = n1201 ^ n1147 ^ 1'b0 ;
  assign n1203 = n1202 ^ n760 ^ x8 ;
  assign n1205 = n673 ^ n283 ^ x247 ;
  assign n1206 = n1205 ^ n867 ^ 1'b0 ;
  assign n1207 = n880 & n1206 ;
  assign n1204 = n1116 ^ n337 ^ x160 ;
  assign n1208 = n1207 ^ n1204 ^ x11 ;
  assign n1210 = ~n288 & n394 ;
  assign n1211 = ~n369 & n1210 ;
  assign n1212 = ( n879 & n940 ) | ( n879 & n1211 ) | ( n940 & n1211 ) ;
  assign n1209 = x59 & ~n992 ;
  assign n1213 = n1212 ^ n1209 ^ 1'b0 ;
  assign n1214 = ~n423 & n699 ;
  assign n1215 = n1214 ^ n567 ^ 1'b0 ;
  assign n1216 = n1215 ^ n1165 ^ n756 ;
  assign n1219 = n366 ^ x92 ^ x61 ;
  assign n1220 = n1219 ^ x254 ^ x180 ;
  assign n1217 = ( x208 & x218 ) | ( x208 & n998 ) | ( x218 & n998 ) ;
  assign n1218 = n1217 ^ n496 ^ n495 ;
  assign n1221 = n1220 ^ n1218 ^ n576 ;
  assign n1224 = n798 ^ n394 ^ x210 ;
  assign n1222 = ~n516 & n1155 ;
  assign n1223 = n1222 ^ n1205 ^ 1'b0 ;
  assign n1225 = n1224 ^ n1223 ^ n879 ;
  assign n1226 = ( n557 & n635 ) | ( n557 & n1225 ) | ( n635 & n1225 ) ;
  assign n1227 = n436 ^ x169 ^ x161 ;
  assign n1228 = n953 ^ n551 ^ n271 ;
  assign n1229 = ~n1227 & n1228 ;
  assign n1230 = n739 ^ x55 ^ 1'b0 ;
  assign n1231 = x122 & ~n1230 ;
  assign n1232 = n276 ^ x39 ^ 1'b0 ;
  assign n1233 = ~n502 & n1232 ;
  assign n1240 = n660 ^ n288 ^ x0 ;
  assign n1237 = x149 & n476 ;
  assign n1238 = n1237 ^ x61 ^ 1'b0 ;
  assign n1239 = x88 & ~n1238 ;
  assign n1241 = n1240 ^ n1239 ^ 1'b0 ;
  assign n1234 = n809 ^ x63 ^ 1'b0 ;
  assign n1235 = ~n680 & n1234 ;
  assign n1236 = n1235 ^ n685 ^ x0 ;
  assign n1242 = n1241 ^ n1236 ^ n698 ;
  assign n1243 = n1233 & ~n1242 ;
  assign n1244 = n1243 ^ x203 ^ 1'b0 ;
  assign n1245 = n304 & n1244 ;
  assign n1246 = ( n382 & n1231 ) | ( n382 & n1245 ) | ( n1231 & n1245 ) ;
  assign n1247 = n1246 ^ n529 ^ 1'b0 ;
  assign n1248 = n1229 | n1247 ;
  assign n1251 = x237 & n457 ;
  assign n1252 = n1251 ^ n426 ^ 1'b0 ;
  assign n1253 = n1252 ^ x226 ^ x45 ;
  assign n1249 = ( x50 & n416 ) | ( x50 & ~n736 ) | ( n416 & ~n736 ) ;
  assign n1250 = ( x101 & ~n1144 ) | ( x101 & n1249 ) | ( ~n1144 & n1249 ) ;
  assign n1254 = n1253 ^ n1250 ^ n1199 ;
  assign n1255 = ( ~x1 & x115 ) | ( ~x1 & n709 ) | ( x115 & n709 ) ;
  assign n1256 = x156 & n1255 ;
  assign n1260 = n544 | n644 ;
  assign n1261 = x19 | n1260 ;
  assign n1257 = ( ~n342 & n536 ) | ( ~n342 & n998 ) | ( n536 & n998 ) ;
  assign n1258 = n1257 ^ n522 ^ x253 ;
  assign n1259 = n1258 ^ n937 ^ n319 ;
  assign n1262 = n1261 ^ n1259 ^ n395 ;
  assign n1270 = n365 ^ x137 ^ 1'b0 ;
  assign n1267 = n390 | n800 ;
  assign n1268 = x142 | n1267 ;
  assign n1269 = n1268 ^ n613 ^ x230 ;
  assign n1271 = n1270 ^ n1269 ^ n324 ;
  assign n1263 = n1224 ^ n600 ^ x51 ;
  assign n1264 = ( ~n725 & n799 ) | ( ~n725 & n1263 ) | ( n799 & n1263 ) ;
  assign n1265 = n827 & n1264 ;
  assign n1266 = ~n1133 & n1265 ;
  assign n1272 = n1271 ^ n1266 ^ n818 ;
  assign n1277 = n1102 ^ n315 ^ 1'b0 ;
  assign n1278 = ~n578 & n1277 ;
  assign n1279 = n1278 ^ x242 ^ x114 ;
  assign n1284 = n491 ^ x191 ^ x95 ;
  assign n1283 = ( x28 & ~x197 ) | ( x28 & n423 ) | ( ~x197 & n423 ) ;
  assign n1280 = n276 ^ x89 ^ x47 ;
  assign n1281 = ( ~x21 & x56 ) | ( ~x21 & n626 ) | ( x56 & n626 ) ;
  assign n1282 = ( ~x96 & n1280 ) | ( ~x96 & n1281 ) | ( n1280 & n1281 ) ;
  assign n1285 = n1284 ^ n1283 ^ n1282 ;
  assign n1286 = n1279 | n1285 ;
  assign n1287 = n807 | n1286 ;
  assign n1288 = n1287 ^ x71 ^ 1'b0 ;
  assign n1273 = n267 & ~n667 ;
  assign n1274 = n1273 ^ n437 ^ 1'b0 ;
  assign n1275 = n1274 ^ n1180 ^ n656 ;
  assign n1276 = ( n407 & ~n1162 ) | ( n407 & n1275 ) | ( ~n1162 & n1275 ) ;
  assign n1289 = n1288 ^ n1276 ^ n1145 ;
  assign n1290 = ( ~x37 & x199 ) | ( ~x37 & n457 ) | ( x199 & n457 ) ;
  assign n1291 = ( n1169 & n1226 ) | ( n1169 & n1290 ) | ( n1226 & n1290 ) ;
  assign n1292 = n1291 ^ n798 ^ n533 ;
  assign n1293 = n1292 ^ n1092 ^ n518 ;
  assign n1298 = ( x64 & x70 ) | ( x64 & ~n304 ) | ( x70 & ~n304 ) ;
  assign n1296 = ( ~x226 & n391 ) | ( ~x226 & n735 ) | ( n391 & n735 ) ;
  assign n1297 = n1296 ^ n914 ^ n675 ;
  assign n1299 = n1298 ^ n1297 ^ x109 ;
  assign n1294 = n1098 ^ n324 ^ x145 ;
  assign n1295 = n1294 ^ n857 ^ 1'b0 ;
  assign n1300 = n1299 ^ n1295 ^ 1'b0 ;
  assign n1301 = n624 | n1300 ;
  assign n1302 = n1301 ^ n861 ^ x49 ;
  assign n1303 = n451 ^ n286 ^ x109 ;
  assign n1304 = ( ~n880 & n1022 ) | ( ~n880 & n1303 ) | ( n1022 & n1303 ) ;
  assign n1305 = ( x87 & x181 ) | ( x87 & ~n320 ) | ( x181 & ~n320 ) ;
  assign n1306 = n1305 ^ n401 ^ x29 ;
  assign n1307 = ( ~x143 & n384 ) | ( ~x143 & n1306 ) | ( n384 & n1306 ) ;
  assign n1308 = ( ~n330 & n714 ) | ( ~n330 & n1172 ) | ( n714 & n1172 ) ;
  assign n1312 = n287 ^ x201 ^ x111 ;
  assign n1313 = n1312 ^ n724 ^ x11 ;
  assign n1309 = x232 & ~n801 ;
  assign n1310 = ~x218 & n1309 ;
  assign n1311 = n327 & ~n1310 ;
  assign n1314 = n1313 ^ n1311 ^ 1'b0 ;
  assign n1315 = n440 ^ n379 ^ x116 ;
  assign n1316 = ~n1314 & n1315 ;
  assign n1317 = n1316 ^ n1091 ^ n422 ;
  assign n1318 = n500 | n923 ;
  assign n1331 = x183 ^ x147 ^ x142 ;
  assign n1329 = ( x81 & x127 ) | ( x81 & ~n509 ) | ( x127 & ~n509 ) ;
  assign n1330 = n287 & n1329 ;
  assign n1332 = n1331 ^ n1330 ^ 1'b0 ;
  assign n1333 = ( n410 & ~n426 ) | ( n410 & n1149 ) | ( ~n426 & n1149 ) ;
  assign n1334 = ( n823 & n1332 ) | ( n823 & ~n1333 ) | ( n1332 & ~n1333 ) ;
  assign n1324 = ( x173 & n710 ) | ( x173 & ~n1236 ) | ( n710 & ~n1236 ) ;
  assign n1325 = ~n926 & n1324 ;
  assign n1326 = n1325 ^ n768 ^ n319 ;
  assign n1327 = ~x152 & n1263 ;
  assign n1328 = ~n1326 & n1327 ;
  assign n1319 = ( x4 & ~x246 ) | ( x4 & n422 ) | ( ~x246 & n422 ) ;
  assign n1320 = x145 & ~n1157 ;
  assign n1321 = n562 & ~n1320 ;
  assign n1322 = ( ~x220 & n1319 ) | ( ~x220 & n1321 ) | ( n1319 & n1321 ) ;
  assign n1323 = n1322 ^ n342 ^ x111 ;
  assign n1335 = n1334 ^ n1328 ^ n1323 ;
  assign n1336 = n1117 ^ n922 ^ n743 ;
  assign n1339 = n340 ^ x62 ^ x61 ;
  assign n1337 = n505 ^ x209 ^ x72 ;
  assign n1338 = ( x29 & x181 ) | ( x29 & n1337 ) | ( x181 & n1337 ) ;
  assign n1340 = n1339 ^ n1338 ^ x2 ;
  assign n1341 = x227 & ~n1340 ;
  assign n1342 = n1336 & n1341 ;
  assign n1343 = ( x225 & n278 ) | ( x225 & ~n951 ) | ( n278 & ~n951 ) ;
  assign n1344 = n1343 ^ n1074 ^ n947 ;
  assign n1345 = n440 & ~n1344 ;
  assign n1346 = ( x149 & n1342 ) | ( x149 & ~n1345 ) | ( n1342 & ~n1345 ) ;
  assign n1347 = ( x13 & n557 ) | ( x13 & n849 ) | ( n557 & n849 ) ;
  assign n1348 = n1078 ^ x20 ^ 1'b0 ;
  assign n1349 = n1347 & ~n1348 ;
  assign n1350 = ~n964 & n1202 ;
  assign n1351 = n1350 ^ n1228 ^ 1'b0 ;
  assign n1352 = n596 ^ n502 ^ n279 ;
  assign n1353 = n1352 ^ n1126 ^ 1'b0 ;
  assign n1354 = x200 & n364 ;
  assign n1355 = n1354 ^ n390 ^ 1'b0 ;
  assign n1356 = n1355 ^ n568 ^ x119 ;
  assign n1357 = n1356 ^ n806 ^ n760 ;
  assign n1358 = x152 & n838 ;
  assign n1359 = n960 & n1358 ;
  assign n1360 = n1359 ^ n822 ^ n710 ;
  assign n1361 = n1360 ^ n730 ^ x177 ;
  assign n1362 = ( n1353 & n1357 ) | ( n1353 & n1361 ) | ( n1357 & n1361 ) ;
  assign n1363 = n399 ^ x231 ^ x13 ;
  assign n1364 = ( ~x228 & n1357 ) | ( ~x228 & n1363 ) | ( n1357 & n1363 ) ;
  assign n1390 = ( x32 & ~n286 ) | ( x32 & n471 ) | ( ~n286 & n471 ) ;
  assign n1391 = n1390 ^ x88 ^ x70 ;
  assign n1392 = n1391 ^ n760 ^ n457 ;
  assign n1393 = ( x191 & ~n904 ) | ( x191 & n1392 ) | ( ~n904 & n1392 ) ;
  assign n1382 = ( ~x166 & x253 ) | ( ~x166 & n1130 ) | ( x253 & n1130 ) ;
  assign n1383 = n1382 ^ n974 ^ n580 ;
  assign n1384 = ( x233 & n790 ) | ( x233 & ~n852 ) | ( n790 & ~n852 ) ;
  assign n1385 = ( ~n308 & n518 ) | ( ~n308 & n1384 ) | ( n518 & n1384 ) ;
  assign n1386 = ( n815 & ~n1383 ) | ( n815 & n1385 ) | ( ~n1383 & n1385 ) ;
  assign n1370 = n552 ^ n339 ^ x252 ;
  assign n1371 = ( x91 & ~x198 ) | ( x91 & n958 ) | ( ~x198 & n958 ) ;
  assign n1372 = n1371 ^ n384 ^ x31 ;
  assign n1373 = ( x44 & n698 ) | ( x44 & n1372 ) | ( n698 & n1372 ) ;
  assign n1374 = n1373 ^ n968 ^ n583 ;
  assign n1375 = x56 & x164 ;
  assign n1376 = n1375 ^ x110 ^ 1'b0 ;
  assign n1377 = ( n511 & n659 ) | ( n511 & ~n1376 ) | ( n659 & ~n1376 ) ;
  assign n1378 = ( x21 & x75 ) | ( x21 & ~x223 ) | ( x75 & ~x223 ) ;
  assign n1379 = n1378 ^ n1313 ^ x218 ;
  assign n1380 = ( n1218 & n1377 ) | ( n1218 & n1379 ) | ( n1377 & n1379 ) ;
  assign n1381 = ( n1370 & n1374 ) | ( n1370 & ~n1380 ) | ( n1374 & ~n1380 ) ;
  assign n1365 = ( x45 & x168 ) | ( x45 & ~n539 ) | ( x168 & ~n539 ) ;
  assign n1366 = n1365 ^ n367 ^ x251 ;
  assign n1367 = n320 ^ x224 ^ x139 ;
  assign n1368 = n1220 & ~n1367 ;
  assign n1369 = ~n1366 & n1368 ;
  assign n1387 = n1386 ^ n1381 ^ n1369 ;
  assign n1388 = x61 & x114 ;
  assign n1389 = ~n1387 & n1388 ;
  assign n1394 = n1393 ^ n1389 ^ 1'b0 ;
  assign n1395 = n533 ^ n530 ^ 1'b0 ;
  assign n1421 = n265 ^ x190 ^ 1'b0 ;
  assign n1422 = n558 & n1421 ;
  assign n1399 = ( x12 & ~n923 ) | ( x12 & n946 ) | ( ~n923 & n946 ) ;
  assign n1401 = n637 ^ n342 ^ 1'b0 ;
  assign n1402 = ~n260 & n1401 ;
  assign n1403 = n1402 ^ n1163 ^ 1'b0 ;
  assign n1404 = n339 & n1403 ;
  assign n1400 = ~n643 & n1033 ;
  assign n1405 = n1404 ^ n1400 ^ 1'b0 ;
  assign n1406 = ( n393 & ~n1399 ) | ( n393 & n1405 ) | ( ~n1399 & n1405 ) ;
  assign n1398 = x53 | n275 ;
  assign n1407 = n1406 ^ n1398 ^ n633 ;
  assign n1397 = ( x254 & n315 ) | ( x254 & n608 ) | ( n315 & n608 ) ;
  assign n1408 = n1407 ^ n1397 ^ n1191 ;
  assign n1411 = ( ~x33 & n302 ) | ( ~x33 & n875 ) | ( n302 & n875 ) ;
  assign n1412 = n1411 ^ x7 ^ 1'b0 ;
  assign n1413 = x39 & n1412 ;
  assign n1414 = n1413 ^ x77 ^ 1'b0 ;
  assign n1409 = n1044 | n1283 ;
  assign n1410 = n830 & ~n1409 ;
  assign n1415 = n1414 ^ n1410 ^ 1'b0 ;
  assign n1416 = ~n377 & n1415 ;
  assign n1417 = n1416 ^ n589 ^ 1'b0 ;
  assign n1418 = n1149 & n1417 ;
  assign n1419 = ( ~n1056 & n1408 ) | ( ~n1056 & n1418 ) | ( n1408 & n1418 ) ;
  assign n1420 = n1419 ^ n1411 ^ 1'b0 ;
  assign n1423 = n1422 ^ n1420 ^ 1'b0 ;
  assign n1396 = x124 & ~n278 ;
  assign n1424 = n1423 ^ n1396 ^ 1'b0 ;
  assign n1425 = ( n399 & n517 ) | ( n399 & ~n1424 ) | ( n517 & ~n1424 ) ;
  assign n1426 = n1425 ^ n312 ^ 1'b0 ;
  assign n1427 = n1395 & n1426 ;
  assign n1438 = n653 ^ n578 ^ x160 ;
  assign n1437 = ( ~x34 & x198 ) | ( ~x34 & n339 ) | ( x198 & n339 ) ;
  assign n1432 = ( x66 & n528 ) | ( x66 & ~n552 ) | ( n528 & ~n552 ) ;
  assign n1433 = x195 & n730 ;
  assign n1434 = ~n1432 & n1433 ;
  assign n1428 = n1002 ^ x141 ^ x120 ;
  assign n1429 = n1105 ^ x187 ^ x186 ;
  assign n1430 = n1429 ^ x226 ^ x41 ;
  assign n1431 = ( x159 & ~n1428 ) | ( x159 & n1430 ) | ( ~n1428 & n1430 ) ;
  assign n1435 = n1434 ^ n1431 ^ x55 ;
  assign n1436 = ~n307 & n1435 ;
  assign n1439 = n1438 ^ n1437 ^ n1436 ;
  assign n1441 = x167 & ~n479 ;
  assign n1440 = ( ~x181 & n436 ) | ( ~x181 & n1233 ) | ( n436 & n1233 ) ;
  assign n1442 = n1441 ^ n1440 ^ n292 ;
  assign n1443 = ( n313 & n326 ) | ( n313 & ~n1442 ) | ( n326 & ~n1442 ) ;
  assign n1444 = ( n1305 & n1439 ) | ( n1305 & ~n1443 ) | ( n1439 & ~n1443 ) ;
  assign n1460 = ( ~n339 & n471 ) | ( ~n339 & n579 ) | ( n471 & n579 ) ;
  assign n1461 = n1460 ^ n844 ^ n440 ;
  assign n1462 = n1461 ^ n1339 ^ n1105 ;
  assign n1458 = n518 & ~n1180 ;
  assign n1459 = n1458 ^ n365 ^ 1'b0 ;
  assign n1463 = n1462 ^ n1459 ^ n718 ;
  assign n1464 = n1463 ^ n655 ^ n440 ;
  assign n1452 = n541 ^ n532 ^ 1'b0 ;
  assign n1453 = n307 & n1452 ;
  assign n1454 = ( n885 & ~n928 ) | ( n885 & n1370 ) | ( ~n928 & n1370 ) ;
  assign n1455 = n1454 ^ n369 ^ x149 ;
  assign n1456 = ( ~n313 & n1453 ) | ( ~n313 & n1455 ) | ( n1453 & n1455 ) ;
  assign n1445 = ( x187 & n364 ) | ( x187 & ~n379 ) | ( n364 & ~n379 ) ;
  assign n1446 = n1445 ^ n751 ^ x41 ;
  assign n1447 = n823 ^ n500 ^ n341 ;
  assign n1448 = ( ~n906 & n1184 ) | ( ~n906 & n1447 ) | ( n1184 & n1447 ) ;
  assign n1449 = x208 & ~n1448 ;
  assign n1450 = n411 & n1449 ;
  assign n1451 = n1446 & n1450 ;
  assign n1457 = n1456 ^ n1451 ^ n851 ;
  assign n1465 = n1464 ^ n1457 ^ n778 ;
  assign n1466 = ~n946 & n1465 ;
  assign n1467 = n1444 & n1466 ;
  assign n1468 = n326 & ~n689 ;
  assign n1469 = n569 & n1468 ;
  assign n1470 = ( n1268 & n1399 ) | ( n1268 & n1469 ) | ( n1399 & n1469 ) ;
  assign n1471 = ( ~x19 & x110 ) | ( ~x19 & x159 ) | ( x110 & x159 ) ;
  assign n1472 = x190 & n1083 ;
  assign n1473 = ~n1215 & n1472 ;
  assign n1474 = n346 & n1473 ;
  assign n1475 = ( ~n662 & n1471 ) | ( ~n662 & n1474 ) | ( n1471 & n1474 ) ;
  assign n1476 = n1356 ^ n1183 ^ n316 ;
  assign n1477 = n579 ^ n271 ^ x59 ;
  assign n1478 = ( n340 & n737 ) | ( n340 & n1477 ) | ( n737 & n1477 ) ;
  assign n1479 = n1478 ^ n555 ^ n311 ;
  assign n1480 = x80 & ~n1479 ;
  assign n1481 = n1480 ^ n396 ^ 1'b0 ;
  assign n1482 = n1476 & n1481 ;
  assign n1483 = n1183 ^ x121 ^ 1'b0 ;
  assign n1486 = ( n556 & n587 ) | ( n556 & ~n851 ) | ( n587 & ~n851 ) ;
  assign n1484 = ( x15 & x55 ) | ( x15 & ~n1207 ) | ( x55 & ~n1207 ) ;
  assign n1485 = ( n430 & ~n858 ) | ( n430 & n1484 ) | ( ~n858 & n1484 ) ;
  assign n1487 = n1486 ^ n1485 ^ x222 ;
  assign n1488 = ~n536 & n890 ;
  assign n1489 = n1488 ^ x164 ^ 1'b0 ;
  assign n1490 = n1489 ^ n742 ^ 1'b0 ;
  assign n1491 = n1487 & ~n1490 ;
  assign n1492 = ( n1066 & ~n1483 ) | ( n1066 & n1491 ) | ( ~n1483 & n1491 ) ;
  assign n1500 = ~n337 & n725 ;
  assign n1493 = ( x42 & n323 ) | ( x42 & ~n619 ) | ( n323 & ~n619 ) ;
  assign n1494 = ~n409 & n448 ;
  assign n1495 = n1494 ^ n737 ^ 1'b0 ;
  assign n1496 = ( x17 & ~x171 ) | ( x17 & n629 ) | ( ~x171 & n629 ) ;
  assign n1497 = ( x43 & n1071 ) | ( x43 & ~n1496 ) | ( n1071 & ~n1496 ) ;
  assign n1498 = n1495 & ~n1497 ;
  assign n1499 = ~n1493 & n1498 ;
  assign n1501 = n1500 ^ n1499 ^ 1'b0 ;
  assign n1502 = ( ~x159 & n356 ) | ( ~x159 & n1501 ) | ( n356 & n1501 ) ;
  assign n1503 = ( n396 & n415 ) | ( n396 & n1255 ) | ( n415 & n1255 ) ;
  assign n1510 = n466 ^ x61 ^ x32 ;
  assign n1511 = ( x59 & n1461 ) | ( x59 & n1510 ) | ( n1461 & n1510 ) ;
  assign n1512 = ( x230 & n571 ) | ( x230 & n1511 ) | ( n571 & n1511 ) ;
  assign n1513 = n671 ^ n654 ^ 1'b0 ;
  assign n1514 = n561 | n1513 ;
  assign n1515 = ( x167 & ~n706 ) | ( x167 & n1514 ) | ( ~n706 & n1514 ) ;
  assign n1516 = n1263 & n1515 ;
  assign n1517 = ~n487 & n1516 ;
  assign n1518 = ( n305 & n1512 ) | ( n305 & ~n1517 ) | ( n1512 & ~n1517 ) ;
  assign n1507 = x235 ^ x202 ^ x88 ;
  assign n1504 = ( n272 & n604 ) | ( n272 & n876 ) | ( n604 & n876 ) ;
  assign n1505 = ( ~n424 & n775 ) | ( ~n424 & n1504 ) | ( n775 & n1504 ) ;
  assign n1506 = n606 | n1505 ;
  assign n1508 = n1507 ^ n1506 ^ 1'b0 ;
  assign n1509 = ( n893 & ~n1255 ) | ( n893 & n1508 ) | ( ~n1255 & n1508 ) ;
  assign n1519 = n1518 ^ n1509 ^ n1274 ;
  assign n1522 = ( x74 & n368 ) | ( x74 & ~n431 ) | ( n368 & ~n431 ) ;
  assign n1523 = ( n660 & ~n912 ) | ( n660 & n1522 ) | ( ~n912 & n1522 ) ;
  assign n1532 = n707 ^ n359 ^ x103 ;
  assign n1533 = ( x150 & ~n898 ) | ( x150 & n1532 ) | ( ~n898 & n1532 ) ;
  assign n1530 = ( x88 & n265 ) | ( x88 & ~n477 ) | ( n265 & ~n477 ) ;
  assign n1524 = n362 & n607 ;
  assign n1525 = n1524 ^ n431 ^ 1'b0 ;
  assign n1526 = n1525 ^ x35 ^ 1'b0 ;
  assign n1527 = n377 | n1526 ;
  assign n1528 = ( n911 & n1162 ) | ( n911 & n1527 ) | ( n1162 & n1527 ) ;
  assign n1529 = ( n306 & n1113 ) | ( n306 & ~n1528 ) | ( n1113 & ~n1528 ) ;
  assign n1531 = n1530 ^ n1529 ^ n1097 ;
  assign n1534 = n1533 ^ n1531 ^ n1006 ;
  assign n1535 = ( n1012 & n1523 ) | ( n1012 & ~n1534 ) | ( n1523 & ~n1534 ) ;
  assign n1520 = ( n546 & n784 ) | ( n546 & ~n1306 ) | ( n784 & ~n1306 ) ;
  assign n1521 = x18 & ~n1520 ;
  assign n1536 = n1535 ^ n1521 ^ 1'b0 ;
  assign n1537 = n1312 ^ n793 ^ x199 ;
  assign n1538 = ( x69 & n733 ) | ( x69 & ~n1537 ) | ( n733 & ~n1537 ) ;
  assign n1539 = n1538 ^ n931 ^ x71 ;
  assign n1540 = n569 | n1153 ;
  assign n1541 = n1540 ^ x199 ^ 1'b0 ;
  assign n1542 = ~n604 & n695 ;
  assign n1543 = n1542 ^ n262 ^ 1'b0 ;
  assign n1544 = ( ~n856 & n1541 ) | ( ~n856 & n1543 ) | ( n1541 & n1543 ) ;
  assign n1545 = n1211 ^ n661 ^ n604 ;
  assign n1546 = n946 ^ n655 ^ x185 ;
  assign n1547 = n1546 ^ n295 ^ 1'b0 ;
  assign n1548 = n1547 ^ x210 ^ 1'b0 ;
  assign n1549 = n1545 | n1548 ;
  assign n1550 = ~n823 & n1242 ;
  assign n1551 = ( n1140 & ~n1143 ) | ( n1140 & n1550 ) | ( ~n1143 & n1550 ) ;
  assign n1563 = n1170 ^ n710 ^ 1'b0 ;
  assign n1564 = n559 & n1563 ;
  assign n1562 = n620 ^ n256 ^ x187 ;
  assign n1558 = ( ~x61 & x146 ) | ( ~x61 & n367 ) | ( x146 & n367 ) ;
  assign n1559 = n1558 ^ n694 ^ 1'b0 ;
  assign n1557 = ( ~x96 & n474 ) | ( ~x96 & n876 ) | ( n474 & n876 ) ;
  assign n1554 = ( x104 & n405 ) | ( x104 & n957 ) | ( n405 & n957 ) ;
  assign n1555 = n1554 ^ n906 ^ n672 ;
  assign n1553 = n1486 ^ n1016 ^ n588 ;
  assign n1556 = n1555 ^ n1553 ^ 1'b0 ;
  assign n1560 = n1559 ^ n1557 ^ n1556 ;
  assign n1552 = n610 ^ x146 ^ 1'b0 ;
  assign n1561 = n1560 ^ n1552 ^ 1'b0 ;
  assign n1565 = n1564 ^ n1562 ^ n1561 ;
  assign n1566 = x238 & ~n397 ;
  assign n1573 = ( x68 & n480 ) | ( x68 & ~n707 ) | ( n480 & ~n707 ) ;
  assign n1567 = n1252 ^ n552 ^ x113 ;
  assign n1568 = n1567 ^ n710 ^ n528 ;
  assign n1569 = n831 ^ n501 ^ 1'b0 ;
  assign n1570 = n1569 ^ x202 ^ 1'b0 ;
  assign n1571 = n1568 | n1570 ;
  assign n1572 = n1571 ^ n1380 ^ n401 ;
  assign n1574 = n1573 ^ n1572 ^ 1'b0 ;
  assign n1575 = n1574 ^ n400 ^ x231 ;
  assign n1576 = ( n359 & ~n1293 ) | ( n359 & n1575 ) | ( ~n1293 & n1575 ) ;
  assign n1577 = n671 ^ n583 ^ x16 ;
  assign n1578 = n1339 & ~n1407 ;
  assign n1579 = n1195 & n1578 ;
  assign n1580 = x59 & n1579 ;
  assign n1581 = ( n1349 & n1577 ) | ( n1349 & ~n1580 ) | ( n1577 & ~n1580 ) ;
  assign n1582 = x167 & ~n422 ;
  assign n1585 = n720 ^ n469 ^ x104 ;
  assign n1583 = ( x34 & n368 ) | ( x34 & n860 ) | ( n368 & n860 ) ;
  assign n1584 = x9 & n1583 ;
  assign n1586 = n1585 ^ n1584 ^ 1'b0 ;
  assign n1587 = ( n653 & ~n1582 ) | ( n653 & n1586 ) | ( ~n1582 & n1586 ) ;
  assign n1588 = n862 & ~n1587 ;
  assign n1589 = n949 & ~n1553 ;
  assign n1590 = n1589 ^ n1440 ^ 1'b0 ;
  assign n1591 = ( x4 & ~x149 ) | ( x4 & x192 ) | ( ~x149 & x192 ) ;
  assign n1592 = n1591 ^ n1204 ^ x65 ;
  assign n1593 = n642 | n1592 ;
  assign n1594 = n1593 ^ n1582 ^ 1'b0 ;
  assign n1597 = n766 ^ n334 ^ x167 ;
  assign n1598 = n1597 ^ n1043 ^ 1'b0 ;
  assign n1595 = n839 ^ x84 ^ 1'b0 ;
  assign n1596 = ( n326 & ~n688 ) | ( n326 & n1595 ) | ( ~n688 & n1595 ) ;
  assign n1599 = n1598 ^ n1596 ^ x11 ;
  assign n1602 = n790 ^ x200 ^ x109 ;
  assign n1603 = n361 & n1602 ;
  assign n1604 = n1603 ^ x237 ^ 1'b0 ;
  assign n1600 = ( x175 & n583 ) | ( x175 & n769 ) | ( n583 & n769 ) ;
  assign n1601 = ( n457 & ~n1073 ) | ( n457 & n1600 ) | ( ~n1073 & n1600 ) ;
  assign n1605 = n1604 ^ n1601 ^ n966 ;
  assign n1606 = n629 ^ x251 ^ 1'b0 ;
  assign n1607 = n1606 ^ n1191 ^ 1'b0 ;
  assign n1608 = n1554 & n1607 ;
  assign n1609 = ( n462 & n1605 ) | ( n462 & ~n1608 ) | ( n1605 & ~n1608 ) ;
  assign n1610 = ( n1594 & n1599 ) | ( n1594 & n1609 ) | ( n1599 & n1609 ) ;
  assign n1618 = n1527 ^ n965 ^ n857 ;
  assign n1619 = ( n521 & ~n777 ) | ( n521 & n1618 ) | ( ~n777 & n1618 ) ;
  assign n1611 = ( ~x251 & n379 ) | ( ~x251 & n752 ) | ( n379 & n752 ) ;
  assign n1612 = n1477 ^ x123 ^ x115 ;
  assign n1613 = n1612 ^ n931 ^ x23 ;
  assign n1614 = n1613 ^ n1071 ^ x69 ;
  assign n1615 = n1141 & ~n1614 ;
  assign n1616 = ~x22 & n1615 ;
  assign n1617 = ( ~x81 & n1611 ) | ( ~x81 & n1616 ) | ( n1611 & n1616 ) ;
  assign n1620 = n1619 ^ n1617 ^ n426 ;
  assign n1621 = ( x24 & n683 ) | ( x24 & ~n947 ) | ( n683 & ~n947 ) ;
  assign n1625 = ( n1025 & n1479 ) | ( n1025 & ~n1496 ) | ( n1479 & ~n1496 ) ;
  assign n1626 = n1625 ^ n328 ^ 1'b0 ;
  assign n1623 = n1275 ^ n541 ^ n366 ;
  assign n1624 = n1623 ^ n436 ^ n430 ;
  assign n1622 = n1009 ^ n713 ^ n490 ;
  assign n1627 = n1626 ^ n1624 ^ n1622 ;
  assign n1628 = n693 & n698 ;
  assign n1629 = n564 & n1628 ;
  assign n1630 = ( x17 & n441 ) | ( x17 & n634 ) | ( n441 & n634 ) ;
  assign n1631 = n571 ^ x168 ^ x82 ;
  assign n1632 = ( ~n552 & n1630 ) | ( ~n552 & n1631 ) | ( n1630 & n1631 ) ;
  assign n1633 = n407 ^ x80 ^ 1'b0 ;
  assign n1634 = n1632 & n1633 ;
  assign n1635 = ( n1170 & n1629 ) | ( n1170 & ~n1634 ) | ( n1629 & ~n1634 ) ;
  assign n1636 = n981 ^ n970 ^ n608 ;
  assign n1647 = ( x39 & x101 ) | ( x39 & ~x185 ) | ( x101 & ~x185 ) ;
  assign n1645 = ( x68 & x158 ) | ( x68 & n775 ) | ( x158 & n775 ) ;
  assign n1646 = n1645 ^ n1622 ^ n725 ;
  assign n1637 = ( x96 & ~x251 ) | ( x96 & n874 ) | ( ~x251 & n874 ) ;
  assign n1639 = n1127 ^ n327 ^ x146 ;
  assign n1640 = ~n998 & n1639 ;
  assign n1641 = ~x123 & n1640 ;
  assign n1638 = n537 & ~n597 ;
  assign n1642 = n1641 ^ n1638 ^ n1010 ;
  assign n1643 = x33 & n1642 ;
  assign n1644 = ~n1637 & n1643 ;
  assign n1648 = n1647 ^ n1646 ^ n1644 ;
  assign n1649 = n1567 ^ x184 ^ x3 ;
  assign n1650 = n424 ^ n280 ^ 1'b0 ;
  assign n1651 = n511 | n1650 ;
  assign n1652 = ( n966 & n1649 ) | ( n966 & ~n1651 ) | ( n1649 & ~n1651 ) ;
  assign n1653 = n468 | n1652 ;
  assign n1654 = n389 & ~n1653 ;
  assign n1655 = n874 & n1579 ;
  assign n1656 = n809 ^ n505 ^ x111 ;
  assign n1657 = ( ~n960 & n1655 ) | ( ~n960 & n1656 ) | ( n1655 & n1656 ) ;
  assign n1658 = ~n549 & n1657 ;
  assign n1659 = n1658 ^ n312 ^ 1'b0 ;
  assign n1660 = ( n1092 & ~n1122 ) | ( n1092 & n1515 ) | ( ~n1122 & n1515 ) ;
  assign n1661 = n1079 & ~n1340 ;
  assign n1662 = n1661 ^ x32 ^ 1'b0 ;
  assign n1663 = n1662 ^ n1087 ^ x2 ;
  assign n1664 = ( x172 & n1004 ) | ( x172 & n1663 ) | ( n1004 & n1663 ) ;
  assign n1665 = n1006 ^ n359 ^ x168 ;
  assign n1666 = x100 & x167 ;
  assign n1669 = n621 ^ x121 ^ 1'b0 ;
  assign n1667 = n806 ^ n567 ^ x185 ;
  assign n1668 = n369 & ~n1667 ;
  assign n1670 = n1669 ^ n1668 ^ 1'b0 ;
  assign n1671 = ( x95 & ~x231 ) | ( x95 & n1274 ) | ( ~x231 & n1274 ) ;
  assign n1672 = n1670 & ~n1671 ;
  assign n1673 = n367 & n1672 ;
  assign n1674 = ( n356 & n593 ) | ( n356 & n1673 ) | ( n593 & n1673 ) ;
  assign n1675 = ( n689 & n1666 ) | ( n689 & n1674 ) | ( n1666 & n1674 ) ;
  assign n1676 = n1675 ^ n1553 ^ x147 ;
  assign n1677 = ( n1658 & ~n1665 ) | ( n1658 & n1676 ) | ( ~n1665 & n1676 ) ;
  assign n1678 = ( n1660 & n1664 ) | ( n1660 & n1677 ) | ( n1664 & n1677 ) ;
  assign n1679 = n369 & n1469 ;
  assign n1680 = n423 ^ x108 ^ x10 ;
  assign n1681 = n472 & ~n1579 ;
  assign n1682 = ~n1680 & n1681 ;
  assign n1683 = x109 & n869 ;
  assign n1684 = n1380 & n1683 ;
  assign n1685 = ( x178 & n1682 ) | ( x178 & ~n1684 ) | ( n1682 & ~n1684 ) ;
  assign n1686 = ( ~n519 & n1679 ) | ( ~n519 & n1685 ) | ( n1679 & n1685 ) ;
  assign n1692 = n1568 ^ n725 ^ x100 ;
  assign n1688 = x11 & n264 ;
  assign n1689 = ~n1199 & n1688 ;
  assign n1690 = ( n461 & ~n719 ) | ( n461 & n1689 ) | ( ~n719 & n1689 ) ;
  assign n1687 = n569 | n1145 ;
  assign n1691 = n1690 ^ n1687 ^ 1'b0 ;
  assign n1693 = n1692 ^ n1691 ^ n659 ;
  assign n1694 = ( x19 & ~x129 ) | ( x19 & x238 ) | ( ~x129 & x238 ) ;
  assign n1695 = n1478 | n1694 ;
  assign n1696 = ( x102 & ~n1174 ) | ( x102 & n1695 ) | ( ~n1174 & n1695 ) ;
  assign n1697 = ( ~x52 & x75 ) | ( ~x52 & n263 ) | ( x75 & n263 ) ;
  assign n1698 = x114 & ~n441 ;
  assign n1699 = n1698 ^ n1562 ^ n517 ;
  assign n1700 = ( n339 & n1697 ) | ( n339 & ~n1699 ) | ( n1697 & ~n1699 ) ;
  assign n1705 = n1057 ^ x160 ^ 1'b0 ;
  assign n1702 = n1002 | n1113 ;
  assign n1703 = n1702 ^ x9 ^ 1'b0 ;
  assign n1704 = n1703 ^ n341 ^ x26 ;
  assign n1701 = n1587 ^ n1196 ^ n939 ;
  assign n1706 = n1705 ^ n1704 ^ n1701 ;
  assign n1713 = n1043 ^ x61 ^ x49 ;
  assign n1710 = n517 ^ x89 ^ 1'b0 ;
  assign n1709 = ( ~n1434 & n1469 ) | ( ~n1434 & n1586 ) | ( n1469 & n1586 ) ;
  assign n1707 = n1614 ^ n1445 ^ n373 ;
  assign n1708 = n1707 ^ n1454 ^ 1'b0 ;
  assign n1711 = n1710 ^ n1709 ^ n1708 ;
  assign n1712 = n1711 ^ n566 ^ x14 ;
  assign n1714 = n1713 ^ n1712 ^ 1'b0 ;
  assign n1715 = n710 ^ x65 ^ x13 ;
  assign n1724 = n379 ^ x123 ^ x105 ;
  assign n1725 = ( n330 & n521 ) | ( n330 & n1724 ) | ( n521 & n1724 ) ;
  assign n1726 = ~n1568 & n1725 ;
  assign n1727 = ( n367 & n1523 ) | ( n367 & n1726 ) | ( n1523 & n1726 ) ;
  assign n1718 = n1008 ^ n936 ^ 1'b0 ;
  assign n1719 = n1168 & n1718 ;
  assign n1720 = n1719 ^ n478 ^ 1'b0 ;
  assign n1721 = ~n323 & n1720 ;
  assign n1722 = n1721 ^ n488 ^ x213 ;
  assign n1716 = n310 & ~n900 ;
  assign n1717 = ( n1150 & n1568 ) | ( n1150 & n1716 ) | ( n1568 & n1716 ) ;
  assign n1723 = n1722 ^ n1719 ^ n1717 ;
  assign n1728 = n1727 ^ n1723 ^ 1'b0 ;
  assign n1729 = n1715 | n1728 ;
  assign n1731 = n355 ^ n305 ^ x210 ;
  assign n1732 = n1731 ^ n866 ^ 1'b0 ;
  assign n1733 = ~n334 & n1732 ;
  assign n1730 = n979 ^ n368 ^ 1'b0 ;
  assign n1734 = n1733 ^ n1730 ^ n1253 ;
  assign n1738 = n1484 ^ n904 ^ x132 ;
  assign n1735 = n308 & ~n1514 ;
  assign n1736 = n1735 ^ x201 ^ 1'b0 ;
  assign n1737 = ( n858 & ~n1296 ) | ( n858 & n1736 ) | ( ~n1296 & n1736 ) ;
  assign n1739 = n1738 ^ n1737 ^ n880 ;
  assign n1740 = n911 & ~n1081 ;
  assign n1741 = n1740 ^ x237 ^ 1'b0 ;
  assign n1742 = n610 ^ x174 ^ x2 ;
  assign n1743 = ( x219 & ~n448 ) | ( x219 & n947 ) | ( ~n448 & n947 ) ;
  assign n1744 = n1742 & n1743 ;
  assign n1745 = n1744 ^ n952 ^ n561 ;
  assign n1746 = n820 ^ n396 ^ x174 ;
  assign n1747 = n1746 ^ n779 ^ n665 ;
  assign n1748 = ( x161 & n575 ) | ( x161 & ~n898 ) | ( n575 & ~n898 ) ;
  assign n1749 = ( ~n866 & n1095 ) | ( ~n866 & n1748 ) | ( n1095 & n1748 ) ;
  assign n1750 = n1749 ^ x51 ^ 1'b0 ;
  assign n1751 = n1747 | n1750 ;
  assign n1752 = n646 ^ x87 ^ x73 ;
  assign n1753 = n1752 ^ n1493 ^ n552 ;
  assign n1755 = n1193 ^ n409 ^ x9 ;
  assign n1756 = ( n279 & ~n1116 ) | ( n279 & n1755 ) | ( ~n1116 & n1755 ) ;
  assign n1757 = ( ~x75 & n660 ) | ( ~x75 & n1756 ) | ( n660 & n1756 ) ;
  assign n1754 = n1337 ^ n1044 ^ 1'b0 ;
  assign n1758 = n1757 ^ n1754 ^ n558 ;
  assign n1759 = n1753 & n1758 ;
  assign n1768 = ( x169 & ~x235 ) | ( x169 & n308 ) | ( ~x235 & n308 ) ;
  assign n1764 = x40 & x226 ;
  assign n1765 = n1764 ^ n384 ^ 1'b0 ;
  assign n1761 = n727 & ~n907 ;
  assign n1760 = ( ~x79 & n648 ) | ( ~x79 & n793 ) | ( n648 & n793 ) ;
  assign n1762 = n1761 ^ n1760 ^ 1'b0 ;
  assign n1763 = n306 | n1762 ;
  assign n1766 = n1765 ^ n1763 ^ n775 ;
  assign n1767 = n1766 ^ n1512 ^ x240 ;
  assign n1769 = n1768 ^ n1767 ^ n670 ;
  assign n1770 = n1632 ^ n424 ^ x248 ;
  assign n1771 = n1680 ^ n530 ^ x244 ;
  assign n1772 = n1591 ^ n452 ^ 1'b0 ;
  assign n1773 = ~n1771 & n1772 ;
  assign n1774 = ( ~n790 & n1770 ) | ( ~n790 & n1773 ) | ( n1770 & n1773 ) ;
  assign n1775 = ~n1769 & n1774 ;
  assign n1776 = n994 ^ x216 ^ x2 ;
  assign n1777 = ( n400 & n1181 ) | ( n400 & ~n1532 ) | ( n1181 & ~n1532 ) ;
  assign n1778 = ( n547 & ~n986 ) | ( n547 & n1777 ) | ( ~n986 & n1777 ) ;
  assign n1779 = ( n332 & ~n1518 ) | ( n332 & n1778 ) | ( ~n1518 & n1778 ) ;
  assign n1791 = n476 ^ n432 ^ x45 ;
  assign n1792 = n1791 ^ n810 ^ n656 ;
  assign n1788 = n594 | n1595 ;
  assign n1789 = n1788 ^ x199 ^ 1'b0 ;
  assign n1790 = ( ~n651 & n1510 ) | ( ~n651 & n1789 ) | ( n1510 & n1789 ) ;
  assign n1793 = n1792 ^ n1790 ^ 1'b0 ;
  assign n1785 = n1432 ^ n1083 ^ n313 ;
  assign n1786 = n1638 | n1785 ;
  assign n1787 = n920 | n1786 ;
  assign n1781 = n541 ^ n338 ^ x232 ;
  assign n1782 = n1781 ^ n1733 ^ n733 ;
  assign n1783 = n1782 ^ n692 ^ x165 ;
  assign n1780 = n464 & n523 ;
  assign n1784 = n1783 ^ n1780 ^ n1727 ;
  assign n1794 = n1793 ^ n1787 ^ n1784 ;
  assign n1795 = n887 ^ n782 ^ n498 ;
  assign n1796 = n1795 ^ n1562 ^ n705 ;
  assign n1799 = n1656 ^ x247 ^ 1'b0 ;
  assign n1800 = n1382 | n1799 ;
  assign n1797 = n1441 ^ n1332 ^ n516 ;
  assign n1798 = n1797 ^ n899 ^ x49 ;
  assign n1801 = n1800 ^ n1798 ^ n390 ;
  assign n1802 = ( ~x110 & n838 ) | ( ~x110 & n1801 ) | ( n838 & n1801 ) ;
  assign n1803 = ( ~x46 & x49 ) | ( ~x46 & x148 ) | ( x49 & x148 ) ;
  assign n1804 = n1803 ^ n929 ^ n337 ;
  assign n1805 = ( ~n442 & n1249 ) | ( ~n442 & n1804 ) | ( n1249 & n1804 ) ;
  assign n1806 = ~n1648 & n1805 ;
  assign n1810 = ( n700 & n1161 ) | ( n700 & n1184 ) | ( n1161 & n1184 ) ;
  assign n1807 = n501 ^ n476 ^ x72 ;
  assign n1808 = ~n1511 & n1807 ;
  assign n1809 = n1808 ^ n1071 ^ n382 ;
  assign n1811 = n1810 ^ n1809 ^ n1174 ;
  assign n1816 = n1781 ^ n832 ^ n653 ;
  assign n1812 = n635 ^ n479 ^ x37 ;
  assign n1813 = n1592 ^ n1367 ^ x51 ;
  assign n1814 = ( n581 & n1812 ) | ( n581 & ~n1813 ) | ( n1812 & ~n1813 ) ;
  assign n1815 = n1814 ^ n1594 ^ x2 ;
  assign n1817 = n1816 ^ n1815 ^ n1769 ;
  assign n1818 = n1181 | n1299 ;
  assign n1819 = n1817 & ~n1818 ;
  assign n1824 = n1665 ^ n1145 ^ n569 ;
  assign n1820 = x185 & n1412 ;
  assign n1821 = n1820 ^ x67 ^ 1'b0 ;
  assign n1822 = n541 ^ n338 ^ x50 ;
  assign n1823 = ( ~n1010 & n1821 ) | ( ~n1010 & n1822 ) | ( n1821 & n1822 ) ;
  assign n1825 = n1824 ^ n1823 ^ n964 ;
  assign n1829 = ( x251 & n371 ) | ( x251 & ~n378 ) | ( n371 & ~n378 ) ;
  assign n1827 = n965 ^ n747 ^ x101 ;
  assign n1826 = ( n954 & n956 ) | ( n954 & n1144 ) | ( n956 & n1144 ) ;
  assign n1828 = n1827 ^ n1826 ^ n1325 ;
  assign n1830 = n1829 ^ n1828 ^ n1249 ;
  assign n1831 = ( n1598 & n1719 ) | ( n1598 & ~n1830 ) | ( n1719 & ~n1830 ) ;
  assign n1832 = n1016 ^ n277 ^ x223 ;
  assign n1834 = x224 | n733 ;
  assign n1833 = n675 ^ n290 ^ 1'b0 ;
  assign n1835 = n1834 ^ n1833 ^ x44 ;
  assign n1836 = n916 | n1631 ;
  assign n1837 = n1836 ^ n1568 ^ n299 ;
  assign n1838 = n1837 ^ n954 ^ x58 ;
  assign n1845 = ( x60 & n434 ) | ( x60 & n613 ) | ( n434 & n613 ) ;
  assign n1840 = ( ~x17 & x143 ) | ( ~x17 & n260 ) | ( x143 & n260 ) ;
  assign n1841 = ( ~x70 & n580 ) | ( ~x70 & n1840 ) | ( n580 & n1840 ) ;
  assign n1839 = n1611 ^ n1598 ^ n318 ;
  assign n1842 = n1841 ^ n1839 ^ n962 ;
  assign n1843 = n1842 ^ n380 ^ 1'b0 ;
  assign n1844 = n1797 & ~n1843 ;
  assign n1846 = n1845 ^ n1844 ^ n1783 ;
  assign n1855 = n281 ^ x113 ^ 1'b0 ;
  assign n1856 = ~n651 & n1855 ;
  assign n1857 = n1856 ^ n1532 ^ n699 ;
  assign n1847 = n538 ^ x213 ^ x189 ;
  assign n1849 = x188 ^ x107 ^ x95 ;
  assign n1850 = ( n633 & n985 ) | ( n633 & ~n1849 ) | ( n985 & ~n1849 ) ;
  assign n1851 = ( ~x192 & n1316 ) | ( ~x192 & n1850 ) | ( n1316 & n1850 ) ;
  assign n1852 = ( n339 & ~n680 ) | ( n339 & n1851 ) | ( ~n680 & n1851 ) ;
  assign n1848 = n1587 ^ n549 ^ n321 ;
  assign n1853 = n1852 ^ n1848 ^ 1'b0 ;
  assign n1854 = n1847 | n1853 ;
  assign n1858 = n1857 ^ n1854 ^ 1'b0 ;
  assign n1859 = ( ~n321 & n840 ) | ( ~n321 & n1333 ) | ( n840 & n1333 ) ;
  assign n1860 = n720 ^ n593 ^ x50 ;
  assign n1861 = n552 & ~n1294 ;
  assign n1862 = n1860 & n1861 ;
  assign n1868 = n594 ^ n408 ^ x94 ;
  assign n1867 = ( x31 & n725 ) | ( x31 & ~n743 ) | ( n725 & ~n743 ) ;
  assign n1865 = ( x114 & n631 ) | ( x114 & n710 ) | ( n631 & n710 ) ;
  assign n1866 = ( ~n302 & n690 ) | ( ~n302 & n1865 ) | ( n690 & n1865 ) ;
  assign n1869 = n1868 ^ n1867 ^ n1866 ;
  assign n1870 = ( n392 & n940 ) | ( n392 & ~n1869 ) | ( n940 & ~n1869 ) ;
  assign n1863 = n1182 & n1753 ;
  assign n1864 = ( ~n642 & n1850 ) | ( ~n642 & n1863 ) | ( n1850 & n1863 ) ;
  assign n1871 = n1870 ^ n1864 ^ n986 ;
  assign n1872 = ( n851 & n1198 ) | ( n851 & n1871 ) | ( n1198 & n1871 ) ;
  assign n1880 = x38 & n469 ;
  assign n1881 = n1880 ^ n258 ^ 1'b0 ;
  assign n1873 = ( x183 & n536 ) | ( x183 & n822 ) | ( n536 & n822 ) ;
  assign n1874 = x1 & x88 ;
  assign n1875 = ~n1453 & n1874 ;
  assign n1876 = ( n797 & n1873 ) | ( n797 & n1875 ) | ( n1873 & n1875 ) ;
  assign n1877 = ( n330 & n888 ) | ( n330 & ~n1876 ) | ( n888 & ~n1876 ) ;
  assign n1878 = n1499 ^ n678 ^ x14 ;
  assign n1879 = ( n1797 & ~n1877 ) | ( n1797 & n1878 ) | ( ~n1877 & n1878 ) ;
  assign n1882 = n1881 ^ n1879 ^ n695 ;
  assign n1883 = ( n1082 & n1872 ) | ( n1082 & n1882 ) | ( n1872 & n1882 ) ;
  assign n1884 = x96 & x232 ;
  assign n1885 = ~x237 & n1884 ;
  assign n1886 = ( n833 & n1497 ) | ( n833 & ~n1885 ) | ( n1497 & ~n1885 ) ;
  assign n1887 = n725 ^ n545 ^ n408 ;
  assign n1888 = n1887 ^ n1098 ^ n810 ;
  assign n1889 = ( ~n509 & n904 ) | ( ~n509 & n1313 ) | ( n904 & n1313 ) ;
  assign n1890 = n406 ^ n371 ^ 1'b0 ;
  assign n1891 = n1890 ^ n1018 ^ n448 ;
  assign n1892 = n1891 ^ n941 ^ 1'b0 ;
  assign n1893 = n522 | n1892 ;
  assign n1894 = n1893 ^ x175 ^ x67 ;
  assign n1895 = ( n580 & n1889 ) | ( n580 & ~n1894 ) | ( n1889 & ~n1894 ) ;
  assign n1896 = ~n311 & n1895 ;
  assign n1899 = ( x170 & ~n293 ) | ( x170 & n1568 ) | ( ~n293 & n1568 ) ;
  assign n1897 = n1036 ^ n789 ^ 1'b0 ;
  assign n1898 = n1897 ^ n1478 ^ n1085 ;
  assign n1900 = n1899 ^ n1898 ^ n1731 ;
  assign n1903 = ( ~n315 & n373 ) | ( ~n315 & n975 ) | ( n373 & n975 ) ;
  assign n1904 = n1903 ^ n1558 ^ n1477 ;
  assign n1901 = ( x228 & ~n1382 ) | ( x228 & n1473 ) | ( ~n1382 & n1473 ) ;
  assign n1902 = ( ~n397 & n946 ) | ( ~n397 & n1901 ) | ( n946 & n1901 ) ;
  assign n1905 = n1904 ^ n1902 ^ n271 ;
  assign n1906 = x19 & ~n396 ;
  assign n1907 = ~n1905 & n1906 ;
  assign n1908 = ( x170 & n914 ) | ( x170 & n1907 ) | ( n914 & n1907 ) ;
  assign n1913 = n654 & ~n1792 ;
  assign n1914 = ~n1660 & n1913 ;
  assign n1915 = ( ~n766 & n1765 ) | ( ~n766 & n1914 ) | ( n1765 & n1914 ) ;
  assign n1909 = ( x237 & n736 ) | ( x237 & n775 ) | ( n736 & n775 ) ;
  assign n1910 = n1856 ^ n1139 ^ n696 ;
  assign n1911 = ( n529 & ~n1909 ) | ( n529 & n1910 ) | ( ~n1909 & n1910 ) ;
  assign n1912 = ( n1110 & n1770 ) | ( n1110 & ~n1911 ) | ( n1770 & ~n1911 ) ;
  assign n1916 = n1915 ^ n1912 ^ 1'b0 ;
  assign n1921 = n1112 ^ n1082 ^ n420 ;
  assign n1922 = n1921 ^ n1689 ^ n1669 ;
  assign n1923 = n1922 ^ n1315 ^ n705 ;
  assign n1924 = n1923 ^ n1710 ^ n887 ;
  assign n1917 = x196 & ~n1840 ;
  assign n1918 = n810 & n1917 ;
  assign n1919 = n1918 ^ n1379 ^ n287 ;
  assign n1920 = ( n1135 & n1166 ) | ( n1135 & n1919 ) | ( n1166 & n1919 ) ;
  assign n1925 = n1924 ^ n1920 ^ x200 ;
  assign n1926 = n1925 ^ n613 ^ x61 ;
  assign n1927 = ( x75 & ~x119 ) | ( x75 & n519 ) | ( ~x119 & n519 ) ;
  assign n1928 = n980 ^ n918 ^ x54 ;
  assign n1929 = x161 & ~n680 ;
  assign n1930 = n1929 ^ n345 ^ 1'b0 ;
  assign n1931 = n1754 & ~n1930 ;
  assign n1932 = n1928 & n1931 ;
  assign n1936 = n1002 ^ n724 ^ n587 ;
  assign n1937 = ( x26 & n1841 ) | ( x26 & n1936 ) | ( n1841 & n1936 ) ;
  assign n1938 = ( x55 & ~n432 ) | ( x55 & n1937 ) | ( ~n432 & n1937 ) ;
  assign n1934 = n624 | n1841 ;
  assign n1935 = n689 & ~n1934 ;
  assign n1939 = n1938 ^ n1935 ^ x220 ;
  assign n1933 = n911 & ~n1592 ;
  assign n1940 = n1939 ^ n1933 ^ 1'b0 ;
  assign n1941 = n1940 ^ n927 ^ x195 ;
  assign n1943 = n1695 ^ n1019 ^ n898 ;
  assign n1942 = ( x171 & n554 ) | ( x171 & ~n1069 ) | ( n554 & ~n1069 ) ;
  assign n1944 = n1943 ^ n1942 ^ n912 ;
  assign n1951 = n1899 ^ n990 ^ n744 ;
  assign n1945 = ( n490 & n1139 ) | ( n490 & ~n1738 ) | ( n1139 & ~n1738 ) ;
  assign n1946 = ( n642 & n1047 ) | ( n642 & n1149 ) | ( n1047 & n1149 ) ;
  assign n1947 = n299 | n737 ;
  assign n1948 = n1946 | n1947 ;
  assign n1949 = ~n357 & n1948 ;
  assign n1950 = n1945 & n1949 ;
  assign n1952 = n1951 ^ n1950 ^ n576 ;
  assign n1953 = n807 | n1952 ;
  assign n1959 = x18 & n582 ;
  assign n1956 = n832 ^ x184 ^ x83 ;
  assign n1957 = ( n809 & ~n1319 ) | ( n809 & n1956 ) | ( ~n1319 & n1956 ) ;
  assign n1954 = ( x240 & x245 ) | ( x240 & ~n1943 ) | ( x245 & ~n1943 ) ;
  assign n1955 = x150 & ~n1954 ;
  assign n1958 = n1957 ^ n1955 ^ x180 ;
  assign n1960 = n1959 ^ n1958 ^ n1742 ;
  assign n1963 = n1808 ^ n464 ^ x110 ;
  assign n1961 = ( ~x149 & n506 ) | ( ~x149 & n877 ) | ( n506 & n877 ) ;
  assign n1962 = ( x21 & ~n1305 ) | ( x21 & n1961 ) | ( ~n1305 & n1961 ) ;
  assign n1964 = n1963 ^ n1962 ^ n308 ;
  assign n1965 = ( n857 & ~n1738 ) | ( n857 & n1964 ) | ( ~n1738 & n1964 ) ;
  assign n1966 = n295 & n303 ;
  assign n1967 = n623 & n1966 ;
  assign n1968 = n1967 ^ x183 ^ x64 ;
  assign n1969 = ~n1169 & n1968 ;
  assign n1970 = n367 & n1969 ;
  assign n1971 = n1970 ^ n1778 ^ n1406 ;
  assign n1972 = ( ~n1338 & n1499 ) | ( ~n1338 & n1971 ) | ( n1499 & n1971 ) ;
  assign n1973 = ( ~n333 & n1220 ) | ( ~n333 & n1972 ) | ( n1220 & n1972 ) ;
  assign n1974 = n1973 ^ n688 ^ 1'b0 ;
  assign n1975 = n1965 & n1974 ;
  assign n1976 = ~x12 & n391 ;
  assign n1977 = n333 | n1976 ;
  assign n1978 = ( n321 & n822 ) | ( n321 & n1977 ) | ( n822 & n1977 ) ;
  assign n1979 = ( n392 & n635 ) | ( n392 & n1792 ) | ( n635 & n1792 ) ;
  assign n1980 = n1979 ^ n1483 ^ n1303 ;
  assign n1981 = n1980 ^ n1963 ^ n608 ;
  assign n1982 = n1978 | n1981 ;
  assign n1983 = n1982 ^ x217 ^ 1'b0 ;
  assign n1984 = n1753 ^ n1207 ^ n753 ;
  assign n1985 = n1767 ^ n410 ^ 1'b0 ;
  assign n1986 = n1489 ^ n737 ^ n389 ;
  assign n1987 = n1986 ^ x218 ^ x37 ;
  assign n1988 = ( ~n1010 & n1985 ) | ( ~n1010 & n1987 ) | ( n1985 & n1987 ) ;
  assign n1998 = n514 & n1020 ;
  assign n1999 = ~n1438 & n1998 ;
  assign n1993 = n1639 ^ n1398 ^ n1331 ;
  assign n1992 = x224 & n267 ;
  assign n1994 = n1993 ^ n1992 ^ 1'b0 ;
  assign n1995 = n523 & ~n567 ;
  assign n1996 = ~n897 & n1995 ;
  assign n1997 = ( x3 & ~n1994 ) | ( x3 & n1996 ) | ( ~n1994 & n1996 ) ;
  assign n1989 = n845 ^ n832 ^ n323 ;
  assign n1990 = ( n703 & ~n745 ) | ( n703 & n1989 ) | ( ~n745 & n1989 ) ;
  assign n1991 = ( n1064 & ~n1682 ) | ( n1064 & n1990 ) | ( ~n1682 & n1990 ) ;
  assign n2000 = n1999 ^ n1997 ^ n1991 ;
  assign n2001 = n2000 ^ n529 ^ 1'b0 ;
  assign n2002 = n1346 & n2001 ;
  assign n2003 = n1909 ^ n1416 ^ n1133 ;
  assign n2004 = ( x138 & n406 ) | ( x138 & ~n742 ) | ( n406 & ~n742 ) ;
  assign n2005 = ( ~x86 & n1103 ) | ( ~x86 & n1128 ) | ( n1103 & n1128 ) ;
  assign n2006 = n2005 ^ n1830 ^ 1'b0 ;
  assign n2018 = n1475 ^ n949 ^ n548 ;
  assign n2008 = ( x220 & n332 ) | ( x220 & n446 ) | ( n332 & n446 ) ;
  assign n2007 = x188 & x235 ;
  assign n2009 = n2008 ^ n2007 ^ 1'b0 ;
  assign n2010 = n2009 ^ n1434 ^ n782 ;
  assign n2011 = n2010 ^ n894 ^ 1'b0 ;
  assign n2012 = n328 & n2011 ;
  assign n2013 = x190 & n2012 ;
  assign n2014 = n814 & n2013 ;
  assign n2015 = ( n623 & ~n822 ) | ( n623 & n2014 ) | ( ~n822 & n2014 ) ;
  assign n2016 = ~n372 & n2015 ;
  assign n2017 = n2016 ^ n887 ^ x182 ;
  assign n2019 = n2018 ^ n2017 ^ 1'b0 ;
  assign n2020 = x20 & n2019 ;
  assign n2021 = x78 & n2020 ;
  assign n2022 = n1444 & n2021 ;
  assign n2026 = n558 | n866 ;
  assign n2027 = n2026 ^ n1220 ^ x245 ;
  assign n2024 = x213 ^ x51 ^ 1'b0 ;
  assign n2023 = ( x121 & n492 ) | ( x121 & n1238 ) | ( n492 & n1238 ) ;
  assign n2025 = n2024 ^ n2023 ^ n1164 ;
  assign n2028 = n2027 ^ n2025 ^ 1'b0 ;
  assign n2029 = n2028 ^ n1848 ^ n1199 ;
  assign n2030 = ( ~n425 & n1016 ) | ( ~n425 & n1591 ) | ( n1016 & n1591 ) ;
  assign n2031 = n2030 ^ n846 ^ x18 ;
  assign n2032 = n2031 ^ n1432 ^ 1'b0 ;
  assign n2033 = n1901 ^ n1447 ^ n828 ;
  assign n2034 = ( x250 & n1382 ) | ( x250 & ~n2033 ) | ( n1382 & ~n2033 ) ;
  assign n2035 = ( n1352 & n2032 ) | ( n1352 & n2034 ) | ( n2032 & n2034 ) ;
  assign n2036 = ( x131 & ~n286 ) | ( x131 & n751 ) | ( ~n286 & n751 ) ;
  assign n2037 = ( x54 & ~n706 ) | ( x54 & n2036 ) | ( ~n706 & n2036 ) ;
  assign n2038 = n1343 ^ n1042 ^ x17 ;
  assign n2039 = ( n1444 & ~n1830 ) | ( n1444 & n2038 ) | ( ~n1830 & n2038 ) ;
  assign n2045 = n448 ^ n368 ^ 1'b0 ;
  assign n2046 = ~n720 & n2045 ;
  assign n2047 = ~n389 & n1084 ;
  assign n2048 = n2047 ^ x110 ^ 1'b0 ;
  assign n2049 = ( ~n1139 & n2046 ) | ( ~n1139 & n2048 ) | ( n2046 & n2048 ) ;
  assign n2040 = ( ~n1199 & n1631 ) | ( ~n1199 & n1641 ) | ( n1631 & n1641 ) ;
  assign n2041 = n2040 ^ n1795 ^ n1724 ;
  assign n2042 = ( n373 & ~n826 ) | ( n373 & n2041 ) | ( ~n826 & n2041 ) ;
  assign n2043 = n2042 ^ n588 ^ n301 ;
  assign n2044 = n824 & ~n2043 ;
  assign n2050 = n2049 ^ n2044 ^ 1'b0 ;
  assign n2052 = n492 ^ n405 ^ x189 ;
  assign n2051 = ( ~x143 & x186 ) | ( ~x143 & n1921 ) | ( x186 & n1921 ) ;
  assign n2053 = n2052 ^ n2051 ^ 1'b0 ;
  assign n2054 = n1098 & n2053 ;
  assign n2055 = n1332 ^ n912 ^ 1'b0 ;
  assign n2056 = x24 & ~n2055 ;
  assign n2057 = ~n705 & n2056 ;
  assign n2058 = n964 & n2057 ;
  assign n2059 = n1186 ^ x157 ^ 1'b0 ;
  assign n2060 = ( x252 & ~n1754 ) | ( x252 & n2059 ) | ( ~n1754 & n2059 ) ;
  assign n2061 = ~n2058 & n2060 ;
  assign n2062 = ~n2054 & n2061 ;
  assign n2063 = ~n1161 & n1942 ;
  assign n2064 = n1178 | n2063 ;
  assign n2065 = n2064 ^ n1868 ^ x115 ;
  assign n2066 = n906 ^ n688 ^ n529 ;
  assign n2067 = ( n1238 & n1530 ) | ( n1238 & ~n2066 ) | ( n1530 & ~n2066 ) ;
  assign n2073 = ( ~n320 & n922 ) | ( ~n320 & n1155 ) | ( n922 & n1155 ) ;
  assign n2071 = n1337 ^ n321 ^ 1'b0 ;
  assign n2069 = n998 ^ n546 ^ 1'b0 ;
  assign n2070 = ~n2036 & n2069 ;
  assign n2068 = ( x90 & n409 ) | ( x90 & ~n907 ) | ( n409 & ~n907 ) ;
  assign n2072 = n2071 ^ n2070 ^ n2068 ;
  assign n2074 = n2073 ^ n2072 ^ n546 ;
  assign n2075 = n2073 ^ n388 ^ 1'b0 ;
  assign n2076 = n669 & ~n2075 ;
  assign n2077 = n310 | n2076 ;
  assign n2078 = n2036 ^ n931 ^ 1'b0 ;
  assign n2079 = x37 & n580 ;
  assign n2080 = ~n2078 & n2079 ;
  assign n2081 = ( n1985 & n2032 ) | ( n1985 & n2080 ) | ( n2032 & n2080 ) ;
  assign n2082 = x81 & n1038 ;
  assign n2083 = n1648 & n2082 ;
  assign n2087 = n294 ^ x210 ^ x25 ;
  assign n2086 = x213 & n1591 ;
  assign n2088 = n2087 ^ n2086 ^ 1'b0 ;
  assign n2089 = ( x31 & x150 ) | ( x31 & n2088 ) | ( x150 & n2088 ) ;
  assign n2090 = n2089 ^ n493 ^ n487 ;
  assign n2084 = x24 | n288 ;
  assign n2085 = n1068 & n2084 ;
  assign n2091 = n2090 ^ n2085 ^ 1'b0 ;
  assign n2092 = n2091 ^ n953 ^ n436 ;
  assign n2093 = n569 | n744 ;
  assign n2094 = n772 & ~n2093 ;
  assign n2095 = ( ~n580 & n996 ) | ( ~n580 & n1967 ) | ( n996 & n1967 ) ;
  assign n2096 = n2084 ^ n783 ^ 1'b0 ;
  assign n2097 = ( n597 & n2095 ) | ( n597 & n2096 ) | ( n2095 & n2096 ) ;
  assign n2098 = n1183 ^ n775 ^ x191 ;
  assign n2105 = ( x221 & n1021 ) | ( x221 & n1034 ) | ( n1021 & n1034 ) ;
  assign n2100 = ~x182 & x242 ;
  assign n2099 = n962 ^ n927 ^ 1'b0 ;
  assign n2101 = n2100 ^ n2099 ^ n617 ;
  assign n2102 = ( n397 & n425 ) | ( n397 & ~n538 ) | ( n425 & ~n538 ) ;
  assign n2103 = ( x119 & n1258 ) | ( x119 & n2102 ) | ( n1258 & n2102 ) ;
  assign n2104 = ( n1393 & n2101 ) | ( n1393 & ~n2103 ) | ( n2101 & ~n2103 ) ;
  assign n2106 = n2105 ^ n2104 ^ 1'b0 ;
  assign n2107 = ( ~x229 & n831 ) | ( ~x229 & n1263 ) | ( n831 & n1263 ) ;
  assign n2108 = ( ~x147 & x152 ) | ( ~x147 & n678 ) | ( x152 & n678 ) ;
  assign n2109 = ( n604 & ~n2107 ) | ( n604 & n2108 ) | ( ~n2107 & n2108 ) ;
  assign n2110 = ( n427 & n1194 ) | ( n427 & n1486 ) | ( n1194 & n1486 ) ;
  assign n2111 = n2110 ^ n1198 ^ n998 ;
  assign n2112 = n310 | n2111 ;
  assign n2113 = n2112 ^ n1952 ^ n412 ;
  assign n2114 = n1814 ^ n695 ^ x60 ;
  assign n2137 = ( x50 & ~n906 ) | ( x50 & n1331 ) | ( ~n906 & n1331 ) ;
  assign n2138 = n2137 ^ n1199 ^ x153 ;
  assign n2134 = ( n612 & n846 ) | ( n612 & n1020 ) | ( n846 & n1020 ) ;
  assign n2135 = ( ~n893 & n1268 ) | ( ~n893 & n2134 ) | ( n1268 & n2134 ) ;
  assign n2130 = n1204 & n1928 ;
  assign n2131 = ( x228 & n1080 ) | ( x228 & ~n2130 ) | ( n1080 & ~n2130 ) ;
  assign n2132 = ( n531 & ~n777 ) | ( n531 & n2131 ) | ( ~n777 & n2131 ) ;
  assign n2133 = n2132 ^ n1367 ^ n838 ;
  assign n2115 = ( x24 & x104 ) | ( x24 & ~n501 ) | ( x104 & ~n501 ) ;
  assign n2116 = n582 & ~n1460 ;
  assign n2117 = ~n2115 & n2116 ;
  assign n2118 = n673 ^ x234 ^ 1'b0 ;
  assign n2119 = ~n2117 & n2118 ;
  assign n2120 = n1407 | n1780 ;
  assign n2121 = x14 & n2120 ;
  assign n2122 = ~n2119 & n2121 ;
  assign n2123 = n760 ^ n569 ^ 1'b0 ;
  assign n2124 = n327 & n2123 ;
  assign n2125 = n485 & n2124 ;
  assign n2126 = ( x225 & n346 ) | ( x225 & n1919 ) | ( n346 & n1919 ) ;
  assign n2127 = ( n2122 & n2125 ) | ( n2122 & ~n2126 ) | ( n2125 & ~n2126 ) ;
  assign n2128 = ~n940 & n1648 ;
  assign n2129 = n2127 & n2128 ;
  assign n2136 = n2135 ^ n2133 ^ n2129 ;
  assign n2139 = n2138 ^ n2136 ^ 1'b0 ;
  assign n2140 = n2114 | n2139 ;
  assign n2141 = n1493 ^ n681 ^ n342 ;
  assign n2142 = n1956 ^ n1001 ^ n482 ;
  assign n2143 = ( ~x136 & n303 ) | ( ~x136 & n2142 ) | ( n303 & n2142 ) ;
  assign n2144 = n2143 ^ n904 ^ 1'b0 ;
  assign n2145 = n727 & n2144 ;
  assign n2146 = n2145 ^ n542 ^ 1'b0 ;
  assign n2147 = ( n1605 & ~n2141 ) | ( n1605 & n2146 ) | ( ~n2141 & n2146 ) ;
  assign n2148 = ( ~n293 & n1608 ) | ( ~n293 & n2147 ) | ( n1608 & n2147 ) ;
  assign n2149 = n1575 & ~n1763 ;
  assign n2150 = n2149 ^ n1057 ^ 1'b0 ;
  assign n2151 = ~n839 & n1734 ;
  assign n2152 = n2151 ^ n442 ^ x173 ;
  assign n2153 = ( n562 & n810 ) | ( n562 & n1781 ) | ( n810 & n1781 ) ;
  assign n2154 = ( n335 & n338 ) | ( n335 & ~n568 ) | ( n338 & ~n568 ) ;
  assign n2155 = n588 ^ x35 ^ 1'b0 ;
  assign n2156 = ( n434 & n2154 ) | ( n434 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = ( n700 & n732 ) | ( n700 & ~n2156 ) | ( n732 & ~n2156 ) ;
  assign n2158 = ~n2153 & n2157 ;
  assign n2159 = n2158 ^ n331 ^ 1'b0 ;
  assign n2160 = n704 ^ x176 ^ 1'b0 ;
  assign n2161 = n352 | n2160 ;
  assign n2162 = n2161 ^ x68 ^ 1'b0 ;
  assign n2163 = n1066 | n2161 ;
  assign n2164 = n575 & ~n2163 ;
  assign n2165 = ( n282 & ~n1041 ) | ( n282 & n2164 ) | ( ~n1041 & n2164 ) ;
  assign n2166 = n2162 | n2165 ;
  assign n2167 = n2159 & ~n2166 ;
  assign n2169 = n1567 ^ n1113 ^ 1'b0 ;
  assign n2170 = x125 | n2169 ;
  assign n2171 = n2170 ^ n1611 ^ 1'b0 ;
  assign n2172 = ( ~n486 & n1722 ) | ( ~n486 & n2171 ) | ( n1722 & n2171 ) ;
  assign n2168 = x149 & ~n528 ;
  assign n2173 = n2172 ^ n2168 ^ x118 ;
  assign n2176 = n747 ^ x243 ^ x168 ;
  assign n2174 = n1619 ^ n1601 ^ n610 ;
  assign n2175 = n2174 ^ n1866 ^ n1061 ;
  assign n2177 = n2176 ^ n2175 ^ n488 ;
  assign n2178 = n2177 ^ n1063 ^ 1'b0 ;
  assign n2179 = n1710 ^ x83 ^ x53 ;
  assign n2180 = n375 | n2179 ;
  assign n2181 = x211 & n1163 ;
  assign n2182 = n1792 & n2181 ;
  assign n2183 = ( ~n632 & n727 ) | ( ~n632 & n2182 ) | ( n727 & n2182 ) ;
  assign n2184 = n1328 ^ n1135 ^ 1'b0 ;
  assign n2185 = n2183 & ~n2184 ;
  assign n2186 = n262 & n2185 ;
  assign n2187 = n2186 ^ n943 ^ 1'b0 ;
  assign n2188 = ( n328 & ~n440 ) | ( n328 & n1046 ) | ( ~n440 & n1046 ) ;
  assign n2189 = n1155 ^ x184 ^ 1'b0 ;
  assign n2190 = n1233 & n2189 ;
  assign n2191 = ( x191 & ~n2188 ) | ( x191 & n2190 ) | ( ~n2188 & n2190 ) ;
  assign n2192 = n1012 ^ n771 ^ n437 ;
  assign n2193 = n2192 ^ n270 ^ 1'b0 ;
  assign n2194 = n1021 ^ n290 ^ 1'b0 ;
  assign n2195 = n2194 ^ n957 ^ 1'b0 ;
  assign n2196 = n406 & n2195 ;
  assign n2197 = ( ~n637 & n1697 ) | ( ~n637 & n2196 ) | ( n1697 & n2196 ) ;
  assign n2198 = n1106 & ~n2197 ;
  assign n2199 = n2198 ^ n2073 ^ 1'b0 ;
  assign n2200 = n828 ^ n701 ^ x224 ;
  assign n2201 = ( n361 & n565 ) | ( n361 & n2200 ) | ( n565 & n2200 ) ;
  assign n2202 = n1511 ^ n696 ^ n521 ;
  assign n2203 = n1159 & n1923 ;
  assign n2204 = n1662 & n2203 ;
  assign n2205 = n2204 ^ n1507 ^ n676 ;
  assign n2206 = ( n571 & ~n2202 ) | ( n571 & n2205 ) | ( ~n2202 & n2205 ) ;
  assign n2207 = n2201 & ~n2206 ;
  assign n2208 = n2207 ^ n1596 ^ 1'b0 ;
  assign n2209 = ( ~n1631 & n1790 ) | ( ~n1631 & n2191 ) | ( n1790 & n2191 ) ;
  assign n2222 = n283 ^ x200 ^ x102 ;
  assign n2210 = ( x233 & n642 ) | ( x233 & n831 ) | ( n642 & n831 ) ;
  assign n2211 = n1220 ^ n488 ^ x166 ;
  assign n2212 = n2211 ^ n1032 ^ n401 ;
  assign n2219 = n1149 ^ n423 ^ n279 ;
  assign n2216 = n1533 ^ n1223 ^ n1182 ;
  assign n2213 = n1373 ^ n976 ^ n514 ;
  assign n2214 = ~n1546 & n2213 ;
  assign n2215 = n2214 ^ n725 ^ 1'b0 ;
  assign n2217 = n2216 ^ n2215 ^ n1597 ;
  assign n2218 = ( x18 & ~n742 ) | ( x18 & n2217 ) | ( ~n742 & n2217 ) ;
  assign n2220 = n2219 ^ n2218 ^ n2103 ;
  assign n2221 = ( n2210 & ~n2212 ) | ( n2210 & n2220 ) | ( ~n2212 & n2220 ) ;
  assign n2223 = n2222 ^ n2221 ^ n1670 ;
  assign n2224 = ( ~n929 & n994 ) | ( ~n929 & n1967 ) | ( n994 & n1967 ) ;
  assign n2225 = x40 & ~n2224 ;
  assign n2226 = n2225 ^ n932 ^ n635 ;
  assign n2227 = ( n335 & n540 ) | ( n335 & ~n1112 ) | ( n540 & ~n1112 ) ;
  assign n2228 = n2227 ^ n339 ^ 1'b0 ;
  assign n2229 = n929 ^ n746 ^ n411 ;
  assign n2230 = x88 & ~x113 ;
  assign n2231 = ( n265 & n1572 ) | ( n265 & ~n1698 ) | ( n1572 & ~n1698 ) ;
  assign n2232 = ( n1001 & n2230 ) | ( n1001 & ~n2231 ) | ( n2230 & ~n2231 ) ;
  assign n2233 = x225 & n477 ;
  assign n2234 = ( n2229 & n2232 ) | ( n2229 & ~n2233 ) | ( n2232 & ~n2233 ) ;
  assign n2235 = ( n777 & n1601 ) | ( n777 & n2234 ) | ( n1601 & n2234 ) ;
  assign n2236 = x1 & n652 ;
  assign n2237 = n2236 ^ x210 ^ 1'b0 ;
  assign n2238 = n2237 ^ n543 ^ n320 ;
  assign n2239 = ( n460 & n811 ) | ( n460 & n1223 ) | ( n811 & n1223 ) ;
  assign n2240 = n2238 & ~n2239 ;
  assign n2245 = n1478 ^ n810 ^ x242 ;
  assign n2246 = n2245 ^ n1043 ^ n721 ;
  assign n2241 = n1157 ^ n1103 ^ n582 ;
  assign n2242 = n2241 ^ n2172 ^ n800 ;
  assign n2243 = ( n1004 & n1771 ) | ( n1004 & ~n1897 ) | ( n1771 & ~n1897 ) ;
  assign n2244 = n2242 | n2243 ;
  assign n2247 = n2246 ^ n2244 ^ n359 ;
  assign n2248 = n1436 ^ n1088 ^ n971 ;
  assign n2251 = n1812 ^ n1207 ^ n703 ;
  assign n2269 = n2251 ^ x226 ^ x70 ;
  assign n2270 = n2269 ^ n1841 ^ 1'b0 ;
  assign n2271 = n981 | n2270 ;
  assign n2249 = n330 & n714 ;
  assign n2250 = ~n1122 & n2249 ;
  assign n2252 = n983 ^ x59 ^ 1'b0 ;
  assign n2253 = n2251 | n2252 ;
  assign n2254 = ( x121 & n2194 ) | ( x121 & n2253 ) | ( n2194 & n2253 ) ;
  assign n2255 = ( n1371 & ~n2250 ) | ( n1371 & n2254 ) | ( ~n2250 & n2254 ) ;
  assign n2256 = ( ~x185 & n504 ) | ( ~x185 & n866 ) | ( n504 & n866 ) ;
  assign n2257 = ( n1495 & n1970 ) | ( n1495 & n2256 ) | ( n1970 & n2256 ) ;
  assign n2258 = ( n468 & n1347 ) | ( n468 & n1780 ) | ( n1347 & n1780 ) ;
  assign n2259 = ~n954 & n2258 ;
  assign n2260 = n2259 ^ n1849 ^ 1'b0 ;
  assign n2261 = ( n1258 & n2257 ) | ( n1258 & n2260 ) | ( n2257 & n2260 ) ;
  assign n2262 = ( x87 & ~n509 ) | ( x87 & n1347 ) | ( ~n509 & n1347 ) ;
  assign n2263 = ( n579 & n1102 ) | ( n579 & ~n1725 ) | ( n1102 & ~n1725 ) ;
  assign n2264 = n2263 ^ n661 ^ 1'b0 ;
  assign n2265 = n339 & ~n2264 ;
  assign n2266 = n2265 ^ n1344 ^ 1'b0 ;
  assign n2267 = n2262 & ~n2266 ;
  assign n2268 = ( n2255 & ~n2261 ) | ( n2255 & n2267 ) | ( ~n2261 & n2267 ) ;
  assign n2272 = n2271 ^ n2268 ^ n576 ;
  assign n2273 = n446 ^ x148 ^ x117 ;
  assign n2274 = ~n455 & n2273 ;
  assign n2275 = n2274 ^ n286 ^ 1'b0 ;
  assign n2282 = n1384 ^ n785 ^ 1'b0 ;
  assign n2283 = x148 & ~n2282 ;
  assign n2284 = n2009 ^ n1125 ^ 1'b0 ;
  assign n2285 = n2283 & ~n2284 ;
  assign n2276 = n968 ^ n521 ^ 1'b0 ;
  assign n2277 = n2255 ^ n1989 ^ 1'b0 ;
  assign n2278 = n1392 | n2277 ;
  assign n2279 = n2278 ^ n1166 ^ 1'b0 ;
  assign n2280 = ~n2276 & n2279 ;
  assign n2281 = n1790 & n2280 ;
  assign n2286 = n2285 ^ n2281 ^ 1'b0 ;
  assign n2287 = ( ~n1174 & n2275 ) | ( ~n1174 & n2286 ) | ( n2275 & n2286 ) ;
  assign n2288 = n883 & n2273 ;
  assign n2289 = n2288 ^ x172 ^ 1'b0 ;
  assign n2290 = ( n405 & ~n2169 ) | ( n405 & n2289 ) | ( ~n2169 & n2289 ) ;
  assign n2291 = ( ~n1371 & n1574 ) | ( ~n1371 & n2046 ) | ( n1574 & n2046 ) ;
  assign n2292 = ( ~n814 & n1382 ) | ( ~n814 & n2291 ) | ( n1382 & n2291 ) ;
  assign n2293 = n1114 ^ n612 ^ 1'b0 ;
  assign n2294 = n2293 ^ n1429 ^ n370 ;
  assign n2295 = ( n410 & n824 ) | ( n410 & n847 ) | ( n824 & n847 ) ;
  assign n2296 = n2295 ^ n1352 ^ x134 ;
  assign n2297 = ( n565 & n2294 ) | ( n565 & ~n2296 ) | ( n2294 & ~n2296 ) ;
  assign n2298 = ( ~n2038 & n2292 ) | ( ~n2038 & n2297 ) | ( n2292 & n2297 ) ;
  assign n2299 = n1441 & ~n2089 ;
  assign n2300 = n1515 ^ n1185 ^ n286 ;
  assign n2301 = n2300 ^ n1752 ^ x38 ;
  assign n2302 = n753 ^ n743 ^ n420 ;
  assign n2303 = ( n655 & n1528 ) | ( n655 & ~n2302 ) | ( n1528 & ~n2302 ) ;
  assign n2304 = ( n1809 & ~n2301 ) | ( n1809 & n2303 ) | ( ~n2301 & n2303 ) ;
  assign n2305 = n2074 ^ n1520 ^ n494 ;
  assign n2309 = ( n287 & n506 ) | ( n287 & ~n1296 ) | ( n506 & ~n1296 ) ;
  assign n2310 = n2309 ^ n841 ^ n523 ;
  assign n2311 = n2310 ^ n1808 ^ n687 ;
  assign n2308 = n947 ^ n343 ^ x159 ;
  assign n2306 = x189 & n869 ;
  assign n2307 = n2306 ^ x251 ^ 1'b0 ;
  assign n2312 = n2311 ^ n2308 ^ n2307 ;
  assign n2317 = n546 ^ x27 ^ 1'b0 ;
  assign n2318 = n2317 ^ n956 ^ n952 ;
  assign n2313 = n1463 ^ n987 ^ x232 ;
  assign n2314 = ~n692 & n2313 ;
  assign n2315 = n2314 ^ n733 ^ 1'b0 ;
  assign n2316 = n1366 & n2315 ;
  assign n2319 = n2318 ^ n2316 ^ n654 ;
  assign n2320 = ( ~n348 & n1631 ) | ( ~n348 & n1999 ) | ( n1631 & n1999 ) ;
  assign n2321 = n1528 | n2320 ;
  assign n2322 = n1948 | n2321 ;
  assign n2323 = n377 ^ x144 ^ 1'b0 ;
  assign n2324 = ( x119 & ~n2102 ) | ( x119 & n2323 ) | ( ~n2102 & n2323 ) ;
  assign n2325 = n2324 ^ n2172 ^ n1553 ;
  assign n2326 = ( n313 & n792 ) | ( n313 & ~n856 ) | ( n792 & ~n856 ) ;
  assign n2328 = ( x38 & n1283 ) | ( x38 & n1344 ) | ( n1283 & n1344 ) ;
  assign n2327 = n1745 & ~n1898 ;
  assign n2329 = n2328 ^ n2327 ^ 1'b0 ;
  assign n2330 = n1746 & n2329 ;
  assign n2331 = n1604 ^ n1562 ^ n1105 ;
  assign n2332 = n1419 ^ n1185 ^ n642 ;
  assign n2333 = ( x212 & ~n505 ) | ( x212 & n1180 ) | ( ~n505 & n1180 ) ;
  assign n2334 = x205 ^ x194 ^ x108 ;
  assign n2335 = n2334 ^ n2217 ^ n548 ;
  assign n2336 = n2335 ^ n1386 ^ n975 ;
  assign n2337 = n893 & n1362 ;
  assign n2338 = ( ~n1583 & n2336 ) | ( ~n1583 & n2337 ) | ( n2336 & n2337 ) ;
  assign n2339 = ( n905 & n2333 ) | ( n905 & ~n2338 ) | ( n2333 & ~n2338 ) ;
  assign n2340 = n1930 ^ x139 ^ 1'b0 ;
  assign n2341 = x58 & ~n2340 ;
  assign n2342 = n1384 ^ n607 ^ x149 ;
  assign n2343 = n2342 ^ n323 ^ x100 ;
  assign n2344 = n2343 ^ n1165 ^ n461 ;
  assign n2352 = n727 ^ n528 ^ n484 ;
  assign n2349 = x140 & n574 ;
  assign n2350 = ( n539 & n716 ) | ( n539 & n2349 ) | ( n716 & n2349 ) ;
  assign n2345 = ( ~x17 & n384 ) | ( ~x17 & n1268 ) | ( n384 & n1268 ) ;
  assign n2346 = ~n663 & n2345 ;
  assign n2347 = n665 & n2346 ;
  assign n2348 = n2347 ^ n541 ^ n502 ;
  assign n2351 = n2350 ^ n2348 ^ n1731 ;
  assign n2353 = n2352 ^ n2351 ^ 1'b0 ;
  assign n2354 = n2344 & ~n2353 ;
  assign n2355 = n498 & n1829 ;
  assign n2356 = n2355 ^ n747 ^ 1'b0 ;
  assign n2357 = n491 ^ x124 ^ 1'b0 ;
  assign n2358 = x27 & ~n2357 ;
  assign n2359 = n2358 ^ n2119 ^ 1'b0 ;
  assign n2360 = x31 & n2359 ;
  assign n2361 = ~x112 & n2360 ;
  assign n2362 = n2361 ^ n1684 ^ n1385 ;
  assign n2363 = n1611 ^ n771 ^ 1'b0 ;
  assign n2364 = ( n715 & n1878 ) | ( n715 & n2363 ) | ( n1878 & n2363 ) ;
  assign n2365 = ( n2356 & ~n2362 ) | ( n2356 & n2364 ) | ( ~n2362 & n2364 ) ;
  assign n2366 = n2365 ^ n1883 ^ n710 ;
  assign n2367 = ( n1440 & n1991 ) | ( n1440 & n2311 ) | ( n1991 & n2311 ) ;
  assign n2368 = ( ~x30 & n621 ) | ( ~x30 & n716 ) | ( n621 & n716 ) ;
  assign n2369 = ( n768 & n2367 ) | ( n768 & ~n2368 ) | ( n2367 & ~n2368 ) ;
  assign n2370 = n814 | n1372 ;
  assign n2371 = n1840 & ~n2370 ;
  assign n2372 = ( n518 & n1240 ) | ( n518 & n2371 ) | ( n1240 & n2371 ) ;
  assign n2374 = n555 ^ x235 ^ x91 ;
  assign n2373 = x110 & x166 ;
  assign n2375 = n2374 ^ n2373 ^ 1'b0 ;
  assign n2376 = n1299 | n2375 ;
  assign n2377 = n331 & ~n2376 ;
  assign n2378 = ~x249 & n2377 ;
  assign n2379 = n2378 ^ n1482 ^ n1159 ;
  assign n2380 = n2379 ^ n1724 ^ 1'b0 ;
  assign n2381 = ~n2372 & n2380 ;
  assign n2382 = n569 | n1199 ;
  assign n2383 = n1001 ^ n390 ^ n384 ;
  assign n2384 = ( n311 & ~n2324 ) | ( n311 & n2383 ) | ( ~n2324 & n2383 ) ;
  assign n2385 = ( ~n544 & n2382 ) | ( ~n544 & n2384 ) | ( n2382 & n2384 ) ;
  assign n2386 = x188 & x228 ;
  assign n2387 = ( n505 & n1032 ) | ( n505 & ~n2386 ) | ( n1032 & ~n2386 ) ;
  assign n2388 = n297 ^ n286 ^ x252 ;
  assign n2389 = ( ~x101 & n2078 ) | ( ~x101 & n2388 ) | ( n2078 & n2388 ) ;
  assign n2390 = n452 & ~n704 ;
  assign n2391 = ~n548 & n2390 ;
  assign n2392 = ( n1445 & n2389 ) | ( n1445 & ~n2391 ) | ( n2389 & ~n2391 ) ;
  assign n2402 = n1789 & ~n2137 ;
  assign n2400 = n1324 ^ n321 ^ 1'b0 ;
  assign n2401 = ( x46 & ~n338 ) | ( x46 & n2400 ) | ( ~n338 & n2400 ) ;
  assign n2393 = ( n335 & n1045 ) | ( n335 & ~n2101 ) | ( n1045 & ~n2101 ) ;
  assign n2394 = n2393 ^ n1583 ^ x245 ;
  assign n2395 = ( n304 & n701 ) | ( n304 & n931 ) | ( n701 & n931 ) ;
  assign n2396 = ( ~n342 & n1015 ) | ( ~n342 & n1157 ) | ( n1015 & n1157 ) ;
  assign n2397 = n2396 ^ n375 ^ n324 ;
  assign n2398 = ~n2395 & n2397 ;
  assign n2399 = ~n2394 & n2398 ;
  assign n2403 = n2402 ^ n2401 ^ n2399 ;
  assign n2404 = n2403 ^ n1377 ^ 1'b0 ;
  assign n2406 = ( x46 & n595 ) | ( x46 & ~n2384 ) | ( n595 & ~n2384 ) ;
  assign n2405 = n377 | n1450 ;
  assign n2407 = n2406 ^ n2405 ^ n1957 ;
  assign n2408 = ( x223 & ~n804 ) | ( x223 & n1597 ) | ( ~n804 & n1597 ) ;
  assign n2409 = n2084 ^ n1692 ^ 1'b0 ;
  assign n2410 = ~n1914 & n2409 ;
  assign n2411 = ~n855 & n2170 ;
  assign n2412 = n522 & n2411 ;
  assign n2413 = ( n2408 & ~n2410 ) | ( n2408 & n2412 ) | ( ~n2410 & n2412 ) ;
  assign n2414 = ( x45 & ~n403 ) | ( x45 & n1363 ) | ( ~n403 & n1363 ) ;
  assign n2415 = ( x101 & ~n1387 ) | ( x101 & n2414 ) | ( ~n1387 & n2414 ) ;
  assign n2416 = n2415 ^ n2178 ^ n2099 ;
  assign n2417 = n1555 ^ n666 ^ x94 ;
  assign n2418 = n661 & n1290 ;
  assign n2419 = ~n2095 & n2418 ;
  assign n2420 = n2419 ^ n1484 ^ 1'b0 ;
  assign n2421 = n2420 ^ n923 ^ n480 ;
  assign n2422 = n2421 ^ n1927 ^ x216 ;
  assign n2423 = ( ~n415 & n2417 ) | ( ~n415 & n2422 ) | ( n2417 & n2422 ) ;
  assign n2424 = n724 & ~n2257 ;
  assign n2425 = n1785 ^ n1016 ^ n838 ;
  assign n2426 = n774 | n2425 ;
  assign n2427 = ( n296 & n785 ) | ( n296 & ~n2426 ) | ( n785 & ~n2426 ) ;
  assign n2428 = ( x132 & n2424 ) | ( x132 & n2427 ) | ( n2424 & n2427 ) ;
  assign n2436 = n652 & n1914 ;
  assign n2437 = ( x175 & ~n2201 ) | ( x175 & n2436 ) | ( ~n2201 & n2436 ) ;
  assign n2429 = n2410 ^ n1503 ^ 1'b0 ;
  assign n2432 = n1175 ^ n776 ^ x64 ;
  assign n2430 = ( ~n826 & n1193 ) | ( ~n826 & n1935 ) | ( n1193 & n1935 ) ;
  assign n2431 = ( n915 & n1727 ) | ( n915 & ~n2430 ) | ( n1727 & ~n2430 ) ;
  assign n2433 = n2432 ^ n2431 ^ n345 ;
  assign n2434 = n2300 | n2433 ;
  assign n2435 = n2429 | n2434 ;
  assign n2438 = n2437 ^ n2435 ^ 1'b0 ;
  assign n2439 = n642 | n2438 ;
  assign n2440 = n1972 ^ n1663 ^ 1'b0 ;
  assign n2441 = n502 ^ n501 ^ 1'b0 ;
  assign n2442 = n2441 ^ n1406 ^ n822 ;
  assign n2443 = n2442 ^ n1800 ^ n1116 ;
  assign n2444 = n1558 ^ n1469 ^ n577 ;
  assign n2445 = n1597 ^ n594 ^ n525 ;
  assign n2446 = n1419 | n2445 ;
  assign n2447 = ( n2443 & ~n2444 ) | ( n2443 & n2446 ) | ( ~n2444 & n2446 ) ;
  assign n2448 = ( n1938 & n2440 ) | ( n1938 & ~n2447 ) | ( n2440 & ~n2447 ) ;
  assign n2449 = n842 | n2024 ;
  assign n2450 = n1112 | n2449 ;
  assign n2451 = n2450 ^ n912 ^ n756 ;
  assign n2455 = x199 ^ x178 ^ x132 ;
  assign n2453 = n583 ^ n440 ^ x163 ;
  assign n2452 = ( ~n748 & n1081 ) | ( ~n748 & n1090 ) | ( n1081 & n1090 ) ;
  assign n2454 = n2453 ^ n2452 ^ n951 ;
  assign n2456 = n2455 ^ n2454 ^ n1041 ;
  assign n2457 = ( n1174 & ~n1243 ) | ( n1174 & n2456 ) | ( ~n1243 & n2456 ) ;
  assign n2458 = n1049 & n2457 ;
  assign n2459 = n1873 ^ n1324 ^ n1227 ;
  assign n2460 = n2459 ^ n1909 ^ n1316 ;
  assign n2461 = n2155 ^ n1694 ^ 1'b0 ;
  assign n2462 = n2253 | n2461 ;
  assign n2463 = n556 & ~n2462 ;
  assign n2464 = ~n2460 & n2463 ;
  assign n2465 = ( x196 & ~n894 ) | ( x196 & n1774 ) | ( ~n894 & n1774 ) ;
  assign n2466 = n2465 ^ n1872 ^ 1'b0 ;
  assign n2467 = n1491 | n1571 ;
  assign n2468 = n2467 ^ n2171 ^ n1965 ;
  assign n2469 = ( ~n689 & n895 ) | ( ~n689 & n1836 ) | ( n895 & n1836 ) ;
  assign n2470 = n2469 ^ n487 ^ 1'b0 ;
  assign n2471 = n1233 & n2470 ;
  assign n2476 = n1829 ^ x33 ^ 1'b0 ;
  assign n2472 = n2046 ^ n397 ^ 1'b0 ;
  assign n2473 = n2472 ^ n904 ^ x142 ;
  assign n2474 = ( x206 & ~n829 ) | ( x206 & n936 ) | ( ~n829 & n936 ) ;
  assign n2475 = ( n1700 & n2473 ) | ( n1700 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2477 = n2476 ^ n2475 ^ n1063 ;
  assign n2480 = ( n1313 & ~n1411 ) | ( n1313 & n1704 ) | ( ~n1411 & n1704 ) ;
  assign n2478 = n1605 ^ n583 ^ 1'b0 ;
  assign n2479 = n2478 ^ n2415 ^ n1696 ;
  assign n2481 = n2480 ^ n2479 ^ n632 ;
  assign n2482 = ( x162 & n267 ) | ( x162 & ~n1904 ) | ( n267 & ~n1904 ) ;
  assign n2484 = n480 & n824 ;
  assign n2483 = n2348 ^ n445 ^ n414 ;
  assign n2485 = n2484 ^ n2483 ^ x156 ;
  assign n2486 = n2485 ^ n2396 ^ n604 ;
  assign n2487 = n1956 & ~n2486 ;
  assign n2488 = ( n855 & n2482 ) | ( n855 & ~n2487 ) | ( n2482 & ~n2487 ) ;
  assign n2495 = ( x26 & n1318 ) | ( x26 & n1406 ) | ( n1318 & n1406 ) ;
  assign n2489 = x45 & x81 ;
  assign n2490 = n2489 ^ n501 ^ 1'b0 ;
  assign n2492 = n1461 ^ x213 ^ x87 ;
  assign n2491 = n1377 ^ n1053 ^ n556 ;
  assign n2493 = n2492 ^ n2491 ^ 1'b0 ;
  assign n2494 = ( n654 & n2490 ) | ( n654 & ~n2493 ) | ( n2490 & ~n2493 ) ;
  assign n2496 = n2495 ^ n2494 ^ 1'b0 ;
  assign n2497 = n2481 ^ n1043 ^ 1'b0 ;
  assign n2498 = n284 & ~n1059 ;
  assign n2499 = ( n1093 & n1326 ) | ( n1093 & n2498 ) | ( n1326 & n2498 ) ;
  assign n2500 = ( x20 & n1241 ) | ( x20 & ~n2499 ) | ( n1241 & ~n2499 ) ;
  assign n2501 = ( ~n267 & n622 ) | ( ~n267 & n2500 ) | ( n622 & n2500 ) ;
  assign n2502 = ( x68 & ~n1261 ) | ( x68 & n1757 ) | ( ~n1261 & n1757 ) ;
  assign n2503 = n1903 ^ n1546 ^ 1'b0 ;
  assign n2504 = n1263 & ~n2503 ;
  assign n2505 = ( n1704 & n2502 ) | ( n1704 & n2504 ) | ( n2502 & n2504 ) ;
  assign n2506 = n2395 ^ n600 ^ n575 ;
  assign n2507 = n2506 ^ n500 ^ x193 ;
  assign n2510 = ( ~x40 & x55 ) | ( ~x40 & x73 ) | ( x55 & x73 ) ;
  assign n2508 = x85 & ~n410 ;
  assign n2509 = n1461 & n2508 ;
  assign n2511 = n2510 ^ n2509 ^ 1'b0 ;
  assign n2512 = ( n2078 & n2507 ) | ( n2078 & ~n2511 ) | ( n2507 & ~n2511 ) ;
  assign n2513 = ~n940 & n2512 ;
  assign n2514 = ~n2505 & n2513 ;
  assign n2517 = ( x63 & ~n496 ) | ( x63 & n2117 ) | ( ~n496 & n2117 ) ;
  assign n2518 = n2517 ^ x227 ^ x107 ;
  assign n2515 = n1669 ^ n779 ^ n769 ;
  assign n2516 = ( n1495 & ~n1604 ) | ( n1495 & n2515 ) | ( ~n1604 & n2515 ) ;
  assign n2519 = n2518 ^ n2516 ^ x45 ;
  assign n2523 = ( n895 & ~n1153 ) | ( n895 & n1822 ) | ( ~n1153 & n1822 ) ;
  assign n2520 = n1224 ^ n1006 ^ x131 ;
  assign n2521 = n752 & n2520 ;
  assign n2522 = ( ~n881 & n997 ) | ( ~n881 & n2521 ) | ( n997 & n2521 ) ;
  assign n2524 = n2523 ^ n2522 ^ n1751 ;
  assign n2529 = n1904 & n2102 ;
  assign n2530 = n2529 ^ n895 ^ 1'b0 ;
  assign n2527 = n412 ^ n320 ^ n276 ;
  assign n2525 = n806 ^ n661 ^ x121 ;
  assign n2526 = ( ~x46 & n1522 ) | ( ~x46 & n2525 ) | ( n1522 & n2525 ) ;
  assign n2528 = n2527 ^ n2526 ^ n1085 ;
  assign n2531 = n2530 ^ n2528 ^ 1'b0 ;
  assign n2532 = n2531 ^ n1944 ^ 1'b0 ;
  assign n2533 = n625 & n2532 ;
  assign n2534 = n1053 ^ n566 ^ 1'b0 ;
  assign n2535 = n829 & ~n2534 ;
  assign n2536 = n2535 ^ n1301 ^ n686 ;
  assign n2537 = n2324 ^ n1518 ^ x168 ;
  assign n2538 = ( n2174 & n2523 ) | ( n2174 & n2537 ) | ( n2523 & n2537 ) ;
  assign n2554 = ( n722 & ~n1254 ) | ( n722 & n1785 ) | ( ~n1254 & n1785 ) ;
  assign n2539 = n897 ^ n441 ^ 1'b0 ;
  assign n2540 = ( ~n293 & n439 ) | ( ~n293 & n2539 ) | ( n439 & n2539 ) ;
  assign n2547 = x102 & x171 ;
  assign n2548 = ~n2527 & n2547 ;
  assign n2549 = n1507 | n2155 ;
  assign n2550 = n2445 | n2549 ;
  assign n2551 = ( n686 & n2548 ) | ( n686 & ~n2550 ) | ( n2548 & ~n2550 ) ;
  assign n2541 = n1155 ^ n362 ^ x52 ;
  assign n2542 = n2012 ^ n482 ^ n436 ;
  assign n2543 = ( ~n1546 & n2170 ) | ( ~n1546 & n2542 ) | ( n2170 & n2542 ) ;
  assign n2544 = n2543 ^ n1996 ^ 1'b0 ;
  assign n2545 = ( n1529 & n1857 ) | ( n1529 & ~n1924 ) | ( n1857 & ~n1924 ) ;
  assign n2546 = ( n2541 & ~n2544 ) | ( n2541 & n2545 ) | ( ~n2544 & n2545 ) ;
  assign n2552 = n2551 ^ n2546 ^ 1'b0 ;
  assign n2553 = ~n2540 & n2552 ;
  assign n2555 = n2554 ^ n2553 ^ n1638 ;
  assign n2556 = n2350 ^ n1164 ^ x99 ;
  assign n2557 = ( n599 & n2296 ) | ( n599 & n2556 ) | ( n2296 & n2556 ) ;
  assign n2558 = n2388 ^ n1379 ^ n973 ;
  assign n2559 = ~n815 & n2558 ;
  assign n2560 = ( n541 & n2557 ) | ( n541 & n2559 ) | ( n2557 & n2559 ) ;
  assign n2561 = ( n969 & ~n2555 ) | ( n969 & n2560 ) | ( ~n2555 & n2560 ) ;
  assign n2562 = ~n1517 & n1736 ;
  assign n2563 = n1897 ^ n1840 ^ 1'b0 ;
  assign n2564 = n2563 ^ n1325 ^ n1103 ;
  assign n2569 = x38 | n1551 ;
  assign n2565 = n1667 ^ n282 ^ x110 ;
  assign n2566 = ( x73 & n295 ) | ( x73 & n2565 ) | ( n295 & n2565 ) ;
  assign n2567 = ( n1266 & ~n2005 ) | ( n1266 & n2566 ) | ( ~n2005 & n2566 ) ;
  assign n2568 = ( n518 & n833 ) | ( n518 & ~n2567 ) | ( n833 & ~n2567 ) ;
  assign n2570 = n2569 ^ n2568 ^ n1736 ;
  assign n2571 = ( ~n1991 & n2564 ) | ( ~n1991 & n2570 ) | ( n2564 & n2570 ) ;
  assign n2572 = n2571 ^ n895 ^ x146 ;
  assign n2573 = n1111 ^ n1059 ^ 1'b0 ;
  assign n2574 = n2455 | n2573 ;
  assign n2575 = ( ~x141 & n1543 ) | ( ~x141 & n1986 ) | ( n1543 & n1986 ) ;
  assign n2576 = n1111 ^ n319 ^ 1'b0 ;
  assign n2577 = n1852 ^ n957 ^ x247 ;
  assign n2578 = ( x13 & n2028 ) | ( x13 & n2577 ) | ( n2028 & n2577 ) ;
  assign n2579 = x152 & n2578 ;
  assign n2580 = n1342 & n2579 ;
  assign n2581 = ( x181 & n411 ) | ( x181 & ~n1258 ) | ( n411 & ~n1258 ) ;
  assign n2582 = n2581 ^ n1448 ^ n688 ;
  assign n2583 = n1899 ^ n544 ^ n346 ;
  assign n2584 = n2583 ^ n1157 ^ 1'b0 ;
  assign n2585 = ~n2582 & n2584 ;
  assign n2586 = n1994 ^ n1117 ^ 1'b0 ;
  assign n2587 = n2586 ^ n1823 ^ n1425 ;
  assign n2593 = ( n517 & ~n530 ) | ( n517 & n859 ) | ( ~n530 & n859 ) ;
  assign n2594 = ~n2210 & n2593 ;
  assign n2592 = n1646 ^ n619 ^ n275 ;
  assign n2595 = n2594 ^ n2592 ^ n2260 ;
  assign n2588 = n601 ^ n370 ^ x132 ;
  assign n2589 = ( n368 & ~n426 ) | ( n368 & n2588 ) | ( ~n426 & n2588 ) ;
  assign n2590 = ( x157 & n532 ) | ( x157 & n1798 ) | ( n532 & n1798 ) ;
  assign n2591 = ( n388 & n2589 ) | ( n388 & n2590 ) | ( n2589 & n2590 ) ;
  assign n2596 = n2595 ^ n2591 ^ n1371 ;
  assign n2597 = ( n486 & ~n2150 ) | ( n486 & n2413 ) | ( ~n2150 & n2413 ) ;
  assign n2598 = n1496 ^ n427 ^ x212 ;
  assign n2599 = n2598 ^ n892 ^ x254 ;
  assign n2600 = ( x7 & ~n849 ) | ( x7 & n2599 ) | ( ~n849 & n2599 ) ;
  assign n2601 = n2312 & ~n2600 ;
  assign n2608 = ~x79 & n1246 ;
  assign n2609 = n2608 ^ x41 ^ 1'b0 ;
  assign n2606 = n621 ^ n308 ^ x222 ;
  assign n2605 = ( n545 & ~n992 ) | ( n545 & n1155 ) | ( ~n992 & n1155 ) ;
  assign n2602 = ( ~n710 & n797 ) | ( ~n710 & n1414 ) | ( n797 & n1414 ) ;
  assign n2603 = n2602 ^ n2179 ^ 1'b0 ;
  assign n2604 = x123 & n2603 ;
  assign n2607 = n2606 ^ n2605 ^ n2604 ;
  assign n2610 = n2609 ^ n2607 ^ n937 ;
  assign n2611 = n2610 ^ n2294 ^ 1'b0 ;
  assign n2612 = n2601 | n2611 ;
  assign n2613 = n1887 ^ n1613 ^ 1'b0 ;
  assign n2614 = x24 & n422 ;
  assign n2615 = n2614 ^ x65 ^ 1'b0 ;
  assign n2616 = n2615 ^ n877 ^ x131 ;
  assign n2617 = n2616 ^ n1495 ^ x59 ;
  assign n2618 = n2617 ^ n2108 ^ n1370 ;
  assign n2619 = n2618 ^ n1315 ^ n315 ;
  assign n2620 = n2619 ^ n2244 ^ n1700 ;
  assign n2621 = n777 | n1586 ;
  assign n2622 = x151 | n2621 ;
  assign n2623 = ( n617 & ~n766 ) | ( n617 & n2622 ) | ( ~n766 & n2622 ) ;
  assign n2624 = n2510 ^ x59 ^ 1'b0 ;
  assign n2625 = n2623 & n2624 ;
  assign n2626 = ( ~x236 & n1936 ) | ( ~x236 & n2625 ) | ( n1936 & n2625 ) ;
  assign n2629 = ( x2 & x73 ) | ( x2 & ~x122 ) | ( x73 & ~x122 ) ;
  assign n2627 = ( ~n258 & n689 ) | ( ~n258 & n997 ) | ( n689 & n997 ) ;
  assign n2628 = ( ~n1255 & n2153 ) | ( ~n1255 & n2627 ) | ( n2153 & n2627 ) ;
  assign n2630 = n2629 ^ n2628 ^ n1332 ;
  assign n2631 = x243 & ~n884 ;
  assign n2632 = ( x2 & x29 ) | ( x2 & n575 ) | ( x29 & n575 ) ;
  assign n2633 = n2632 ^ n354 ^ x190 ;
  assign n2634 = n1909 | n2633 ;
  assign n2635 = n2084 | n2634 ;
  assign n2636 = n2635 ^ n637 ^ 1'b0 ;
  assign n2637 = ( n1053 & ~n2631 ) | ( n1053 & n2636 ) | ( ~n2631 & n2636 ) ;
  assign n2638 = ( n2626 & n2630 ) | ( n2626 & n2637 ) | ( n2630 & n2637 ) ;
  assign n2639 = n1856 ^ x24 ^ 1'b0 ;
  assign n2640 = x152 & n2639 ;
  assign n2654 = ( n452 & n815 ) | ( n452 & n1310 ) | ( n815 & n1310 ) ;
  assign n2655 = n2654 ^ n1824 ^ n929 ;
  assign n2645 = x51 ^ x9 ^ 1'b0 ;
  assign n2646 = n2645 ^ n1689 ^ x214 ;
  assign n2647 = ( n342 & n2348 ) | ( n342 & ~n2646 ) | ( n2348 & ~n2646 ) ;
  assign n2648 = n1313 ^ n306 ^ 1'b0 ;
  assign n2649 = n343 | n2648 ;
  assign n2650 = n453 & n1264 ;
  assign n2651 = n2650 ^ n294 ^ 1'b0 ;
  assign n2652 = ~n2649 & n2651 ;
  assign n2653 = n2647 & n2652 ;
  assign n2641 = n1841 ^ n1530 ^ n453 ;
  assign n2642 = n1410 ^ n487 ^ 1'b0 ;
  assign n2643 = n1840 | n2642 ;
  assign n2644 = n2641 & ~n2643 ;
  assign n2656 = n2655 ^ n2653 ^ n2644 ;
  assign n2657 = x127 & x155 ;
  assign n2658 = ~x167 & n2657 ;
  assign n2659 = n2658 ^ n1945 ^ 1'b0 ;
  assign n2660 = n2659 ^ n1443 ^ x99 ;
  assign n2661 = n2660 ^ n914 ^ x174 ;
  assign n2664 = n1278 ^ n1039 ^ x144 ;
  assign n2663 = ( n1525 & n1707 ) | ( n1525 & ~n2211 ) | ( n1707 & ~n2211 ) ;
  assign n2665 = n2664 ^ n2663 ^ n1186 ;
  assign n2662 = ~x0 & n920 ;
  assign n2666 = n2665 ^ n2662 ^ n2088 ;
  assign n2667 = n1850 ^ n575 ^ x26 ;
  assign n2668 = n2667 ^ n1783 ^ n422 ;
  assign n2669 = ( ~n946 & n2383 ) | ( ~n946 & n2668 ) | ( n2383 & n2668 ) ;
  assign n2672 = ( n888 & ~n993 ) | ( n888 & n2032 ) | ( ~n993 & n2032 ) ;
  assign n2673 = n711 & n1060 ;
  assign n2674 = ~n918 & n2673 ;
  assign n2675 = x37 & ~n2674 ;
  assign n2676 = ~n2672 & n2675 ;
  assign n2670 = ( n341 & ~n1383 ) | ( n341 & n2646 ) | ( ~n1383 & n2646 ) ;
  assign n2671 = n2670 ^ n1854 ^ n526 ;
  assign n2677 = n2676 ^ n2671 ^ n359 ;
  assign n2678 = n1591 & ~n1989 ;
  assign n2679 = ~x247 & n2678 ;
  assign n2680 = n1889 & n2679 ;
  assign n2681 = ( ~n1595 & n1825 ) | ( ~n1595 & n2680 ) | ( n1825 & n2680 ) ;
  assign n2682 = n2681 ^ n2261 ^ n367 ;
  assign n2687 = n964 ^ x242 ^ 1'b0 ;
  assign n2683 = n2616 ^ n590 ^ 1'b0 ;
  assign n2684 = n857 & n2683 ;
  assign n2685 = n1828 ^ x108 ^ 1'b0 ;
  assign n2686 = n2684 & ~n2685 ;
  assign n2688 = n2687 ^ n2686 ^ n2336 ;
  assign n2692 = n1791 ^ n1434 ^ n447 ;
  assign n2693 = n2692 ^ n1077 ^ n1073 ;
  assign n2689 = ~n305 & n768 ;
  assign n2690 = ~n2336 & n2689 ;
  assign n2691 = ( x114 & n2009 ) | ( x114 & ~n2690 ) | ( n2009 & ~n2690 ) ;
  assign n2694 = n2693 ^ n2691 ^ n400 ;
  assign n2706 = n1215 ^ n1091 ^ n348 ;
  assign n2709 = ( ~x41 & x46 ) | ( ~x41 & n279 ) | ( x46 & n279 ) ;
  assign n2707 = n1074 ^ n949 ^ n368 ;
  assign n2708 = ( x55 & n881 ) | ( x55 & ~n2707 ) | ( n881 & ~n2707 ) ;
  assign n2710 = n2709 ^ n2708 ^ n518 ;
  assign n2711 = ( n2265 & ~n2706 ) | ( n2265 & n2710 ) | ( ~n2706 & n2710 ) ;
  assign n2700 = n2622 ^ n1477 ^ n923 ;
  assign n2701 = n1029 ^ n529 ^ x108 ;
  assign n2702 = n1036 | n2701 ;
  assign n2703 = n2702 ^ n1595 ^ 1'b0 ;
  assign n2704 = n2165 & ~n2703 ;
  assign n2705 = ( n2122 & n2700 ) | ( n2122 & ~n2704 ) | ( n2700 & ~n2704 ) ;
  assign n2695 = n394 & n1710 ;
  assign n2696 = n2695 ^ n982 ^ 1'b0 ;
  assign n2697 = n800 ^ n583 ^ x140 ;
  assign n2698 = n2697 ^ n669 ^ x25 ;
  assign n2699 = ( n1182 & ~n2696 ) | ( n1182 & n2698 ) | ( ~n2696 & n2698 ) ;
  assign n2712 = n2711 ^ n2705 ^ n2699 ;
  assign n2713 = n2511 ^ n1952 ^ n1899 ;
  assign n2714 = ( ~n441 & n1964 ) | ( ~n441 & n2146 ) | ( n1964 & n2146 ) ;
  assign n2715 = n922 ^ n265 ^ x115 ;
  assign n2716 = ( n406 & n2491 ) | ( n406 & n2715 ) | ( n2491 & n2715 ) ;
  assign n2719 = x179 & n1530 ;
  assign n2720 = n2719 ^ x135 ^ 1'b0 ;
  assign n2717 = n1332 & ~n1571 ;
  assign n2718 = n2717 ^ n549 ^ n409 ;
  assign n2721 = n2720 ^ n2718 ^ 1'b0 ;
  assign n2722 = ( n350 & n2716 ) | ( n350 & ~n2721 ) | ( n2716 & ~n2721 ) ;
  assign n2723 = n2089 ^ x120 ^ 1'b0 ;
  assign n2724 = n2078 ^ n1914 ^ n1130 ;
  assign n2725 = ( ~n2194 & n2556 ) | ( ~n2194 & n2724 ) | ( n2556 & n2724 ) ;
  assign n2726 = ( n380 & ~n434 ) | ( n380 & n1278 ) | ( ~n434 & n1278 ) ;
  assign n2727 = ( n281 & ~n574 ) | ( n281 & n689 ) | ( ~n574 & n689 ) ;
  assign n2728 = ( n608 & n1083 ) | ( n608 & n1139 ) | ( n1083 & n1139 ) ;
  assign n2729 = ( n1318 & n2727 ) | ( n1318 & n2728 ) | ( n2727 & n2728 ) ;
  assign n2730 = ( ~n1379 & n2726 ) | ( ~n1379 & n2729 ) | ( n2726 & n2729 ) ;
  assign n2731 = ( n2723 & n2725 ) | ( n2723 & ~n2730 ) | ( n2725 & ~n2730 ) ;
  assign n2732 = ( ~x169 & n596 ) | ( ~x169 & n661 ) | ( n596 & n661 ) ;
  assign n2733 = ( n394 & ~n874 ) | ( n394 & n2732 ) | ( ~n874 & n2732 ) ;
  assign n2734 = ( n359 & n2176 ) | ( n359 & n2733 ) | ( n2176 & n2733 ) ;
  assign n2735 = n2539 ^ n1057 ^ 1'b0 ;
  assign n2736 = n1703 & n2735 ;
  assign n2737 = ~n2348 & n2736 ;
  assign n2738 = n2737 ^ n968 ^ x202 ;
  assign n2739 = ~n2734 & n2738 ;
  assign n2740 = ~n2431 & n2739 ;
  assign n2741 = n453 & n2740 ;
  assign n2742 = n2349 ^ n1018 ^ 1'b0 ;
  assign n2743 = n983 | n2742 ;
  assign n2744 = n2743 ^ n1558 ^ 1'b0 ;
  assign n2745 = x7 & ~n2156 ;
  assign n2746 = ~n2026 & n2745 ;
  assign n2747 = ( n831 & ~n957 ) | ( n831 & n2746 ) | ( ~n957 & n2746 ) ;
  assign n2757 = n532 | n1021 ;
  assign n2758 = n2757 ^ n1617 ^ n838 ;
  assign n2752 = x207 | n794 ;
  assign n2749 = n2317 ^ n788 ^ 1'b0 ;
  assign n2750 = x64 & n2749 ;
  assign n2748 = x48 & n696 ;
  assign n2751 = n2750 ^ n2748 ^ 1'b0 ;
  assign n2753 = n2752 ^ n2751 ^ n2701 ;
  assign n2754 = x218 & ~n1383 ;
  assign n2755 = n2753 & n2754 ;
  assign n2756 = n2755 ^ n2375 ^ n380 ;
  assign n2759 = n2758 ^ n2756 ^ n2414 ;
  assign n2760 = n1007 & ~n1618 ;
  assign n2761 = n890 & n1886 ;
  assign n2762 = ~n2760 & n2761 ;
  assign n2763 = ( ~n387 & n2759 ) | ( ~n387 & n2762 ) | ( n2759 & n2762 ) ;
  assign n2770 = n373 ^ x96 ^ x24 ;
  assign n2771 = ~n541 & n1144 ;
  assign n2772 = n2770 & n2771 ;
  assign n2773 = n2772 ^ n1461 ^ n1430 ;
  assign n2767 = n1065 ^ n637 ^ 1'b0 ;
  assign n2768 = n1356 & ~n2767 ;
  assign n2764 = n1133 & ~n2507 ;
  assign n2765 = ( x176 & ~n1644 ) | ( x176 & n2564 ) | ( ~n1644 & n2564 ) ;
  assign n2766 = ( x31 & n2764 ) | ( x31 & ~n2765 ) | ( n2764 & ~n2765 ) ;
  assign n2769 = n2768 ^ n2766 ^ 1'b0 ;
  assign n2774 = n2773 ^ n2769 ^ 1'b0 ;
  assign n2775 = ( n736 & n1241 ) | ( n736 & n1478 ) | ( n1241 & n1478 ) ;
  assign n2776 = ( n1557 & n1665 ) | ( n1557 & ~n2775 ) | ( n1665 & ~n2775 ) ;
  assign n2777 = ~n2490 & n2628 ;
  assign n2778 = n2776 & ~n2777 ;
  assign n2779 = n2778 ^ n1533 ^ 1'b0 ;
  assign n2780 = ( x215 & ~n2760 ) | ( x215 & n2779 ) | ( ~n2760 & n2779 ) ;
  assign n2783 = n1282 ^ x189 ^ 1'b0 ;
  assign n2781 = n876 & ~n1928 ;
  assign n2782 = n2781 ^ n706 ^ 1'b0 ;
  assign n2784 = n2783 ^ n2782 ^ n2220 ;
  assign n2785 = n459 ^ x129 ^ 1'b0 ;
  assign n2786 = n2164 | n2785 ;
  assign n2787 = n2773 ^ n2510 ^ n1025 ;
  assign n2788 = n1060 & n2787 ;
  assign n2789 = n2786 & n2788 ;
  assign n2799 = n956 ^ n760 ^ n295 ;
  assign n2800 = n2799 ^ x126 ^ 1'b0 ;
  assign n2795 = n585 ^ x232 ^ x117 ;
  assign n2796 = n600 & n959 ;
  assign n2797 = ~n2795 & n2796 ;
  assign n2798 = n877 & ~n2797 ;
  assign n2801 = n2800 ^ n2798 ^ 1'b0 ;
  assign n2793 = n403 & n797 ;
  assign n2794 = n2793 ^ x192 ^ 1'b0 ;
  assign n2802 = n2801 ^ n2794 ^ n1316 ;
  assign n2790 = ( n307 & n805 ) | ( n307 & n1850 ) | ( n805 & n1850 ) ;
  assign n2791 = n2636 & n2790 ;
  assign n2792 = n855 | n2791 ;
  assign n2803 = n2802 ^ n2792 ^ 1'b0 ;
  assign n2804 = n2056 ^ n594 ^ 1'b0 ;
  assign n2805 = ( n304 & n2800 ) | ( n304 & n2804 ) | ( n2800 & n2804 ) ;
  assign n2806 = n1248 & ~n2805 ;
  assign n2807 = ( n2789 & n2803 ) | ( n2789 & n2806 ) | ( n2803 & n2806 ) ;
  assign n2809 = ( x148 & n999 ) | ( x148 & ~n1568 ) | ( n999 & ~n1568 ) ;
  assign n2808 = ( n1204 & n1893 ) | ( n1204 & ~n1942 ) | ( n1893 & ~n1942 ) ;
  assign n2810 = n2809 ^ n2808 ^ n1639 ;
  assign n2811 = n2807 & n2810 ;
  assign n2822 = n1849 ^ n1224 ^ 1'b0 ;
  assign n2823 = n373 & n2822 ;
  assign n2821 = n771 ^ n705 ^ n395 ;
  assign n2818 = n593 ^ n406 ^ x213 ;
  assign n2819 = n1360 ^ n1024 ^ n377 ;
  assign n2820 = ( x62 & n2818 ) | ( x62 & ~n2819 ) | ( n2818 & ~n2819 ) ;
  assign n2824 = n2823 ^ n2821 ^ n2820 ;
  assign n2817 = x38 & ~n2372 ;
  assign n2825 = n2824 ^ n2817 ^ 1'b0 ;
  assign n2812 = ( n626 & ~n1069 ) | ( n626 & n1848 ) | ( ~n1069 & n1848 ) ;
  assign n2814 = ( ~n602 & n811 ) | ( ~n602 & n1631 ) | ( n811 & n1631 ) ;
  assign n2813 = n1445 & n2087 ;
  assign n2815 = n2814 ^ n2813 ^ 1'b0 ;
  assign n2816 = ( n966 & n2812 ) | ( n966 & n2815 ) | ( n2812 & n2815 ) ;
  assign n2826 = n2825 ^ n2816 ^ n2447 ;
  assign n2828 = ( n431 & n724 ) | ( n431 & ~n939 ) | ( n724 & ~n939 ) ;
  assign n2829 = ( n319 & ~n371 ) | ( n319 & n1365 ) | ( ~n371 & n1365 ) ;
  assign n2830 = ( n2804 & n2828 ) | ( n2804 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = n2830 ^ n1961 ^ 1'b0 ;
  assign n2827 = ( x14 & ~n1397 ) | ( x14 & n1760 ) | ( ~n1397 & n1760 ) ;
  assign n2832 = n2831 ^ n2827 ^ n1382 ;
  assign n2833 = ( ~n800 & n1645 ) | ( ~n800 & n1978 ) | ( n1645 & n1978 ) ;
  assign n2884 = n953 ^ x251 ^ 1'b0 ;
  assign n2885 = ( ~x236 & n2087 ) | ( ~x236 & n2884 ) | ( n2087 & n2884 ) ;
  assign n2881 = n641 & n2350 ;
  assign n2882 = ( ~n640 & n1140 ) | ( ~n640 & n2881 ) | ( n1140 & n2881 ) ;
  assign n2883 = n2882 ^ n1533 ^ n1144 ;
  assign n2886 = n2885 ^ n2883 ^ x175 ;
  assign n2869 = ( n356 & n495 ) | ( n356 & ~n822 ) | ( n495 & ~n822 ) ;
  assign n2870 = n2727 ^ n1755 ^ n1220 ;
  assign n2871 = ( n299 & ~n2869 ) | ( n299 & n2870 ) | ( ~n2869 & n2870 ) ;
  assign n2872 = x67 & ~n2871 ;
  assign n2873 = n2872 ^ n672 ^ 1'b0 ;
  assign n2875 = ( ~x118 & n407 ) | ( ~x118 & n455 ) | ( n407 & n455 ) ;
  assign n2876 = ( n521 & n1241 ) | ( n521 & ~n2875 ) | ( n1241 & ~n2875 ) ;
  assign n2877 = n2876 ^ n1463 ^ n1279 ;
  assign n2874 = ( x111 & ~n1199 ) | ( x111 & n1454 ) | ( ~n1199 & n1454 ) ;
  assign n2878 = n2877 ^ n2874 ^ n810 ;
  assign n2879 = n2873 & ~n2878 ;
  assign n2867 = ( x150 & n426 ) | ( x150 & n1359 ) | ( n426 & n1359 ) ;
  assign n2862 = n1056 & n1970 ;
  assign n2863 = n2432 ^ n2082 ^ n889 ;
  assign n2864 = ( ~n970 & n2862 ) | ( ~n970 & n2863 ) | ( n2862 & n2863 ) ;
  assign n2865 = n2864 ^ n1285 ^ n876 ;
  assign n2866 = n842 | n2865 ;
  assign n2868 = n2867 ^ n2866 ^ 1'b0 ;
  assign n2880 = n2879 ^ n2868 ^ n790 ;
  assign n2834 = ( n815 & ~n1381 ) | ( n815 & n2617 ) | ( ~n1381 & n2617 ) ;
  assign n2835 = ( n359 & n642 ) | ( n359 & n2834 ) | ( n642 & n2834 ) ;
  assign n2836 = ~n828 & n2835 ;
  assign n2856 = ( x87 & ~n1242 ) | ( x87 & n1336 ) | ( ~n1242 & n1336 ) ;
  assign n2857 = n2856 ^ n748 ^ x181 ;
  assign n2858 = ( ~x250 & n1980 ) | ( ~x250 & n2857 ) | ( n1980 & n2857 ) ;
  assign n2859 = n2858 ^ x39 ^ 1'b0 ;
  assign n2854 = n928 ^ n874 ^ x12 ;
  assign n2855 = n2237 & ~n2854 ;
  assign n2837 = n853 & ~n2388 ;
  assign n2838 = n2837 ^ n1173 ^ 1'b0 ;
  assign n2847 = x15 & ~n639 ;
  assign n2848 = ~n1305 & n2847 ;
  assign n2846 = ( n544 & n629 ) | ( n544 & ~n855 ) | ( n629 & ~n855 ) ;
  assign n2849 = n2848 ^ n2846 ^ x90 ;
  assign n2844 = ( ~x60 & x84 ) | ( ~x60 & n1170 ) | ( x84 & n1170 ) ;
  assign n2845 = n2844 ^ n1006 ^ n947 ;
  assign n2850 = n2849 ^ n2845 ^ 1'b0 ;
  assign n2851 = n2850 ^ n1675 ^ n1039 ;
  assign n2839 = ( ~x25 & n362 ) | ( ~x25 & n1279 ) | ( n362 & n1279 ) ;
  assign n2840 = ( n295 & n1320 ) | ( n295 & n2839 ) | ( n1320 & n2839 ) ;
  assign n2841 = n1047 ^ n910 ^ n601 ;
  assign n2842 = n2841 ^ n321 ^ x163 ;
  assign n2843 = ( ~n1883 & n2840 ) | ( ~n1883 & n2842 ) | ( n2840 & n2842 ) ;
  assign n2852 = n2851 ^ n2843 ^ x118 ;
  assign n2853 = ( n747 & ~n2838 ) | ( n747 & n2852 ) | ( ~n2838 & n2852 ) ;
  assign n2860 = n2859 ^ n2855 ^ n2853 ;
  assign n2861 = ( n1282 & ~n2836 ) | ( n1282 & n2860 ) | ( ~n2836 & n2860 ) ;
  assign n2887 = n2886 ^ n2880 ^ n2861 ;
  assign n2888 = n2887 ^ n876 ^ 1'b0 ;
  assign n2889 = ~n1042 & n2888 ;
  assign n2890 = n539 & ~n1032 ;
  assign n2891 = n2890 ^ n1255 ^ 1'b0 ;
  assign n2892 = n2638 ^ n874 ^ 1'b0 ;
  assign n2895 = n2275 ^ n1161 ^ 1'b0 ;
  assign n2893 = n537 & ~n788 ;
  assign n2894 = n2893 ^ n1508 ^ 1'b0 ;
  assign n2896 = n2895 ^ n2894 ^ x153 ;
  assign n2897 = n2868 ^ n466 ^ n448 ;
  assign n2898 = ( n854 & ~n1389 ) | ( n854 & n2897 ) | ( ~n1389 & n2897 ) ;
  assign n2901 = ( x98 & ~n613 ) | ( x98 & n1393 ) | ( ~n613 & n1393 ) ;
  assign n2899 = n2509 ^ x236 ^ x174 ;
  assign n2900 = ~n2175 & n2899 ;
  assign n2902 = n2901 ^ n2900 ^ n2509 ;
  assign n2903 = n2632 ^ n1946 ^ n824 ;
  assign n2904 = n1763 ^ n623 ^ x210 ;
  assign n2905 = ( n885 & ~n2192 ) | ( n885 & n2904 ) | ( ~n2192 & n2904 ) ;
  assign n2906 = ( n2879 & n2903 ) | ( n2879 & n2905 ) | ( n2903 & n2905 ) ;
  assign n2907 = n1117 ^ n772 ^ x170 ;
  assign n2908 = x157 & ~n2907 ;
  assign n2909 = n2908 ^ n1760 ^ 1'b0 ;
  assign n2910 = ( n1753 & n2906 ) | ( n1753 & ~n2909 ) | ( n2906 & ~n2909 ) ;
  assign n2911 = ( n318 & n626 ) | ( n318 & ~n2910 ) | ( n626 & ~n2910 ) ;
  assign n2912 = ( x78 & n436 ) | ( x78 & n857 ) | ( n436 & n857 ) ;
  assign n2913 = n980 & n2101 ;
  assign n2914 = ~n276 & n2913 ;
  assign n2916 = ( n965 & ~n1780 ) | ( n965 & n2076 ) | ( ~n1780 & n2076 ) ;
  assign n2917 = n2916 ^ n2716 ^ n1254 ;
  assign n2915 = ~n1143 & n1451 ;
  assign n2918 = n2917 ^ n2915 ^ 1'b0 ;
  assign n2919 = ( n2912 & n2914 ) | ( n2912 & n2918 ) | ( n2914 & n2918 ) ;
  assign n2920 = ( ~n658 & n1221 ) | ( ~n658 & n1669 ) | ( n1221 & n1669 ) ;
  assign n2921 = ( n655 & n1807 ) | ( n655 & ~n1970 ) | ( n1807 & ~n1970 ) ;
  assign n2922 = ( ~n1705 & n1963 ) | ( ~n1705 & n2134 ) | ( n1963 & n2134 ) ;
  assign n2923 = ( x35 & n2921 ) | ( x35 & ~n2922 ) | ( n2921 & ~n2922 ) ;
  assign n2924 = n1656 ^ n1399 ^ 1'b0 ;
  assign n2925 = n1447 & ~n2924 ;
  assign n2926 = ( ~n852 & n2923 ) | ( ~n852 & n2925 ) | ( n2923 & n2925 ) ;
  assign n2927 = ( n2919 & n2920 ) | ( n2919 & ~n2926 ) | ( n2920 & ~n2926 ) ;
  assign n2929 = n845 ^ n633 ^ 1'b0 ;
  assign n2930 = ( x38 & n2041 ) | ( x38 & ~n2929 ) | ( n2041 & ~n2929 ) ;
  assign n2928 = n2710 ^ n1755 ^ n1451 ;
  assign n2931 = n2930 ^ n2928 ^ n1438 ;
  assign n2932 = n2931 ^ n2776 ^ n2760 ;
  assign n2947 = n1922 ^ n1532 ^ 1'b0 ;
  assign n2943 = n2350 ^ n1781 ^ 1'b0 ;
  assign n2944 = n2943 ^ n2808 ^ 1'b0 ;
  assign n2945 = ~n1106 & n2944 ;
  assign n2946 = n2945 ^ n1916 ^ n963 ;
  assign n2933 = ( ~n545 & n2066 ) | ( ~n545 & n2629 ) | ( n2066 & n2629 ) ;
  assign n2937 = ( n379 & n2382 ) | ( n379 & ~n2445 ) | ( n2382 & ~n2445 ) ;
  assign n2938 = ( x244 & n341 ) | ( x244 & ~n2937 ) | ( n341 & ~n2937 ) ;
  assign n2935 = n2089 ^ n1113 ^ n403 ;
  assign n2936 = ( n326 & n800 ) | ( n326 & n2935 ) | ( n800 & n2935 ) ;
  assign n2934 = ( x212 & n670 ) | ( x212 & ~n2084 ) | ( n670 & ~n2084 ) ;
  assign n2939 = n2938 ^ n2936 ^ n2934 ;
  assign n2940 = ( n926 & n1369 ) | ( n926 & n2939 ) | ( n1369 & n2939 ) ;
  assign n2941 = n1567 & ~n2940 ;
  assign n2942 = ~n2933 & n2941 ;
  assign n2948 = n2947 ^ n2946 ^ n2942 ;
  assign n2970 = ( ~n377 & n1001 ) | ( ~n377 & n1008 ) | ( n1001 & n1008 ) ;
  assign n2969 = ~n830 & n934 ;
  assign n2971 = n2970 ^ n2969 ^ 1'b0 ;
  assign n2967 = n2309 ^ n1084 ^ n530 ;
  assign n2968 = ( n1752 & n2273 ) | ( n1752 & n2967 ) | ( n2273 & n2967 ) ;
  assign n2949 = ( x33 & n760 ) | ( x33 & n1585 ) | ( n760 & n1585 ) ;
  assign n2950 = ( x218 & n1863 ) | ( x218 & n2949 ) | ( n1863 & n2949 ) ;
  assign n2951 = n2582 | n2950 ;
  assign n2964 = n1644 ^ n996 ^ x11 ;
  assign n2952 = n340 ^ x141 ^ 1'b0 ;
  assign n2953 = x77 | n2294 ;
  assign n2954 = n2953 ^ n1680 ^ n1647 ;
  assign n2955 = x116 & ~n1036 ;
  assign n2956 = ~x115 & n2955 ;
  assign n2957 = n2956 ^ n1392 ^ n614 ;
  assign n2958 = n2957 ^ n1587 ^ 1'b0 ;
  assign n2959 = x56 & ~n2958 ;
  assign n2960 = ( x246 & ~n1574 ) | ( x246 & n2959 ) | ( ~n1574 & n2959 ) ;
  assign n2961 = x138 & n2665 ;
  assign n2962 = ~n2960 & n2961 ;
  assign n2963 = ( ~n2952 & n2954 ) | ( ~n2952 & n2962 ) | ( n2954 & n2962 ) ;
  assign n2965 = n2964 ^ n2963 ^ 1'b0 ;
  assign n2966 = n2951 & n2965 ;
  assign n2972 = n2971 ^ n2968 ^ n2966 ;
  assign n2981 = n1027 ^ n443 ^ n331 ;
  assign n2979 = n682 ^ n482 ^ n271 ;
  assign n2975 = n749 ^ n728 ^ x231 ;
  assign n2978 = n2975 ^ n2775 ^ n827 ;
  assign n2976 = ( n526 & n685 ) | ( n526 & n2975 ) | ( n685 & n2975 ) ;
  assign n2977 = n2976 ^ n2430 ^ n710 ;
  assign n2980 = n2979 ^ n2978 ^ n2977 ;
  assign n2982 = n2981 ^ n2980 ^ n2227 ;
  assign n2973 = ( ~n1514 & n1781 ) | ( ~n1514 & n2227 ) | ( n1781 & n2227 ) ;
  assign n2974 = ~n1515 & n2973 ;
  assign n2983 = n2982 ^ n2974 ^ n2137 ;
  assign n2984 = n820 ^ n651 ^ x112 ;
  assign n2985 = n2984 ^ n2768 ^ n951 ;
  assign n2986 = n2870 ^ n1061 ^ 1'b0 ;
  assign n2987 = n2985 & ~n2986 ;
  assign n2988 = n1887 ^ n1455 ^ n1065 ;
  assign n2989 = n2987 & n2988 ;
  assign n2990 = n2989 ^ n1141 ^ 1'b0 ;
  assign n2991 = ~n494 & n2990 ;
  assign n2992 = ( ~n2114 & n2983 ) | ( ~n2114 & n2991 ) | ( n2983 & n2991 ) ;
  assign n2993 = n1598 ^ n1383 ^ x122 ;
  assign n2994 = n1532 ^ n486 ^ 1'b0 ;
  assign n2995 = n566 | n1139 ;
  assign n2996 = x236 | n2995 ;
  assign n2997 = n892 ^ n581 ^ 1'b0 ;
  assign n2998 = n621 | n2997 ;
  assign n2999 = n2998 ^ n798 ^ 1'b0 ;
  assign n3000 = n987 | n2999 ;
  assign n3001 = n2996 & n3000 ;
  assign n3002 = ( n1812 & n2994 ) | ( n1812 & n3001 ) | ( n2994 & n3001 ) ;
  assign n3003 = ( n1667 & n2993 ) | ( n1667 & ~n3002 ) | ( n2993 & ~n3002 ) ;
  assign n3004 = n1396 ^ n1083 ^ n260 ;
  assign n3005 = ( x237 & ~n2538 ) | ( x237 & n3004 ) | ( ~n2538 & n3004 ) ;
  assign n3006 = n1946 ^ n1476 ^ n1337 ;
  assign n3007 = n3006 ^ n2210 ^ n1168 ;
  assign n3008 = n3007 ^ n1595 ^ x90 ;
  assign n3009 = n2056 & n3008 ;
  assign n3010 = n3009 ^ n2901 ^ 1'b0 ;
  assign n3011 = n3010 ^ n2987 ^ n480 ;
  assign n3028 = n1814 ^ n1435 ^ n485 ;
  assign n3027 = n923 ^ n884 ^ n413 ;
  assign n3029 = n3028 ^ n3027 ^ n996 ;
  assign n3030 = n720 ^ n572 ^ 1'b0 ;
  assign n3031 = n2867 & n3030 ;
  assign n3032 = n270 & n3031 ;
  assign n3033 = n3029 & n3032 ;
  assign n3034 = n3033 ^ n2864 ^ n1156 ;
  assign n3023 = x167 ^ x79 ^ 1'b0 ;
  assign n3024 = x106 & n3023 ;
  assign n3025 = ~n742 & n3024 ;
  assign n3021 = n587 | n1243 ;
  assign n3022 = ( n270 & n842 ) | ( n270 & ~n3021 ) | ( n842 & ~n3021 ) ;
  assign n3016 = n890 | n1031 ;
  assign n3017 = n1033 & ~n3016 ;
  assign n3018 = n3017 ^ n1451 ^ 1'b0 ;
  assign n3019 = ( n1253 & ~n2015 ) | ( n1253 & n3018 ) | ( ~n2015 & n3018 ) ;
  assign n3020 = ( n1074 & n1806 ) | ( n1074 & n3019 ) | ( n1806 & n3019 ) ;
  assign n3026 = n3025 ^ n3022 ^ n3020 ;
  assign n3014 = n579 | n1860 ;
  assign n3012 = ( ~n319 & n926 ) | ( ~n319 & n1363 ) | ( n926 & n1363 ) ;
  assign n3013 = ( x197 & ~n272 ) | ( x197 & n3012 ) | ( ~n272 & n3012 ) ;
  assign n3015 = n3014 ^ n3013 ^ n1552 ;
  assign n3035 = n3034 ^ n3026 ^ n3015 ;
  assign n3041 = n505 & n2241 ;
  assign n3042 = n1523 ^ n1195 ^ n345 ;
  assign n3043 = ~n3041 & n3042 ;
  assign n3044 = n3043 ^ n811 ^ 1'b0 ;
  assign n3036 = n1381 ^ x167 ^ 1'b0 ;
  assign n3037 = x67 & n3036 ;
  assign n3038 = n3037 ^ n1907 ^ 1'b0 ;
  assign n3039 = n1005 & ~n3038 ;
  assign n3040 = n3039 ^ x90 ^ 1'b0 ;
  assign n3045 = n3044 ^ n3040 ^ 1'b0 ;
  assign n3047 = ( n579 & ~n594 ) | ( n579 & n1120 ) | ( ~n594 & n1120 ) ;
  assign n3048 = n3047 ^ x218 ^ 1'b0 ;
  assign n3046 = ~n579 & n2856 ;
  assign n3049 = n3048 ^ n3046 ^ 1'b0 ;
  assign n3050 = n620 ^ x81 ^ 1'b0 ;
  assign n3051 = n3050 ^ n2488 ^ n1079 ;
  assign n3054 = n2768 ^ x38 ^ 1'b0 ;
  assign n3055 = n3054 ^ n2812 ^ 1'b0 ;
  assign n3052 = ( n280 & ~n898 ) | ( n280 & n1730 ) | ( ~n898 & n1730 ) ;
  assign n3053 = ( n345 & n977 ) | ( n345 & n3052 ) | ( n977 & n3052 ) ;
  assign n3056 = n3055 ^ n3053 ^ n2387 ;
  assign n3077 = ( n966 & n2383 ) | ( n966 & n2510 ) | ( n2383 & n2510 ) ;
  assign n3078 = n1746 & n3077 ;
  assign n3066 = n804 ^ n451 ^ n283 ;
  assign n3067 = n597 ^ n553 ^ 1'b0 ;
  assign n3068 = n1585 & n3067 ;
  assign n3069 = ~x174 & n3068 ;
  assign n3072 = n1168 ^ n345 ^ x4 ;
  assign n3070 = ~n1157 & n2323 ;
  assign n3071 = n3070 ^ n1263 ^ 1'b0 ;
  assign n3073 = n3072 ^ n3071 ^ n1133 ;
  assign n3074 = ( n465 & n3069 ) | ( n465 & n3073 ) | ( n3069 & n3073 ) ;
  assign n3075 = ( ~n1406 & n3066 ) | ( ~n1406 & n3074 ) | ( n3066 & n3074 ) ;
  assign n3076 = n3075 ^ n2844 ^ x201 ;
  assign n3079 = n3078 ^ n3076 ^ x183 ;
  assign n3057 = ~n284 & n676 ;
  assign n3058 = ( n472 & ~n606 ) | ( n472 & n3057 ) | ( ~n606 & n3057 ) ;
  assign n3059 = n452 & n1161 ;
  assign n3060 = n3059 ^ x121 ^ 1'b0 ;
  assign n3061 = n1507 ^ x230 ^ 1'b0 ;
  assign n3062 = n3061 ^ n2838 ^ 1'b0 ;
  assign n3063 = n2766 & ~n3062 ;
  assign n3064 = ( n997 & n3060 ) | ( n997 & ~n3063 ) | ( n3060 & ~n3063 ) ;
  assign n3065 = ( ~n1743 & n3058 ) | ( ~n1743 & n3064 ) | ( n3058 & n3064 ) ;
  assign n3080 = n3079 ^ n3065 ^ x125 ;
  assign n3081 = x195 & n743 ;
  assign n3082 = ~n1149 & n3081 ;
  assign n3083 = n3077 ^ n335 ^ 1'b0 ;
  assign n3084 = n3083 ^ n3028 ^ n1107 ;
  assign n3085 = n3082 & n3084 ;
  assign n3086 = n2607 ^ n1199 ^ n559 ;
  assign n3087 = n2975 ^ n2790 ^ x162 ;
  assign n3088 = ( ~n659 & n845 ) | ( ~n659 & n3087 ) | ( n845 & n3087 ) ;
  assign n3089 = n2801 | n3088 ;
  assign n3090 = ( ~n2265 & n2565 ) | ( ~n2265 & n3089 ) | ( n2565 & n3089 ) ;
  assign n3091 = x16 & x165 ;
  assign n3092 = n3091 ^ n522 ^ 1'b0 ;
  assign n3093 = ( n1123 & n1379 ) | ( n1123 & ~n3092 ) | ( n1379 & ~n3092 ) ;
  assign n3094 = ( n1751 & n2630 ) | ( n1751 & n3093 ) | ( n2630 & n3093 ) ;
  assign n3095 = ( n392 & n2339 ) | ( n392 & n3094 ) | ( n2339 & n3094 ) ;
  assign n3096 = n1374 ^ n1298 ^ n479 ;
  assign n3097 = ( n1304 & ~n1481 ) | ( n1304 & n2093 ) | ( ~n1481 & n2093 ) ;
  assign n3098 = ( ~n1279 & n2617 ) | ( ~n1279 & n3097 ) | ( n2617 & n3097 ) ;
  assign n3099 = n1769 | n3098 ;
  assign n3100 = n3099 ^ n2676 ^ 1'b0 ;
  assign n3101 = n296 & ~n2009 ;
  assign n3102 = n3100 & n3101 ;
  assign n3103 = n3096 | n3102 ;
  assign n3104 = n1405 ^ n745 ^ n362 ;
  assign n3105 = n3104 ^ n874 ^ x125 ;
  assign n3106 = n3105 ^ n2317 ^ n374 ;
  assign n3107 = n3106 ^ n1164 ^ 1'b0 ;
  assign n3108 = n2862 ^ n2048 ^ n898 ;
  assign n3109 = ( n778 & n1042 ) | ( n778 & ~n1849 ) | ( n1042 & ~n1849 ) ;
  assign n3110 = ( n2663 & ~n2906 ) | ( n2663 & n3109 ) | ( ~n2906 & n3109 ) ;
  assign n3111 = n2209 ^ n964 ^ n625 ;
  assign n3112 = x119 | n1595 ;
  assign n3113 = n3112 ^ n2681 ^ n1595 ;
  assign n3117 = n2153 ^ n1231 ^ n1143 ;
  assign n3118 = n3117 ^ n1278 ^ n514 ;
  assign n3115 = n1753 ^ n683 ^ n544 ;
  assign n3114 = n957 ^ n313 ^ x114 ;
  assign n3116 = n3115 ^ n3114 ^ n812 ;
  assign n3119 = n3118 ^ n3116 ^ n3026 ;
  assign n3120 = ( x13 & n408 ) | ( x13 & ~n2211 ) | ( n408 & ~n2211 ) ;
  assign n3121 = x128 & ~n3120 ;
  assign n3122 = n3121 ^ n1534 ^ 1'b0 ;
  assign n3123 = n2483 ^ n500 ^ x201 ;
  assign n3124 = ~n1551 & n2886 ;
  assign n3125 = n1344 ^ n1211 ^ 1'b0 ;
  assign n3126 = n727 & n3125 ;
  assign n3127 = ( n3123 & n3124 ) | ( n3123 & n3126 ) | ( n3124 & n3126 ) ;
  assign n3128 = ~n981 & n3127 ;
  assign n3141 = n1865 ^ n1591 ^ n1527 ;
  assign n3142 = ( n1107 & n1220 ) | ( n1107 & n3141 ) | ( n1220 & n3141 ) ;
  assign n3143 = n2293 ^ n972 ^ 1'b0 ;
  assign n3144 = ( x34 & n3142 ) | ( x34 & ~n3143 ) | ( n3142 & ~n3143 ) ;
  assign n3129 = n2383 ^ n778 ^ n740 ;
  assign n3130 = ( ~x217 & n648 ) | ( ~x217 & n3129 ) | ( n648 & n3129 ) ;
  assign n3131 = ( ~x93 & n384 ) | ( ~x93 & n2952 ) | ( n384 & n2952 ) ;
  assign n3132 = n3131 ^ x19 ^ 1'b0 ;
  assign n3133 = ~n1868 & n3132 ;
  assign n3134 = ( n1649 & n3130 ) | ( n1649 & ~n3133 ) | ( n3130 & ~n3133 ) ;
  assign n3135 = n1252 | n3134 ;
  assign n3136 = n2527 | n3135 ;
  assign n3137 = ( ~n297 & n363 ) | ( ~n297 & n1928 ) | ( n363 & n1928 ) ;
  assign n3138 = n3137 ^ n2867 ^ n1875 ;
  assign n3139 = n3138 ^ n2897 ^ n359 ;
  assign n3140 = n3136 & ~n3139 ;
  assign n3145 = n3144 ^ n3140 ^ 1'b0 ;
  assign n3146 = ( ~n579 & n826 ) | ( ~n579 & n2395 ) | ( n826 & n2395 ) ;
  assign n3147 = ( ~n704 & n1619 ) | ( ~n704 & n3146 ) | ( n1619 & n3146 ) ;
  assign n3148 = ( x154 & n473 ) | ( x154 & ~n3147 ) | ( n473 & ~n3147 ) ;
  assign n3158 = ~n997 & n2352 ;
  assign n3149 = n897 ^ n629 ^ n263 ;
  assign n3150 = ~n1071 & n1612 ;
  assign n3151 = ( x154 & n3149 ) | ( x154 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3153 = ( x223 & n1408 ) | ( x223 & n2093 ) | ( n1408 & n2093 ) ;
  assign n3154 = ( x181 & n849 ) | ( x181 & n2217 ) | ( n849 & n2217 ) ;
  assign n3155 = ( n1048 & n3153 ) | ( n1048 & n3154 ) | ( n3153 & n3154 ) ;
  assign n3152 = n1724 ^ n1533 ^ n582 ;
  assign n3156 = n3155 ^ n3152 ^ 1'b0 ;
  assign n3157 = n3151 & ~n3156 ;
  assign n3159 = n3158 ^ n3157 ^ n2982 ;
  assign n3160 = ( ~n1616 & n2107 ) | ( ~n1616 & n2680 ) | ( n2107 & n2680 ) ;
  assign n3161 = n2327 | n3160 ;
  assign n3162 = n3159 & ~n3161 ;
  assign n3163 = ( n2005 & n2605 ) | ( n2005 & n2857 ) | ( n2605 & n2857 ) ;
  assign n3164 = x239 & ~n1840 ;
  assign n3165 = ~n3163 & n3164 ;
  assign n3166 = n1482 ^ n571 ^ 1'b0 ;
  assign n3167 = ( n2733 & n2949 ) | ( n2733 & ~n3166 ) | ( n2949 & ~n3166 ) ;
  assign n3171 = n350 & n1226 ;
  assign n3172 = n3171 ^ n1852 ^ 1'b0 ;
  assign n3168 = n1149 ^ n611 ^ x5 ;
  assign n3169 = ( x198 & ~n852 ) | ( x198 & n3168 ) | ( ~n852 & n3168 ) ;
  assign n3170 = n3169 ^ n770 ^ x210 ;
  assign n3173 = n3172 ^ n3170 ^ n1503 ;
  assign n3191 = n1573 ^ n552 ^ 1'b0 ;
  assign n3188 = n931 ^ x213 ^ x17 ;
  assign n3189 = n3188 ^ n2542 ^ 1'b0 ;
  assign n3190 = n3189 ^ n1144 ^ n696 ;
  assign n3174 = n2250 ^ x34 ^ 1'b0 ;
  assign n3185 = n3129 ^ n2609 ^ 1'b0 ;
  assign n3175 = n1019 ^ n259 ^ 1'b0 ;
  assign n3176 = n2520 & n3175 ;
  assign n3177 = ( ~n1189 & n3041 ) | ( ~n1189 & n3176 ) | ( n3041 & n3176 ) ;
  assign n3178 = ~n1558 & n1667 ;
  assign n3179 = n2058 | n3088 ;
  assign n3180 = n3178 & ~n3179 ;
  assign n3181 = n1810 ^ n778 ^ n368 ;
  assign n3182 = n3181 ^ n2504 ^ 1'b0 ;
  assign n3183 = ( ~n3177 & n3180 ) | ( ~n3177 & n3182 ) | ( n3180 & n3182 ) ;
  assign n3184 = n1012 | n3183 ;
  assign n3186 = n3185 ^ n3184 ^ 1'b0 ;
  assign n3187 = n3174 | n3186 ;
  assign n3192 = n3191 ^ n3190 ^ n3187 ;
  assign n3193 = n2081 ^ n767 ^ x172 ;
  assign n3194 = n3193 ^ n849 ^ 1'b0 ;
  assign n3195 = n3174 ^ n1993 ^ n334 ;
  assign n3196 = n3028 ^ n1246 ^ n954 ;
  assign n3197 = ( ~n1155 & n1261 ) | ( ~n1155 & n3196 ) | ( n1261 & n3196 ) ;
  assign n3198 = n590 & n607 ;
  assign n3199 = n733 & n3198 ;
  assign n3207 = n1312 ^ x6 ^ 1'b0 ;
  assign n3205 = ( x33 & n1220 ) | ( x33 & n1405 ) | ( n1220 & n1405 ) ;
  assign n3200 = n1112 ^ n1019 ^ x23 ;
  assign n3201 = x197 & ~n665 ;
  assign n3202 = n766 & n3201 ;
  assign n3203 = n3202 ^ n1631 ^ x242 ;
  assign n3204 = ( n1508 & n3200 ) | ( n1508 & n3203 ) | ( n3200 & n3203 ) ;
  assign n3206 = n3205 ^ n3204 ^ n894 ;
  assign n3208 = n3207 ^ n3206 ^ n455 ;
  assign n3209 = n2096 ^ n1618 ^ n1156 ;
  assign n3210 = n3209 ^ n2942 ^ n1677 ;
  assign n3211 = ( n760 & ~n1716 ) | ( n760 & n2027 ) | ( ~n1716 & n2027 ) ;
  assign n3212 = ( x105 & ~n401 ) | ( x105 & n531 ) | ( ~n401 & n531 ) ;
  assign n3213 = ( n525 & ~n2241 ) | ( n525 & n3212 ) | ( ~n2241 & n3212 ) ;
  assign n3214 = ( n821 & ~n1986 ) | ( n821 & n3213 ) | ( ~n1986 & n3213 ) ;
  assign n3215 = ( ~x239 & n2544 ) | ( ~x239 & n3214 ) | ( n2544 & n3214 ) ;
  assign n3216 = ( x207 & n829 ) | ( x207 & ~n1631 ) | ( n829 & ~n1631 ) ;
  assign n3217 = n528 & n3216 ;
  assign n3218 = n3217 ^ n1065 ^ 1'b0 ;
  assign n3219 = n3218 ^ n1638 ^ 1'b0 ;
  assign n3220 = ~n3215 & n3219 ;
  assign n3221 = n3220 ^ n2934 ^ 1'b0 ;
  assign n3222 = ( ~n2196 & n3211 ) | ( ~n2196 & n3221 ) | ( n3211 & n3221 ) ;
  assign n3230 = ~n565 & n727 ;
  assign n3223 = n1689 ^ n1505 ^ 1'b0 ;
  assign n3224 = x152 ^ x72 ^ 1'b0 ;
  assign n3225 = n3224 ^ n1791 ^ n691 ;
  assign n3226 = n3225 ^ n2095 ^ 1'b0 ;
  assign n3227 = n3223 & ~n3226 ;
  assign n3228 = n827 & ~n1333 ;
  assign n3229 = ~n3227 & n3228 ;
  assign n3231 = n3230 ^ n3229 ^ n2446 ;
  assign n3232 = x226 & n611 ;
  assign n3233 = n3232 ^ n715 ^ 1'b0 ;
  assign n3234 = n1856 & n3233 ;
  assign n3235 = n1312 ^ x133 ^ x95 ;
  assign n3236 = n3235 ^ n1087 ^ n387 ;
  assign n3237 = n3236 ^ x236 ^ 1'b0 ;
  assign n3238 = n3237 ^ n1013 ^ 1'b0 ;
  assign n3239 = n3234 & n3238 ;
  assign n3240 = ~n3131 & n3223 ;
  assign n3241 = n3240 ^ n1103 ^ 1'b0 ;
  assign n3242 = n3241 ^ n2002 ^ 1'b0 ;
  assign n3243 = ( n303 & n951 ) | ( n303 & ~n3242 ) | ( n951 & ~n3242 ) ;
  assign n3244 = n566 ^ n565 ^ x235 ;
  assign n3245 = n852 & ~n2828 ;
  assign n3246 = n3245 ^ n2495 ^ x222 ;
  assign n3247 = ( x203 & ~n713 ) | ( x203 & n1411 ) | ( ~n713 & n1411 ) ;
  assign n3248 = ( ~n1956 & n3246 ) | ( ~n1956 & n3247 ) | ( n3246 & n3247 ) ;
  assign n3261 = n2071 ^ n1968 ^ n1438 ;
  assign n3262 = ( n1313 & n1595 ) | ( n1313 & ~n3261 ) | ( n1595 & ~n3261 ) ;
  assign n3259 = ( x108 & ~n485 ) | ( x108 & n1155 ) | ( ~n485 & n1155 ) ;
  assign n3260 = n3259 ^ n2819 ^ 1'b0 ;
  assign n3250 = n1255 ^ n1184 ^ 1'b0 ;
  assign n3249 = n1365 & ~n2764 ;
  assign n3251 = n3250 ^ n3249 ^ x154 ;
  assign n3252 = n1053 ^ n672 ^ 1'b0 ;
  assign n3253 = n2764 & ~n3252 ;
  assign n3254 = n2981 ^ n1812 ^ n1088 ;
  assign n3255 = n3254 ^ n1231 ^ x59 ;
  assign n3256 = n2933 & n3255 ;
  assign n3257 = ~n3253 & n3256 ;
  assign n3258 = ( n1217 & n3251 ) | ( n1217 & n3257 ) | ( n3251 & n3257 ) ;
  assign n3263 = n3262 ^ n3260 ^ n3258 ;
  assign n3264 = x31 | n2938 ;
  assign n3265 = ( n853 & ~n1942 ) | ( n853 & n2976 ) | ( ~n1942 & n2976 ) ;
  assign n3266 = n1125 & n3075 ;
  assign n3267 = ( n2339 & n3265 ) | ( n2339 & ~n3266 ) | ( n3265 & ~n3266 ) ;
  assign n3269 = n2775 ^ n405 ^ x130 ;
  assign n3271 = n3269 ^ n926 ^ n311 ;
  assign n3272 = n3271 ^ n906 ^ 1'b0 ;
  assign n3268 = n1924 ^ n1453 ^ n727 ;
  assign n3270 = n3269 ^ n3268 ^ n377 ;
  assign n3273 = n3272 ^ n3270 ^ 1'b0 ;
  assign n3274 = n3267 | n3273 ;
  assign n3275 = n2518 ^ n1207 ^ x183 ;
  assign n3276 = x247 & ~n522 ;
  assign n3277 = ~n505 & n3276 ;
  assign n3278 = ( x101 & ~n2084 ) | ( x101 & n3277 ) | ( ~n2084 & n3277 ) ;
  assign n3279 = ( n313 & ~n3275 ) | ( n313 & n3278 ) | ( ~n3275 & n3278 ) ;
  assign n3280 = ~n1424 & n1587 ;
  assign n3281 = n3280 ^ n1308 ^ 1'b0 ;
  assign n3282 = n985 ^ n778 ^ 1'b0 ;
  assign n3288 = ( ~n1865 & n1870 ) | ( ~n1865 & n2358 ) | ( n1870 & n2358 ) ;
  assign n3289 = n3288 ^ x166 ^ x10 ;
  assign n3286 = n2787 ^ n2633 ^ 1'b0 ;
  assign n3287 = n2556 & n3286 ;
  assign n3290 = n3289 ^ n3287 ^ n1045 ;
  assign n3283 = n912 ^ n823 ^ 1'b0 ;
  assign n3284 = n1774 & n3283 ;
  assign n3285 = n1172 & n3284 ;
  assign n3291 = n3290 ^ n3285 ^ 1'b0 ;
  assign n3292 = n3282 & n3291 ;
  assign n3293 = n373 ^ x60 ^ x32 ;
  assign n3294 = n2478 | n3293 ;
  assign n3295 = n3294 ^ n1749 ^ n918 ;
  assign n3296 = ( n790 & n1175 ) | ( n790 & n1538 ) | ( n1175 & n1538 ) ;
  assign n3297 = n3296 ^ n1461 ^ x190 ;
  assign n3302 = n2078 & ~n2867 ;
  assign n3303 = ( n654 & n1943 ) | ( n654 & n3302 ) | ( n1943 & n3302 ) ;
  assign n3298 = ~n678 & n2012 ;
  assign n3299 = n1632 ^ n1469 ^ 1'b0 ;
  assign n3300 = n964 | n3299 ;
  assign n3301 = ( n342 & n3298 ) | ( n342 & ~n3300 ) | ( n3298 & ~n3300 ) ;
  assign n3304 = n3303 ^ n3301 ^ 1'b0 ;
  assign n3307 = n1235 & n1591 ;
  assign n3308 = n3307 ^ n997 ^ 1'b0 ;
  assign n3305 = ( n396 & n922 ) | ( n396 & n1316 ) | ( n922 & n1316 ) ;
  assign n3306 = ( x212 & n521 ) | ( x212 & ~n3305 ) | ( n521 & ~n3305 ) ;
  assign n3309 = n3308 ^ n3306 ^ n301 ;
  assign n3310 = x152 & ~n3309 ;
  assign n3311 = ~n3011 & n3310 ;
  assign n3319 = n3211 ^ n1821 ^ n1546 ;
  assign n3312 = x87 & x151 ;
  assign n3313 = n2904 & n3312 ;
  assign n3316 = n2408 ^ n2200 ^ x127 ;
  assign n3315 = n1523 ^ n445 ^ x225 ;
  assign n3314 = ( ~x135 & n622 ) | ( ~x135 & n1773 ) | ( n622 & n1773 ) ;
  assign n3317 = n3316 ^ n3315 ^ n3314 ;
  assign n3318 = ( n882 & ~n3313 ) | ( n882 & n3317 ) | ( ~n3313 & n3317 ) ;
  assign n3320 = n3319 ^ n3318 ^ n3074 ;
  assign n3321 = n3320 ^ n2491 ^ n1285 ;
  assign n3322 = n3321 ^ n2909 ^ n2628 ;
  assign n3323 = n296 ^ x213 ^ 1'b0 ;
  assign n3324 = n1339 & n3323 ;
  assign n3325 = n3324 ^ n2383 ^ 1'b0 ;
  assign n3326 = n1044 | n3325 ;
  assign n3327 = n1410 ^ n410 ^ 1'b0 ;
  assign n3328 = n655 & n3327 ;
  assign n3329 = ( ~n2957 & n3326 ) | ( ~n2957 & n3328 ) | ( n3326 & n3328 ) ;
  assign n3330 = x161 & n1441 ;
  assign n3331 = n1270 & n3330 ;
  assign n3332 = n3331 ^ n3015 ^ n1131 ;
  assign n3333 = n982 & ~n2601 ;
  assign n3334 = ( n1747 & n1800 ) | ( n1747 & ~n1994 ) | ( n1800 & ~n1994 ) ;
  assign n3335 = n3334 ^ n1999 ^ n1857 ;
  assign n3336 = ( x69 & ~n2114 ) | ( x69 & n2514 ) | ( ~n2114 & n2514 ) ;
  assign n3337 = n3336 ^ n2245 ^ n1677 ;
  assign n3339 = n2941 ^ n2544 ^ 1'b0 ;
  assign n3338 = ~n2375 & n3220 ;
  assign n3340 = n3339 ^ n3338 ^ 1'b0 ;
  assign n3341 = ( n615 & n1782 ) | ( n615 & n1891 ) | ( n1782 & n1891 ) ;
  assign n3342 = ( n690 & n2110 ) | ( n690 & n3341 ) | ( n2110 & n3341 ) ;
  assign n3343 = n3342 ^ n3096 ^ 1'b0 ;
  assign n3354 = n465 & ~n1682 ;
  assign n3353 = n2318 ^ n1879 ^ 1'b0 ;
  assign n3352 = x79 & n2130 ;
  assign n3355 = n3354 ^ n3353 ^ n3352 ;
  assign n3356 = ( n538 & n2628 ) | ( n538 & n3355 ) | ( n2628 & n3355 ) ;
  assign n3357 = ( n1829 & ~n2500 ) | ( n1829 & n3356 ) | ( ~n2500 & n3356 ) ;
  assign n3345 = n1061 ^ n982 ^ n574 ;
  assign n3346 = x59 & ~n1828 ;
  assign n3347 = n408 & n3346 ;
  assign n3348 = n3347 ^ n1323 ^ n430 ;
  assign n3349 = n3348 ^ n2777 ^ n782 ;
  assign n3350 = ( n1318 & n3345 ) | ( n1318 & n3349 ) | ( n3345 & n3349 ) ;
  assign n3351 = n2493 & ~n3350 ;
  assign n3358 = n3357 ^ n3351 ^ 1'b0 ;
  assign n3344 = n539 & n610 ;
  assign n3359 = n3358 ^ n3344 ^ 1'b0 ;
  assign n3360 = n2291 ^ n1410 ^ n1069 ;
  assign n3364 = ( ~x221 & n503 ) | ( ~x221 & n1824 ) | ( n503 & n1824 ) ;
  assign n3361 = ( ~n448 & n666 ) | ( ~n448 & n2300 ) | ( n666 & n2300 ) ;
  assign n3362 = n3361 ^ n1511 ^ 1'b0 ;
  assign n3363 = n626 & n3362 ;
  assign n3365 = n3364 ^ n3363 ^ n1798 ;
  assign n3366 = n2660 & n3365 ;
  assign n3367 = n3360 & n3366 ;
  assign n3370 = ( x188 & n1386 ) | ( x188 & ~n2629 ) | ( n1386 & ~n2629 ) ;
  assign n3371 = ( x179 & n400 ) | ( x179 & ~n548 ) | ( n400 & ~n548 ) ;
  assign n3372 = ( ~n491 & n3370 ) | ( ~n491 & n3371 ) | ( n3370 & n3371 ) ;
  assign n3368 = n1473 ^ n1284 ^ n418 ;
  assign n3369 = ( n2983 & n3236 ) | ( n2983 & n3368 ) | ( n3236 & n3368 ) ;
  assign n3373 = n3372 ^ n3369 ^ n971 ;
  assign n3374 = n722 & ~n1848 ;
  assign n3377 = ~n595 & n1956 ;
  assign n3375 = n2625 ^ x95 ^ 1'b0 ;
  assign n3376 = n3375 ^ n1921 ^ n364 ;
  assign n3378 = n3377 ^ n3376 ^ n3214 ;
  assign n3382 = n1090 ^ n564 ^ 1'b0 ;
  assign n3383 = n2012 & n3382 ;
  assign n3380 = n2070 ^ n345 ^ x229 ;
  assign n3381 = n1073 & ~n3380 ;
  assign n3384 = n3383 ^ n3381 ^ 1'b0 ;
  assign n3379 = n318 & n2209 ;
  assign n3385 = n3384 ^ n3379 ^ 1'b0 ;
  assign n3387 = n2799 ^ x109 ^ 1'b0 ;
  assign n3386 = n1280 ^ n810 ^ n337 ;
  assign n3388 = n3387 ^ n3386 ^ n715 ;
  assign n3389 = ~n651 & n1552 ;
  assign n3390 = n1976 & n3389 ;
  assign n3391 = n2154 & n3390 ;
  assign n3392 = ( n495 & n1585 ) | ( n495 & n1594 ) | ( n1585 & n1594 ) ;
  assign n3393 = n2430 | n2976 ;
  assign n3394 = n3392 & ~n3393 ;
  assign n3395 = ( n761 & ~n1489 ) | ( n761 & n3394 ) | ( ~n1489 & n3394 ) ;
  assign n3396 = ( n3388 & ~n3391 ) | ( n3388 & n3395 ) | ( ~n3391 & n3395 ) ;
  assign n3400 = n2929 ^ n1363 ^ n388 ;
  assign n3401 = n3400 ^ n2400 ^ n590 ;
  assign n3397 = n2358 ^ n1134 ^ x191 ;
  assign n3398 = n1897 ^ n341 ^ n286 ;
  assign n3399 = ( ~n823 & n3397 ) | ( ~n823 & n3398 ) | ( n3397 & n3398 ) ;
  assign n3402 = n3401 ^ n3399 ^ x152 ;
  assign n3403 = n2106 ^ n1602 ^ n1369 ;
  assign n3404 = n734 ^ n395 ^ x151 ;
  assign n3405 = ( n773 & n2865 ) | ( n773 & ~n3404 ) | ( n2865 & ~n3404 ) ;
  assign n3406 = n1806 & ~n3405 ;
  assign n3407 = n3406 ^ n3115 ^ n768 ;
  assign n3408 = ( n457 & ~n988 ) | ( n457 & n2875 ) | ( ~n988 & n2875 ) ;
  assign n3409 = ( n876 & n3067 ) | ( n876 & n3408 ) | ( n3067 & n3408 ) ;
  assign n3410 = n3409 ^ n2895 ^ n829 ;
  assign n3411 = n1179 & ~n2814 ;
  assign n3412 = ~n3410 & n3411 ;
  assign n3413 = ( x16 & n694 ) | ( x16 & ~n1104 ) | ( n694 & ~n1104 ) ;
  assign n3414 = ( x151 & n1110 ) | ( x151 & ~n1185 ) | ( n1110 & ~n1185 ) ;
  assign n3415 = x134 & ~n1748 ;
  assign n3416 = n3415 ^ n1477 ^ 1'b0 ;
  assign n3417 = ( x68 & n2667 ) | ( x68 & ~n3416 ) | ( n2667 & ~n3416 ) ;
  assign n3418 = n3417 ^ n1198 ^ x118 ;
  assign n3419 = ~n3414 & n3418 ;
  assign n3420 = ( n1907 & ~n3033 ) | ( n1907 & n3419 ) | ( ~n3033 & n3419 ) ;
  assign n3431 = n3168 ^ n1808 ^ n1065 ;
  assign n3432 = n474 & ~n3431 ;
  assign n3433 = ~n962 & n3432 ;
  assign n3424 = n1742 ^ n555 ^ 1'b0 ;
  assign n3425 = n3191 & n3424 ;
  assign n3426 = n729 | n998 ;
  assign n3427 = n3426 ^ x111 ^ 1'b0 ;
  assign n3428 = ( ~n295 & n2881 ) | ( ~n295 & n3427 ) | ( n2881 & n3427 ) ;
  assign n3429 = ( n1599 & n3425 ) | ( n1599 & n3428 ) | ( n3425 & n3428 ) ;
  assign n3421 = n965 ^ n486 ^ x247 ;
  assign n3422 = n3421 ^ n1105 ^ n670 ;
  assign n3423 = n2543 & ~n3422 ;
  assign n3430 = n3429 ^ n3423 ^ 1'b0 ;
  assign n3434 = n3433 ^ n3430 ^ n2857 ;
  assign n3435 = n3315 & ~n3434 ;
  assign n3436 = ( ~x61 & n1634 ) | ( ~x61 & n2222 ) | ( n1634 & n2222 ) ;
  assign n3437 = ( n2406 & ~n2759 ) | ( n2406 & n3436 ) | ( ~n2759 & n3436 ) ;
  assign n3438 = ~n3049 & n3437 ;
  assign n3439 = ~x208 & n3438 ;
  assign n3440 = ~n1200 & n1370 ;
  assign n3441 = n3440 ^ n365 ^ 1'b0 ;
  assign n3442 = ~n3016 & n3441 ;
  assign n3443 = n1475 & n3442 ;
  assign n3444 = n2126 ^ n948 ^ n879 ;
  assign n3445 = n1527 ^ n1412 ^ n383 ;
  assign n3446 = ( n1412 & n2659 ) | ( n1412 & n3445 ) | ( n2659 & n3445 ) ;
  assign n3447 = ( n753 & n2994 ) | ( n753 & ~n3446 ) | ( n2994 & ~n3446 ) ;
  assign n3453 = n775 ^ n753 ^ x236 ;
  assign n3454 = n3453 ^ n971 ^ x106 ;
  assign n3448 = n962 ^ x102 ^ x80 ;
  assign n3449 = n3448 ^ n564 ^ 1'b0 ;
  assign n3450 = x25 & n3449 ;
  assign n3451 = n3450 ^ x196 ^ x154 ;
  assign n3452 = n1021 & ~n3451 ;
  assign n3455 = n3454 ^ n3452 ^ 1'b0 ;
  assign n3456 = n448 & ~n1656 ;
  assign n3457 = n1863 ^ n283 ^ 1'b0 ;
  assign n3458 = n392 & n3457 ;
  assign n3459 = n3458 ^ n2623 ^ n2402 ;
  assign n3460 = n480 | n3459 ;
  assign n3461 = n3456 | n3460 ;
  assign n3462 = ~n3455 & n3461 ;
  assign n3463 = n2646 ^ n2473 ^ x73 ;
  assign n3464 = ( n478 & ~n2197 ) | ( n478 & n3463 ) | ( ~n2197 & n3463 ) ;
  assign n3466 = n1291 & ~n1618 ;
  assign n3467 = n3466 ^ n370 ^ 1'b0 ;
  assign n3465 = n1155 & n2311 ;
  assign n3468 = n3467 ^ n3465 ^ 1'b0 ;
  assign n3469 = n3468 ^ n1528 ^ n1030 ;
  assign n3470 = ( n283 & n3444 ) | ( n283 & n3469 ) | ( n3444 & n3469 ) ;
  assign n3471 = ( n610 & n732 ) | ( n610 & n2665 ) | ( n732 & n2665 ) ;
  assign n3472 = n3471 ^ n1272 ^ n948 ;
  assign n3473 = ( n844 & ~n2627 ) | ( n844 & n3472 ) | ( ~n2627 & n3472 ) ;
  assign n3476 = n1840 ^ n966 ^ x13 ;
  assign n3474 = ( x217 & ~n1008 ) | ( x217 & n2566 ) | ( ~n1008 & n2566 ) ;
  assign n3475 = n1138 & n3474 ;
  assign n3477 = n3476 ^ n3475 ^ 1'b0 ;
  assign n3480 = n1626 ^ n844 ^ 1'b0 ;
  assign n3478 = n2382 ^ n1334 ^ 1'b0 ;
  assign n3479 = ( n1188 & n1714 ) | ( n1188 & ~n3478 ) | ( n1714 & ~n3478 ) ;
  assign n3481 = n3480 ^ n3479 ^ n2041 ;
  assign n3482 = ( n1189 & n2386 ) | ( n1189 & n2620 ) | ( n2386 & n2620 ) ;
  assign n3483 = ( n2325 & n3481 ) | ( n2325 & n3482 ) | ( n3481 & n3482 ) ;
  assign n3484 = ( x77 & ~x114 ) | ( x77 & n1996 ) | ( ~x114 & n1996 ) ;
  assign n3485 = n562 & ~n1009 ;
  assign n3486 = ~n3250 & n3485 ;
  assign n3487 = ( ~n2134 & n3484 ) | ( ~n2134 & n3486 ) | ( n3484 & n3486 ) ;
  assign n3489 = n805 & n2386 ;
  assign n3490 = ~n2828 & n3489 ;
  assign n3491 = n3490 ^ n1386 ^ n1010 ;
  assign n3492 = n3491 ^ n2504 ^ 1'b0 ;
  assign n3488 = n3007 ^ n2830 ^ n2606 ;
  assign n3493 = n3492 ^ n3488 ^ n1908 ;
  assign n3494 = n1326 & n3493 ;
  assign n3495 = ( n2173 & n3264 ) | ( n2173 & n3494 ) | ( n3264 & n3494 ) ;
  assign n3497 = n3212 ^ n1217 ^ x145 ;
  assign n3496 = ( n923 & n1699 ) | ( n923 & ~n2738 ) | ( n1699 & ~n2738 ) ;
  assign n3498 = n3497 ^ n3496 ^ 1'b0 ;
  assign n3499 = n652 & n2311 ;
  assign n3500 = n3499 ^ n2975 ^ 1'b0 ;
  assign n3501 = n3500 ^ n1644 ^ n1218 ;
  assign n3502 = x65 & ~n3501 ;
  assign n3503 = n1658 & n3502 ;
  assign n3504 = n2210 ^ n597 ^ n343 ;
  assign n3505 = n1899 ^ n798 ^ n324 ;
  assign n3506 = n3505 ^ n1398 ^ n596 ;
  assign n3507 = ( n1220 & n3504 ) | ( n1220 & ~n3506 ) | ( n3504 & ~n3506 ) ;
  assign n3508 = ~n1376 & n3453 ;
  assign n3509 = n1102 & n3508 ;
  assign n3510 = n3509 ^ n1132 ^ 1'b0 ;
  assign n3511 = x160 & ~n3510 ;
  assign n3512 = n2097 ^ n1475 ^ 1'b0 ;
  assign n3520 = ( n805 & ~n811 ) | ( n805 & n1912 ) | ( ~n811 & n1912 ) ;
  assign n3513 = n425 & ~n620 ;
  assign n3514 = n3513 ^ x195 ^ 1'b0 ;
  assign n3515 = n933 | n3514 ;
  assign n3516 = n3515 ^ n1392 ^ 1'b0 ;
  assign n3517 = n3516 ^ n3294 ^ n2378 ;
  assign n3518 = n1402 & n2311 ;
  assign n3519 = n3517 & n3518 ;
  assign n3521 = n3520 ^ n3519 ^ n521 ;
  assign n3522 = n2760 ^ n720 ^ 1'b0 ;
  assign n3523 = ( x50 & ~n2967 ) | ( x50 & n3522 ) | ( ~n2967 & n3522 ) ;
  assign n3524 = n3523 ^ x73 ^ 1'b0 ;
  assign n3525 = n3524 ^ n772 ^ x161 ;
  assign n3526 = n3392 ^ n2939 ^ 1'b0 ;
  assign n3527 = n1523 ^ n1161 ^ 1'b0 ;
  assign n3528 = n2293 & n3527 ;
  assign n3529 = ~n352 & n840 ;
  assign n3530 = ~x130 & n3529 ;
  assign n3531 = n3530 ^ n2956 ^ n1885 ;
  assign n3532 = n3287 ^ n1742 ^ n482 ;
  assign n3533 = ( n3528 & ~n3531 ) | ( n3528 & n3532 ) | ( ~n3531 & n3532 ) ;
  assign n3534 = n1890 ^ n1455 ^ n1178 ;
  assign n3535 = ( x92 & x193 ) | ( x92 & n280 ) | ( x193 & n280 ) ;
  assign n3536 = n3535 ^ n3314 ^ 1'b0 ;
  assign n3537 = n3534 & n3536 ;
  assign n3538 = n3537 ^ n3410 ^ 1'b0 ;
  assign n3539 = ( ~n286 & n644 ) | ( ~n286 & n1923 ) | ( n644 & n1923 ) ;
  assign n3540 = n2067 & ~n3539 ;
  assign n3541 = ~n1431 & n3540 ;
  assign n3542 = n1127 ^ n304 ^ n277 ;
  assign n3543 = ( x186 & ~n800 ) | ( x186 & n2716 ) | ( ~n800 & n2716 ) ;
  assign n3544 = n3542 & ~n3543 ;
  assign n3545 = ( n441 & n829 ) | ( n441 & ~n2459 ) | ( n829 & ~n2459 ) ;
  assign n3546 = ( ~x244 & n523 ) | ( ~x244 & n640 ) | ( n523 & n640 ) ;
  assign n3547 = n3546 ^ x236 ^ 1'b0 ;
  assign n3548 = n3547 ^ n2541 ^ n2221 ;
  assign n3549 = ( n317 & n3545 ) | ( n317 & n3548 ) | ( n3545 & n3548 ) ;
  assign n3550 = ( n2297 & n3544 ) | ( n2297 & ~n3549 ) | ( n3544 & ~n3549 ) ;
  assign n3551 = ( n3359 & n3541 ) | ( n3359 & n3550 ) | ( n3541 & n3550 ) ;
  assign n3552 = n2406 ^ n795 ^ 1'b0 ;
  assign n3553 = ( ~n1651 & n2862 ) | ( ~n1651 & n3552 ) | ( n2862 & n3552 ) ;
  assign n3576 = ( x44 & n769 ) | ( x44 & ~n2071 ) | ( n769 & ~n2071 ) ;
  assign n3577 = n459 ^ x183 ^ x42 ;
  assign n3578 = ( n637 & ~n1045 ) | ( n637 & n3577 ) | ( ~n1045 & n3577 ) ;
  assign n3579 = ( n922 & n3576 ) | ( n922 & n3578 ) | ( n3576 & n3578 ) ;
  assign n3570 = ~n862 & n1573 ;
  assign n3571 = n3570 ^ n555 ^ 1'b0 ;
  assign n3572 = n1137 & n3571 ;
  assign n3567 = n772 ^ x204 ^ 1'b0 ;
  assign n3568 = n1514 | n3567 ;
  assign n3569 = n3568 ^ n2809 ^ 1'b0 ;
  assign n3555 = ~n316 & n666 ;
  assign n3556 = n3555 ^ n1338 ^ 1'b0 ;
  assign n3557 = n3556 ^ n1157 ^ n705 ;
  assign n3554 = ( n1188 & ~n2649 ) | ( n1188 & n2667 ) | ( ~n2649 & n2667 ) ;
  assign n3558 = n3557 ^ n3554 ^ x135 ;
  assign n3559 = ( n356 & n1043 ) | ( n356 & ~n1536 ) | ( n1043 & ~n1536 ) ;
  assign n3564 = n441 ^ n428 ^ x130 ;
  assign n3560 = ( x35 & n737 ) | ( x35 & n2349 ) | ( n737 & n2349 ) ;
  assign n3561 = n3560 ^ n643 ^ x141 ;
  assign n3562 = n3561 ^ n1087 ^ n719 ;
  assign n3563 = n3562 ^ n2710 ^ n1834 ;
  assign n3565 = n3564 ^ n3563 ^ n2179 ;
  assign n3566 = ( n3558 & n3559 ) | ( n3558 & ~n3565 ) | ( n3559 & ~n3565 ) ;
  assign n3573 = n3572 ^ n3569 ^ n3566 ;
  assign n3574 = ( n980 & n1953 ) | ( n980 & ~n2728 ) | ( n1953 & ~n2728 ) ;
  assign n3575 = n3573 & n3574 ;
  assign n3580 = n3579 ^ n3575 ^ 1'b0 ;
  assign n3581 = ( n2096 & ~n2330 ) | ( n2096 & n2420 ) | ( ~n2330 & n2420 ) ;
  assign n3582 = n3557 ^ n2566 ^ n1730 ;
  assign n3583 = n3582 ^ n3547 ^ x33 ;
  assign n3584 = ( ~n457 & n2084 ) | ( ~n457 & n3583 ) | ( n2084 & n3583 ) ;
  assign n3586 = n805 & ~n2885 ;
  assign n3587 = n3586 ^ n1809 ^ 1'b0 ;
  assign n3585 = ( n704 & n1993 ) | ( n704 & n3098 ) | ( n1993 & n3098 ) ;
  assign n3588 = n3587 ^ n3585 ^ n932 ;
  assign n3589 = ( x232 & n1989 ) | ( x232 & n3588 ) | ( n1989 & n3588 ) ;
  assign n3590 = n3589 ^ n1963 ^ n1258 ;
  assign n3591 = ( ~n2006 & n3584 ) | ( ~n2006 & n3590 ) | ( n3584 & n3590 ) ;
  assign n3592 = ~n2752 & n2815 ;
  assign n3593 = ( n2554 & n2846 ) | ( n2554 & ~n3592 ) | ( n2846 & ~n3592 ) ;
  assign n3594 = n3593 ^ n3111 ^ n1572 ;
  assign n3595 = ( x237 & ~n1291 ) | ( x237 & n2213 ) | ( ~n1291 & n2213 ) ;
  assign n3596 = n3151 & n3595 ;
  assign n3597 = n1486 & n3596 ;
  assign n3598 = ( x4 & n1184 ) | ( x4 & ~n2038 ) | ( n1184 & ~n2038 ) ;
  assign n3599 = ( n1117 & n2183 ) | ( n1117 & n3598 ) | ( n2183 & n3598 ) ;
  assign n3621 = ( ~n784 & n815 ) | ( ~n784 & n1655 ) | ( n815 & n1655 ) ;
  assign n3605 = ( ~n558 & n1554 ) | ( ~n558 & n1865 ) | ( n1554 & n1865 ) ;
  assign n3607 = n271 & ~n1218 ;
  assign n3608 = n3607 ^ n385 ^ 1'b0 ;
  assign n3609 = ~n1005 & n3608 ;
  assign n3606 = ( x132 & n823 ) | ( x132 & ~n1749 ) | ( n823 & ~n1749 ) ;
  assign n3610 = n3609 ^ n3606 ^ n1373 ;
  assign n3611 = x131 & n3610 ;
  assign n3612 = n3611 ^ n3421 ^ 1'b0 ;
  assign n3613 = n3605 & ~n3612 ;
  assign n3614 = x120 & n2499 ;
  assign n3615 = x171 & n3614 ;
  assign n3616 = n3615 ^ n2551 ^ 1'b0 ;
  assign n3617 = n2008 ^ n1406 ^ n306 ;
  assign n3618 = ( n1138 & n1223 ) | ( n1138 & n3617 ) | ( n1223 & n3617 ) ;
  assign n3619 = n3144 & ~n3618 ;
  assign n3620 = ( n3613 & ~n3616 ) | ( n3613 & n3619 ) | ( ~n3616 & n3619 ) ;
  assign n3602 = n2131 & n2183 ;
  assign n3603 = n3602 ^ n958 ^ 1'b0 ;
  assign n3600 = n1900 ^ n929 ^ 1'b0 ;
  assign n3601 = n2334 | n3600 ;
  assign n3604 = n3603 ^ n3601 ^ n2759 ;
  assign n3622 = n3621 ^ n3620 ^ n3604 ;
  assign n3623 = ( n288 & n743 ) | ( n288 & ~n866 ) | ( n743 & ~n866 ) ;
  assign n3624 = n3623 ^ n655 ^ n392 ;
  assign n3625 = n1296 ^ n596 ^ 1'b0 ;
  assign n3626 = n1406 ^ x105 ^ 1'b0 ;
  assign n3627 = n2821 & ~n3626 ;
  assign n3628 = ( n283 & n735 ) | ( n283 & n2770 ) | ( n735 & n2770 ) ;
  assign n3629 = ( n1196 & ~n2442 ) | ( n1196 & n3628 ) | ( ~n2442 & n3628 ) ;
  assign n3630 = ( ~n1384 & n2971 ) | ( ~n1384 & n3629 ) | ( n2971 & n3629 ) ;
  assign n3631 = n2653 ^ n1666 ^ x172 ;
  assign n3632 = ( ~n858 & n1670 ) | ( ~n858 & n2772 ) | ( n1670 & n2772 ) ;
  assign n3634 = n980 ^ n539 ^ n512 ;
  assign n3635 = n3634 ^ n985 ^ x224 ;
  assign n3636 = x148 & n622 ;
  assign n3637 = ( x120 & ~n336 ) | ( x120 & n1223 ) | ( ~n336 & n1223 ) ;
  assign n3638 = ( n3635 & n3636 ) | ( n3635 & n3637 ) | ( n3636 & n3637 ) ;
  assign n3633 = ( ~x142 & n1435 ) | ( ~x142 & n2294 ) | ( n1435 & n2294 ) ;
  assign n3639 = n3638 ^ n3633 ^ 1'b0 ;
  assign n3640 = n3639 ^ n1836 ^ 1'b0 ;
  assign n3641 = n3640 ^ n1748 ^ n779 ;
  assign n3643 = n2111 | n2589 ;
  assign n3644 = n1402 | n3643 ;
  assign n3645 = ( n730 & ~n1939 ) | ( n730 & n2772 ) | ( ~n1939 & n2772 ) ;
  assign n3646 = n3645 ^ n1731 ^ x204 ;
  assign n3647 = n2894 ^ n2201 ^ 1'b0 ;
  assign n3648 = ~n3646 & n3647 ;
  assign n3649 = ( n2183 & n3644 ) | ( n2183 & ~n3648 ) | ( n3644 & ~n3648 ) ;
  assign n3642 = ( n2250 & n2471 ) | ( n2250 & ~n3428 ) | ( n2471 & ~n3428 ) ;
  assign n3650 = n3649 ^ n3642 ^ 1'b0 ;
  assign n3651 = n2453 ^ n1782 ^ n1428 ;
  assign n3652 = ( ~n437 & n494 ) | ( ~n437 & n3651 ) | ( n494 & n3651 ) ;
  assign n3653 = n3652 ^ n724 ^ 1'b0 ;
  assign n3654 = n3392 ^ n1897 ^ 1'b0 ;
  assign n3655 = ( ~n1630 & n1649 ) | ( ~n1630 & n3654 ) | ( n1649 & n3654 ) ;
  assign n3656 = n410 ^ x184 ^ 1'b0 ;
  assign n3657 = n2243 | n3656 ;
  assign n3658 = n3657 ^ n1146 ^ 1'b0 ;
  assign n3659 = n3658 ^ n3497 ^ n552 ;
  assign n3660 = ( n2433 & n3655 ) | ( n2433 & ~n3659 ) | ( n3655 & ~n3659 ) ;
  assign n3662 = ( n498 & n932 ) | ( n498 & n2869 ) | ( n932 & n2869 ) ;
  assign n3661 = ( x111 & n466 ) | ( x111 & n1174 ) | ( n466 & n1174 ) ;
  assign n3663 = n3662 ^ n3661 ^ n1479 ;
  assign n3664 = ( x76 & n341 ) | ( x76 & ~n439 ) | ( n341 & ~n439 ) ;
  assign n3666 = n286 & ~n317 ;
  assign n3667 = n3666 ^ n909 ^ 1'b0 ;
  assign n3668 = ( n2202 & ~n2602 ) | ( n2202 & n3667 ) | ( ~n2602 & n3667 ) ;
  assign n3669 = n3668 ^ n632 ^ 1'b0 ;
  assign n3665 = n947 & ~n1197 ;
  assign n3670 = n3669 ^ n3665 ^ 1'b0 ;
  assign n3671 = ( ~x9 & n801 ) | ( ~x9 & n3670 ) | ( n801 & n3670 ) ;
  assign n3672 = n2443 | n2782 ;
  assign n3673 = ( n1882 & n2070 ) | ( n1882 & n3037 ) | ( n2070 & n3037 ) ;
  assign n3674 = ( x30 & n3672 ) | ( x30 & ~n3673 ) | ( n3672 & ~n3673 ) ;
  assign n3675 = n3636 ^ n2137 ^ n1510 ;
  assign n3676 = ( n558 & n1132 ) | ( n558 & n3675 ) | ( n1132 & n3675 ) ;
  assign n3677 = n486 & ~n2862 ;
  assign n3678 = n3677 ^ n2356 ^ 1'b0 ;
  assign n3679 = ( n506 & ~n928 ) | ( n506 & n3223 ) | ( ~n928 & n3223 ) ;
  assign n3680 = n3678 & n3679 ;
  assign n3681 = n2112 & ~n3680 ;
  assign n3682 = ( n963 & n1619 ) | ( n963 & n2335 ) | ( n1619 & n2335 ) ;
  assign n3683 = n1746 & n2849 ;
  assign n3684 = ~n845 & n3683 ;
  assign n3685 = ~n3682 & n3684 ;
  assign n3686 = ( n503 & ~n1166 ) | ( n503 & n3685 ) | ( ~n1166 & n3685 ) ;
  assign n3687 = n1128 ^ n305 ^ x137 ;
  assign n3688 = n1422 & n1596 ;
  assign n3689 = ~n647 & n3688 ;
  assign n3690 = n3687 & n3689 ;
  assign n3691 = n2215 ^ n965 ^ n525 ;
  assign n3692 = ~n1336 & n2145 ;
  assign n3693 = n3692 ^ n3037 ^ 1'b0 ;
  assign n3694 = n3585 ^ n2907 ^ n1081 ;
  assign n3695 = ( n3287 & ~n3693 ) | ( n3287 & n3694 ) | ( ~n3693 & n3694 ) ;
  assign n3696 = ( n1948 & n2842 ) | ( n1948 & ~n3695 ) | ( n2842 & ~n3695 ) ;
  assign n3697 = n2070 ^ n1305 ^ x55 ;
  assign n3698 = n1495 | n2704 ;
  assign n3699 = n3698 ^ n1898 ^ 1'b0 ;
  assign n3700 = ( n1696 & ~n2197 ) | ( n1696 & n3400 ) | ( ~n2197 & n3400 ) ;
  assign n3701 = ( ~n288 & n290 ) | ( ~n288 & n533 ) | ( n290 & n533 ) ;
  assign n3702 = ( n776 & n1342 ) | ( n776 & n3701 ) | ( n1342 & n3701 ) ;
  assign n3706 = n688 ^ x180 ^ 1'b0 ;
  assign n3704 = x161 & n1227 ;
  assign n3705 = n3704 ^ n1961 ^ 1'b0 ;
  assign n3707 = n3706 ^ n3705 ^ n2374 ;
  assign n3708 = n3707 ^ n3514 ^ 1'b0 ;
  assign n3703 = n1943 ^ n1529 ^ 1'b0 ;
  assign n3709 = n3708 ^ n3703 ^ 1'b0 ;
  assign n3710 = ( n781 & n811 ) | ( n781 & n2227 ) | ( n811 & n2227 ) ;
  assign n3711 = n2122 ^ n1293 ^ 1'b0 ;
  assign n3712 = n3710 | n3711 ;
  assign n3713 = n3712 ^ n2548 ^ 1'b0 ;
  assign n3714 = ( n3702 & ~n3709 ) | ( n3702 & n3713 ) | ( ~n3709 & n3713 ) ;
  assign n3715 = n2911 ^ n1147 ^ 1'b0 ;
  assign n3716 = ~n495 & n3474 ;
  assign n3717 = n3715 & n3716 ;
  assign n3718 = ( x160 & n908 ) | ( x160 & n2633 ) | ( n908 & n2633 ) ;
  assign n3719 = n3718 ^ n2978 ^ n1314 ;
  assign n3720 = ( n2272 & n3241 ) | ( n2272 & n3719 ) | ( n3241 & n3719 ) ;
  assign n3721 = ( x140 & ~n2646 ) | ( x140 & n3720 ) | ( ~n2646 & n3720 ) ;
  assign n3722 = n3543 ^ n2384 ^ x187 ;
  assign n3723 = n2206 | n3318 ;
  assign n3724 = n3723 ^ n1779 ^ 1'b0 ;
  assign n3727 = ( x61 & x108 ) | ( x61 & ~n1182 ) | ( x108 & ~n1182 ) ;
  assign n3725 = n2979 ^ n1136 ^ 1'b0 ;
  assign n3726 = n3725 ^ n1543 ^ n620 ;
  assign n3728 = n3727 ^ n3726 ^ n728 ;
  assign n3729 = n3728 ^ n3623 ^ n547 ;
  assign n3739 = n3093 ^ n1422 ^ n701 ;
  assign n3740 = n3458 ^ x222 ^ 1'b0 ;
  assign n3741 = n3739 & n3740 ;
  assign n3730 = ~n2967 & n3235 ;
  assign n3731 = n3041 & n3730 ;
  assign n3732 = ( x165 & n256 ) | ( x165 & ~n1840 ) | ( n256 & ~n1840 ) ;
  assign n3734 = ~n1085 & n3572 ;
  assign n3735 = n3072 & n3734 ;
  assign n3733 = n2255 ^ n1749 ^ 1'b0 ;
  assign n3736 = n3735 ^ n3733 ^ x175 ;
  assign n3737 = ( n3308 & n3732 ) | ( n3308 & ~n3736 ) | ( n3732 & ~n3736 ) ;
  assign n3738 = n3731 & n3737 ;
  assign n3742 = n3741 ^ n3738 ^ 1'b0 ;
  assign n3743 = ( ~x141 & n676 ) | ( ~x141 & n818 ) | ( n676 & n818 ) ;
  assign n3744 = ( x203 & n1253 ) | ( x203 & ~n3743 ) | ( n1253 & ~n3743 ) ;
  assign n3745 = n3744 ^ n3639 ^ n2172 ;
  assign n3755 = n2875 ^ n2119 ^ n1215 ;
  assign n3752 = ( x161 & n385 ) | ( x161 & n2073 ) | ( n385 & n2073 ) ;
  assign n3751 = n663 | n2791 ;
  assign n3753 = n3752 ^ n3751 ^ 1'b0 ;
  assign n3748 = x59 & ~n1791 ;
  assign n3749 = n3748 ^ n321 ^ 1'b0 ;
  assign n3750 = ( n957 & n1733 ) | ( n957 & n3749 ) | ( n1733 & n3749 ) ;
  assign n3754 = n3753 ^ n3750 ^ n673 ;
  assign n3756 = n3755 ^ n3754 ^ n1504 ;
  assign n3747 = ( x149 & n1976 ) | ( x149 & n2219 ) | ( n1976 & n2219 ) ;
  assign n3746 = n2700 ^ n770 ^ n561 ;
  assign n3757 = n3756 ^ n3747 ^ n3746 ;
  assign n3758 = n3757 ^ n2974 ^ n1751 ;
  assign n3759 = n2944 ^ n2544 ^ 1'b0 ;
  assign n3760 = n2834 | n3759 ;
  assign n3761 = n346 | n1501 ;
  assign n3762 = n487 & n1182 ;
  assign n3763 = n3762 ^ n2052 ^ 1'b0 ;
  assign n3764 = n2609 | n2808 ;
  assign n3769 = ( x94 & ~x203 ) | ( x94 & n2441 ) | ( ~x203 & n2441 ) ;
  assign n3770 = n3769 ^ n1455 ^ n675 ;
  assign n3765 = ( n279 & n631 ) | ( n279 & n876 ) | ( n631 & n876 ) ;
  assign n3766 = ( n1127 & n3037 ) | ( n1127 & ~n3765 ) | ( n3037 & ~n3765 ) ;
  assign n3767 = n3766 ^ n2831 ^ x9 ;
  assign n3768 = n3767 ^ n1479 ^ n997 ;
  assign n3771 = n3770 ^ n3768 ^ n2491 ;
  assign n3772 = n3771 ^ n3543 ^ n1050 ;
  assign n3773 = ( n3331 & n3764 ) | ( n3331 & n3772 ) | ( n3764 & n3772 ) ;
  assign n3774 = ( n394 & n1218 ) | ( n394 & ~n1686 ) | ( n1218 & ~n1686 ) ;
  assign n3775 = n2964 & ~n3774 ;
  assign n3776 = ~n1846 & n3775 ;
  assign n3777 = n1463 & n3490 ;
  assign n3780 = ( x31 & n592 ) | ( x31 & n2408 ) | ( n592 & n2408 ) ;
  assign n3781 = ( n952 & ~n2706 ) | ( n952 & n3780 ) | ( ~n2706 & n3780 ) ;
  assign n3782 = n405 & n3608 ;
  assign n3783 = ( n1664 & n3781 ) | ( n1664 & n3782 ) | ( n3781 & n3782 ) ;
  assign n3778 = n3668 ^ n3578 ^ n722 ;
  assign n3779 = n3778 ^ n730 ^ n379 ;
  assign n3784 = n3783 ^ n3779 ^ n3151 ;
  assign n3785 = ( n2559 & n3178 ) | ( n2559 & ~n3784 ) | ( n3178 & ~n3784 ) ;
  assign n3786 = ( ~n2996 & n3777 ) | ( ~n2996 & n3785 ) | ( n3777 & n3785 ) ;
  assign n3787 = n3786 ^ n1739 ^ 1'b0 ;
  assign n3788 = ( n373 & ~n1690 ) | ( n373 & n2959 ) | ( ~n1690 & n2959 ) ;
  assign n3789 = ( ~x81 & n472 ) | ( ~x81 & n3788 ) | ( n472 & n3788 ) ;
  assign n3790 = ( n826 & n2835 ) | ( n826 & n3789 ) | ( n2835 & n3789 ) ;
  assign n3791 = n3790 ^ n982 ^ n292 ;
  assign n3793 = n596 ^ n430 ^ n332 ;
  assign n3792 = ( n1320 & n2388 ) | ( n1320 & n3605 ) | ( n2388 & n3605 ) ;
  assign n3794 = n3793 ^ n3792 ^ x247 ;
  assign n3795 = n3794 ^ n1754 ^ 1'b0 ;
  assign n3796 = n3795 ^ n1205 ^ 1'b0 ;
  assign n3797 = n735 ^ x51 ^ 1'b0 ;
  assign n3798 = ( n1080 & n2664 ) | ( n1080 & ~n3797 ) | ( n2664 & ~n3797 ) ;
  assign n3799 = ( x10 & n729 ) | ( x10 & ~n784 ) | ( n729 & ~n784 ) ;
  assign n3800 = n3799 ^ n2231 ^ n346 ;
  assign n3801 = ~n1550 & n3800 ;
  assign n3802 = ( x246 & n3798 ) | ( x246 & ~n3801 ) | ( n3798 & ~n3801 ) ;
  assign n3806 = x236 & ~n2716 ;
  assign n3807 = ~n405 & n3806 ;
  assign n3803 = x244 | n1299 ;
  assign n3804 = n3803 ^ n3060 ^ 1'b0 ;
  assign n3805 = n2790 & ~n3804 ;
  assign n3808 = n3807 ^ n3805 ^ n2928 ;
  assign n3809 = n375 & ~n1499 ;
  assign n3810 = n3809 ^ n2959 ^ 1'b0 ;
  assign n3811 = n3810 ^ n1881 ^ n1754 ;
  assign n3812 = n511 & n3811 ;
  assign n3813 = n1986 ^ n1041 ^ n425 ;
  assign n3814 = n3813 ^ n2921 ^ n2693 ;
  assign n3815 = n3812 | n3814 ;
  assign n3816 = n1423 & ~n3815 ;
  assign n3817 = n567 | n595 ;
  assign n3818 = n3816 & ~n3817 ;
  assign n3819 = n1784 ^ n1263 ^ 1'b0 ;
  assign n3820 = n2388 ^ n1952 ^ n352 ;
  assign n3821 = n3819 | n3820 ;
  assign n3822 = n632 & ~n3821 ;
  assign n3823 = ( n582 & ~n982 ) | ( n582 & n1711 ) | ( ~n982 & n1711 ) ;
  assign n3824 = n3305 ^ n866 ^ n647 ;
  assign n3825 = n3824 ^ n1961 ^ n1699 ;
  assign n3826 = ( x237 & ~n3823 ) | ( x237 & n3825 ) | ( ~n3823 & n3825 ) ;
  assign n3832 = ~n770 & n2787 ;
  assign n3833 = n1500 & n3832 ;
  assign n3830 = ( n1950 & ~n2062 ) | ( n1950 & n2773 ) | ( ~n2062 & n2773 ) ;
  assign n3831 = ( n2296 & ~n2302 ) | ( n2296 & n3830 ) | ( ~n2302 & n3830 ) ;
  assign n3827 = ~n529 & n3528 ;
  assign n3828 = n3827 ^ n3610 ^ 1'b0 ;
  assign n3829 = n1246 & ~n3828 ;
  assign n3834 = n3833 ^ n3831 ^ n3829 ;
  assign n3835 = n327 | n912 ;
  assign n3836 = n2525 ^ x249 ^ 1'b0 ;
  assign n3837 = n3836 ^ n1761 ^ n607 ;
  assign n3838 = ( ~n1657 & n3835 ) | ( ~n1657 & n3837 ) | ( n3835 & n3837 ) ;
  assign n3843 = ( n1552 & n1862 ) | ( n1552 & n2836 ) | ( n1862 & n2836 ) ;
  assign n3839 = ( ~n1052 & n1359 ) | ( ~n1052 & n2984 ) | ( n1359 & n2984 ) ;
  assign n3840 = n3839 ^ n3268 ^ n1594 ;
  assign n3841 = ( n1768 & n3659 ) | ( n1768 & ~n3840 ) | ( n3659 & ~n3840 ) ;
  assign n3842 = n2917 & n3841 ;
  assign n3844 = n3843 ^ n3842 ^ 1'b0 ;
  assign n3845 = ( n2522 & ~n3838 ) | ( n2522 & n3844 ) | ( ~n3838 & n3844 ) ;
  assign n3846 = n1527 ^ n621 ^ x189 ;
  assign n3847 = n1761 ^ n305 ^ x1 ;
  assign n3848 = ( n1142 & n1160 ) | ( n1142 & n3847 ) | ( n1160 & n3847 ) ;
  assign n3849 = ( ~n711 & n2693 ) | ( ~n711 & n3651 ) | ( n2693 & n3651 ) ;
  assign n3850 = n3848 & ~n3849 ;
  assign n3851 = n3846 & n3850 ;
  assign n3852 = ~n1349 & n2105 ;
  assign n3853 = n3852 ^ n2868 ^ n514 ;
  assign n3854 = n3851 | n3853 ;
  assign n3855 = ( n1505 & n1557 ) | ( n1505 & ~n2730 ) | ( n1557 & ~n2730 ) ;
  assign n3856 = n3855 ^ n820 ^ 1'b0 ;
  assign n3857 = n2750 ^ n1572 ^ n647 ;
  assign n3858 = n1972 | n3857 ;
  assign n3859 = n690 | n3858 ;
  assign n3861 = ( n287 & ~n1039 ) | ( n287 & n2238 ) | ( ~n1039 & n2238 ) ;
  assign n3860 = n3705 ^ n1869 ^ x152 ;
  assign n3862 = n3861 ^ n3860 ^ n875 ;
  assign n3863 = ( ~n987 & n3859 ) | ( ~n987 & n3862 ) | ( n3859 & n3862 ) ;
  assign n3864 = n1730 ^ n1671 ^ n463 ;
  assign n3865 = n3864 ^ n1989 ^ n505 ;
  assign n3866 = n3865 ^ x251 ^ 1'b0 ;
  assign n3867 = ( n2760 & ~n3863 ) | ( n2760 & n3866 ) | ( ~n3863 & n3866 ) ;
  assign n3868 = n3867 ^ x42 ^ 1'b0 ;
  assign n3869 = n1836 & ~n3868 ;
  assign n3871 = n3347 ^ n1280 ^ 1'b0 ;
  assign n3870 = n3235 ^ n1364 ^ n1191 ;
  assign n3872 = n3871 ^ n3870 ^ n279 ;
  assign n3875 = ( ~n428 & n1467 ) | ( ~n428 & n2465 ) | ( n1467 & n2465 ) ;
  assign n3876 = n3875 ^ n2384 ^ n299 ;
  assign n3873 = n3793 ^ n2444 ^ x85 ;
  assign n3874 = ( n2273 & n2864 ) | ( n2273 & n3873 ) | ( n2864 & n3873 ) ;
  assign n3877 = n3876 ^ n3874 ^ n1447 ;
  assign n3879 = n3368 ^ n2697 ^ n1044 ;
  assign n3880 = n2556 & n3879 ;
  assign n3878 = n2455 ^ n1126 ^ x33 ;
  assign n3881 = n3880 ^ n3878 ^ 1'b0 ;
  assign n3882 = n2101 & n3881 ;
  assign n3883 = ( ~n1411 & n1602 ) | ( ~n1411 & n3882 ) | ( n1602 & n3882 ) ;
  assign n3884 = n2978 ^ n852 ^ n569 ;
  assign n3885 = ( x35 & n2786 ) | ( x35 & ~n3884 ) | ( n2786 & ~n3884 ) ;
  assign n3886 = n3072 ^ n1391 ^ 1'b0 ;
  assign n3887 = n2435 & n3886 ;
  assign n3888 = n2649 | n3887 ;
  assign n3889 = ( x158 & x197 ) | ( x158 & ~n3888 ) | ( x197 & ~n3888 ) ;
  assign n3890 = ~n1656 & n2984 ;
  assign n3891 = n3890 ^ n3739 ^ 1'b0 ;
  assign n3892 = n3891 ^ n3542 ^ n1612 ;
  assign n3896 = n1353 & ~n2720 ;
  assign n3897 = n3896 ^ n2662 ^ 1'b0 ;
  assign n3895 = n1332 & ~n3050 ;
  assign n3898 = n3897 ^ n3895 ^ 1'b0 ;
  assign n3893 = ~n1708 & n2553 ;
  assign n3894 = ( n2779 & ~n3547 ) | ( n2779 & n3893 ) | ( ~n3547 & n3893 ) ;
  assign n3899 = n3898 ^ n3894 ^ n415 ;
  assign n3900 = ( ~n3889 & n3892 ) | ( ~n3889 & n3899 ) | ( n3892 & n3899 ) ;
  assign n3901 = ( n1227 & n1857 ) | ( n1227 & n3347 ) | ( n1857 & n3347 ) ;
  assign n3902 = ( ~n1962 & n3614 ) | ( ~n1962 & n3901 ) | ( n3614 & n3901 ) ;
  assign n3906 = n2848 ^ n1968 ^ 1'b0 ;
  assign n3907 = ( n375 & n2238 ) | ( n375 & ~n3906 ) | ( n2238 & ~n3906 ) ;
  assign n3908 = ( n3357 & ~n3847 ) | ( n3357 & n3907 ) | ( ~n3847 & n3907 ) ;
  assign n3903 = n927 ^ n636 ^ 1'b0 ;
  assign n3904 = n3671 | n3903 ;
  assign n3905 = n1238 | n3904 ;
  assign n3909 = n3908 ^ n3905 ^ 1'b0 ;
  assign n3917 = n2245 ^ n1804 ^ n1493 ;
  assign n3912 = n295 ^ x239 ^ 1'b0 ;
  assign n3913 = x33 & n3912 ;
  assign n3914 = n3578 ^ n2760 ^ 1'b0 ;
  assign n3915 = ~n2361 & n3914 ;
  assign n3916 = ( n3516 & n3913 ) | ( n3516 & n3915 ) | ( n3913 & n3915 ) ;
  assign n3918 = n3917 ^ n3916 ^ n413 ;
  assign n3910 = n2170 ^ n1464 ^ 1'b0 ;
  assign n3911 = ( n2538 & ~n3322 ) | ( n2538 & n3910 ) | ( ~n3322 & n3910 ) ;
  assign n3919 = n3918 ^ n3911 ^ n1144 ;
  assign n3920 = n2437 ^ n1075 ^ x172 ;
  assign n3921 = ~n422 & n2447 ;
  assign n3922 = ( ~n854 & n1560 ) | ( ~n854 & n3921 ) | ( n1560 & n3921 ) ;
  assign n3931 = n3154 ^ n1604 ^ 1'b0 ;
  assign n3932 = n1149 & ~n3931 ;
  assign n3927 = ( x215 & n1013 ) | ( x215 & n2491 ) | ( n1013 & n2491 ) ;
  assign n3928 = ( n1302 & n1592 ) | ( n1302 & n1864 ) | ( n1592 & n1864 ) ;
  assign n3929 = n1393 | n3928 ;
  assign n3930 = ( n2043 & ~n3927 ) | ( n2043 & n3929 ) | ( ~n3927 & n3929 ) ;
  assign n3923 = n1083 ^ n980 ^ n492 ;
  assign n3924 = ( ~n721 & n947 ) | ( ~n721 & n1177 ) | ( n947 & n1177 ) ;
  assign n3925 = ( n1774 & n2108 ) | ( n1774 & n3275 ) | ( n2108 & n3275 ) ;
  assign n3926 = ( n3923 & n3924 ) | ( n3923 & ~n3925 ) | ( n3924 & ~n3925 ) ;
  assign n3933 = n3932 ^ n3930 ^ n3926 ;
  assign n3934 = n3922 & ~n3933 ;
  assign n3935 = n3920 & n3934 ;
  assign n3937 = n566 | n1389 ;
  assign n3936 = ( x126 & ~x141 ) | ( x126 & n1878 ) | ( ~x141 & n1878 ) ;
  assign n3938 = n3937 ^ n3936 ^ n1085 ;
  assign n3945 = n2567 ^ n2014 ^ 1'b0 ;
  assign n3943 = n3431 ^ n1761 ^ 1'b0 ;
  assign n3944 = n2384 | n3943 ;
  assign n3946 = n3945 ^ n3944 ^ 1'b0 ;
  assign n3947 = n3946 ^ n3644 ^ n2301 ;
  assign n3948 = x77 | n3947 ;
  assign n3940 = ( n920 & n1496 ) | ( n920 & n1562 ) | ( n1496 & n1562 ) ;
  assign n3939 = n2959 ^ n992 ^ n956 ;
  assign n3941 = n3940 ^ n3939 ^ n1986 ;
  assign n3942 = n3941 ^ n2255 ^ x75 ;
  assign n3949 = n3948 ^ n3942 ^ n1030 ;
  assign n3950 = n3066 ^ n1440 ^ n1282 ;
  assign n3951 = n3950 ^ n400 ^ 1'b0 ;
  assign n3952 = ( ~n1944 & n3949 ) | ( ~n1944 & n3951 ) | ( n3949 & n3951 ) ;
  assign n3953 = n355 & ~n544 ;
  assign n3954 = ~x142 & n3953 ;
  assign n3955 = n3954 ^ n1849 ^ 1'b0 ;
  assign n3956 = ( x10 & n2851 ) | ( x10 & ~n3701 ) | ( n2851 & ~n3701 ) ;
  assign n3957 = n715 & n3741 ;
  assign n3958 = ( ~x21 & n2902 ) | ( ~x21 & n3957 ) | ( n2902 & n3957 ) ;
  assign n3959 = ( n1050 & n2188 ) | ( n1050 & n2943 ) | ( n2188 & n2943 ) ;
  assign n3960 = n3959 ^ n2656 ^ x132 ;
  assign n3961 = n1147 ^ x91 ^ 1'b0 ;
  assign n3964 = ( n1946 & n2670 ) | ( n1946 & ~n2867 ) | ( n2670 & ~n2867 ) ;
  assign n3962 = n703 ^ n509 ^ n377 ;
  assign n3963 = ( n859 & ~n1288 ) | ( n859 & n3962 ) | ( ~n1288 & n3962 ) ;
  assign n3965 = n3964 ^ n3963 ^ n3317 ;
  assign n3966 = n3965 ^ x124 ^ 1'b0 ;
  assign n3967 = ( n1695 & n3961 ) | ( n1695 & ~n3966 ) | ( n3961 & ~n3966 ) ;
  assign n3968 = n1549 ^ n1465 ^ n898 ;
  assign n3971 = n1943 ^ n1525 ^ x199 ;
  assign n3969 = n390 | n2161 ;
  assign n3970 = ( n986 & ~n1408 ) | ( n986 & n3969 ) | ( ~n1408 & n3969 ) ;
  assign n3972 = n3971 ^ n3970 ^ n428 ;
  assign n3973 = n3972 ^ n1854 ^ x37 ;
  assign n3974 = n2197 | n3973 ;
  assign n3975 = n3968 | n3974 ;
  assign n3976 = ( n283 & n424 ) | ( n283 & ~n1135 ) | ( n424 & ~n1135 ) ;
  assign n3977 = n964 & n3976 ;
  assign n3978 = n3977 ^ n3634 ^ 1'b0 ;
  assign n3979 = ( x75 & ~n1538 ) | ( x75 & n2735 ) | ( ~n1538 & n2735 ) ;
  assign n3980 = ( ~n3192 & n3978 ) | ( ~n3192 & n3979 ) | ( n3978 & n3979 ) ;
  assign n3981 = ( n2504 & n2848 ) | ( n2504 & n2880 ) | ( n2848 & n2880 ) ;
  assign n3982 = n2056 ^ n646 ^ n503 ;
  assign n3983 = n3982 ^ n1291 ^ n1114 ;
  assign n3984 = ( n2040 & n3981 ) | ( n2040 & n3983 ) | ( n3981 & n3983 ) ;
  assign n3985 = n1058 & n1915 ;
  assign n3986 = x205 & n1767 ;
  assign n3987 = n3985 & n3986 ;
  assign n3988 = n1324 ^ n1202 ^ n665 ;
  assign n3989 = n3988 ^ n1946 ^ n1794 ;
  assign n3990 = n636 & ~n3989 ;
  assign n3991 = n3990 ^ n1948 ^ 1'b0 ;
  assign n3992 = x180 & ~n636 ;
  assign n3993 = n3992 ^ n2104 ^ 1'b0 ;
  assign n4009 = n1378 ^ n1040 ^ 1'b0 ;
  assign n3999 = n966 ^ n633 ^ x162 ;
  assign n4000 = ( n696 & n1169 ) | ( n696 & ~n3999 ) | ( n1169 & ~n3999 ) ;
  assign n4005 = ( n567 & n1106 ) | ( n567 & n3560 ) | ( n1106 & n3560 ) ;
  assign n4001 = n540 & n649 ;
  assign n4002 = ~n3093 & n4001 ;
  assign n4003 = ( n1102 & n1195 ) | ( n1102 & ~n4002 ) | ( n1195 & ~n4002 ) ;
  assign n4004 = n4003 ^ n3380 ^ 1'b0 ;
  assign n4006 = n4005 ^ n4004 ^ n2067 ;
  assign n4007 = ( ~n504 & n3021 ) | ( ~n504 & n4006 ) | ( n3021 & n4006 ) ;
  assign n4008 = ( n2962 & ~n4000 ) | ( n2962 & n4007 ) | ( ~n4000 & n4007 ) ;
  assign n3994 = ( n472 & ~n851 ) | ( n472 & n1316 ) | ( ~n851 & n1316 ) ;
  assign n3995 = n1473 ^ x212 ^ 1'b0 ;
  assign n3996 = ( x190 & n1638 ) | ( x190 & ~n2293 ) | ( n1638 & ~n2293 ) ;
  assign n3997 = ( n2804 & n3995 ) | ( n2804 & ~n3996 ) | ( n3995 & ~n3996 ) ;
  assign n3998 = ( n788 & n3994 ) | ( n788 & ~n3997 ) | ( n3994 & ~n3997 ) ;
  assign n4010 = n4009 ^ n4008 ^ n3998 ;
  assign n4011 = n2737 ^ n2157 ^ n1736 ;
  assign n4019 = ( ~n1363 & n1591 ) | ( ~n1363 & n1655 ) | ( n1591 & n1655 ) ;
  assign n4020 = n2099 ^ n1371 ^ n393 ;
  assign n4021 = ( ~n1471 & n2024 ) | ( ~n1471 & n4020 ) | ( n2024 & n4020 ) ;
  assign n4022 = n3606 ^ n654 ^ 1'b0 ;
  assign n4023 = ~n3041 & n4022 ;
  assign n4024 = ( ~n4019 & n4021 ) | ( ~n4019 & n4023 ) | ( n4021 & n4023 ) ;
  assign n4017 = n3427 ^ n899 ^ x93 ;
  assign n4015 = n1655 ^ n641 ^ 1'b0 ;
  assign n4013 = n1805 ^ n867 ^ 1'b0 ;
  assign n4014 = n1242 | n4013 ;
  assign n4016 = n4015 ^ n4014 ^ n2335 ;
  assign n4018 = n4017 ^ n4016 ^ n3365 ;
  assign n4012 = ( x212 & n693 ) | ( x212 & ~n1243 ) | ( n693 & ~n1243 ) ;
  assign n4025 = n4024 ^ n4018 ^ n4012 ;
  assign n4026 = ( n315 & n2485 ) | ( n315 & ~n2606 ) | ( n2485 & ~n2606 ) ;
  assign n4027 = n4026 ^ n2845 ^ n1224 ;
  assign n4028 = n4027 ^ n2879 ^ n1604 ;
  assign n4029 = n4028 ^ n3111 ^ n1460 ;
  assign n4030 = n1241 ^ n1216 ^ n783 ;
  assign n4031 = ( n2319 & n3743 ) | ( n2319 & ~n4030 ) | ( n3743 & ~n4030 ) ;
  assign n4032 = ( ~n2130 & n4029 ) | ( ~n2130 & n4031 ) | ( n4029 & n4031 ) ;
  assign n4033 = ( n4011 & ~n4025 ) | ( n4011 & n4032 ) | ( ~n4025 & n4032 ) ;
  assign n4034 = n3759 ^ n1625 ^ n757 ;
  assign n4035 = n4034 ^ n3981 ^ x98 ;
  assign n4036 = n2647 ^ n1105 ^ n505 ;
  assign n4037 = n4036 ^ n2895 ^ 1'b0 ;
  assign n4038 = n2109 ^ n766 ^ x77 ;
  assign n4039 = ( n436 & n447 ) | ( n436 & n2558 ) | ( n447 & n2558 ) ;
  assign n4040 = n2014 ^ n1459 ^ 1'b0 ;
  assign n4041 = n4040 ^ n3490 ^ 1'b0 ;
  assign n4042 = n2527 & n4041 ;
  assign n4043 = n4042 ^ n2482 ^ n1418 ;
  assign n4044 = ( n1907 & n2638 ) | ( n1907 & ~n4043 ) | ( n2638 & ~n4043 ) ;
  assign n4045 = n2448 ^ n2095 ^ n1547 ;
  assign n4046 = n941 & n4045 ;
  assign n4047 = n4046 ^ n2210 ^ 1'b0 ;
  assign n4049 = n2150 ^ n982 ^ x196 ;
  assign n4048 = n480 ^ n439 ^ x11 ;
  assign n4050 = n4049 ^ n4048 ^ 1'b0 ;
  assign n4051 = n2228 ^ n2196 ^ n1567 ;
  assign n4052 = n3083 ^ n333 ^ 1'b0 ;
  assign n4053 = n4051 & ~n4052 ;
  assign n4054 = n1182 & n2830 ;
  assign n4055 = n4054 ^ n2743 ^ 1'b0 ;
  assign n4056 = ( n1359 & n4053 ) | ( n1359 & n4055 ) | ( n4053 & n4055 ) ;
  assign n4062 = n3727 ^ n3468 ^ n2977 ;
  assign n4063 = n1363 ^ x186 ^ x152 ;
  assign n4064 = n3277 ^ n1194 ^ n956 ;
  assign n4065 = n3253 & ~n4064 ;
  assign n4066 = ~n4063 & n4065 ;
  assign n4067 = n1135 & ~n4066 ;
  assign n4068 = n901 & n4067 ;
  assign n4069 = n3619 | n4068 ;
  assign n4070 = n4062 & ~n4069 ;
  assign n4059 = n3054 ^ n2138 ^ n2134 ;
  assign n4058 = x218 & n622 ;
  assign n4060 = n4059 ^ n4058 ^ 1'b0 ;
  assign n4057 = n3752 ^ n2589 ^ n2500 ;
  assign n4061 = n4060 ^ n4057 ^ n804 ;
  assign n4071 = n4070 ^ n4061 ^ n2289 ;
  assign n4080 = ( n313 & n2881 ) | ( n313 & ~n3057 ) | ( n2881 & ~n3057 ) ;
  assign n4075 = n1592 ^ n1071 ^ x226 ;
  assign n4076 = x17 & ~n4075 ;
  assign n4077 = ~n517 & n4076 ;
  assign n4072 = ( n1161 & ~n2769 ) | ( n1161 & n4066 ) | ( ~n2769 & n4066 ) ;
  assign n4073 = n2776 ^ n2572 ^ n1474 ;
  assign n4074 = ( n3968 & n4072 ) | ( n3968 & ~n4073 ) | ( n4072 & ~n4073 ) ;
  assign n4078 = n4077 ^ n4074 ^ n2868 ;
  assign n4079 = ( n1871 & n2359 ) | ( n1871 & ~n4078 ) | ( n2359 & ~n4078 ) ;
  assign n4081 = n4080 ^ n4079 ^ n3255 ;
  assign n4091 = ( ~n2492 & n2850 ) | ( ~n2492 & n3007 ) | ( n2850 & n3007 ) ;
  assign n4086 = n1250 & n2717 ;
  assign n4087 = n4086 ^ n1384 ^ 1'b0 ;
  assign n4088 = ( n1204 & n3007 ) | ( n1204 & ~n4087 ) | ( n3007 & ~n4087 ) ;
  assign n4083 = n653 ^ x190 ^ 1'b0 ;
  assign n4084 = n3725 & n4083 ;
  assign n4082 = n2096 ^ n813 ^ x67 ;
  assign n4085 = n4084 ^ n4082 ^ 1'b0 ;
  assign n4089 = n4088 ^ n4085 ^ n2027 ;
  assign n4090 = n4089 ^ n736 ^ x116 ;
  assign n4092 = n4091 ^ n4090 ^ n3685 ;
  assign n4093 = n1881 ^ n1405 ^ 1'b0 ;
  assign n4094 = n2435 ^ n923 ^ n567 ;
  assign n4095 = ( ~n1280 & n4093 ) | ( ~n1280 & n4094 ) | ( n4093 & n4094 ) ;
  assign n4096 = n409 ^ x12 ^ 1'b0 ;
  assign n4097 = n4096 ^ n2857 ^ n1708 ;
  assign n4098 = ( n3429 & n3593 ) | ( n3429 & ~n4097 ) | ( n3593 & ~n4097 ) ;
  assign n4104 = ( n2036 & ~n2848 ) | ( n2036 & n3545 ) | ( ~n2848 & n3545 ) ;
  assign n4100 = n1125 ^ n1017 ^ x178 ;
  assign n4099 = ( n565 & ~n2790 ) | ( n565 & n3505 ) | ( ~n2790 & n3505 ) ;
  assign n4101 = n4100 ^ n4099 ^ n1159 ;
  assign n4102 = n4101 ^ n3250 ^ 1'b0 ;
  assign n4103 = n2142 & ~n4102 ;
  assign n4105 = n4104 ^ n4103 ^ n3873 ;
  assign n4106 = n2901 ^ n983 ^ 1'b0 ;
  assign n4107 = ~n256 & n4106 ;
  assign n4108 = ( n587 & n2323 ) | ( n587 & n3861 ) | ( n2323 & n3861 ) ;
  assign n4109 = ( n733 & n4107 ) | ( n733 & n4108 ) | ( n4107 & n4108 ) ;
  assign n4110 = n4109 ^ n1384 ^ n270 ;
  assign n4111 = n4110 ^ n2417 ^ n959 ;
  assign n4112 = n1736 ^ x131 ^ 1'b0 ;
  assign n4113 = x19 & ~n4112 ;
  assign n4114 = n4113 ^ n2455 ^ x25 ;
  assign n4115 = ~n2452 & n4114 ;
  assign n4116 = n3316 ^ n2940 ^ n2706 ;
  assign n4117 = n2641 ^ n1429 ^ n739 ;
  assign n4118 = n4117 ^ n2630 ^ n585 ;
  assign n4119 = n3937 ^ n1870 ^ x135 ;
  assign n4120 = n288 & ~n4119 ;
  assign n4121 = n4120 ^ x29 ^ 1'b0 ;
  assign n4122 = n648 ^ n546 ^ x178 ;
  assign n4123 = x138 & ~n1331 ;
  assign n4124 = ~x160 & n4123 ;
  assign n4125 = n4124 ^ n704 ^ 1'b0 ;
  assign n4126 = x128 & n4125 ;
  assign n4127 = n4126 ^ n4096 ^ n1170 ;
  assign n4128 = ( n3044 & n3592 ) | ( n3044 & n4127 ) | ( n3592 & n4127 ) ;
  assign n4134 = ( x56 & n323 ) | ( x56 & ~n715 ) | ( n323 & ~n715 ) ;
  assign n4135 = ( ~n621 & n3392 ) | ( ~n621 & n4134 ) | ( n3392 & n4134 ) ;
  assign n4133 = ( n631 & n1767 ) | ( n631 & n3136 ) | ( n1767 & n3136 ) ;
  assign n4130 = ( n972 & n1724 ) | ( n972 & ~n2703 ) | ( n1724 & ~n2703 ) ;
  assign n4131 = n4130 ^ n3626 ^ n3105 ;
  assign n4129 = ( ~n814 & n1798 ) | ( ~n814 & n2473 ) | ( n1798 & n2473 ) ;
  assign n4132 = n4131 ^ n4129 ^ n3589 ;
  assign n4136 = n4135 ^ n4133 ^ n4132 ;
  assign n4137 = n4136 ^ n2460 ^ x230 ;
  assign n4138 = ( n4122 & ~n4128 ) | ( n4122 & n4137 ) | ( ~n4128 & n4137 ) ;
  assign n4139 = ~n4121 & n4138 ;
  assign n4140 = n3617 & n4139 ;
  assign n4141 = ( ~n1419 & n4118 ) | ( ~n1419 & n4140 ) | ( n4118 & n4140 ) ;
  assign n4145 = ( ~n940 & n1690 ) | ( ~n940 & n2507 ) | ( n1690 & n2507 ) ;
  assign n4146 = n4145 ^ n1018 ^ x121 ;
  assign n4142 = ( n1323 & ~n3254 ) | ( n1323 & n3331 ) | ( ~n3254 & n3331 ) ;
  assign n4143 = ( n855 & n1631 ) | ( n855 & n4142 ) | ( n1631 & n4142 ) ;
  assign n4144 = n2565 | n4143 ;
  assign n4147 = n4146 ^ n4144 ^ 1'b0 ;
  assign n4148 = n1573 ^ n897 ^ x69 ;
  assign n4155 = n3467 ^ n3102 ^ x39 ;
  assign n4156 = n4155 ^ n2535 ^ n2303 ;
  assign n4157 = n4156 ^ n3291 ^ 1'b0 ;
  assign n4158 = ( x225 & n3054 ) | ( x225 & ~n4157 ) | ( n3054 & ~n4157 ) ;
  assign n4149 = n1325 | n2956 ;
  assign n4150 = ( x194 & ~n475 ) | ( x194 & n1580 ) | ( ~n475 & n1580 ) ;
  assign n4151 = ( n3363 & n4149 ) | ( n3363 & ~n4150 ) | ( n4149 & ~n4150 ) ;
  assign n4152 = n4151 ^ n1935 ^ 1'b0 ;
  assign n4153 = ( n1984 & n2901 ) | ( n1984 & n4152 ) | ( n2901 & n4152 ) ;
  assign n4154 = n299 | n4153 ;
  assign n4159 = n4158 ^ n4154 ^ 1'b0 ;
  assign n4172 = ( x81 & n294 ) | ( x81 & ~n296 ) | ( n294 & ~n296 ) ;
  assign n4173 = ~n1337 & n2582 ;
  assign n4174 = n4173 ^ n2359 ^ 1'b0 ;
  assign n4175 = n4172 | n4174 ;
  assign n4176 = n3646 & ~n4175 ;
  assign n4177 = ( ~x140 & n1975 ) | ( ~x140 & n3410 ) | ( n1975 & n3410 ) ;
  assign n4178 = ( n1975 & n4176 ) | ( n1975 & n4177 ) | ( n4176 & n4177 ) ;
  assign n4160 = n2703 ^ n2628 ^ x107 ;
  assign n4161 = ( n548 & n2278 ) | ( n548 & ~n4160 ) | ( n2278 & ~n4160 ) ;
  assign n4162 = n4161 ^ n2879 ^ n770 ;
  assign n4163 = ( n775 & n1399 ) | ( n775 & ~n1885 ) | ( n1399 & ~n1885 ) ;
  assign n4164 = n4163 ^ n2309 ^ n623 ;
  assign n4165 = n4164 ^ n2543 ^ n2516 ;
  assign n4166 = n836 ^ n602 ^ n500 ;
  assign n4167 = ( n868 & n3629 ) | ( n868 & n4166 ) | ( n3629 & n4166 ) ;
  assign n4168 = n2715 ^ n410 ^ x251 ;
  assign n4169 = ~n1186 & n4168 ;
  assign n4170 = ( n4165 & ~n4167 ) | ( n4165 & n4169 ) | ( ~n4167 & n4169 ) ;
  assign n4171 = n4162 & ~n4170 ;
  assign n4179 = n4178 ^ n4171 ^ 1'b0 ;
  assign n4180 = ( n654 & n729 ) | ( n654 & n1224 ) | ( n729 & n1224 ) ;
  assign n4181 = n4180 ^ n1808 ^ 1'b0 ;
  assign n4182 = n4181 ^ n981 ^ 1'b0 ;
  assign n4183 = ( ~n576 & n1461 ) | ( ~n576 & n2301 ) | ( n1461 & n2301 ) ;
  assign n4184 = n1898 ^ n1112 ^ n1080 ;
  assign n4185 = n3354 & n4184 ;
  assign n4186 = n4183 & n4185 ;
  assign n4187 = ( ~n495 & n1629 ) | ( ~n495 & n1976 ) | ( n1629 & n1976 ) ;
  assign n4188 = ( n3094 & n3598 ) | ( n3094 & n4187 ) | ( n3598 & n4187 ) ;
  assign n4189 = ( ~n4182 & n4186 ) | ( ~n4182 & n4188 ) | ( n4186 & n4188 ) ;
  assign n4190 = n4189 ^ n2601 ^ n1291 ;
  assign n4191 = n4142 ^ n2671 ^ n2083 ;
  assign n4192 = n4191 ^ n275 ^ 1'b0 ;
  assign n4195 = n3294 ^ n2140 ^ n1839 ;
  assign n4193 = n387 ^ x198 ^ 1'b0 ;
  assign n4194 = n2637 & ~n4193 ;
  assign n4196 = n4195 ^ n4194 ^ n1103 ;
  assign n4197 = n1845 ^ n1224 ^ n543 ;
  assign n4198 = n3543 ^ n2842 ^ n872 ;
  assign n4199 = n4197 & ~n4198 ;
  assign n4200 = n3534 ^ n2119 ^ n1717 ;
  assign n4201 = ~n3857 & n4200 ;
  assign n4202 = n4201 ^ n3669 ^ 1'b0 ;
  assign n4203 = n1836 & ~n4202 ;
  assign n4204 = x191 & n747 ;
  assign n4205 = n2542 ^ n1867 ^ n1083 ;
  assign n4206 = ( x97 & n639 ) | ( x97 & ~n4205 ) | ( n639 & ~n4205 ) ;
  assign n4207 = ( n2605 & ~n2853 ) | ( n2605 & n4206 ) | ( ~n2853 & n4206 ) ;
  assign n4208 = ( n412 & n4204 ) | ( n412 & ~n4207 ) | ( n4204 & ~n4207 ) ;
  assign n4209 = ( ~n3269 & n3998 ) | ( ~n3269 & n4208 ) | ( n3998 & n4208 ) ;
  assign n4210 = ( n944 & n2090 ) | ( n944 & ~n2852 ) | ( n2090 & ~n2852 ) ;
  assign n4212 = n3564 ^ x118 ^ 1'b0 ;
  assign n4211 = n2089 ^ n259 ^ 1'b0 ;
  assign n4213 = n4212 ^ n4211 ^ n1938 ;
  assign n4214 = ( n2600 & n4210 ) | ( n2600 & ~n4213 ) | ( n4210 & ~n4213 ) ;
  assign n4215 = n4214 ^ n2935 ^ n1091 ;
  assign n4216 = ~n671 & n1075 ;
  assign n4217 = ( n813 & ~n1716 ) | ( n813 & n4216 ) | ( ~n1716 & n4216 ) ;
  assign n4218 = ( n401 & ~n954 ) | ( n401 & n1092 ) | ( ~n954 & n1092 ) ;
  assign n4219 = n4218 ^ n2998 ^ 1'b0 ;
  assign n4220 = n4219 ^ n3812 ^ 1'b0 ;
  assign n4221 = ~n4217 & n4220 ;
  assign n4222 = n3530 ^ n334 ^ x206 ;
  assign n4223 = n400 ^ n354 ^ 1'b0 ;
  assign n4224 = ( n3733 & ~n4222 ) | ( n3733 & n4223 ) | ( ~n4222 & n4223 ) ;
  assign n4232 = n2738 & ~n2993 ;
  assign n4233 = n4232 ^ n2594 ^ 1'b0 ;
  assign n4234 = n4233 ^ n779 ^ n559 ;
  assign n4228 = n689 ^ n634 ^ 1'b0 ;
  assign n4229 = n1834 & ~n4228 ;
  assign n4230 = n4229 ^ n2865 ^ n2630 ;
  assign n4231 = ( n1026 & n4100 ) | ( n1026 & ~n4230 ) | ( n4100 & ~n4230 ) ;
  assign n4225 = ~n260 & n936 ;
  assign n4226 = n4225 ^ n2903 ^ 1'b0 ;
  assign n4227 = n4226 ^ n940 ^ n538 ;
  assign n4235 = n4234 ^ n4231 ^ n4227 ;
  assign n4236 = ( n1063 & ~n2027 ) | ( n1063 & n3143 ) | ( ~n2027 & n3143 ) ;
  assign n4237 = ( n743 & ~n2316 ) | ( n743 & n4236 ) | ( ~n2316 & n4236 ) ;
  assign n4238 = ( ~n2589 & n2720 ) | ( ~n2589 & n4237 ) | ( n2720 & n4237 ) ;
  assign n4239 = ( n3672 & n3687 ) | ( n3672 & ~n4238 ) | ( n3687 & ~n4238 ) ;
  assign n4245 = ( ~n1471 & n2005 ) | ( ~n1471 & n3250 ) | ( n2005 & n3250 ) ;
  assign n4244 = n3395 | n4130 ;
  assign n4240 = n1642 & n1863 ;
  assign n4241 = n4240 ^ n1131 ^ 1'b0 ;
  assign n4242 = n4241 ^ n2721 ^ n1286 ;
  assign n4243 = ( n722 & n3200 ) | ( n722 & ~n4242 ) | ( n3200 & ~n4242 ) ;
  assign n4246 = n4245 ^ n4244 ^ n4243 ;
  assign n4247 = n2491 ^ n1754 ^ n554 ;
  assign n4248 = x149 & n4247 ;
  assign n4249 = n4248 ^ n1425 ^ 1'b0 ;
  assign n4250 = ( n1465 & n2194 ) | ( n1465 & ~n2197 ) | ( n2194 & ~n2197 ) ;
  assign n4251 = ( n2310 & n2831 ) | ( n2310 & n3686 ) | ( n2831 & n3686 ) ;
  assign n4253 = ( n407 & n1784 ) | ( n407 & n2567 ) | ( n1784 & n2567 ) ;
  assign n4252 = n3610 ^ n3568 ^ n2180 ;
  assign n4254 = n4253 ^ n4252 ^ n3243 ;
  assign n4255 = n4254 ^ n3831 ^ n1939 ;
  assign n4258 = x7 & n3756 ;
  assign n4256 = ( x171 & ~n2350 ) | ( x171 & n2605 ) | ( ~n2350 & n2605 ) ;
  assign n4257 = ( n1229 & n2094 ) | ( n1229 & n4256 ) | ( n2094 & n4256 ) ;
  assign n4259 = n4258 ^ n4257 ^ 1'b0 ;
  assign n4260 = x152 & ~n4259 ;
  assign n4261 = n2231 ^ x194 ^ x166 ;
  assign n4262 = n2769 | n4261 ;
  assign n4263 = n698 & n915 ;
  assign n4264 = ~n666 & n4263 ;
  assign n4265 = ( n2851 & ~n4179 ) | ( n2851 & n4264 ) | ( ~n4179 & n4264 ) ;
  assign n4266 = n2838 ^ n1634 ^ 1'b0 ;
  assign n4267 = x12 & n4266 ;
  assign n4268 = n803 & n4267 ;
  assign n4269 = n4268 ^ n1105 ^ 1'b0 ;
  assign n4270 = n3893 ^ n2183 ^ 1'b0 ;
  assign n4271 = n1376 & n4270 ;
  assign n4272 = n681 ^ n294 ^ 1'b0 ;
  assign n4273 = ( n353 & ~n2875 ) | ( n353 & n3196 ) | ( ~n2875 & n3196 ) ;
  assign n4274 = ( n1170 & ~n2939 ) | ( n1170 & n4253 ) | ( ~n2939 & n4253 ) ;
  assign n4275 = ( n4231 & n4273 ) | ( n4231 & ~n4274 ) | ( n4273 & ~n4274 ) ;
  assign n4276 = ( n338 & n4272 ) | ( n338 & ~n4275 ) | ( n4272 & ~n4275 ) ;
  assign n4277 = n2713 ^ n1205 ^ x25 ;
  assign n4278 = n4066 & n4277 ;
  assign n4279 = n4278 ^ x64 ^ 1'b0 ;
  assign n4280 = n3705 & n4279 ;
  assign n4281 = n2459 ^ n2312 ^ x82 ;
  assign n4282 = n4281 ^ n1250 ^ n680 ;
  assign n4283 = n2038 ^ n1605 ^ n1039 ;
  assign n4284 = n3044 & ~n4283 ;
  assign n4285 = n4284 ^ n1050 ^ 1'b0 ;
  assign n4286 = ( n1175 & ~n2701 ) | ( n1175 & n2857 ) | ( ~n2701 & n2857 ) ;
  assign n4287 = ( n3275 & n4285 ) | ( n3275 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4288 = n2078 ^ n1541 ^ 1'b0 ;
  assign n4289 = n1753 & n3004 ;
  assign n4290 = n2664 & ~n4289 ;
  assign n4291 = n1132 & ~n2248 ;
  assign n4292 = n4291 ^ n1262 ^ 1'b0 ;
  assign n4293 = n3326 ^ n1814 ^ n1390 ;
  assign n4294 = n2516 ^ n1812 ^ x145 ;
  assign n4295 = ( n3328 & ~n3454 ) | ( n3328 & n4294 ) | ( ~n3454 & n4294 ) ;
  assign n4296 = ( n320 & n1225 ) | ( n320 & n1747 ) | ( n1225 & n1747 ) ;
  assign n4297 = n1692 & n4296 ;
  assign n4298 = n4297 ^ n1246 ^ 1'b0 ;
  assign n4299 = n766 | n1111 ;
  assign n4300 = ( n752 & ~n2115 ) | ( n752 & n2966 ) | ( ~n2115 & n2966 ) ;
  assign n4301 = ( n4298 & ~n4299 ) | ( n4298 & n4300 ) | ( ~n4299 & n4300 ) ;
  assign n4302 = n4301 ^ n3178 ^ 1'b0 ;
  assign n4303 = n4295 & n4302 ;
  assign n4304 = n1518 ^ n914 ^ n270 ;
  assign n4305 = ( n495 & n620 ) | ( n495 & ~n1266 ) | ( n620 & ~n1266 ) ;
  assign n4306 = n4305 ^ n696 ^ n350 ;
  assign n4307 = n661 ^ x103 ^ x96 ;
  assign n4308 = ( n4304 & n4306 ) | ( n4304 & n4307 ) | ( n4306 & n4307 ) ;
  assign n4309 = ( n374 & ~n745 ) | ( n374 & n944 ) | ( ~n745 & n944 ) ;
  assign n4310 = ( n2718 & ~n3778 ) | ( n2718 & n4309 ) | ( ~n3778 & n4309 ) ;
  assign n4311 = n4310 ^ n2257 ^ x248 ;
  assign n4312 = ( n2564 & n4308 ) | ( n2564 & n4311 ) | ( n4308 & n4311 ) ;
  assign n4313 = n3028 ^ n2686 ^ n1464 ;
  assign n4314 = ( n2147 & ~n2734 ) | ( n2147 & n3476 ) | ( ~n2734 & n3476 ) ;
  assign n4315 = ( n869 & n1487 ) | ( n869 & n2400 ) | ( n1487 & n2400 ) ;
  assign n4316 = n905 & ~n1408 ;
  assign n4317 = ~n3319 & n4316 ;
  assign n4318 = n4317 ^ n649 ^ 1'b0 ;
  assign n4319 = ( n3753 & n4315 ) | ( n3753 & ~n4318 ) | ( n4315 & ~n4318 ) ;
  assign n4320 = ( n4313 & ~n4314 ) | ( n4313 & n4319 ) | ( ~n4314 & n4319 ) ;
  assign n4326 = n3546 ^ n732 ^ 1'b0 ;
  assign n4327 = n611 & n4326 ;
  assign n4328 = ( ~n844 & n2232 ) | ( ~n844 & n4327 ) | ( n2232 & n4327 ) ;
  assign n4324 = ( n1408 & n1881 ) | ( n1408 & n3287 ) | ( n1881 & n3287 ) ;
  assign n4325 = ( n882 & ~n3990 ) | ( n882 & n4324 ) | ( ~n3990 & n4324 ) ;
  assign n4322 = n4229 ^ n1956 ^ n1842 ;
  assign n4321 = n4267 ^ n1257 ^ 1'b0 ;
  assign n4323 = n4322 ^ n4321 ^ n2358 ;
  assign n4329 = n4328 ^ n4325 ^ n4323 ;
  assign n4330 = ( ~x17 & n2010 ) | ( ~x17 & n2068 ) | ( n2010 & n2068 ) ;
  assign n4331 = n2114 | n4330 ;
  assign n4332 = n4331 ^ n1568 ^ 1'b0 ;
  assign n4333 = n4332 ^ n2782 ^ n1714 ;
  assign n4334 = ( n479 & n2119 ) | ( n479 & ~n3889 ) | ( n2119 & ~n3889 ) ;
  assign n4335 = n2395 ^ n1854 ^ n1178 ;
  assign n4336 = ( n1097 & n3921 ) | ( n1097 & n4335 ) | ( n3921 & n4335 ) ;
  assign n4337 = ~n1067 & n2786 ;
  assign n4338 = ( n625 & ~n2641 ) | ( n625 & n4337 ) | ( ~n2641 & n4337 ) ;
  assign n4339 = n904 & ~n4338 ;
  assign n4340 = ~n3087 & n4339 ;
  assign n4341 = ( ~n3733 & n3861 ) | ( ~n3733 & n4340 ) | ( n3861 & n4340 ) ;
  assign n4342 = n4341 ^ n2887 ^ 1'b0 ;
  assign n4343 = n4336 & n4342 ;
  assign n4344 = ( n4030 & n4334 ) | ( n4030 & n4343 ) | ( n4334 & n4343 ) ;
  assign n4346 = n3130 ^ n1667 ^ 1'b0 ;
  assign n4347 = ~n1828 & n4346 ;
  assign n4345 = x238 | n3864 ;
  assign n4348 = n4347 ^ n4345 ^ n968 ;
  assign n4349 = ( n1352 & ~n3331 ) | ( n1352 & n4348 ) | ( ~n3331 & n4348 ) ;
  assign n4350 = ( n330 & n823 ) | ( n330 & n2192 ) | ( n823 & n2192 ) ;
  assign n4351 = n1264 & ~n2240 ;
  assign n4352 = n4350 | n4351 ;
  assign n4366 = ( n687 & n1256 ) | ( n687 & n3265 ) | ( n1256 & n3265 ) ;
  assign n4353 = ~n1040 & n2251 ;
  assign n4354 = ( n1999 & n2809 ) | ( n1999 & n4353 ) | ( n2809 & n4353 ) ;
  assign n4355 = n2237 ^ n436 ^ 1'b0 ;
  assign n4358 = ( x67 & ~n369 ) | ( x67 & n966 ) | ( ~n369 & n966 ) ;
  assign n4357 = n3514 ^ n2099 ^ n359 ;
  assign n4356 = n2723 ^ n2089 ^ n1785 ;
  assign n4359 = n4358 ^ n4357 ^ n4356 ;
  assign n4360 = ( n4354 & n4355 ) | ( n4354 & ~n4359 ) | ( n4355 & ~n4359 ) ;
  assign n4361 = ( x197 & n2680 ) | ( x197 & ~n4360 ) | ( n2680 & ~n4360 ) ;
  assign n4362 = n3785 ^ n2097 ^ n1558 ;
  assign n4363 = n1447 & ~n4362 ;
  assign n4364 = ~n3262 & n4363 ;
  assign n4365 = ( ~n2197 & n4361 ) | ( ~n2197 & n4364 ) | ( n4361 & n4364 ) ;
  assign n4367 = n4366 ^ n4365 ^ 1'b0 ;
  assign n4368 = n1868 | n4367 ;
  assign n4369 = ( n854 & n1755 ) | ( n854 & n4368 ) | ( n1755 & n4368 ) ;
  assign n4370 = n3137 ^ x57 ^ 1'b0 ;
  assign n4371 = n735 & ~n1713 ;
  assign n4372 = n4371 ^ n1317 ^ x116 ;
  assign n4373 = ( ~n1919 & n2849 ) | ( ~n1919 & n4130 ) | ( n2849 & n4130 ) ;
  assign n4374 = ( ~n1546 & n3892 ) | ( ~n1546 & n4373 ) | ( n3892 & n4373 ) ;
  assign n4375 = ( n716 & n1580 ) | ( n716 & n4099 ) | ( n1580 & n4099 ) ;
  assign n4376 = ( n2165 & ~n2437 ) | ( n2165 & n2485 ) | ( ~n2437 & n2485 ) ;
  assign n4377 = ~n1808 & n4376 ;
  assign n4378 = n4377 ^ n1102 ^ 1'b0 ;
  assign n4379 = ( n2331 & n4375 ) | ( n2331 & n4378 ) | ( n4375 & n4378 ) ;
  assign n4380 = n3215 ^ n2475 ^ 1'b0 ;
  assign n4381 = n4379 & ~n4380 ;
  assign n4382 = n4381 ^ n3766 ^ x142 ;
  assign n4383 = n2850 ^ x183 ^ 1'b0 ;
  assign n4384 = n1712 | n3536 ;
  assign n4385 = n3606 ^ n3265 ^ 1'b0 ;
  assign n4386 = ( n4383 & n4384 ) | ( n4383 & ~n4385 ) | ( n4384 & ~n4385 ) ;
  assign n4387 = n1715 ^ n1173 ^ 1'b0 ;
  assign n4388 = n614 & n4387 ;
  assign n4389 = ( ~x98 & x207 ) | ( ~x98 & n4388 ) | ( x207 & n4388 ) ;
  assign n4390 = n4389 ^ n547 ^ 1'b0 ;
  assign n4391 = n4386 & n4390 ;
  assign n4393 = n2923 ^ x220 ^ 1'b0 ;
  assign n4394 = n1404 & n4393 ;
  assign n4392 = n4217 ^ n1276 ^ n756 ;
  assign n4395 = n4394 ^ n4392 ^ 1'b0 ;
  assign n4396 = n4395 ^ n2237 ^ n1221 ;
  assign n4397 = ( n2063 & n4085 ) | ( n2063 & ~n4396 ) | ( n4085 & ~n4396 ) ;
  assign n4398 = x25 | n1605 ;
  assign n4402 = n1921 & n2406 ;
  assign n4403 = n529 & n4402 ;
  assign n4399 = ( ~n1366 & n2250 ) | ( ~n1366 & n2687 ) | ( n2250 & n2687 ) ;
  assign n4400 = n3137 | n4399 ;
  assign n4401 = n4109 | n4400 ;
  assign n4404 = n4403 ^ n4401 ^ n3029 ;
  assign n4405 = ( x130 & x212 ) | ( x130 & ~n1815 ) | ( x212 & ~n1815 ) ;
  assign n4406 = n4405 ^ n3701 ^ n1920 ;
  assign n4407 = ~n973 & n4406 ;
  assign n4411 = ~n500 & n4304 ;
  assign n4409 = ( n1191 & n1253 ) | ( n1191 & n1705 ) | ( n1253 & n1705 ) ;
  assign n4408 = n356 & n1967 ;
  assign n4410 = n4409 ^ n4408 ^ n713 ;
  assign n4412 = n4411 ^ n4410 ^ n861 ;
  assign n4413 = n4412 ^ n4321 ^ n1075 ;
  assign n4414 = n2631 ^ n891 ^ 1'b0 ;
  assign n4415 = ( n1647 & ~n2801 ) | ( n1647 & n4338 ) | ( ~n2801 & n4338 ) ;
  assign n4416 = n1856 ^ n445 ^ 1'b0 ;
  assign n4417 = n4415 | n4416 ;
  assign n4418 = ( n1418 & n4414 ) | ( n1418 & n4417 ) | ( n4414 & n4417 ) ;
  assign n4419 = n1464 ^ x163 ^ 1'b0 ;
  assign n4420 = n4419 ^ n3500 ^ n1200 ;
  assign n4421 = ( n1238 & ~n2451 ) | ( n1238 & n3841 ) | ( ~n2451 & n3841 ) ;
  assign n4427 = n1940 ^ n1770 ^ n732 ;
  assign n4428 = n4427 ^ n703 ^ x252 ;
  assign n4422 = ( n1169 & ~n1600 ) | ( n1169 & n1865 ) | ( ~n1600 & n1865 ) ;
  assign n4423 = n2227 | n4422 ;
  assign n4424 = n2593 ^ x72 ^ x26 ;
  assign n4425 = n4424 ^ n3056 ^ n1392 ;
  assign n4426 = ( n3926 & ~n4423 ) | ( n3926 & n4425 ) | ( ~n4423 & n4425 ) ;
  assign n4429 = n4428 ^ n4426 ^ n506 ;
  assign n4444 = n3749 ^ n2582 ^ n1583 ;
  assign n4445 = n4444 ^ n1253 ^ 1'b0 ;
  assign n4446 = n1634 & n4445 ;
  assign n4447 = n4446 ^ n3405 ^ n2358 ;
  assign n4448 = ( ~x55 & n307 ) | ( ~x55 & n4447 ) | ( n307 & n4447 ) ;
  assign n4430 = ( n582 & ~n977 ) | ( n582 & n1845 ) | ( ~n977 & n1845 ) ;
  assign n4431 = n4430 ^ n3212 ^ n914 ;
  assign n4439 = ( ~x214 & n794 ) | ( ~x214 & n2070 ) | ( n794 & n2070 ) ;
  assign n4432 = ( ~x142 & x203 ) | ( ~x142 & n1181 ) | ( x203 & n1181 ) ;
  assign n4433 = ( n642 & ~n964 ) | ( n642 & n4432 ) | ( ~n964 & n4432 ) ;
  assign n4434 = n4433 ^ n846 ^ x40 ;
  assign n4435 = n528 & n734 ;
  assign n4436 = n4435 ^ n1573 ^ 1'b0 ;
  assign n4437 = ( n2871 & n4434 ) | ( n2871 & ~n4436 ) | ( n4434 & ~n4436 ) ;
  assign n4438 = ~n2825 & n4437 ;
  assign n4440 = n4439 ^ n4438 ^ 1'b0 ;
  assign n4441 = ( n518 & n951 ) | ( n518 & n4440 ) | ( n951 & n4440 ) ;
  assign n4442 = ~n4431 & n4441 ;
  assign n4443 = ~n3724 & n4442 ;
  assign n4449 = n4448 ^ n4443 ^ 1'b0 ;
  assign n4450 = n1560 & ~n4449 ;
  assign n4463 = n2929 ^ n1597 ^ n784 ;
  assign n4451 = n2399 | n2900 ;
  assign n4452 = n4451 ^ n2849 ^ 1'b0 ;
  assign n4455 = n2782 ^ n2324 ^ n397 ;
  assign n4456 = n977 & ~n4455 ;
  assign n4457 = n4456 ^ n1268 ^ 1'b0 ;
  assign n4458 = ( n699 & n2626 ) | ( n699 & ~n4457 ) | ( n2626 & ~n4457 ) ;
  assign n4459 = ( x236 & n2692 ) | ( x236 & ~n4458 ) | ( n2692 & ~n4458 ) ;
  assign n4453 = ~x75 & n505 ;
  assign n4454 = n4453 ^ n3106 ^ n2626 ;
  assign n4460 = n4459 ^ n4454 ^ 1'b0 ;
  assign n4461 = n4460 ^ n2976 ^ 1'b0 ;
  assign n4462 = n4452 & n4461 ;
  assign n4464 = n4463 ^ n4462 ^ 1'b0 ;
  assign n4465 = ( ~n528 & n3750 ) | ( ~n528 & n4122 ) | ( n3750 & n4122 ) ;
  assign n4466 = ( ~n556 & n1316 ) | ( ~n556 & n4465 ) | ( n1316 & n4465 ) ;
  assign n4467 = ( n785 & n1296 ) | ( n785 & n3079 ) | ( n1296 & n3079 ) ;
  assign n4468 = ( n1033 & n3057 ) | ( n1033 & n3170 ) | ( n3057 & n3170 ) ;
  assign n4469 = ( ~x38 & n1976 ) | ( ~x38 & n2120 ) | ( n1976 & n2120 ) ;
  assign n4470 = n1501 ^ n1030 ^ 1'b0 ;
  assign n4471 = n472 & n4470 ;
  assign n4472 = ( ~n1854 & n4469 ) | ( ~n1854 & n4471 ) | ( n4469 & n4471 ) ;
  assign n4477 = ~n794 & n1146 ;
  assign n4478 = ~x126 & n4477 ;
  assign n4475 = n1937 ^ n1566 ^ 1'b0 ;
  assign n4476 = ~n1594 & n4475 ;
  assign n4473 = n2747 ^ n552 ^ n312 ;
  assign n4474 = n403 & n4473 ;
  assign n4479 = n4478 ^ n4476 ^ n4474 ;
  assign n4480 = n308 & n1495 ;
  assign n4481 = n660 & n4480 ;
  assign n4482 = ( ~n2102 & n3136 ) | ( ~n2102 & n4481 ) | ( n3136 & n4481 ) ;
  assign n4483 = n784 & ~n2005 ;
  assign n4484 = n1312 & n4483 ;
  assign n4485 = n4484 ^ n4359 ^ n1207 ;
  assign n4486 = n1284 & ~n1919 ;
  assign n4487 = n4485 & n4486 ;
  assign n4488 = ( n2895 & ~n4482 ) | ( n2895 & n4487 ) | ( ~n4482 & n4487 ) ;
  assign n4489 = ~n698 & n1284 ;
  assign n4492 = n540 ^ x128 ^ 1'b0 ;
  assign n4493 = x49 & n4492 ;
  assign n4494 = ( n2590 & ~n3315 ) | ( n2590 & n4493 ) | ( ~n3315 & n4493 ) ;
  assign n4495 = n4494 ^ n2316 ^ 1'b0 ;
  assign n4496 = n1644 | n4495 ;
  assign n4490 = n413 ^ x39 ^ 1'b0 ;
  assign n4491 = n1133 & ~n4490 ;
  assign n4497 = n4496 ^ n4491 ^ n2000 ;
  assign n4498 = ( n613 & n4489 ) | ( n613 & n4497 ) | ( n4489 & n4497 ) ;
  assign n4499 = n2150 & n4366 ;
  assign n4500 = n4499 ^ n1514 ^ 1'b0 ;
  assign n4501 = n3490 ^ n894 ^ 1'b0 ;
  assign n4502 = n2815 & ~n4501 ;
  assign n4503 = n4502 ^ n3163 ^ n1534 ;
  assign n4504 = n753 ^ n630 ^ 1'b0 ;
  assign n4505 = n1606 & ~n4504 ;
  assign n4506 = ( ~n2243 & n3454 ) | ( ~n2243 & n4505 ) | ( n3454 & n4505 ) ;
  assign n4507 = n601 | n999 ;
  assign n4508 = n2790 | n4507 ;
  assign n4515 = n3445 ^ n2665 ^ n1492 ;
  assign n4510 = n3241 & n4168 ;
  assign n4511 = n4510 ^ x90 ^ 1'b0 ;
  assign n4512 = n688 | n4511 ;
  assign n4509 = ( n343 & n2041 ) | ( n343 & n2867 ) | ( n2041 & n2867 ) ;
  assign n4513 = n4512 ^ n4509 ^ n692 ;
  assign n4514 = ~n3204 & n4513 ;
  assign n4516 = n4515 ^ n4514 ^ 1'b0 ;
  assign n4517 = ( n4155 & ~n4508 ) | ( n4155 & n4516 ) | ( ~n4508 & n4516 ) ;
  assign n4518 = n4517 ^ n3281 ^ 1'b0 ;
  assign n4519 = n1758 & ~n3837 ;
  assign n4520 = n4519 ^ n3077 ^ 1'b0 ;
  assign n4521 = n1924 ^ n784 ^ x171 ;
  assign n4522 = n3578 & n4521 ;
  assign n4523 = n4522 ^ n2291 ^ 1'b0 ;
  assign n4524 = ( n840 & ~n4520 ) | ( n840 & n4523 ) | ( ~n4520 & n4523 ) ;
  assign n4525 = n4524 ^ n3208 ^ n3064 ;
  assign n4526 = n3298 ^ n2706 ^ n2568 ;
  assign n4527 = n4526 ^ n893 ^ 1'b0 ;
  assign n4528 = n1984 & ~n4527 ;
  assign n4529 = n3784 ^ n1822 ^ 1'b0 ;
  assign n4530 = ( n393 & ~n1168 ) | ( n393 & n2606 ) | ( ~n1168 & n2606 ) ;
  assign n4531 = n3345 ^ n2823 ^ n1829 ;
  assign n4532 = n4124 | n4531 ;
  assign n4533 = n4532 ^ n2981 ^ 1'b0 ;
  assign n4534 = ( n4179 & n4530 ) | ( n4179 & ~n4533 ) | ( n4530 & ~n4533 ) ;
  assign n4535 = ( ~n1937 & n1960 ) | ( ~n1937 & n3726 ) | ( n1960 & n3726 ) ;
  assign n4536 = n1810 ^ n1558 ^ x0 ;
  assign n4537 = ( ~n817 & n2427 ) | ( ~n817 & n4536 ) | ( n2427 & n4536 ) ;
  assign n4538 = ( n2432 & n3355 ) | ( n2432 & ~n4537 ) | ( n3355 & ~n4537 ) ;
  assign n4539 = ( n4311 & n4535 ) | ( n4311 & n4538 ) | ( n4535 & n4538 ) ;
  assign n4540 = n4539 ^ n4415 ^ n1896 ;
  assign n4541 = n1645 ^ n1448 ^ n1197 ;
  assign n4542 = n2476 & ~n4541 ;
  assign n4543 = ~n3614 & n4542 ;
  assign n4548 = n2082 ^ n629 ^ 1'b0 ;
  assign n4549 = n900 | n4548 ;
  assign n4550 = ( n1476 & ~n2553 ) | ( n1476 & n4549 ) | ( ~n2553 & n4549 ) ;
  assign n4544 = ( n1778 & n2159 ) | ( n1778 & ~n2981 ) | ( n2159 & ~n2981 ) ;
  assign n4545 = n4544 ^ n4108 ^ n2294 ;
  assign n4546 = ( ~n2444 & n4066 ) | ( ~n2444 & n4545 ) | ( n4066 & n4545 ) ;
  assign n4547 = n4546 ^ n3218 ^ n632 ;
  assign n4551 = n4550 ^ n4547 ^ 1'b0 ;
  assign n4552 = ( ~n1153 & n1725 ) | ( ~n1153 & n2256 ) | ( n1725 & n2256 ) ;
  assign n4553 = n4552 ^ n525 ^ 1'b0 ;
  assign n4554 = ( n4543 & ~n4551 ) | ( n4543 & n4553 ) | ( ~n4551 & n4553 ) ;
  assign n4555 = n2324 ^ n1322 ^ 1'b0 ;
  assign n4556 = n1569 | n4555 ;
  assign n4557 = ( n1463 & ~n3944 ) | ( n1463 & n4556 ) | ( ~n3944 & n4556 ) ;
  assign n4558 = n4557 ^ n1848 ^ n1637 ;
  assign n4559 = ( ~n901 & n1369 ) | ( ~n901 & n2382 ) | ( n1369 & n2382 ) ;
  assign n4560 = ( n2172 & n3516 ) | ( n2172 & n4559 ) | ( n3516 & n4559 ) ;
  assign n4561 = ( n552 & ~n4558 ) | ( n552 & n4560 ) | ( ~n4558 & n4560 ) ;
  assign n4565 = ( n620 & ~n923 ) | ( n620 & n1155 ) | ( ~n923 & n1155 ) ;
  assign n4566 = ( n1444 & ~n2901 ) | ( n1444 & n4565 ) | ( ~n2901 & n4565 ) ;
  assign n4562 = ( n708 & n1873 ) | ( n708 & ~n2107 ) | ( n1873 & ~n2107 ) ;
  assign n4563 = n4562 ^ n3176 ^ n2772 ;
  assign n4564 = ( n1246 & n1562 ) | ( n1246 & ~n4563 ) | ( n1562 & ~n4563 ) ;
  assign n4567 = n4566 ^ n4564 ^ n2022 ;
  assign n4568 = ( n987 & ~n1314 ) | ( n987 & n4567 ) | ( ~n1314 & n4567 ) ;
  assign n4569 = n1365 ^ n1015 ^ x175 ;
  assign n4570 = ( x0 & ~n3528 ) | ( x0 & n4569 ) | ( ~n3528 & n4569 ) ;
  assign n4571 = n1626 | n2943 ;
  assign n4572 = ( n1573 & n2291 ) | ( n1573 & ~n4520 ) | ( n2291 & ~n4520 ) ;
  assign n4573 = ~n931 & n3544 ;
  assign n4574 = ( ~n2735 & n4572 ) | ( ~n2735 & n4573 ) | ( n4572 & n4573 ) ;
  assign n4575 = ( n1394 & ~n4571 ) | ( n1394 & n4574 ) | ( ~n4571 & n4574 ) ;
  assign n4577 = x18 & ~n1486 ;
  assign n4578 = ( n1288 & n1656 ) | ( n1288 & ~n4577 ) | ( n1656 & ~n4577 ) ;
  assign n4576 = n2686 ^ n1396 ^ n271 ;
  assign n4579 = n4578 ^ n4576 ^ 1'b0 ;
  assign n4580 = n2632 ^ n792 ^ n326 ;
  assign n4581 = n3750 ^ n1996 ^ n302 ;
  assign n4582 = n4581 ^ n3778 ^ n2456 ;
  assign n4583 = n4580 & ~n4582 ;
  assign n4584 = n588 | n680 ;
  assign n4585 = n3533 | n4584 ;
  assign n4586 = n4585 ^ n3725 ^ n1085 ;
  assign n4587 = n827 & n1302 ;
  assign n4588 = n4587 ^ n3041 ^ 1'b0 ;
  assign n4602 = n2956 ^ n1032 ^ 1'b0 ;
  assign n4603 = n391 & n4602 ;
  assign n4604 = ( ~n1155 & n2243 ) | ( ~n1155 & n4603 ) | ( n2243 & n4603 ) ;
  assign n4605 = ( n667 & n2030 ) | ( n667 & n4604 ) | ( n2030 & n4604 ) ;
  assign n4596 = n1797 ^ n846 ^ x12 ;
  assign n4599 = n2459 ^ n1550 ^ n615 ;
  assign n4597 = ( x13 & n463 ) | ( x13 & n1707 ) | ( n463 & n1707 ) ;
  assign n4598 = n4597 ^ n2773 ^ 1'b0 ;
  assign n4600 = n4599 ^ n4598 ^ n4310 ;
  assign n4601 = ( n1406 & n4596 ) | ( n1406 & n4600 ) | ( n4596 & n4600 ) ;
  assign n4606 = n4605 ^ n4601 ^ n1491 ;
  assign n4589 = ( n1355 & ~n1733 ) | ( n1355 & n3129 ) | ( ~n1733 & n3129 ) ;
  assign n4590 = ( n2571 & n4571 ) | ( n2571 & n4589 ) | ( n4571 & n4589 ) ;
  assign n4591 = ~n482 & n891 ;
  assign n4592 = n4591 ^ n3505 ^ 1'b0 ;
  assign n4593 = n1053 & ~n4592 ;
  assign n4594 = n4593 ^ n4020 ^ 1'b0 ;
  assign n4595 = ~n4590 & n4594 ;
  assign n4607 = n4606 ^ n4595 ^ x77 ;
  assign n4608 = n532 & ~n2643 ;
  assign n4609 = ( ~x193 & n374 ) | ( ~x193 & n4608 ) | ( n374 & n4608 ) ;
  assign n4610 = ( n2869 & n4149 ) | ( n2869 & n4609 ) | ( n4149 & n4609 ) ;
  assign n4611 = ~n1778 & n2691 ;
  assign n4612 = ~n1834 & n4611 ;
  assign n4613 = n4612 ^ n3004 ^ x61 ;
  assign n4614 = ( ~n2583 & n4610 ) | ( ~n2583 & n4613 ) | ( n4610 & n4613 ) ;
  assign n4615 = n2231 ^ n1963 ^ 1'b0 ;
  assign n4616 = n1431 & ~n4615 ;
  assign n4617 = n873 & n4164 ;
  assign n4618 = n315 & n4617 ;
  assign n4619 = n3678 ^ n2854 ^ 1'b0 ;
  assign n4620 = ~n4618 & n4619 ;
  assign n4621 = n4620 ^ n1208 ^ 1'b0 ;
  assign n4622 = n4616 & n4621 ;
  assign n4623 = ( n1040 & n1427 ) | ( n1040 & n3713 ) | ( n1427 & n3713 ) ;
  assign n4626 = ~n396 & n3788 ;
  assign n4627 = n4626 ^ n3638 ^ n1749 ;
  assign n4628 = n985 ^ n842 ^ n681 ;
  assign n4629 = ( n296 & n4627 ) | ( n296 & ~n4628 ) | ( n4627 & ~n4628 ) ;
  assign n4624 = ( ~n1047 & n1281 ) | ( ~n1047 & n4075 ) | ( n1281 & n4075 ) ;
  assign n4625 = n4624 ^ n2738 ^ x167 ;
  assign n4630 = n4629 ^ n4625 ^ 1'b0 ;
  assign n4631 = n2294 ^ n897 ^ 1'b0 ;
  assign n4632 = ( x234 & ~n2697 ) | ( x234 & n3246 ) | ( ~n2697 & n3246 ) ;
  assign n4633 = ( ~n1217 & n4631 ) | ( ~n1217 & n4632 ) | ( n4631 & n4632 ) ;
  assign n4641 = n4366 ^ n3626 ^ n1651 ;
  assign n4642 = n4641 ^ n3530 ^ n748 ;
  assign n4639 = n3864 ^ n3361 ^ n706 ;
  assign n4637 = ( x181 & x191 ) | ( x181 & n1238 ) | ( x191 & n1238 ) ;
  assign n4634 = n1446 & n3087 ;
  assign n4635 = n4634 ^ n722 ^ 1'b0 ;
  assign n4636 = ( n1315 & n4218 ) | ( n1315 & ~n4635 ) | ( n4218 & ~n4635 ) ;
  assign n4638 = n4637 ^ n4636 ^ n3878 ;
  assign n4640 = n4639 ^ n4638 ^ x17 ;
  assign n4643 = n4642 ^ n4640 ^ n3249 ;
  assign n4644 = n939 ^ n880 ^ x196 ;
  assign n4645 = n4644 ^ n3317 ^ 1'b0 ;
  assign n4646 = n1567 & n4645 ;
  assign n4647 = ( n695 & ~n1976 ) | ( n695 & n2367 ) | ( ~n1976 & n2367 ) ;
  assign n4648 = n2217 ^ n1165 ^ n1138 ;
  assign n4649 = n654 & n4648 ;
  assign n4650 = n4649 ^ n2863 ^ 1'b0 ;
  assign n4651 = n4650 ^ n1116 ^ n752 ;
  assign n4652 = ( x14 & n3837 ) | ( x14 & n4651 ) | ( n3837 & n4651 ) ;
  assign n4653 = ( x207 & n468 ) | ( x207 & n1294 ) | ( n468 & n1294 ) ;
  assign n4654 = n4653 ^ n2159 ^ n1107 ;
  assign n4655 = n1905 ^ n1080 ^ 1'b0 ;
  assign n4656 = ( ~n4122 & n4654 ) | ( ~n4122 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = ( n1269 & n4652 ) | ( n1269 & n4656 ) | ( n4652 & n4656 ) ;
  assign n4658 = ( ~n2557 & n3861 ) | ( ~n2557 & n4481 ) | ( n3861 & n4481 ) ;
  assign n4659 = ( ~x139 & n827 ) | ( ~x139 & n3022 ) | ( n827 & n3022 ) ;
  assign n4660 = n577 & ~n1737 ;
  assign n4661 = n4660 ^ n3422 ^ 1'b0 ;
  assign n4662 = n4661 ^ n915 ^ x77 ;
  assign n4663 = ( x126 & ~n2604 ) | ( x126 & n3096 ) | ( ~n2604 & n3096 ) ;
  assign n4664 = ( n340 & n2715 ) | ( n340 & n4663 ) | ( n2715 & n4663 ) ;
  assign n4665 = ( n973 & ~n2720 ) | ( n973 & n4664 ) | ( ~n2720 & n4664 ) ;
  assign n4666 = ( n2218 & n2725 ) | ( n2218 & ~n4665 ) | ( n2725 & ~n4665 ) ;
  assign n4667 = ( ~n4659 & n4662 ) | ( ~n4659 & n4666 ) | ( n4662 & n4666 ) ;
  assign n4668 = ( n2090 & n4658 ) | ( n2090 & ~n4667 ) | ( n4658 & ~n4667 ) ;
  assign n4669 = n4353 ^ n3214 ^ n431 ;
  assign n4677 = ( x140 & ~n1377 ) | ( x140 & n4107 ) | ( ~n1377 & n4107 ) ;
  assign n4675 = n4469 ^ n1664 ^ x133 ;
  assign n4676 = n3824 & ~n4675 ;
  assign n4670 = n3120 ^ n2954 ^ n495 ;
  assign n4671 = ( ~n999 & n2087 ) | ( ~n999 & n3733 ) | ( n2087 & n3733 ) ;
  assign n4672 = n2070 & n4671 ;
  assign n4673 = n3204 & n4672 ;
  assign n4674 = ( n891 & n4670 ) | ( n891 & ~n4673 ) | ( n4670 & ~n4673 ) ;
  assign n4678 = n4677 ^ n4676 ^ n4674 ;
  assign n4679 = n3224 & ~n4678 ;
  assign n4680 = n1387 & ~n4549 ;
  assign n4681 = n3808 & n4680 ;
  assign n4688 = ~n400 & n829 ;
  assign n4684 = n1697 ^ n1079 ^ x173 ;
  assign n4682 = n3595 ^ x232 ^ 1'b0 ;
  assign n4683 = ~n1945 & n4682 ;
  assign n4685 = n4684 ^ n4683 ^ n2446 ;
  assign n4686 = n4685 ^ n1839 ^ x189 ;
  assign n4687 = ( x20 & n1876 ) | ( x20 & ~n4686 ) | ( n1876 & ~n4686 ) ;
  assign n4689 = n4688 ^ n4687 ^ n4034 ;
  assign n4705 = n3237 | n4599 ;
  assign n4690 = n1930 ^ n640 ^ x30 ;
  assign n4691 = n3769 ^ n316 ^ 1'b0 ;
  assign n4692 = n2700 & n4691 ;
  assign n4693 = ( n2087 & n4690 ) | ( n2087 & n4692 ) | ( n4690 & n4692 ) ;
  assign n4694 = n4693 ^ n4597 ^ n2795 ;
  assign n4695 = ( x83 & n1951 ) | ( x83 & ~n2839 ) | ( n1951 & ~n2839 ) ;
  assign n4696 = n4695 ^ n1838 ^ 1'b0 ;
  assign n4697 = n4694 | n4696 ;
  assign n4698 = n3544 ^ n733 ^ n727 ;
  assign n4699 = n4698 ^ n1715 ^ n319 ;
  assign n4700 = n4699 ^ n3029 ^ n2000 ;
  assign n4701 = n1398 & n4700 ;
  assign n4702 = ( ~n966 & n1736 ) | ( ~n966 & n2418 ) | ( n1736 & n2418 ) ;
  assign n4703 = ( n3657 & n4701 ) | ( n3657 & ~n4702 ) | ( n4701 & ~n4702 ) ;
  assign n4704 = ( n1200 & n4697 ) | ( n1200 & ~n4703 ) | ( n4697 & ~n4703 ) ;
  assign n4706 = n4705 ^ n4704 ^ n2945 ;
  assign n4718 = n686 ^ n391 ^ 1'b0 ;
  assign n4707 = x230 & n1656 ;
  assign n4708 = n4707 ^ n823 ^ n283 ;
  assign n4711 = n324 & n3324 ;
  assign n4712 = n1726 & n4711 ;
  assign n4713 = ( n1129 & n3421 ) | ( n1129 & ~n4712 ) | ( n3421 & ~n4712 ) ;
  assign n4714 = ( ~n1437 & n1758 ) | ( ~n1437 & n4713 ) | ( n1758 & n4713 ) ;
  assign n4709 = n602 & ~n4544 ;
  assign n4710 = ~x99 & n4709 ;
  assign n4715 = n4714 ^ n4710 ^ n2842 ;
  assign n4716 = ( n781 & n4708 ) | ( n781 & ~n4715 ) | ( n4708 & ~n4715 ) ;
  assign n4717 = ( n689 & n1453 ) | ( n689 & n4716 ) | ( n1453 & n4716 ) ;
  assign n4719 = n4718 ^ n4717 ^ n761 ;
  assign n4720 = n2420 ^ n453 ^ x71 ;
  assign n4721 = n4283 ^ n3754 ^ n2218 ;
  assign n4722 = ( n3557 & ~n4720 ) | ( n3557 & n4721 ) | ( ~n4720 & n4721 ) ;
  assign n4724 = n4248 ^ n3582 ^ n2536 ;
  assign n4725 = n4724 ^ n2396 ^ 1'b0 ;
  assign n4726 = ( ~n1280 & n3454 ) | ( ~n1280 & n4725 ) | ( n3454 & n4725 ) ;
  assign n4723 = n1005 & ~n3837 ;
  assign n4727 = n4726 ^ n4723 ^ 1'b0 ;
  assign n4728 = n2654 | n4234 ;
  assign n4729 = n4728 ^ n1280 ^ 1'b0 ;
  assign n4730 = ( x107 & n1983 ) | ( x107 & n4729 ) | ( n1983 & n4729 ) ;
  assign n4732 = n1174 ^ n829 ^ n337 ;
  assign n4731 = n3601 ^ n3095 ^ n2556 ;
  assign n4733 = n4732 ^ n4731 ^ n2168 ;
  assign n4734 = ( n606 & ~n1690 ) | ( n606 & n4275 ) | ( ~n1690 & n4275 ) ;
  assign n4735 = n2594 ^ n1306 ^ n732 ;
  assign n4736 = n3954 ^ x249 ^ 1'b0 ;
  assign n4737 = n4735 & ~n4736 ;
  assign n4738 = n4737 ^ x159 ^ x118 ;
  assign n4739 = n950 ^ x85 ^ 1'b0 ;
  assign n4742 = x52 & n1175 ;
  assign n4743 = n4742 ^ x127 ^ 1'b0 ;
  assign n4740 = n2317 | n2799 ;
  assign n4741 = n2482 | n4740 ;
  assign n4744 = n4743 ^ n4741 ^ n1044 ;
  assign n4745 = ( ~n286 & n2550 ) | ( ~n286 & n4744 ) | ( n2550 & n4744 ) ;
  assign n4746 = ( ~n2940 & n4511 ) | ( ~n2940 & n4745 ) | ( n4511 & n4745 ) ;
  assign n4753 = n2027 ^ n1840 ^ 1'b0 ;
  assign n4751 = x62 & ~n1208 ;
  assign n4752 = ~x56 & n4751 ;
  assign n4754 = n4753 ^ n4752 ^ n979 ;
  assign n4747 = n2113 ^ n1335 ^ n1194 ;
  assign n4748 = ( ~x101 & n1140 ) | ( ~x101 & n4533 ) | ( n1140 & n4533 ) ;
  assign n4749 = ( ~n511 & n4747 ) | ( ~n511 & n4748 ) | ( n4747 & n4748 ) ;
  assign n4750 = n3340 & n4749 ;
  assign n4755 = n4754 ^ n4750 ^ 1'b0 ;
  assign n4756 = ( ~n4739 & n4746 ) | ( ~n4739 & n4755 ) | ( n4746 & n4755 ) ;
  assign n4757 = n4151 ^ n1840 ^ n1240 ;
  assign n4758 = n3260 | n4757 ;
  assign n4760 = n1791 ^ n296 ^ 1'b0 ;
  assign n4761 = ( n788 & n2530 ) | ( n788 & n3284 ) | ( n2530 & n3284 ) ;
  assign n4762 = ( n3678 & n3783 ) | ( n3678 & ~n4761 ) | ( n3783 & ~n4761 ) ;
  assign n4763 = ( n689 & n4760 ) | ( n689 & ~n4762 ) | ( n4760 & ~n4762 ) ;
  assign n4759 = ~n1212 & n1591 ;
  assign n4764 = n4763 ^ n4759 ^ x154 ;
  assign n4774 = n1545 ^ n867 ^ n286 ;
  assign n4775 = ( n1856 & n2923 ) | ( n1856 & n4774 ) | ( n2923 & n4774 ) ;
  assign n4766 = n1798 ^ n933 ^ 1'b0 ;
  assign n4767 = n629 & n4766 ;
  assign n4765 = ( n624 & n645 ) | ( n624 & n1684 ) | ( n645 & n1684 ) ;
  assign n4768 = n4767 ^ n4765 ^ n2042 ;
  assign n4769 = n3327 ^ n2649 ^ n1405 ;
  assign n4770 = ( n427 & n1706 ) | ( n427 & ~n4769 ) | ( n1706 & ~n4769 ) ;
  assign n4771 = ( n936 & n4187 ) | ( n936 & n4604 ) | ( n4187 & n4604 ) ;
  assign n4772 = n4771 ^ n3027 ^ n1814 ;
  assign n4773 = ( n4768 & n4770 ) | ( n4768 & n4772 ) | ( n4770 & n4772 ) ;
  assign n4776 = n4775 ^ n4773 ^ 1'b0 ;
  assign n4777 = x166 & n4776 ;
  assign n4780 = n2564 ^ n439 ^ 1'b0 ;
  assign n4778 = ( ~n2587 & n3556 ) | ( ~n2587 & n4552 ) | ( n3556 & n4552 ) ;
  assign n4779 = n4778 ^ n1709 ^ 1'b0 ;
  assign n4781 = n4780 ^ n4779 ^ n1427 ;
  assign n4782 = n1391 ^ n276 ^ 1'b0 ;
  assign n4783 = n970 | n4782 ;
  assign n4784 = ( n272 & n770 ) | ( n272 & ~n2388 ) | ( n770 & ~n2388 ) ;
  assign n4785 = n4784 ^ n2975 ^ x153 ;
  assign n4786 = n4785 ^ n1371 ^ 1'b0 ;
  assign n4787 = ~n3052 & n4786 ;
  assign n4788 = n2060 & n3306 ;
  assign n4789 = ( n4783 & ~n4787 ) | ( n4783 & n4788 ) | ( ~n4787 & n4788 ) ;
  assign n4790 = n3645 & n4314 ;
  assign n4791 = n4789 & n4790 ;
  assign n4792 = n4791 ^ n4730 ^ x32 ;
  assign n4793 = ( n2294 & n2474 ) | ( n2294 & n3706 ) | ( n2474 & n3706 ) ;
  assign n4794 = ( n1771 & ~n4060 ) | ( n1771 & n4793 ) | ( ~n4060 & n4793 ) ;
  assign n4795 = n4794 ^ n2937 ^ n720 ;
  assign n4797 = n1414 ^ n727 ^ 1'b0 ;
  assign n4798 = n4797 ^ n1618 ^ n366 ;
  assign n4796 = n1320 & n2705 ;
  assign n4799 = n4798 ^ n4796 ^ 1'b0 ;
  assign n4801 = n3572 ^ n854 ^ 1'b0 ;
  assign n4802 = n4801 ^ n1897 ^ n1746 ;
  assign n4800 = n2733 | n3065 ;
  assign n4803 = n4802 ^ n4800 ^ 1'b0 ;
  assign n4804 = ( ~n4780 & n4799 ) | ( ~n4780 & n4803 ) | ( n4799 & n4803 ) ;
  assign n4805 = n3087 ^ n1857 ^ 1'b0 ;
  assign n4806 = n1642 & ~n4805 ;
  assign n4807 = n1173 | n1549 ;
  assign n4808 = ( ~n2509 & n4806 ) | ( ~n2509 & n4807 ) | ( n4806 & n4807 ) ;
  assign n4809 = n1022 & ~n4808 ;
  assign n4817 = ~n1504 & n4745 ;
  assign n4810 = ( n428 & ~n1787 ) | ( n428 & n3743 ) | ( ~n1787 & n3743 ) ;
  assign n4811 = n567 | n3422 ;
  assign n4812 = n4811 ^ n619 ^ 1'b0 ;
  assign n4813 = n4812 ^ x233 ^ 1'b0 ;
  assign n4814 = n4810 & n4813 ;
  assign n4815 = n3995 | n4814 ;
  assign n4816 = n4815 ^ n732 ^ 1'b0 ;
  assign n4818 = n4817 ^ n4816 ^ n3157 ;
  assign n4821 = ( ~n2726 & n3069 ) | ( ~n2726 & n4020 ) | ( n3069 & n4020 ) ;
  assign n4822 = ( n814 & n2953 ) | ( n814 & ~n4821 ) | ( n2953 & ~n4821 ) ;
  assign n4819 = n2824 & ~n3939 ;
  assign n4820 = ~x156 & n4819 ;
  assign n4823 = n4822 ^ n4820 ^ n492 ;
  assign n4824 = n4823 ^ n4066 ^ x137 ;
  assign n4825 = n4824 ^ n3392 ^ n1451 ;
  assign n4833 = n380 & n472 ;
  assign n4831 = n1128 & n3205 ;
  assign n4832 = n4831 ^ n3687 ^ 1'b0 ;
  assign n4826 = ~n423 & n2313 ;
  assign n4827 = ~n753 & n4826 ;
  assign n4828 = ( ~n357 & n805 ) | ( ~n357 & n4827 ) | ( n805 & n4827 ) ;
  assign n4829 = ~n606 & n4828 ;
  assign n4830 = ~n2651 & n4829 ;
  assign n4834 = n4833 ^ n4832 ^ n4830 ;
  assign n4835 = ( x254 & n1676 ) | ( x254 & n2302 ) | ( n1676 & n2302 ) ;
  assign n4836 = n4835 ^ n3488 ^ n2396 ;
  assign n4837 = ( ~n2575 & n2703 ) | ( ~n2575 & n4836 ) | ( n2703 & n4836 ) ;
  assign n4838 = ~n1644 & n4837 ;
  assign n4839 = n4838 ^ n2363 ^ 1'b0 ;
  assign n4841 = ~n334 & n2289 ;
  assign n4840 = ( n635 & n1191 ) | ( n635 & ~n3025 ) | ( n1191 & ~n3025 ) ;
  assign n4842 = n4841 ^ n4840 ^ n301 ;
  assign n4846 = ( ~n1042 & n3778 ) | ( ~n1042 & n4708 ) | ( n3778 & n4708 ) ;
  assign n4847 = n2441 ^ x120 ^ x13 ;
  assign n4848 = ~n812 & n4847 ;
  assign n4849 = n4848 ^ n1644 ^ 1'b0 ;
  assign n4850 = n4849 ^ n2362 ^ n1830 ;
  assign n4851 = ( n4130 & n4846 ) | ( n4130 & n4850 ) | ( n4846 & n4850 ) ;
  assign n4843 = ( ~x227 & n2018 ) | ( ~x227 & n3749 ) | ( n2018 & n3749 ) ;
  assign n4844 = ( n1082 & ~n4309 ) | ( n1082 & n4843 ) | ( ~n4309 & n4843 ) ;
  assign n4845 = n4844 ^ n3533 ^ 1'b0 ;
  assign n4852 = n4851 ^ n4845 ^ n4708 ;
  assign n4853 = ( n1734 & n1828 ) | ( n1734 & n3006 ) | ( n1828 & n3006 ) ;
  assign n4854 = n4853 ^ n471 ^ x56 ;
  assign n4855 = n710 & ~n774 ;
  assign n4856 = n4403 & n4855 ;
  assign n4857 = n4181 | n4856 ;
  assign n4858 = n3675 ^ n2412 ^ n632 ;
  assign n4862 = n1939 ^ n1564 ^ 1'b0 ;
  assign n4860 = n2773 ^ n1811 ^ n1723 ;
  assign n4859 = n1216 ^ n732 ^ 1'b0 ;
  assign n4861 = n4860 ^ n4859 ^ n2891 ;
  assign n4863 = n4862 ^ n4861 ^ 1'b0 ;
  assign n4864 = n4863 ^ n1794 ^ n1127 ;
  assign n4873 = ( n1065 & ~n4089 ) | ( n1065 & n4236 ) | ( ~n4089 & n4236 ) ;
  assign n4869 = ( ~n589 & n771 ) | ( ~n589 & n1213 ) | ( n771 & n1213 ) ;
  assign n4870 = n4392 ^ n3225 ^ 1'b0 ;
  assign n4871 = n4869 | n4870 ;
  assign n4866 = n3658 ^ n1435 ^ n1259 ;
  assign n4867 = n4866 ^ n4014 ^ n2780 ;
  assign n4865 = n3726 ^ n2094 ^ 1'b0 ;
  assign n4868 = n4867 ^ n4865 ^ n3916 ;
  assign n4872 = n4871 ^ n4868 ^ n1522 ;
  assign n4874 = n4873 ^ n4872 ^ n4850 ;
  assign n4875 = n4874 ^ n3998 ^ 1'b0 ;
  assign n4876 = n1837 ^ x41 ^ 1'b0 ;
  assign n4877 = ( ~n269 & n2610 ) | ( ~n269 & n4876 ) | ( n2610 & n4876 ) ;
  assign n4878 = n1544 ^ n1539 ^ n924 ;
  assign n4879 = ( n2873 & n4497 ) | ( n2873 & ~n4878 ) | ( n4497 & ~n4878 ) ;
  assign n4882 = n2704 ^ n1360 ^ x240 ;
  assign n4881 = n2441 | n4644 ;
  assign n4883 = n4882 ^ n4881 ^ 1'b0 ;
  assign n4880 = ~n3719 & n4376 ;
  assign n4884 = n4883 ^ n4880 ^ 1'b0 ;
  assign n4891 = n915 ^ n432 ^ n355 ;
  assign n4892 = n4891 ^ n3436 ^ n2543 ;
  assign n4893 = ( n580 & n4423 ) | ( n580 & n4892 ) | ( n4423 & n4892 ) ;
  assign n4894 = n4893 ^ n509 ^ 1'b0 ;
  assign n4885 = n1243 ^ n675 ^ x249 ;
  assign n4886 = n1741 ^ n838 ^ 1'b0 ;
  assign n4887 = n4075 | n4886 ;
  assign n4888 = n1306 & ~n4887 ;
  assign n4889 = ~n2521 & n4888 ;
  assign n4890 = n4885 & ~n4889 ;
  assign n4895 = n4894 ^ n4890 ^ 1'b0 ;
  assign n4896 = n2540 ^ n1215 ^ 1'b0 ;
  assign n4897 = ( ~n4884 & n4895 ) | ( ~n4884 & n4896 ) | ( n4895 & n4896 ) ;
  assign n4898 = ( n4877 & n4879 ) | ( n4877 & n4897 ) | ( n4879 & n4897 ) ;
  assign n4902 = n3654 ^ n800 ^ 1'b0 ;
  assign n4903 = n1624 & n4902 ;
  assign n4904 = ( n1243 & n1781 ) | ( n1243 & n4903 ) | ( n1781 & n4903 ) ;
  assign n4899 = n1606 ^ n1282 ^ 1'b0 ;
  assign n4900 = ( ~n2779 & n3840 ) | ( ~n2779 & n4899 ) | ( n3840 & n4899 ) ;
  assign n4901 = n4900 ^ n3519 ^ n3341 ;
  assign n4905 = n4904 ^ n4901 ^ n1034 ;
  assign n4906 = n3635 ^ n2828 ^ x47 ;
  assign n4907 = ( n1058 & n1286 ) | ( n1058 & n4191 ) | ( n1286 & n4191 ) ;
  assign n4908 = ( n862 & ~n4906 ) | ( n862 & n4907 ) | ( ~n4906 & n4907 ) ;
  assign n4914 = n4714 ^ n3500 ^ x37 ;
  assign n4915 = ( n588 & ~n2876 ) | ( n588 & n3421 ) | ( ~n2876 & n3421 ) ;
  assign n4916 = ( n4063 & ~n4914 ) | ( n4063 & n4915 ) | ( ~n4914 & n4915 ) ;
  assign n4910 = n3388 ^ n2482 ^ n1897 ;
  assign n4909 = n1125 & ~n1333 ;
  assign n4911 = n4910 ^ n4909 ^ 1'b0 ;
  assign n4912 = x140 & n4911 ;
  assign n4913 = n4912 ^ n4406 ^ 1'b0 ;
  assign n4917 = n4916 ^ n4913 ^ n2454 ;
  assign n4925 = n2154 ^ n1987 ^ n718 ;
  assign n4923 = n4430 ^ n521 ^ 1'b0 ;
  assign n4924 = n1616 | n4923 ;
  assign n4926 = n4925 ^ n4924 ^ n859 ;
  assign n4919 = n308 & ~n644 ;
  assign n4918 = n4484 ^ n3621 ^ n824 ;
  assign n4920 = n4919 ^ n4918 ^ n3151 ;
  assign n4921 = ( ~n4247 & n4566 ) | ( ~n4247 & n4920 ) | ( n4566 & n4920 ) ;
  assign n4922 = ( n1246 & ~n1941 ) | ( n1246 & n4921 ) | ( ~n1941 & n4921 ) ;
  assign n4927 = n4926 ^ n4922 ^ 1'b0 ;
  assign n4928 = ~n4917 & n4927 ;
  assign n4946 = n1080 ^ n1074 ^ n342 ;
  assign n4947 = ( n822 & n3057 ) | ( n822 & n4946 ) | ( n3057 & n4946 ) ;
  assign n4948 = n4947 ^ n1404 ^ x60 ;
  assign n4940 = x48 & ~n3944 ;
  assign n4941 = n4940 ^ x81 ^ 1'b0 ;
  assign n4936 = ( n587 & n1031 ) | ( n587 & n2627 ) | ( n1031 & n2627 ) ;
  assign n4937 = ~n1505 & n4936 ;
  assign n4938 = n2056 & n4937 ;
  assign n4939 = n4938 ^ n4172 ^ n1509 ;
  assign n4942 = n4941 ^ n4939 ^ n907 ;
  assign n4934 = ( n1105 & ~n2062 ) | ( n1105 & n2855 ) | ( ~n2062 & n2855 ) ;
  assign n4929 = n1334 | n2900 ;
  assign n4930 = n1264 & n3019 ;
  assign n4931 = ~n469 & n4930 ;
  assign n4932 = n4929 | n4931 ;
  assign n4933 = ( x130 & ~n373 ) | ( x130 & n4932 ) | ( ~n373 & n4932 ) ;
  assign n4935 = n4934 ^ n4933 ^ 1'b0 ;
  assign n4943 = n4942 ^ n4935 ^ n2649 ;
  assign n4944 = n4323 & ~n4943 ;
  assign n4945 = n4944 ^ n320 ^ 1'b0 ;
  assign n4949 = n4948 ^ n4945 ^ n3316 ;
  assign n4950 = n1599 & n2185 ;
  assign n4951 = n3962 & n4950 ;
  assign n4952 = n3379 | n3401 ;
  assign n4953 = n4952 ^ n3557 ^ 1'b0 ;
  assign n4954 = ( n1202 & n3482 ) | ( n1202 & ~n4953 ) | ( n3482 & ~n4953 ) ;
  assign n4955 = ~n4951 & n4954 ;
  assign n4956 = ~n3724 & n4955 ;
  assign n4958 = ( x9 & ~n580 ) | ( x9 & n3463 ) | ( ~n580 & n3463 ) ;
  assign n4957 = ( n387 & n905 ) | ( n387 & ~n1565 ) | ( n905 & ~n1565 ) ;
  assign n4959 = n4958 ^ n4957 ^ n2615 ;
  assign n4965 = ( ~x101 & n1168 ) | ( ~x101 & n3928 ) | ( n1168 & n3928 ) ;
  assign n4960 = n2356 | n2525 ;
  assign n4961 = n4481 ^ n2201 ^ n1128 ;
  assign n4962 = n4961 ^ n3671 ^ n933 ;
  assign n4963 = n4962 ^ n1924 ^ n356 ;
  assign n4964 = n4960 & ~n4963 ;
  assign n4966 = n4965 ^ n4964 ^ 1'b0 ;
  assign n4967 = n2589 ^ n459 ^ 1'b0 ;
  assign n4968 = ~n3390 & n4967 ;
  assign n4969 = n3441 & n4968 ;
  assign n4970 = ~n2089 & n4969 ;
  assign n4971 = n700 & ~n2488 ;
  assign n4972 = n4970 & n4971 ;
  assign n4973 = ( x203 & ~n3056 ) | ( x203 & n3182 ) | ( ~n3056 & n3182 ) ;
  assign n4976 = n2142 ^ n975 ^ 1'b0 ;
  assign n4977 = n4296 & ~n4976 ;
  assign n4978 = n4977 ^ n817 ^ 1'b0 ;
  assign n4979 = n2071 & n4978 ;
  assign n4980 = n4979 ^ n2037 ^ 1'b0 ;
  assign n4974 = n2833 ^ n1865 ^ x174 ;
  assign n4975 = ~n2974 & n4974 ;
  assign n4981 = n4980 ^ n4975 ^ 1'b0 ;
  assign n4982 = ( n1040 & n4973 ) | ( n1040 & n4981 ) | ( n4973 & n4981 ) ;
  assign n4985 = n3067 ^ n1993 ^ n1724 ;
  assign n4986 = n4985 ^ n2830 ^ 1'b0 ;
  assign n4987 = x140 & n4986 ;
  assign n4988 = ( n950 & ~n1583 ) | ( n950 & n4987 ) | ( ~n1583 & n4987 ) ;
  assign n4989 = n4988 ^ n2084 ^ n1575 ;
  assign n4983 = n1676 | n1909 ;
  assign n4984 = n2258 | n4983 ;
  assign n4990 = n4989 ^ n4984 ^ n1256 ;
  assign n4991 = ( x251 & n3028 ) | ( x251 & n4327 ) | ( n3028 & n4327 ) ;
  assign n4992 = n4991 ^ n3066 ^ 1'b0 ;
  assign n4996 = n1352 ^ n1346 ^ x47 ;
  assign n4993 = ( n857 & ~n1571 ) | ( n857 & n2583 ) | ( ~n1571 & n2583 ) ;
  assign n4994 = ( n869 & n4411 ) | ( n869 & ~n4993 ) | ( n4411 & ~n4993 ) ;
  assign n4995 = ( n1595 & n3739 ) | ( n1595 & ~n4994 ) | ( n3739 & ~n4994 ) ;
  assign n4997 = n4996 ^ n4995 ^ n3946 ;
  assign n4998 = ( ~n4990 & n4992 ) | ( ~n4990 & n4997 ) | ( n4992 & n4997 ) ;
  assign n4999 = ( n4972 & n4982 ) | ( n4972 & ~n4998 ) | ( n4982 & ~n4998 ) ;
  assign n5000 = n2877 ^ n2245 ^ x160 ;
  assign n5001 = n5000 ^ n3790 ^ 1'b0 ;
  assign n5002 = n2976 ^ n1794 ^ 1'b0 ;
  assign n5003 = ~n1832 & n5002 ;
  assign n5004 = n2453 ^ n724 ^ x198 ;
  assign n5005 = n2210 | n5004 ;
  assign n5006 = n5005 ^ n2457 ^ 1'b0 ;
  assign n5007 = ~n566 & n5006 ;
  assign n5020 = n3744 ^ n496 ^ 1'b0 ;
  assign n5021 = n3073 ^ n2857 ^ n784 ;
  assign n5022 = ( ~n864 & n5020 ) | ( ~n864 & n5021 ) | ( n5020 & n5021 ) ;
  assign n5011 = x108 & ~n1205 ;
  assign n5012 = ~n517 & n5011 ;
  assign n5013 = ( x104 & n1263 ) | ( x104 & n5012 ) | ( n1263 & n5012 ) ;
  assign n5014 = n5013 ^ n1645 ^ n1283 ;
  assign n5009 = n321 | n2628 ;
  assign n5010 = n1730 | n5009 ;
  assign n5015 = n5014 ^ n5010 ^ 1'b0 ;
  assign n5008 = ( n2399 & ~n2821 ) | ( n2399 & n4108 ) | ( ~n2821 & n4108 ) ;
  assign n5016 = n5015 ^ n5008 ^ n3731 ;
  assign n5017 = n5016 ^ n2949 ^ n554 ;
  assign n5018 = n3144 & ~n5017 ;
  assign n5019 = n5018 ^ n4512 ^ 1'b0 ;
  assign n5023 = n5022 ^ n5019 ^ n3033 ;
  assign n5024 = ( n5003 & ~n5007 ) | ( n5003 & n5023 ) | ( ~n5007 & n5023 ) ;
  assign n5025 = n5024 ^ n1463 ^ 1'b0 ;
  assign n5026 = ( x217 & n1605 ) | ( x217 & ~n3663 ) | ( n1605 & ~n3663 ) ;
  assign n5027 = n2256 | n5026 ;
  assign n5028 = n2067 ^ n1270 ^ n964 ;
  assign n5029 = ( n1768 & ~n4443 ) | ( n1768 & n5028 ) | ( ~n4443 & n5028 ) ;
  assign n5030 = x248 & n2627 ;
  assign n5031 = n5030 ^ n4426 ^ 1'b0 ;
  assign n5032 = ( x38 & ~n3511 ) | ( x38 & n5031 ) | ( ~n3511 & n5031 ) ;
  assign n5033 = n2633 ^ n2113 ^ n412 ;
  assign n5034 = ( n278 & n1561 ) | ( n278 & n3569 ) | ( n1561 & n3569 ) ;
  assign n5035 = n1082 ^ n367 ^ 1'b0 ;
  assign n5036 = n5035 ^ n1885 ^ n790 ;
  assign n5041 = n1103 ^ n535 ^ x141 ;
  assign n5042 = ~n1813 & n5041 ;
  assign n5043 = n5042 ^ n544 ^ 1'b0 ;
  assign n5044 = ( ~x141 & n1320 ) | ( ~x141 & n5043 ) | ( n1320 & n5043 ) ;
  assign n5037 = n3153 ^ n1241 ^ n631 ;
  assign n5038 = n1527 | n5037 ;
  assign n5039 = n5038 ^ n317 ^ 1'b0 ;
  assign n5040 = n5039 ^ n3669 ^ n3302 ;
  assign n5045 = n5044 ^ n5040 ^ n1094 ;
  assign n5046 = n5045 ^ n3354 ^ n2553 ;
  assign n5047 = n5046 ^ x183 ^ 1'b0 ;
  assign n5048 = n1666 & ~n5047 ;
  assign n5049 = ( n5034 & n5036 ) | ( n5034 & n5048 ) | ( n5036 & n5048 ) ;
  assign n5050 = n5049 ^ n4012 ^ n1815 ;
  assign n5051 = n1250 ^ n585 ^ 1'b0 ;
  assign n5052 = n2323 & ~n5051 ;
  assign n5053 = ( ~n682 & n4318 ) | ( ~n682 & n5052 ) | ( n4318 & n5052 ) ;
  assign n5054 = ( n4170 & n5050 ) | ( n4170 & n5053 ) | ( n5050 & n5053 ) ;
  assign n5055 = ( n612 & n1366 ) | ( n612 & ~n4444 ) | ( n1366 & ~n4444 ) ;
  assign n5056 = n5055 ^ n3836 ^ x254 ;
  assign n5057 = ( ~n1744 & n2137 ) | ( ~n1744 & n5056 ) | ( n2137 & n5056 ) ;
  assign n5061 = x55 & n701 ;
  assign n5059 = n4931 ^ n3710 ^ n3261 ;
  assign n5058 = ~n1306 & n4304 ;
  assign n5060 = n5059 ^ n5058 ^ n2758 ;
  assign n5062 = n5061 ^ n5060 ^ n4264 ;
  assign n5063 = n552 & n4785 ;
  assign n5064 = n1198 & n5063 ;
  assign n5065 = ( x167 & ~n5004 ) | ( x167 & n5064 ) | ( ~n5004 & n5064 ) ;
  assign n5066 = ( n1731 & n1747 ) | ( n1731 & n2026 ) | ( n1747 & n2026 ) ;
  assign n5067 = n5066 ^ n2790 ^ 1'b0 ;
  assign n5068 = ( ~n3148 & n3878 ) | ( ~n3148 & n4718 ) | ( n3878 & n4718 ) ;
  assign n5069 = ( n5065 & n5067 ) | ( n5065 & n5068 ) | ( n5067 & n5068 ) ;
  assign n5071 = n4114 ^ n579 ^ 1'b0 ;
  assign n5070 = ( ~n1659 & n3357 ) | ( ~n1659 & n4574 ) | ( n3357 & n4574 ) ;
  assign n5072 = n5071 ^ n5070 ^ n1694 ;
  assign n5073 = n346 | n760 ;
  assign n5074 = n5073 ^ n4172 ^ n1310 ;
  assign n5075 = n5074 ^ n2720 ^ 1'b0 ;
  assign n5076 = x210 & n5075 ;
  assign n5077 = ( n1561 & n3054 ) | ( n1561 & ~n5076 ) | ( n3054 & ~n5076 ) ;
  assign n5078 = n5077 ^ n3443 ^ 1'b0 ;
  assign n5079 = n807 ^ n761 ^ x89 ;
  assign n5080 = ( n4427 & n4793 ) | ( n4427 & n5079 ) | ( n4793 & n5079 ) ;
  assign n5081 = n5080 ^ n3492 ^ n1359 ;
  assign n5082 = ( ~n593 & n2608 ) | ( ~n593 & n3129 ) | ( n2608 & n3129 ) ;
  assign n5083 = ( x204 & ~n757 ) | ( x204 & n5082 ) | ( ~n757 & n5082 ) ;
  assign n5084 = n256 & ~n5083 ;
  assign n5085 = ( n4549 & n4595 ) | ( n4549 & ~n5084 ) | ( n4595 & ~n5084 ) ;
  assign n5088 = ~n1293 & n2949 ;
  assign n5089 = n3750 ^ n1711 ^ n1617 ;
  assign n5090 = ( n3598 & n5088 ) | ( n3598 & ~n5089 ) | ( n5088 & ~n5089 ) ;
  assign n5086 = n1015 ^ n943 ^ n908 ;
  assign n5087 = n3506 & n5086 ;
  assign n5091 = n5090 ^ n5087 ^ n851 ;
  assign n5092 = n5091 ^ n4661 ^ 1'b0 ;
  assign n5093 = n4712 | n5092 ;
  assign n5099 = n518 & ~n1749 ;
  assign n5100 = n5099 ^ n2213 ^ 1'b0 ;
  assign n5101 = n2707 ^ n1895 ^ x40 ;
  assign n5102 = ~n5100 & n5101 ;
  assign n5094 = n4735 ^ n3211 ^ n1370 ;
  assign n5095 = ( n3988 & ~n4132 ) | ( n3988 & n5094 ) | ( ~n4132 & n5094 ) ;
  assign n5096 = n1319 & n5095 ;
  assign n5097 = n5096 ^ n4705 ^ 1'b0 ;
  assign n5098 = ( n3078 & ~n4070 ) | ( n3078 & n5097 ) | ( ~n4070 & n5097 ) ;
  assign n5103 = n5102 ^ n5098 ^ n5093 ;
  assign n5104 = ( ~n1185 & n1428 ) | ( ~n1185 & n4523 ) | ( n1428 & n4523 ) ;
  assign n5105 = n2787 & ~n5104 ;
  assign n5106 = n5105 ^ n2115 ^ 1'b0 ;
  assign n5115 = n1767 ^ n989 ^ n337 ;
  assign n5107 = n4376 ^ x29 ^ 1'b0 ;
  assign n5108 = ( n614 & ~n884 ) | ( n614 & n4798 ) | ( ~n884 & n4798 ) ;
  assign n5109 = n2016 ^ n498 ^ 1'b0 ;
  assign n5110 = n5108 | n5109 ;
  assign n5111 = n5110 ^ n3548 ^ 1'b0 ;
  assign n5112 = n5107 | n5111 ;
  assign n5113 = n3904 | n5112 ;
  assign n5114 = n1765 & ~n5113 ;
  assign n5116 = n5115 ^ n5114 ^ 1'b0 ;
  assign n5117 = ( n1108 & n1760 ) | ( n1108 & n2605 ) | ( n1760 & n2605 ) ;
  assign n5118 = n4364 ^ n3268 ^ n1569 ;
  assign n5119 = n5044 ^ n1486 ^ n287 ;
  assign n5120 = n730 & n5119 ;
  assign n5121 = ~x209 & n5120 ;
  assign n5122 = n5121 ^ n1795 ^ 1'b0 ;
  assign n5123 = n5118 | n5122 ;
  assign n5124 = n5123 ^ n4874 ^ n3606 ;
  assign n5125 = ( ~n840 & n1425 ) | ( ~n840 & n1444 ) | ( n1425 & n1444 ) ;
  assign n5126 = n4166 & ~n5125 ;
  assign n5127 = x240 & n4422 ;
  assign n5128 = ( n3205 & ~n3497 ) | ( n3205 & n5127 ) | ( ~n3497 & n5127 ) ;
  assign n5129 = n5128 ^ n3682 ^ 1'b0 ;
  assign n5130 = n1196 & n5129 ;
  assign n5133 = ( ~x22 & n587 ) | ( ~x22 & n4184 ) | ( n587 & n4184 ) ;
  assign n5131 = n2161 ^ n1943 ^ n525 ;
  assign n5132 = n5131 ^ n4437 ^ n867 ;
  assign n5134 = n5133 ^ n5132 ^ n4158 ;
  assign n5135 = n5134 ^ n915 ^ n486 ;
  assign n5136 = ( n1761 & n5130 ) | ( n1761 & ~n5135 ) | ( n5130 & ~n5135 ) ;
  assign n5137 = ~n541 & n4670 ;
  assign n5138 = ~n3678 & n5137 ;
  assign n5139 = n2230 ^ n1776 ^ x248 ;
  assign n5140 = ( n2218 & n2219 ) | ( n2218 & n5139 ) | ( n2219 & n5139 ) ;
  assign n5141 = n672 | n867 ;
  assign n5142 = n5141 ^ n3718 ^ 1'b0 ;
  assign n5143 = ( n2119 & n2213 ) | ( n2119 & ~n2892 ) | ( n2213 & ~n2892 ) ;
  assign n5144 = n5142 & n5143 ;
  assign n5145 = n1465 & ~n5144 ;
  assign n5152 = ~n1577 & n2495 ;
  assign n5153 = n5152 ^ n4892 ^ x40 ;
  assign n5154 = n5153 ^ n4841 ^ n3801 ;
  assign n5155 = n5154 ^ n1691 ^ n771 ;
  assign n5147 = ( ~n590 & n2401 ) | ( ~n590 & n3542 ) | ( n2401 & n3542 ) ;
  assign n5148 = ( n856 & n3506 ) | ( n856 & ~n5147 ) | ( n3506 & ~n5147 ) ;
  assign n5149 = n2737 ^ n2136 ^ n323 ;
  assign n5150 = n5148 | n5149 ;
  assign n5151 = ( ~x242 & n1921 ) | ( ~x242 & n5150 ) | ( n1921 & n5150 ) ;
  assign n5146 = n415 & ~n704 ;
  assign n5156 = n5155 ^ n5151 ^ n5146 ;
  assign n5157 = ( n430 & n539 ) | ( n430 & ~n549 ) | ( n539 & ~n549 ) ;
  assign n5158 = n5157 ^ n4785 ^ n1351 ;
  assign n5159 = ~n640 & n1594 ;
  assign n5160 = ( n2510 & ~n3812 ) | ( n2510 & n5159 ) | ( ~n3812 & n5159 ) ;
  assign n5161 = n1717 ^ n263 ^ x228 ;
  assign n5162 = ( n1536 & ~n1864 ) | ( n1536 & n5161 ) | ( ~n1864 & n5161 ) ;
  assign n5163 = x57 & ~n5162 ;
  assign n5164 = ~n2195 & n5163 ;
  assign n5165 = n5164 ^ n3741 ^ n3187 ;
  assign n5166 = n746 ^ n539 ^ 1'b0 ;
  assign n5167 = ( n2517 & n2906 ) | ( n2517 & ~n4345 ) | ( n2906 & ~n4345 ) ;
  assign n5168 = n4628 ^ n1543 ^ n292 ;
  assign n5169 = n4840 ^ n2820 ^ n1815 ;
  assign n5170 = ( n3020 & n3537 ) | ( n3020 & ~n5169 ) | ( n3537 & ~n5169 ) ;
  assign n5171 = n5170 ^ n2474 ^ n1961 ;
  assign n5172 = ( n1356 & n5168 ) | ( n1356 & ~n5171 ) | ( n5168 & ~n5171 ) ;
  assign n5175 = ( n1075 & ~n2093 ) | ( n1075 & n2996 ) | ( ~n2093 & n2996 ) ;
  assign n5176 = ( n408 & n3683 ) | ( n408 & ~n5175 ) | ( n3683 & ~n5175 ) ;
  assign n5173 = n295 & n3536 ;
  assign n5174 = ( x172 & n2102 ) | ( x172 & ~n5173 ) | ( n2102 & ~n5173 ) ;
  assign n5177 = n5176 ^ n5174 ^ n2577 ;
  assign n5178 = n4459 ^ n1722 ^ n468 ;
  assign n5179 = x77 & x174 ;
  assign n5180 = n5179 ^ n4688 ^ n2142 ;
  assign n5181 = ( n641 & n5178 ) | ( n641 & ~n5180 ) | ( n5178 & ~n5180 ) ;
  assign n5182 = ( ~n2922 & n5074 ) | ( ~n2922 & n5181 ) | ( n5074 & n5181 ) ;
  assign n5183 = n4019 ^ n3484 ^ n2615 ;
  assign n5184 = ( ~n1815 & n3800 ) | ( ~n1815 & n4785 ) | ( n3800 & n4785 ) ;
  assign n5185 = n5183 & n5184 ;
  assign n5186 = ( n1041 & ~n3015 ) | ( n1041 & n4654 ) | ( ~n3015 & n4654 ) ;
  assign n5187 = n874 & n3151 ;
  assign n5188 = ( ~n384 & n3141 ) | ( ~n384 & n3202 ) | ( n3141 & n3202 ) ;
  assign n5189 = n5188 ^ n3859 ^ 1'b0 ;
  assign n5190 = ( ~n4991 & n5187 ) | ( ~n4991 & n5189 ) | ( n5187 & n5189 ) ;
  assign n5191 = n3848 ^ n1253 ^ 1'b0 ;
  assign n5192 = n3878 ^ n3333 ^ 1'b0 ;
  assign n5194 = n3241 ^ n613 ^ 1'b0 ;
  assign n5195 = n5194 ^ n3577 ^ n1964 ;
  assign n5196 = ~n3035 & n5195 ;
  assign n5193 = n3946 ^ n2031 ^ 1'b0 ;
  assign n5197 = n5196 ^ n5193 ^ 1'b0 ;
  assign n5198 = n1288 & ~n5197 ;
  assign n5199 = n5198 ^ n4504 ^ 1'b0 ;
  assign n5200 = n3152 ^ n1141 ^ n763 ;
  assign n5201 = n3539 ^ n785 ^ 1'b0 ;
  assign n5202 = n5201 ^ n4872 ^ 1'b0 ;
  assign n5203 = n4479 & ~n5202 ;
  assign n5204 = n4787 ^ n1651 ^ 1'b0 ;
  assign n5207 = n4904 ^ n4226 ^ 1'b0 ;
  assign n5208 = n5207 ^ n5017 ^ 1'b0 ;
  assign n5205 = n1871 ^ n549 ^ n286 ;
  assign n5206 = n3523 & n5205 ;
  assign n5209 = n5208 ^ n5206 ^ 1'b0 ;
  assign n5210 = ( ~n2248 & n3621 ) | ( ~n2248 & n5209 ) | ( n3621 & n5209 ) ;
  assign n5211 = ~n5204 & n5210 ;
  assign n5212 = ( n3488 & n3546 ) | ( n3488 & n3765 ) | ( n3546 & n3765 ) ;
  assign n5213 = ~n2930 & n5212 ;
  assign n5214 = n1761 ^ n909 ^ 1'b0 ;
  assign n5218 = ( n2110 & ~n2760 ) | ( n2110 & n3066 ) | ( ~n2760 & n3066 ) ;
  assign n5215 = n4843 ^ n4164 ^ n502 ;
  assign n5216 = n5215 ^ n4675 ^ n4212 ;
  assign n5217 = ( n1129 & n2606 ) | ( n1129 & ~n5216 ) | ( n2606 & ~n5216 ) ;
  assign n5219 = n5218 ^ n5217 ^ n1382 ;
  assign n5220 = ( n1223 & n5214 ) | ( n1223 & n5219 ) | ( n5214 & n5219 ) ;
  assign n5221 = n5220 ^ x184 ^ 1'b0 ;
  assign n5222 = n2033 ^ n1065 ^ n939 ;
  assign n5223 = n5176 ^ n3225 ^ n1113 ;
  assign n5229 = n1863 ^ x16 ^ 1'b0 ;
  assign n5225 = x67 & x146 ;
  assign n5226 = n3560 & n5225 ;
  assign n5227 = n5226 ^ n3797 ^ x71 ;
  assign n5224 = n1873 ^ n1390 ^ n772 ;
  assign n5228 = n5227 ^ n5224 ^ n2933 ;
  assign n5230 = n5229 ^ n5228 ^ 1'b0 ;
  assign n5231 = n3744 ^ n3601 ^ n1058 ;
  assign n5232 = n2531 & n5010 ;
  assign n5233 = n1909 & n5232 ;
  assign n5234 = ( n5230 & ~n5231 ) | ( n5230 & n5233 ) | ( ~n5231 & n5233 ) ;
  assign n5235 = ( n5222 & ~n5223 ) | ( n5222 & n5234 ) | ( ~n5223 & n5234 ) ;
  assign n5236 = ( n3025 & n3129 ) | ( n3025 & ~n4354 ) | ( n3129 & ~n4354 ) ;
  assign n5237 = ( n460 & n2903 ) | ( n460 & ~n5236 ) | ( n2903 & ~n5236 ) ;
  assign n5238 = n5237 ^ n920 ^ n692 ;
  assign n5239 = n424 & ~n5238 ;
  assign n5240 = n4469 & n5239 ;
  assign n5241 = ( n2033 & n2850 ) | ( n2033 & ~n3875 ) | ( n2850 & ~n3875 ) ;
  assign n5242 = n3719 | n5241 ;
  assign n5243 = x178 & ~n3500 ;
  assign n5244 = n2364 ^ n1233 ^ 1'b0 ;
  assign n5245 = n4289 & n5244 ;
  assign n5263 = x101 & n4743 ;
  assign n5264 = n5263 ^ n658 ^ 1'b0 ;
  assign n5260 = n1968 ^ n1386 ^ n667 ;
  assign n5261 = ( n1544 & n2046 ) | ( n1544 & ~n4087 ) | ( n2046 & ~n4087 ) ;
  assign n5262 = ( n3371 & ~n5260 ) | ( n3371 & n5261 ) | ( ~n5260 & n5261 ) ;
  assign n5252 = n2052 ^ n1422 ^ x113 ;
  assign n5253 = n970 & ~n3196 ;
  assign n5254 = n2498 ^ n1709 ^ 1'b0 ;
  assign n5255 = n5253 | n5254 ;
  assign n5256 = n5252 | n5255 ;
  assign n5257 = n5256 ^ n1962 ^ 1'b0 ;
  assign n5250 = ( n413 & n576 ) | ( n413 & ~n1765 ) | ( n576 & ~n1765 ) ;
  assign n5247 = ( x20 & n2957 ) | ( x20 & n3777 ) | ( n2957 & n3777 ) ;
  assign n5248 = ~n689 & n1065 ;
  assign n5249 = ~n5247 & n5248 ;
  assign n5251 = n5250 ^ n5249 ^ n2267 ;
  assign n5258 = n5257 ^ n5251 ^ 1'b0 ;
  assign n5246 = ( n612 & n1225 ) | ( n612 & n1351 ) | ( n1225 & n1351 ) ;
  assign n5259 = n5258 ^ n5246 ^ n2930 ;
  assign n5265 = n5264 ^ n5262 ^ n5259 ;
  assign n5266 = ( n3839 & ~n3940 ) | ( n3839 & n5265 ) | ( ~n3940 & n5265 ) ;
  assign n5270 = ( ~n2170 & n2734 ) | ( ~n2170 & n2795 ) | ( n2734 & n2795 ) ;
  assign n5271 = ( n1999 & ~n2194 ) | ( n1999 & n5270 ) | ( ~n2194 & n5270 ) ;
  assign n5267 = n3605 ^ n1013 ^ x192 ;
  assign n5268 = n5267 ^ n1963 ^ n394 ;
  assign n5269 = n5268 ^ n654 ^ n545 ;
  assign n5272 = n5271 ^ n5269 ^ n3604 ;
  assign n5273 = n5272 ^ n5082 ^ n3169 ;
  assign n5274 = n2697 ^ n1522 ^ 1'b0 ;
  assign n5275 = ( ~n1231 & n1791 ) | ( ~n1231 & n4993 ) | ( n1791 & n4993 ) ;
  assign n5276 = ( n1422 & n5274 ) | ( n1422 & n5275 ) | ( n5274 & n5275 ) ;
  assign n5277 = n5276 ^ n729 ^ n689 ;
  assign n5280 = n328 & ~n1094 ;
  assign n5281 = ~n1830 & n5280 ;
  assign n5278 = n331 | n4937 ;
  assign n5279 = n5278 ^ n4513 ^ x191 ;
  assign n5282 = n5281 ^ n5279 ^ n3822 ;
  assign n5287 = n5073 ^ n2155 ^ n1550 ;
  assign n5288 = ( ~n346 & n3306 ) | ( ~n346 & n5287 ) | ( n3306 & n5287 ) ;
  assign n5285 = n4043 ^ n2743 ^ n496 ;
  assign n5286 = ( ~n1248 & n2542 ) | ( ~n1248 & n5285 ) | ( n2542 & n5285 ) ;
  assign n5283 = ( n1532 & n1635 ) | ( n1532 & n3445 ) | ( n1635 & n3445 ) ;
  assign n5284 = x29 | n5283 ;
  assign n5289 = n5288 ^ n5286 ^ n5284 ;
  assign n5290 = n3127 ^ n2886 ^ x142 ;
  assign n5291 = n5290 ^ n5050 ^ 1'b0 ;
  assign n5292 = n5289 & n5291 ;
  assign n5293 = ~n1866 & n5292 ;
  assign n5294 = ( x86 & n1778 ) | ( x86 & n2506 ) | ( n1778 & n2506 ) ;
  assign n5295 = n2119 ^ n608 ^ 1'b0 ;
  assign n5296 = n5294 | n5295 ;
  assign n5297 = n5296 ^ n1711 ^ n1505 ;
  assign n5298 = n1334 & ~n4563 ;
  assign n5299 = n831 & n5298 ;
  assign n5300 = n840 & n1572 ;
  assign n5301 = ~n2646 & n5300 ;
  assign n5302 = ( ~n3985 & n5299 ) | ( ~n3985 & n5301 ) | ( n5299 & n5301 ) ;
  assign n5309 = n2716 ^ n2546 ^ n1895 ;
  assign n5310 = n5309 ^ n3027 ^ 1'b0 ;
  assign n5304 = n1976 ^ n1968 ^ n1077 ;
  assign n5305 = n891 | n5304 ;
  assign n5306 = n5305 ^ n1320 ^ 1'b0 ;
  assign n5303 = ( ~n1059 & n2964 ) | ( ~n1059 & n3348 ) | ( n2964 & n3348 ) ;
  assign n5307 = n5306 ^ n5303 ^ n2592 ;
  assign n5308 = ( ~n1621 & n3962 ) | ( ~n1621 & n5307 ) | ( n3962 & n5307 ) ;
  assign n5311 = n5310 ^ n5308 ^ 1'b0 ;
  assign n5312 = n1451 ^ n1195 ^ n282 ;
  assign n5313 = n5312 ^ n1525 ^ 1'b0 ;
  assign n5314 = n1395 & n5313 ;
  assign n5315 = n388 & n5314 ;
  assign n5316 = x65 & ~n5315 ;
  assign n5317 = ( ~x126 & n2060 ) | ( ~x126 & n2356 ) | ( n2060 & n2356 ) ;
  assign n5318 = ( x203 & n347 ) | ( x203 & ~n1756 ) | ( n347 & ~n1756 ) ;
  assign n5319 = ( ~n3355 & n4730 ) | ( ~n3355 & n5318 ) | ( n4730 & n5318 ) ;
  assign n5320 = n5319 ^ n1007 ^ 1'b0 ;
  assign n5321 = n5317 | n5320 ;
  assign n5334 = n2848 ^ n503 ^ 1'b0 ;
  assign n5335 = n2292 & ~n5334 ;
  assign n5324 = ( n316 & n3109 ) | ( n316 & ~n4164 ) | ( n3109 & ~n4164 ) ;
  assign n5325 = n4338 ^ n1231 ^ n855 ;
  assign n5326 = n5325 ^ n2349 ^ n1243 ;
  assign n5327 = n5326 ^ n1734 ^ 1'b0 ;
  assign n5328 = ~n5324 & n5327 ;
  assign n5329 = n2260 ^ n1095 ^ n394 ;
  assign n5330 = n5329 ^ n3480 ^ n874 ;
  assign n5331 = n5330 ^ n4110 ^ n1328 ;
  assign n5332 = ( n551 & ~n568 ) | ( n551 & n4064 ) | ( ~n568 & n4064 ) ;
  assign n5333 = ( ~n5328 & n5331 ) | ( ~n5328 & n5332 ) | ( n5331 & n5332 ) ;
  assign n5322 = n1185 ^ n959 ^ x222 ;
  assign n5323 = ~n2391 & n5322 ;
  assign n5336 = n5335 ^ n5333 ^ n5323 ;
  assign n5337 = n3212 ^ n1971 ^ n286 ;
  assign n5338 = n1340 & ~n5337 ;
  assign n5343 = n3562 ^ n1169 ^ n957 ;
  assign n5344 = ( n395 & n2628 ) | ( n395 & ~n5343 ) | ( n2628 & ~n5343 ) ;
  assign n5345 = n5344 ^ n5215 ^ 1'b0 ;
  assign n5346 = n583 | n5345 ;
  assign n5339 = n471 & ~n1595 ;
  assign n5340 = n5339 ^ n1719 ^ n1074 ;
  assign n5341 = ( n1340 & n4553 ) | ( n1340 & n5340 ) | ( n4553 & n5340 ) ;
  assign n5342 = n1791 | n5341 ;
  assign n5347 = n5346 ^ n5342 ^ 1'b0 ;
  assign n5348 = ~n793 & n3270 ;
  assign n5349 = n2107 & n5348 ;
  assign n5350 = n5349 ^ n2253 ^ n1453 ;
  assign n5355 = ( x76 & n1229 ) | ( x76 & ~n1537 ) | ( n1229 & ~n1537 ) ;
  assign n5356 = ~n2786 & n5355 ;
  assign n5357 = n5356 ^ n1335 ^ 1'b0 ;
  assign n5354 = ( ~n1199 & n1680 ) | ( ~n1199 & n2504 ) | ( n1680 & n2504 ) ;
  assign n5358 = n5357 ^ n5354 ^ n1443 ;
  assign n5353 = ( x77 & n334 ) | ( x77 & ~n3505 ) | ( n334 & ~n3505 ) ;
  assign n5351 = n1622 | n5004 ;
  assign n5352 = n1025 | n5351 ;
  assign n5359 = n5358 ^ n5353 ^ n5352 ;
  assign n5360 = n743 & ~n4124 ;
  assign n5361 = n5360 ^ n5039 ^ 1'b0 ;
  assign n5368 = ( n1291 & n1625 ) | ( n1291 & n2484 ) | ( n1625 & n2484 ) ;
  assign n5369 = ( x16 & n2029 ) | ( x16 & n5368 ) | ( n2029 & n5368 ) ;
  assign n5370 = ( n1443 & ~n2255 ) | ( n1443 & n5369 ) | ( ~n2255 & n5369 ) ;
  assign n5362 = n286 & ~n3852 ;
  assign n5363 = n5362 ^ n1882 ^ 1'b0 ;
  assign n5364 = ~n370 & n5363 ;
  assign n5365 = n5364 ^ n2815 ^ 1'b0 ;
  assign n5366 = n1338 & ~n5365 ;
  assign n5367 = n5366 ^ n486 ^ 1'b0 ;
  assign n5371 = n5370 ^ n5367 ^ n1450 ;
  assign n5372 = ~n860 & n5299 ;
  assign n5373 = n5372 ^ n2561 ^ n1859 ;
  assign n5374 = ( n307 & ~n1437 ) | ( n307 & n5373 ) | ( ~n1437 & n5373 ) ;
  assign n5375 = n5374 ^ n1304 ^ 1'b0 ;
  assign n5376 = n5371 & ~n5375 ;
  assign n5377 = ( n3451 & ~n5361 ) | ( n3451 & n5376 ) | ( ~n5361 & n5376 ) ;
  assign n5380 = n3227 & ~n3944 ;
  assign n5378 = ~n1108 & n2859 ;
  assign n5379 = n5378 ^ n1204 ^ 1'b0 ;
  assign n5381 = n5380 ^ n5379 ^ n3223 ;
  assign n5382 = n5055 ^ n4708 ^ n851 ;
  assign n5383 = n5382 ^ n1479 ^ n1435 ;
  assign n5384 = ( x116 & n1879 ) | ( x116 & n5383 ) | ( n1879 & n5383 ) ;
  assign n5385 = n476 & n1535 ;
  assign n5391 = n1511 ^ n693 ^ n666 ;
  assign n5386 = n2637 & ~n3828 ;
  assign n5387 = ~n405 & n5386 ;
  assign n5388 = n1676 ^ n1416 ^ 1'b0 ;
  assign n5389 = ( n2570 & ~n3865 ) | ( n2570 & n5388 ) | ( ~n3865 & n5388 ) ;
  assign n5390 = ( ~n2159 & n5387 ) | ( ~n2159 & n5389 ) | ( n5387 & n5389 ) ;
  assign n5392 = n5391 ^ n5390 ^ 1'b0 ;
  assign n5393 = ~n1981 & n5392 ;
  assign n5394 = ( n1153 & ~n2718 ) | ( n1153 & n3483 ) | ( ~n2718 & n3483 ) ;
  assign n5395 = ~n406 & n5394 ;
  assign n5396 = ( ~x115 & n1352 ) | ( ~x115 & n2563 ) | ( n1352 & n2563 ) ;
  assign n5397 = n5396 ^ x206 ^ 1'b0 ;
  assign n5398 = n4253 & ~n5397 ;
  assign n5399 = n5398 ^ n1657 ^ n881 ;
  assign n5400 = n2963 ^ n985 ^ 1'b0 ;
  assign n5401 = n2916 ^ n2032 ^ n1936 ;
  assign n5402 = n5401 ^ n1641 ^ n604 ;
  assign n5403 = n998 | n5402 ;
  assign n5404 = n2293 & n5403 ;
  assign n5405 = n5404 ^ n3326 ^ 1'b0 ;
  assign n5406 = ( n694 & ~n2739 ) | ( n694 & n3824 ) | ( ~n2739 & n3824 ) ;
  assign n5407 = ( ~n890 & n1155 ) | ( ~n890 & n5406 ) | ( n1155 & n5406 ) ;
  assign n5408 = x12 & n3342 ;
  assign n5409 = ( ~x151 & n1152 ) | ( ~x151 & n5408 ) | ( n1152 & n5408 ) ;
  assign n5410 = n3332 ^ n1552 ^ 1'b0 ;
  assign n5411 = ~n706 & n5410 ;
  assign n5412 = n5411 ^ n2365 ^ 1'b0 ;
  assign n5413 = n5409 & ~n5412 ;
  assign n5414 = ( ~n3893 & n5249 ) | ( ~n3893 & n5413 ) | ( n5249 & n5413 ) ;
  assign n5415 = ( x122 & n1930 ) | ( x122 & n2063 ) | ( n1930 & n2063 ) ;
  assign n5416 = ( x225 & ~n3476 ) | ( x225 & n5415 ) | ( ~n3476 & n5415 ) ;
  assign n5417 = ( n1301 & n2125 ) | ( n1301 & ~n2556 ) | ( n2125 & ~n2556 ) ;
  assign n5418 = ( n1213 & n2476 ) | ( n1213 & n5417 ) | ( n2476 & n5417 ) ;
  assign n5419 = n3654 ^ n3331 ^ n3078 ;
  assign n5420 = ( n1092 & n2206 ) | ( n1092 & n5419 ) | ( n2206 & n5419 ) ;
  assign n5421 = n1835 ^ n580 ^ x2 ;
  assign n5422 = n4710 ^ n1616 ^ n1034 ;
  assign n5423 = n5422 ^ n2556 ^ 1'b0 ;
  assign n5424 = ~n5421 & n5423 ;
  assign n5425 = ( x188 & n643 ) | ( x188 & n1670 ) | ( n643 & n1670 ) ;
  assign n5426 = ( n378 & n475 ) | ( n378 & ~n646 ) | ( n475 & ~n646 ) ;
  assign n5427 = ( n5424 & ~n5425 ) | ( n5424 & n5426 ) | ( ~n5425 & n5426 ) ;
  assign n5428 = n2201 ^ n1497 ^ 1'b0 ;
  assign n5429 = n1062 | n5428 ;
  assign n5430 = ( n2653 & n4671 ) | ( n2653 & ~n5429 ) | ( n4671 & ~n5429 ) ;
  assign n5431 = ~n954 & n1261 ;
  assign n5432 = ~n4801 & n5431 ;
  assign n5433 = n4946 | n5432 ;
  assign n5438 = ( n417 & n1367 ) | ( n417 & n2922 ) | ( n1367 & n2922 ) ;
  assign n5434 = n287 & n2760 ;
  assign n5435 = n5434 ^ x58 ^ 1'b0 ;
  assign n5436 = ~n1813 & n2070 ;
  assign n5437 = ~n5435 & n5436 ;
  assign n5439 = n5438 ^ n5437 ^ 1'b0 ;
  assign n5440 = n2176 ^ x162 ^ 1'b0 ;
  assign n5442 = n1007 & ~n2122 ;
  assign n5441 = n4774 ^ n1999 ^ 1'b0 ;
  assign n5443 = n5442 ^ n5441 ^ n4857 ;
  assign n5448 = ( n491 & n939 ) | ( n491 & n1103 ) | ( n939 & n1103 ) ;
  assign n5449 = n1408 | n5448 ;
  assign n5450 = n3417 | n5449 ;
  assign n5451 = n5450 ^ n3071 ^ 1'b0 ;
  assign n5444 = x63 & n4906 ;
  assign n5445 = n5444 ^ n3147 ^ 1'b0 ;
  assign n5446 = ( n784 & ~n1492 ) | ( n784 & n3266 ) | ( ~n1492 & n3266 ) ;
  assign n5447 = ( n2258 & ~n5445 ) | ( n2258 & n5446 ) | ( ~n5445 & n5446 ) ;
  assign n5452 = n5451 ^ n5447 ^ n2369 ;
  assign n5462 = n3486 ^ n1722 ^ n1390 ;
  assign n5463 = ( n3634 & n4040 ) | ( n3634 & n5462 ) | ( n4040 & n5462 ) ;
  assign n5458 = n1329 ^ n1058 ^ n457 ;
  assign n5459 = n5458 ^ n1404 ^ n1226 ;
  assign n5455 = ~n2424 & n4684 ;
  assign n5456 = n5455 ^ n2378 ^ 1'b0 ;
  assign n5457 = n5456 ^ n4674 ^ n3950 ;
  assign n5460 = n5459 ^ n5457 ^ n982 ;
  assign n5461 = n5460 ^ x235 ^ 1'b0 ;
  assign n5453 = ( x8 & n401 ) | ( x8 & ~n1675 ) | ( n401 & ~n1675 ) ;
  assign n5454 = n5453 ^ n3379 ^ n2764 ;
  assign n5464 = n5463 ^ n5461 ^ n5454 ;
  assign n5465 = ( x113 & n390 ) | ( x113 & n2307 ) | ( n390 & n2307 ) ;
  assign n5466 = n5465 ^ n799 ^ 1'b0 ;
  assign n5467 = n5466 ^ n4530 ^ n2705 ;
  assign n5468 = n3023 ^ n844 ^ 1'b0 ;
  assign n5469 = n4298 | n5297 ;
  assign n5470 = ( ~x204 & n794 ) | ( ~x204 & n820 ) | ( n794 & n820 ) ;
  assign n5471 = n5470 ^ n2979 ^ n2460 ;
  assign n5472 = n1290 & ~n5471 ;
  assign n5473 = n5472 ^ n3215 ^ 1'b0 ;
  assign n5474 = x93 & n879 ;
  assign n5475 = n1975 ^ n760 ^ n487 ;
  assign n5476 = n5475 ^ n3671 ^ n1029 ;
  assign n5477 = ( n969 & n1827 ) | ( n969 & n3200 ) | ( n1827 & n3200 ) ;
  assign n5478 = n2114 | n5477 ;
  assign n5479 = n2179 & ~n5478 ;
  assign n5480 = n5479 ^ n4012 ^ n1883 ;
  assign n5481 = x34 & n437 ;
  assign n5482 = n5481 ^ n2522 ^ 1'b0 ;
  assign n5483 = n5482 ^ n3780 ^ n1155 ;
  assign n5484 = n2481 ^ n1912 ^ 1'b0 ;
  assign n5485 = n5483 & n5484 ;
  assign n5486 = n3777 ^ n1319 ^ n517 ;
  assign n5487 = ( n2095 & n5485 ) | ( n2095 & ~n5486 ) | ( n5485 & ~n5486 ) ;
  assign n5488 = n4239 ^ n3703 ^ 1'b0 ;
  assign n5489 = n5487 & ~n5488 ;
  assign n5492 = n3060 ^ n793 ^ 1'b0 ;
  assign n5493 = n1228 & n5492 ;
  assign n5490 = ~n2251 & n3562 ;
  assign n5491 = n5490 ^ n2848 ^ n859 ;
  assign n5494 = n5493 ^ n5491 ^ n5477 ;
  assign n5495 = ~n1299 & n2402 ;
  assign n5496 = n5495 ^ n5043 ^ 1'b0 ;
  assign n5497 = n5496 ^ n3075 ^ n1821 ;
  assign n5498 = n4283 | n5056 ;
  assign n5499 = ( n5494 & n5497 ) | ( n5494 & ~n5498 ) | ( n5497 & ~n5498 ) ;
  assign n5500 = n4089 ^ n3789 ^ n3151 ;
  assign n5501 = ( n3173 & n4745 ) | ( n3173 & n5500 ) | ( n4745 & n5500 ) ;
  assign n5502 = ( ~n752 & n931 ) | ( ~n752 & n1441 ) | ( n931 & n1441 ) ;
  assign n5503 = n3570 ^ n1166 ^ 1'b0 ;
  assign n5504 = ~n5502 & n5503 ;
  assign n5505 = n4296 ^ n1708 ^ n460 ;
  assign n5506 = n5505 ^ n5257 ^ n3710 ;
  assign n5507 = n5506 ^ n2450 ^ n1208 ;
  assign n5508 = ( ~x27 & n5504 ) | ( ~x27 & n5507 ) | ( n5504 & n5507 ) ;
  assign n5509 = n2254 & n5508 ;
  assign n5510 = ( ~n259 & n854 ) | ( ~n259 & n3067 ) | ( n854 & n3067 ) ;
  assign n5511 = n5510 ^ n3563 ^ n1095 ;
  assign n5512 = n4009 | n4667 ;
  assign n5513 = n1194 ^ x77 ^ 1'b0 ;
  assign n5514 = n863 & n5513 ;
  assign n5515 = ~n1652 & n5514 ;
  assign n5516 = n5515 ^ n2992 ^ 1'b0 ;
  assign n5520 = n2265 & ~n5204 ;
  assign n5521 = n5520 ^ n880 ^ 1'b0 ;
  assign n5517 = n2466 ^ n1187 ^ n996 ;
  assign n5518 = ~n4850 & n5517 ;
  assign n5519 = n5518 ^ n5283 ^ 1'b0 ;
  assign n5522 = n5521 ^ n5519 ^ n3786 ;
  assign n5523 = n5516 & ~n5522 ;
  assign n5524 = ~n3003 & n5523 ;
  assign n5525 = ( n5511 & n5512 ) | ( n5511 & ~n5524 ) | ( n5512 & ~n5524 ) ;
  assign n5528 = n1781 | n2670 ;
  assign n5526 = n1585 ^ n1462 ^ n346 ;
  assign n5527 = n5526 ^ n3608 ^ n393 ;
  assign n5529 = n5528 ^ n5527 ^ n2564 ;
  assign n5530 = n3417 ^ n1212 ^ n526 ;
  assign n5531 = ~n1429 & n3334 ;
  assign n5532 = ( n763 & n5530 ) | ( n763 & n5531 ) | ( n5530 & n5531 ) ;
  assign n5533 = n5529 & ~n5532 ;
  assign n5534 = n5533 ^ n2204 ^ 1'b0 ;
  assign n5535 = n1339 ^ n852 ^ 1'b0 ;
  assign n5536 = ~n3207 & n5535 ;
  assign n5538 = n1649 ^ n1461 ^ n281 ;
  assign n5537 = n1283 ^ x152 ^ 1'b0 ;
  assign n5539 = n5538 ^ n5537 ^ 1'b0 ;
  assign n5540 = ( n487 & ~n5536 ) | ( n487 & n5539 ) | ( ~n5536 & n5539 ) ;
  assign n5542 = n2344 ^ n2308 ^ n1305 ;
  assign n5543 = n5542 ^ n5108 ^ n3678 ;
  assign n5544 = n5543 ^ n4562 ^ x228 ;
  assign n5541 = ( n1371 & n1445 ) | ( n1371 & ~n4238 ) | ( n1445 & ~n4238 ) ;
  assign n5545 = n5544 ^ n5541 ^ n1716 ;
  assign n5546 = n5545 ^ n4493 ^ n4214 ;
  assign n5547 = ( ~n871 & n3260 ) | ( ~n871 & n5546 ) | ( n3260 & n5546 ) ;
  assign n5548 = n1081 | n1582 ;
  assign n5549 = n755 | n5548 ;
  assign n5550 = ( ~n347 & n1392 ) | ( ~n347 & n5549 ) | ( n1392 & n5549 ) ;
  assign n5551 = ( n2769 & n4176 ) | ( n2769 & n5550 ) | ( n4176 & n5550 ) ;
  assign n5552 = ( n3924 & n3976 ) | ( n3924 & ~n4087 ) | ( n3976 & ~n4087 ) ;
  assign n5555 = n2879 ^ n1133 ^ 1'b0 ;
  assign n5553 = n1002 | n3189 ;
  assign n5554 = n3390 & ~n5553 ;
  assign n5556 = n5555 ^ n5554 ^ 1'b0 ;
  assign n5557 = ( n5551 & n5552 ) | ( n5551 & n5556 ) | ( n5552 & n5556 ) ;
  assign n5558 = n2865 ^ n1305 ^ 1'b0 ;
  assign n5565 = ( x178 & ~n2665 ) | ( x178 & n4197 ) | ( ~n2665 & n4197 ) ;
  assign n5563 = n5463 ^ n324 ^ 1'b0 ;
  assign n5564 = n3275 & ~n5563 ;
  assign n5559 = ( n866 & ~n1236 ) | ( n866 & n2707 ) | ( ~n1236 & n2707 ) ;
  assign n5560 = ( n693 & n1236 ) | ( n693 & ~n5559 ) | ( n1236 & ~n5559 ) ;
  assign n5561 = n522 ^ n447 ^ 1'b0 ;
  assign n5562 = n5560 & ~n5561 ;
  assign n5566 = n5565 ^ n5564 ^ n5562 ;
  assign n5567 = ( n2577 & ~n3636 ) | ( n2577 & n5566 ) | ( ~n3636 & n5566 ) ;
  assign n5568 = ~n662 & n5567 ;
  assign n5569 = n1184 | n2615 ;
  assign n5570 = n5569 ^ n3661 ^ 1'b0 ;
  assign n5571 = ( n305 & ~n4685 ) | ( n305 & n5570 ) | ( ~n4685 & n5570 ) ;
  assign n5572 = ( n2987 & n4523 ) | ( n2987 & n5571 ) | ( n4523 & n5571 ) ;
  assign n5574 = ( n531 & n1412 ) | ( n531 & n1997 ) | ( n1412 & n1997 ) ;
  assign n5573 = ( n1191 & n1959 ) | ( n1191 & ~n1977 ) | ( n1959 & ~n1977 ) ;
  assign n5575 = n5574 ^ n5573 ^ n725 ;
  assign n5576 = ( ~x116 & x152 ) | ( ~x116 & n2026 ) | ( x152 & n2026 ) ;
  assign n5577 = ( n773 & n2562 ) | ( n773 & n5576 ) | ( n2562 & n5576 ) ;
  assign n5578 = n5577 ^ n722 ^ 1'b0 ;
  assign n5579 = n4307 ^ n1020 ^ n554 ;
  assign n5580 = n5579 ^ n3203 ^ n286 ;
  assign n5581 = ( n4094 & n5209 ) | ( n4094 & n5580 ) | ( n5209 & n5580 ) ;
  assign n5582 = n1281 ^ n1142 ^ n1007 ;
  assign n5583 = ( n315 & n417 ) | ( n315 & ~n705 ) | ( n417 & ~n705 ) ;
  assign n5584 = ( n2395 & n2668 ) | ( n2395 & n5583 ) | ( n2668 & n5583 ) ;
  assign n5585 = n1662 | n5584 ;
  assign n5586 = n5582 | n5585 ;
  assign n5587 = n5586 ^ n3950 ^ 1'b0 ;
  assign n5588 = ( ~n3082 & n3724 ) | ( ~n3082 & n5587 ) | ( n3724 & n5587 ) ;
  assign n5593 = ( n328 & ~n2243 ) | ( n328 & n3969 ) | ( ~n2243 & n3969 ) ;
  assign n5594 = ~n4763 & n5593 ;
  assign n5595 = n5594 ^ n3916 ^ 1'b0 ;
  assign n5589 = n1053 & n2341 ;
  assign n5590 = n5589 ^ n1007 ^ 1'b0 ;
  assign n5591 = n729 & ~n2351 ;
  assign n5592 = ( n546 & ~n5590 ) | ( n546 & n5591 ) | ( ~n5590 & n5591 ) ;
  assign n5596 = n5595 ^ n5592 ^ n487 ;
  assign n5597 = n5588 & n5596 ;
  assign n5598 = n5597 ^ n1130 ^ 1'b0 ;
  assign n5599 = n1635 & ~n5227 ;
  assign n5600 = n5599 ^ n1105 ^ n960 ;
  assign n5601 = n1726 | n5600 ;
  assign n5602 = ~n1118 & n5601 ;
  assign n5604 = n1930 ^ n412 ^ 1'b0 ;
  assign n5605 = n539 & n5604 ;
  assign n5603 = ( n4383 & ~n4620 ) | ( n4383 & n4626 ) | ( ~n4620 & n4626 ) ;
  assign n5606 = n5605 ^ n5603 ^ n3278 ;
  assign n5607 = ~n5602 & n5606 ;
  assign n5608 = n5607 ^ x240 ^ 1'b0 ;
  assign n5611 = n2705 & ~n3075 ;
  assign n5612 = n5611 ^ n505 ^ 1'b0 ;
  assign n5613 = n5612 ^ n2953 ^ n2029 ;
  assign n5609 = ~n2309 & n2717 ;
  assign n5610 = n5609 ^ n2102 ^ n1130 ;
  assign n5614 = n5613 ^ n5610 ^ n1636 ;
  assign n5615 = n5614 ^ n2699 ^ 1'b0 ;
  assign n5620 = n1990 ^ n1074 ^ x10 ;
  assign n5616 = n2937 ^ n2141 ^ n740 ;
  assign n5617 = n5616 ^ n551 ^ 1'b0 ;
  assign n5618 = n3008 & n5617 ;
  assign n5619 = n5618 ^ n4708 ^ n2309 ;
  assign n5621 = n5620 ^ n5619 ^ n667 ;
  assign n5622 = n5621 ^ n3759 ^ n1932 ;
  assign n5623 = ( n774 & n3736 ) | ( n774 & ~n5622 ) | ( n3736 & ~n5622 ) ;
  assign n5624 = n5623 ^ n2950 ^ n1126 ;
  assign n5625 = n1047 & ~n1380 ;
  assign n5627 = ~n2076 & n3557 ;
  assign n5626 = x164 & n649 ;
  assign n5628 = n5627 ^ n5626 ^ 1'b0 ;
  assign n5629 = n5036 ^ n1809 ^ n1678 ;
  assign n5630 = ( ~n528 & n1686 ) | ( ~n528 & n5629 ) | ( n1686 & n5629 ) ;
  assign n5631 = n5628 & ~n5630 ;
  assign n5632 = ~n5625 & n5631 ;
  assign n5647 = n3606 ^ n340 ^ x181 ;
  assign n5648 = ( x228 & n3397 ) | ( x228 & n3689 ) | ( n3397 & n3689 ) ;
  assign n5649 = n5648 ^ n775 ^ n716 ;
  assign n5650 = ~n1930 & n5649 ;
  assign n5651 = ( n1056 & n5647 ) | ( n1056 & ~n5650 ) | ( n5647 & ~n5650 ) ;
  assign n5652 = ( n1665 & n2326 ) | ( n1665 & n5651 ) | ( n2326 & n5651 ) ;
  assign n5633 = n3131 | n4439 ;
  assign n5634 = n5633 ^ n1175 ^ 1'b0 ;
  assign n5635 = ~n1116 & n1495 ;
  assign n5636 = n718 & n5635 ;
  assign n5637 = ( n1453 & ~n5634 ) | ( n1453 & n5636 ) | ( ~n5634 & n5636 ) ;
  assign n5644 = ( n884 & n1229 ) | ( n884 & n2334 ) | ( n1229 & n2334 ) ;
  assign n5642 = n3271 ^ n2430 ^ 1'b0 ;
  assign n5643 = n3683 & n5642 ;
  assign n5638 = n3628 | n4693 ;
  assign n5639 = n5638 ^ n1422 ^ n964 ;
  assign n5640 = n850 | n1088 ;
  assign n5641 = ( n949 & n5639 ) | ( n949 & ~n5640 ) | ( n5639 & ~n5640 ) ;
  assign n5645 = n5644 ^ n5643 ^ n5641 ;
  assign n5646 = n5637 & n5645 ;
  assign n5653 = n5652 ^ n5646 ^ 1'b0 ;
  assign n5654 = ( ~n3871 & n4237 ) | ( ~n3871 & n4253 ) | ( n4237 & n4253 ) ;
  assign n5655 = n5654 ^ n4150 ^ n1020 ;
  assign n5656 = ( n4513 & ~n5653 ) | ( n4513 & n5655 ) | ( ~n5653 & n5655 ) ;
  assign n5657 = n4877 ^ n2770 ^ n2219 ;
  assign n5658 = n5657 ^ n2441 ^ n399 ;
  assign n5659 = ~n1351 & n2460 ;
  assign n5660 = n975 & n5659 ;
  assign n5661 = ( n696 & ~n1389 ) | ( n696 & n2063 ) | ( ~n1389 & n2063 ) ;
  assign n5662 = n5661 ^ n928 ^ n848 ;
  assign n5663 = ( n1537 & ~n5660 ) | ( n1537 & n5662 ) | ( ~n5660 & n5662 ) ;
  assign n5664 = ( ~n1029 & n2417 ) | ( ~n1029 & n2751 ) | ( n2417 & n2751 ) ;
  assign n5665 = n5664 ^ n3109 ^ n2457 ;
  assign n5666 = n952 | n5665 ;
  assign n5669 = n3037 ^ n601 ^ x236 ;
  assign n5667 = ( n1023 & n1423 ) | ( n1023 & n3726 ) | ( n1423 & n3726 ) ;
  assign n5668 = ( n405 & ~n864 ) | ( n405 & n5667 ) | ( ~n864 & n5667 ) ;
  assign n5670 = n5669 ^ n5668 ^ 1'b0 ;
  assign n5676 = n3214 ^ n2715 ^ x12 ;
  assign n5673 = ( ~n324 & n1845 ) | ( ~n324 & n2126 ) | ( n1845 & n2126 ) ;
  assign n5674 = ( n262 & n3496 ) | ( n262 & n5673 ) | ( n3496 & n5673 ) ;
  assign n5672 = n4981 ^ n2412 ^ n2152 ;
  assign n5675 = n5674 ^ n5672 ^ n5224 ;
  assign n5671 = n3551 ^ n2077 ^ 1'b0 ;
  assign n5677 = n5676 ^ n5675 ^ n5671 ;
  assign n5678 = ( ~n4362 & n5670 ) | ( ~n4362 & n5677 ) | ( n5670 & n5677 ) ;
  assign n5680 = n592 | n3634 ;
  assign n5681 = n2301 | n5680 ;
  assign n5679 = n4739 ^ n1428 ^ 1'b0 ;
  assign n5682 = n5681 ^ n5679 ^ n2643 ;
  assign n5683 = n1050 & ~n1326 ;
  assign n5684 = ( ~x11 & n1596 ) | ( ~x11 & n2338 ) | ( n1596 & n2338 ) ;
  assign n5685 = n4600 | n5684 ;
  assign n5686 = n5683 & n5685 ;
  assign n5687 = n575 ^ n554 ^ 1'b0 ;
  assign n5688 = x182 & ~n5687 ;
  assign n5689 = n5688 ^ n2490 ^ 1'b0 ;
  assign n5690 = n4373 | n5689 ;
  assign n5691 = n3792 ^ n3672 ^ x177 ;
  assign n5692 = ( n2925 & ~n4945 ) | ( n2925 & n5691 ) | ( ~n4945 & n5691 ) ;
  assign n5693 = n3446 ^ n1649 ^ n283 ;
  assign n5694 = ( n446 & ~n619 ) | ( n446 & n5012 ) | ( ~n619 & n5012 ) ;
  assign n5695 = n2684 & n3572 ;
  assign n5696 = n5695 ^ n2143 ^ 1'b0 ;
  assign n5697 = ( n5693 & n5694 ) | ( n5693 & n5696 ) | ( n5694 & n5696 ) ;
  assign n5698 = n1724 & ~n3799 ;
  assign n5699 = ( x218 & ~n3260 ) | ( x218 & n5698 ) | ( ~n3260 & n5698 ) ;
  assign n5700 = ( n1396 & n2686 ) | ( n1396 & ~n5699 ) | ( n2686 & ~n5699 ) ;
  assign n5701 = ~n408 & n5700 ;
  assign n5702 = ( n4313 & n4887 ) | ( n4313 & ~n5701 ) | ( n4887 & ~n5701 ) ;
  assign n5703 = n1522 & ~n5702 ;
  assign n5706 = ( n1461 & n1822 ) | ( n1461 & ~n4812 ) | ( n1822 & ~n4812 ) ;
  assign n5704 = ( x5 & n1594 ) | ( x5 & ~n2849 ) | ( n1594 & ~n2849 ) ;
  assign n5705 = n5704 ^ n5044 ^ n552 ;
  assign n5707 = n5706 ^ n5705 ^ n4427 ;
  assign n5718 = ( ~x109 & n294 ) | ( ~x109 & n2273 ) | ( n294 & n2273 ) ;
  assign n5719 = n5718 ^ n1632 ^ 1'b0 ;
  assign n5714 = n922 & n936 ;
  assign n5715 = ( ~n4685 & n5264 ) | ( ~n4685 & n5714 ) | ( n5264 & n5714 ) ;
  assign n5716 = n5715 ^ n4175 ^ n1238 ;
  assign n5717 = n2304 & ~n5716 ;
  assign n5708 = ~n1078 & n1737 ;
  assign n5709 = ( ~n1522 & n2216 ) | ( ~n1522 & n3142 ) | ( n2216 & n3142 ) ;
  assign n5710 = ( x57 & ~n5708 ) | ( x57 & n5709 ) | ( ~n5708 & n5709 ) ;
  assign n5711 = ( n2970 & n5459 ) | ( n2970 & ~n5710 ) | ( n5459 & ~n5710 ) ;
  assign n5712 = n5711 ^ n3458 ^ n1842 ;
  assign n5713 = ( n2514 & n5294 ) | ( n2514 & ~n5712 ) | ( n5294 & ~n5712 ) ;
  assign n5720 = n5719 ^ n5717 ^ n5713 ;
  assign n5721 = n4042 ^ n3484 ^ n1579 ;
  assign n5722 = ( ~n1487 & n3800 ) | ( ~n1487 & n5721 ) | ( n3800 & n5721 ) ;
  assign n5723 = ~n970 & n5722 ;
  assign n5726 = n557 & n3289 ;
  assign n5727 = n5726 ^ x112 ^ 1'b0 ;
  assign n5728 = ( n457 & ~n4771 ) | ( n457 & n5727 ) | ( ~n4771 & n5727 ) ;
  assign n5724 = n4906 ^ n3008 ^ x72 ;
  assign n5725 = ( n1322 & ~n3133 ) | ( n1322 & n5724 ) | ( ~n3133 & n5724 ) ;
  assign n5729 = n5728 ^ n5725 ^ 1'b0 ;
  assign n5730 = n3732 & ~n5729 ;
  assign n5731 = n5730 ^ n4564 ^ 1'b0 ;
  assign n5732 = n5723 | n5731 ;
  assign n5739 = ( x138 & n281 ) | ( x138 & n1725 ) | ( n281 & n1725 ) ;
  assign n5733 = n4484 ^ x89 ^ 1'b0 ;
  assign n5734 = ( n4661 & n5161 ) | ( n4661 & ~n5733 ) | ( n5161 & ~n5733 ) ;
  assign n5735 = n5016 ^ n1654 ^ 1'b0 ;
  assign n5736 = ( n403 & n1716 ) | ( n403 & ~n3212 ) | ( n1716 & ~n3212 ) ;
  assign n5737 = ( n4685 & n5735 ) | ( n4685 & ~n5736 ) | ( n5735 & ~n5736 ) ;
  assign n5738 = n5734 & n5737 ;
  assign n5740 = n5739 ^ n5738 ^ 1'b0 ;
  assign n5741 = ( ~x12 & n2568 ) | ( ~x12 & n5704 ) | ( n2568 & n5704 ) ;
  assign n5742 = n2260 & n5741 ;
  assign n5743 = n5742 ^ n3353 ^ n1198 ;
  assign n5744 = n5490 ^ n4764 ^ n3443 ;
  assign n5745 = n2998 ^ n2950 ^ n2096 ;
  assign n5746 = ~n1457 & n5745 ;
  assign n5747 = n5746 ^ n1951 ^ 1'b0 ;
  assign n5748 = n5747 ^ n2501 ^ 1'b0 ;
  assign n5749 = ( n1910 & n3659 ) | ( n1910 & n4744 ) | ( n3659 & n4744 ) ;
  assign n5750 = ( n1873 & n5472 ) | ( n1873 & n5749 ) | ( n5472 & n5749 ) ;
  assign n5751 = ( n846 & n5619 ) | ( n846 & ~n5750 ) | ( n5619 & ~n5750 ) ;
  assign n5752 = ( n1768 & ~n2175 ) | ( n1768 & n2945 ) | ( ~n2175 & n2945 ) ;
  assign n5753 = n5752 ^ x138 ^ 1'b0 ;
  assign n5754 = n3744 & n5753 ;
  assign n5755 = n5549 ^ n4173 ^ n3197 ;
  assign n5756 = n5754 | n5755 ;
  assign n5757 = n5756 ^ n2046 ^ n1130 ;
  assign n5758 = n5757 ^ n2311 ^ 1'b0 ;
  assign n5759 = ~n5751 & n5758 ;
  assign n5760 = n3626 ^ n2343 ^ 1'b0 ;
  assign n5761 = n3535 ^ n1293 ^ 1'b0 ;
  assign n5762 = ( n641 & n988 ) | ( n641 & ~n5761 ) | ( n988 & ~n5761 ) ;
  assign n5763 = ~n1863 & n4559 ;
  assign n5764 = ~n3048 & n5763 ;
  assign n5765 = n5764 ^ n707 ^ 1'b0 ;
  assign n5766 = ~n3807 & n5765 ;
  assign n5767 = ( ~n5760 & n5762 ) | ( ~n5760 & n5766 ) | ( n5762 & n5766 ) ;
  assign n5768 = n276 & n5767 ;
  assign n5769 = n5768 ^ x31 ^ 1'b0 ;
  assign n5777 = n2606 ^ n547 ^ x149 ;
  assign n5778 = ( ~n370 & n4629 ) | ( ~n370 & n5777 ) | ( n4629 & n5777 ) ;
  assign n5770 = ( n543 & n1299 ) | ( n543 & n1504 ) | ( n1299 & n1504 ) ;
  assign n5771 = ( n1387 & ~n3790 ) | ( n1387 & n5770 ) | ( ~n3790 & n5770 ) ;
  assign n5773 = n3554 | n4216 ;
  assign n5774 = n5773 ^ n1455 ^ 1'b0 ;
  assign n5772 = ( ~n683 & n4744 ) | ( ~n683 & n5506 ) | ( n4744 & n5506 ) ;
  assign n5775 = n5774 ^ n5772 ^ n4440 ;
  assign n5776 = ( n3060 & n5771 ) | ( n3060 & n5775 ) | ( n5771 & n5775 ) ;
  assign n5779 = n5778 ^ n5776 ^ 1'b0 ;
  assign n5780 = n2661 ^ n2242 ^ n336 ;
  assign n5781 = ~n1595 & n5780 ;
  assign n5782 = n5781 ^ n4773 ^ 1'b0 ;
  assign n5783 = ( ~x135 & n1101 ) | ( ~x135 & n1692 ) | ( n1101 & n1692 ) ;
  assign n5784 = ( n1549 & ~n4059 ) | ( n1549 & n5783 ) | ( ~n4059 & n5783 ) ;
  assign n5785 = n5784 ^ n3052 ^ n2219 ;
  assign n5786 = n4085 ^ n2714 ^ n2407 ;
  assign n5787 = n5786 ^ n2244 ^ n773 ;
  assign n5788 = ( n1465 & n4774 ) | ( n1465 & ~n5787 ) | ( n4774 & ~n5787 ) ;
  assign n5789 = n5788 ^ n1170 ^ 1'b0 ;
  assign n5790 = ~n5785 & n5789 ;
  assign n5791 = n3463 ^ n1858 ^ n340 ;
  assign n5792 = ( n425 & n1939 ) | ( n425 & n2827 ) | ( n1939 & n2827 ) ;
  assign n5793 = ( ~n4053 & n5035 ) | ( ~n4053 & n5792 ) | ( n5035 & n5792 ) ;
  assign n5794 = n3157 ^ n2923 ^ 1'b0 ;
  assign n5795 = ( n1082 & n1323 ) | ( n1082 & n1941 ) | ( n1323 & n1941 ) ;
  assign n5796 = n5795 ^ n5196 ^ n2311 ;
  assign n5797 = x94 | n1428 ;
  assign n5798 = ~n3995 & n5797 ;
  assign n5799 = n5798 ^ n338 ^ 1'b0 ;
  assign n5800 = n5061 ^ n427 ^ x162 ;
  assign n5801 = n818 | n4481 ;
  assign n5802 = ~n1216 & n5801 ;
  assign n5803 = ~n5800 & n5802 ;
  assign n5804 = n1608 & ~n5803 ;
  assign n5805 = n5804 ^ n3823 ^ n1246 ;
  assign n5806 = n4356 ^ n3075 ^ n394 ;
  assign n5807 = n2752 ^ n1282 ^ n1178 ;
  assign n5808 = ( n428 & n1549 ) | ( n428 & ~n5807 ) | ( n1549 & ~n5807 ) ;
  assign n5809 = ~n3875 & n5808 ;
  assign n5810 = n5809 ^ n1727 ^ 1'b0 ;
  assign n5811 = ( n4037 & n5806 ) | ( n4037 & ~n5810 ) | ( n5806 & ~n5810 ) ;
  assign n5812 = ( n3768 & n3824 ) | ( n3768 & n5811 ) | ( n3824 & n5811 ) ;
  assign n5813 = ( n5799 & n5805 ) | ( n5799 & ~n5812 ) | ( n5805 & ~n5812 ) ;
  assign n5815 = ( n3083 & n4187 ) | ( n3083 & ~n5718 ) | ( n4187 & ~n5718 ) ;
  assign n5814 = ( x140 & ~n1636 ) | ( x140 & n2225 ) | ( ~n1636 & n2225 ) ;
  assign n5816 = n5815 ^ n5814 ^ 1'b0 ;
  assign n5817 = n590 & ~n5816 ;
  assign n5818 = n5817 ^ n2656 ^ 1'b0 ;
  assign n5819 = ~n823 & n5818 ;
  assign n5820 = ( n2709 & n2789 ) | ( n2709 & n5380 ) | ( n2789 & n5380 ) ;
  assign n5821 = n3214 ^ n1886 ^ 1'b0 ;
  assign n5822 = n5820 & n5821 ;
  assign n5823 = n5822 ^ n2705 ^ 1'b0 ;
  assign n5824 = n5819 & n5823 ;
  assign n5825 = ~n5317 & n5824 ;
  assign n5826 = ~n1411 & n5825 ;
  assign n5827 = x26 & n1898 ;
  assign n5828 = n5827 ^ n2518 ^ 1'b0 ;
  assign n5829 = n3750 ^ n2564 ^ n1427 ;
  assign n5830 = n5829 ^ n763 ^ 1'b0 ;
  assign n5831 = n5828 & ~n5830 ;
  assign n5832 = ( n4742 & n5022 ) | ( n4742 & n5483 ) | ( n5022 & n5483 ) ;
  assign n5833 = ( n3650 & n5831 ) | ( n3650 & ~n5832 ) | ( n5831 & ~n5832 ) ;
  assign n5837 = n348 & n2959 ;
  assign n5838 = ~x205 & n5837 ;
  assign n5839 = n5838 ^ n5694 ^ n1294 ;
  assign n5834 = ( ~n1692 & n4552 ) | ( ~n1692 & n4810 ) | ( n4552 & n4810 ) ;
  assign n5835 = n4310 | n5665 ;
  assign n5836 = n5834 | n5835 ;
  assign n5840 = n5839 ^ n5836 ^ n1550 ;
  assign n5841 = n4841 ^ n3587 ^ x160 ;
  assign n5842 = n5841 ^ n361 ^ 1'b0 ;
  assign n5843 = n2110 ^ n528 ^ n317 ;
  assign n5844 = n5843 ^ n2255 ^ n1190 ;
  assign n5845 = n5844 ^ n2922 ^ 1'b0 ;
  assign n5846 = n745 ^ n388 ^ n368 ;
  assign n5847 = ~n1502 & n5846 ;
  assign n5848 = ~n4664 & n5847 ;
  assign n5849 = ( ~n632 & n870 ) | ( ~n632 & n3609 ) | ( n870 & n3609 ) ;
  assign n5850 = n5843 ^ n5100 ^ 1'b0 ;
  assign n5851 = n5849 | n5850 ;
  assign n5852 = ( n1120 & n2257 ) | ( n1120 & n5851 ) | ( n2257 & n5851 ) ;
  assign n5853 = ( n5845 & ~n5848 ) | ( n5845 & n5852 ) | ( ~n5848 & n5852 ) ;
  assign n5854 = ( n384 & n5842 ) | ( n384 & n5853 ) | ( n5842 & n5853 ) ;
  assign n5855 = n4444 ^ n1734 ^ x86 ;
  assign n5856 = n5855 ^ n3624 ^ n1294 ;
  assign n5858 = ~n641 & n2295 ;
  assign n5857 = n1611 ^ n1106 ^ x69 ;
  assign n5859 = n5858 ^ n5857 ^ n4520 ;
  assign n5860 = n4734 | n5859 ;
  assign n5861 = n5860 ^ n2835 ^ 1'b0 ;
  assign n5862 = n5861 ^ n5759 ^ n806 ;
  assign n5863 = n1888 | n5845 ;
  assign n5864 = n500 & ~n5863 ;
  assign n5865 = n5864 ^ n2905 ^ n414 ;
  assign n5866 = n5865 ^ n5057 ^ n1918 ;
  assign n5867 = n5866 ^ n3433 ^ 1'b0 ;
  assign n5873 = n1690 ^ n1231 ^ 1'b0 ;
  assign n5870 = n5490 ^ n4596 ^ n1813 ;
  assign n5871 = ~n1328 & n5870 ;
  assign n5868 = n3705 & ~n3985 ;
  assign n5869 = n2891 & n5868 ;
  assign n5872 = n5871 ^ n5869 ^ n5616 ;
  assign n5874 = n5873 ^ n5872 ^ n2084 ;
  assign n5875 = ( n1016 & n2365 ) | ( n1016 & n3569 ) | ( n2365 & n3569 ) ;
  assign n5876 = n5875 ^ n532 ^ 1'b0 ;
  assign n5877 = x190 & n5876 ;
  assign n5878 = ( x214 & ~n297 ) | ( x214 & n428 ) | ( ~n297 & n428 ) ;
  assign n5879 = n5878 ^ n1956 ^ 1'b0 ;
  assign n5880 = ( n3731 & n4168 ) | ( n3731 & ~n5879 ) | ( n4168 & ~n5879 ) ;
  assign n5887 = ( ~x124 & n1460 ) | ( ~x124 & n3316 ) | ( n1460 & n3316 ) ;
  assign n5884 = ( n1756 & n1784 ) | ( n1756 & n5419 ) | ( n1784 & n5419 ) ;
  assign n5885 = n5884 ^ n599 ^ x118 ;
  assign n5883 = n1748 | n4900 ;
  assign n5886 = n5885 ^ n5883 ^ 1'b0 ;
  assign n5881 = n4198 ^ n1497 ^ n810 ;
  assign n5882 = ( n5123 & ~n5764 ) | ( n5123 & n5881 ) | ( ~n5764 & n5881 ) ;
  assign n5888 = n5887 ^ n5886 ^ n5882 ;
  assign n5889 = ( n307 & ~n1627 ) | ( n307 & n5859 ) | ( ~n1627 & n5859 ) ;
  assign n5890 = ( n1180 & ~n5762 ) | ( n1180 & n5889 ) | ( ~n5762 & n5889 ) ;
  assign n5891 = ( ~n3901 & n3995 ) | ( ~n3901 & n5890 ) | ( n3995 & n5890 ) ;
  assign n5892 = ~n923 & n5559 ;
  assign n5893 = ~n2664 & n5892 ;
  assign n5894 = ( x181 & ~n5043 ) | ( x181 & n5893 ) | ( ~n5043 & n5893 ) ;
  assign n5895 = n5894 ^ n1879 ^ n884 ;
  assign n5896 = n5895 ^ n2240 ^ 1'b0 ;
  assign n5897 = n5891 & ~n5896 ;
  assign n5898 = n5694 ^ n4276 ^ n3562 ;
  assign n5899 = ( ~n269 & n1777 ) | ( ~n269 & n4411 ) | ( n1777 & n4411 ) ;
  assign n5907 = n941 & n2679 ;
  assign n5909 = ( n987 & ~n2070 ) | ( n987 & n3268 ) | ( ~n2070 & n3268 ) ;
  assign n5908 = n2721 ^ n1878 ^ n635 ;
  assign n5910 = n5909 ^ n5908 ^ 1'b0 ;
  assign n5911 = ( n2052 & ~n5907 ) | ( n2052 & n5910 ) | ( ~n5907 & n5910 ) ;
  assign n5904 = n4436 ^ n809 ^ 1'b0 ;
  assign n5905 = ( n888 & n2518 ) | ( n888 & ~n5904 ) | ( n2518 & ~n5904 ) ;
  assign n5906 = ( n1026 & n1439 ) | ( n1026 & ~n5905 ) | ( n1439 & ~n5905 ) ;
  assign n5912 = n5911 ^ n5906 ^ x49 ;
  assign n5900 = n3204 ^ n1315 ^ n332 ;
  assign n5901 = n5900 ^ n5734 ^ 1'b0 ;
  assign n5902 = ( x204 & n3021 ) | ( x204 & n5599 ) | ( n3021 & n5599 ) ;
  assign n5903 = ( ~n1397 & n5901 ) | ( ~n1397 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5913 = n5912 ^ n5903 ^ n1522 ;
  assign n5914 = n5913 ^ n2604 ^ 1'b0 ;
  assign n5915 = n3683 & n5914 ;
  assign n5916 = ~n5899 & n5915 ;
  assign n5923 = n801 & ~n1252 ;
  assign n5922 = ( n1114 & n1329 ) | ( n1114 & n1834 ) | ( n1329 & n1834 ) ;
  assign n5924 = n5923 ^ n5922 ^ n1352 ;
  assign n5917 = ( n271 & n432 ) | ( n271 & n2384 ) | ( n432 & n2384 ) ;
  assign n5918 = ( n1165 & n5749 ) | ( n1165 & ~n5917 ) | ( n5749 & ~n5917 ) ;
  assign n5919 = n3989 & n4901 ;
  assign n5920 = n5919 ^ n3333 ^ 1'b0 ;
  assign n5921 = ( ~n1709 & n5918 ) | ( ~n1709 & n5920 ) | ( n5918 & n5920 ) ;
  assign n5925 = n5924 ^ n5921 ^ 1'b0 ;
  assign n5926 = n2625 ^ n2002 ^ n1601 ;
  assign n5927 = ( n1428 & n1920 ) | ( n1428 & ~n5926 ) | ( n1920 & ~n5926 ) ;
  assign n5928 = ~n4899 & n5927 ;
  assign n5929 = n5928 ^ n3278 ^ 1'b0 ;
  assign n5930 = ( n634 & n4647 ) | ( n634 & ~n5929 ) | ( n4647 & ~n5929 ) ;
  assign n5931 = n2176 ^ n2036 ^ n368 ;
  assign n5932 = ~n1406 & n4273 ;
  assign n5933 = n2024 & n5932 ;
  assign n5934 = n1149 & ~n5933 ;
  assign n5935 = n5934 ^ x181 ^ 1'b0 ;
  assign n5942 = n357 | n2382 ;
  assign n5943 = n5942 ^ n1576 ^ 1'b0 ;
  assign n5944 = n5943 ^ n5636 ^ n5301 ;
  assign n5940 = ( ~n415 & n2062 ) | ( ~n415 & n3105 ) | ( n2062 & n3105 ) ;
  assign n5936 = n4325 ^ n2452 ^ 1'b0 ;
  assign n5937 = ~n2938 & n5936 ;
  assign n5938 = n5937 ^ n4989 ^ n793 ;
  assign n5939 = ~n1662 & n5938 ;
  assign n5941 = n5940 ^ n5939 ^ 1'b0 ;
  assign n5945 = n5944 ^ n5941 ^ 1'b0 ;
  assign n5946 = n5935 | n5945 ;
  assign n5947 = n5931 | n5946 ;
  assign n5948 = n5930 | n5947 ;
  assign n5952 = n1018 ^ n973 ^ 1'b0 ;
  assign n5949 = n988 & n1141 ;
  assign n5950 = n2095 & n5949 ;
  assign n5951 = n3284 & ~n5950 ;
  assign n5953 = n5952 ^ n5951 ^ 1'b0 ;
  assign n5954 = ( n397 & ~n557 ) | ( n397 & n5953 ) | ( ~n557 & n5953 ) ;
  assign n5955 = n5954 ^ n559 ^ 1'b0 ;
  assign n5956 = n5688 & n5955 ;
  assign n5957 = n5956 ^ n3966 ^ 1'b0 ;
  assign n5958 = ( n2441 & ~n5067 ) | ( n2441 & n5514 ) | ( ~n5067 & n5514 ) ;
  assign n5959 = n2524 ^ x176 ^ 1'b0 ;
  assign n5960 = n5959 ^ n1981 ^ 1'b0 ;
  assign n5961 = n5958 & n5960 ;
  assign n5962 = n5961 ^ n4648 ^ n4012 ;
  assign n5971 = ( n1847 & n1915 ) | ( n1847 & ~n3014 ) | ( n1915 & ~n3014 ) ;
  assign n5972 = x149 & ~n5971 ;
  assign n5973 = n1902 & n5972 ;
  assign n5974 = n5973 ^ n1989 ^ x118 ;
  assign n5963 = n3353 ^ n2580 ^ n2142 ;
  assign n5964 = n2871 ^ n1072 ^ x72 ;
  assign n5965 = n5964 ^ n3568 ^ n3095 ;
  assign n5966 = ( n1501 & n2156 ) | ( n1501 & ~n4457 ) | ( n2156 & ~n4457 ) ;
  assign n5967 = ~n4354 & n4653 ;
  assign n5968 = n5967 ^ n3826 ^ n2879 ;
  assign n5969 = ( ~n5965 & n5966 ) | ( ~n5965 & n5968 ) | ( n5966 & n5968 ) ;
  assign n5970 = ( ~n2132 & n5963 ) | ( ~n2132 & n5969 ) | ( n5963 & n5969 ) ;
  assign n5975 = n5974 ^ n5970 ^ n2394 ;
  assign n5976 = n4742 ^ n3093 ^ n392 ;
  assign n5977 = n1878 & ~n5976 ;
  assign n5978 = ( ~n952 & n4683 ) | ( ~n952 & n5977 ) | ( n4683 & n5977 ) ;
  assign n5979 = ( n889 & n1539 ) | ( n889 & n1757 ) | ( n1539 & n1757 ) ;
  assign n5980 = n4778 & n5979 ;
  assign n5981 = ( n844 & ~n1909 ) | ( n844 & n2084 ) | ( ~n1909 & n2084 ) ;
  assign n5982 = ( x65 & n671 ) | ( x65 & ~n895 ) | ( n671 & ~n895 ) ;
  assign n5983 = ( ~n1479 & n2276 ) | ( ~n1479 & n5982 ) | ( n2276 & n5982 ) ;
  assign n5984 = ( n1961 & ~n5981 ) | ( n1961 & n5983 ) | ( ~n5981 & n5983 ) ;
  assign n5985 = n373 & n5984 ;
  assign n5986 = n5985 ^ n2541 ^ 1'b0 ;
  assign n5987 = n3860 ^ n1863 ^ n1695 ;
  assign n5988 = n5987 ^ n1241 ^ n448 ;
  assign n5989 = n3583 ^ n1469 ^ 1'b0 ;
  assign n5990 = ~n5988 & n5989 ;
  assign n5991 = ( x233 & n3259 ) | ( x233 & ~n5990 ) | ( n3259 & ~n5990 ) ;
  assign n5992 = n4939 & ~n5372 ;
  assign n5993 = n1423 & n5992 ;
  assign n5994 = ( n5986 & ~n5991 ) | ( n5986 & n5993 ) | ( ~n5991 & n5993 ) ;
  assign n5995 = n5980 | n5994 ;
  assign n5996 = n5978 | n5995 ;
  assign n5997 = n1904 ^ n463 ^ 1'b0 ;
  assign n5998 = n4913 ^ n4523 ^ x70 ;
  assign n5999 = ( n2135 & ~n5997 ) | ( n2135 & n5998 ) | ( ~n5997 & n5998 ) ;
  assign n6000 = n4121 ^ n3965 ^ n2260 ;
  assign n6001 = n2379 | n6000 ;
  assign n6002 = n836 & ~n5800 ;
  assign n6003 = n1370 ^ n273 ^ 1'b0 ;
  assign n6004 = ~n6002 & n6003 ;
  assign n6005 = n1608 ^ x151 ^ 1'b0 ;
  assign n6006 = x241 & n6005 ;
  assign n6007 = ( x171 & n5117 ) | ( x171 & ~n6006 ) | ( n5117 & ~n6006 ) ;
  assign n6008 = n6007 ^ n2107 ^ 1'b0 ;
  assign n6009 = ~n2938 & n6008 ;
  assign n6010 = ( n2430 & n6004 ) | ( n2430 & n6009 ) | ( n6004 & n6009 ) ;
  assign n6011 = ( n3117 & n3566 ) | ( n3117 & ~n4465 ) | ( n3566 & ~n4465 ) ;
  assign n6012 = n2074 | n6011 ;
  assign n6013 = n6010 | n6012 ;
  assign n6014 = n5952 ^ n4747 ^ n3152 ;
  assign n6015 = ( n944 & ~n3483 ) | ( n944 & n5475 ) | ( ~n3483 & n5475 ) ;
  assign n6016 = n4352 & ~n6015 ;
  assign n6017 = n6014 & n6016 ;
  assign n6018 = ( ~n390 & n3766 ) | ( ~n390 & n5050 ) | ( n3766 & n5050 ) ;
  assign n6019 = n5398 & ~n6018 ;
  assign n6020 = ( x42 & x222 ) | ( x42 & n4134 ) | ( x222 & n4134 ) ;
  assign n6021 = n4841 ^ n2540 ^ n1438 ;
  assign n6022 = ( n3609 & n6020 ) | ( n3609 & n6021 ) | ( n6020 & n6021 ) ;
  assign n6025 = ( x54 & ~x134 ) | ( x54 & n2003 ) | ( ~x134 & n2003 ) ;
  assign n6023 = ( n1235 & n2445 ) | ( n1235 & ~n2482 ) | ( n2445 & ~n2482 ) ;
  assign n6024 = ( n1507 & n3400 ) | ( n1507 & n6023 ) | ( n3400 & n6023 ) ;
  assign n6026 = n6025 ^ n6024 ^ n4484 ;
  assign n6027 = ( ~n2691 & n4030 ) | ( ~n2691 & n4836 ) | ( n4030 & n4836 ) ;
  assign n6028 = ( ~n6022 & n6026 ) | ( ~n6022 & n6027 ) | ( n6026 & n6027 ) ;
  assign n6029 = x87 ^ x36 ^ 1'b0 ;
  assign n6030 = ( n1195 & n1276 ) | ( n1195 & ~n3651 ) | ( n1276 & ~n3651 ) ;
  assign n6031 = n3193 ^ n2929 ^ n736 ;
  assign n6032 = n3267 ^ n1839 ^ 1'b0 ;
  assign n6033 = n1514 | n6032 ;
  assign n6034 = ( n4020 & ~n6031 ) | ( n4020 & n6033 ) | ( ~n6031 & n6033 ) ;
  assign n6035 = ( n3774 & n6030 ) | ( n3774 & ~n6034 ) | ( n6030 & ~n6034 ) ;
  assign n6036 = n6035 ^ n5966 ^ x91 ;
  assign n6039 = x18 & ~n3846 ;
  assign n6037 = n5660 ^ n2510 ^ n2459 ;
  assign n6038 = ( n1181 & n3474 ) | ( n1181 & ~n6037 ) | ( n3474 & ~n6037 ) ;
  assign n6040 = n6039 ^ n6038 ^ n2082 ;
  assign n6045 = ~x77 & n1007 ;
  assign n6046 = x224 & ~n641 ;
  assign n6047 = n6045 & n6046 ;
  assign n6041 = n1365 ^ n1117 ^ n645 ;
  assign n6042 = n840 ^ x28 ^ 1'b0 ;
  assign n6043 = n6042 ^ n4987 ^ x208 ;
  assign n6044 = ( ~n548 & n6041 ) | ( ~n548 & n6043 ) | ( n6041 & n6043 ) ;
  assign n6048 = n6047 ^ n6044 ^ 1'b0 ;
  assign n6049 = n2797 & ~n3261 ;
  assign n6050 = ( n1662 & n1834 ) | ( n1662 & ~n6049 ) | ( n1834 & ~n6049 ) ;
  assign n6051 = n6050 ^ n4544 ^ n2006 ;
  assign n6052 = n708 | n1045 ;
  assign n6053 = ~n3947 & n4626 ;
  assign n6054 = ~n597 & n6053 ;
  assign n6055 = n6054 ^ n4641 ^ n2590 ;
  assign n6056 = n6055 ^ n5330 ^ n642 ;
  assign n6057 = n6056 ^ n1814 ^ n1737 ;
  assign n6058 = ( n2570 & n6052 ) | ( n2570 & ~n6057 ) | ( n6052 & ~n6057 ) ;
  assign n6059 = n2431 ^ n752 ^ n505 ;
  assign n6060 = ( n1523 & ~n2664 ) | ( n1523 & n6059 ) | ( ~n2664 & n6059 ) ;
  assign n6061 = n6023 ^ n4547 ^ 1'b0 ;
  assign n6066 = ( n256 & n822 ) | ( n256 & n3701 ) | ( n822 & n3701 ) ;
  assign n6067 = n3971 | n6066 ;
  assign n6062 = ~n752 & n1141 ;
  assign n6063 = ( n1328 & ~n1713 ) | ( n1328 & n6062 ) | ( ~n1713 & n6062 ) ;
  assign n6064 = n6063 ^ n5706 ^ n2674 ;
  assign n6065 = n6020 | n6064 ;
  assign n6068 = n6067 ^ n6065 ^ n4701 ;
  assign n6069 = ( x150 & ~n3142 ) | ( x150 & n6068 ) | ( ~n3142 & n6068 ) ;
  assign n6070 = n6069 ^ n5609 ^ n504 ;
  assign n6071 = n1987 ^ n1040 ^ x130 ;
  assign n6072 = n6071 ^ n3191 ^ n699 ;
  assign n6073 = n6072 ^ n5969 ^ 1'b0 ;
  assign n6075 = n5061 | n5471 ;
  assign n6076 = n3807 & ~n6075 ;
  assign n6077 = n6076 ^ n3621 ^ 1'b0 ;
  assign n6078 = n6077 ^ n1257 ^ 1'b0 ;
  assign n6074 = ( n1270 & n1694 ) | ( n1270 & ~n2031 ) | ( n1694 & ~n2031 ) ;
  assign n6079 = n6078 ^ n6074 ^ n634 ;
  assign n6080 = ( n2846 & n3022 ) | ( n2846 & ~n4857 ) | ( n3022 & ~n4857 ) ;
  assign n6081 = n6080 ^ n3019 ^ n2217 ;
  assign n6082 = ( n2048 & n3509 ) | ( n2048 & ~n5309 ) | ( n3509 & ~n5309 ) ;
  assign n6083 = n6082 ^ n3269 ^ n666 ;
  assign n6084 = ( ~n4410 & n5748 ) | ( ~n4410 & n6083 ) | ( n5748 & n6083 ) ;
  assign n6085 = n295 & n818 ;
  assign n6086 = n2720 & n6085 ;
  assign n6087 = n6086 ^ n5625 ^ n4958 ;
  assign n6088 = n1760 | n5720 ;
  assign n6089 = n6087 & ~n6088 ;
  assign n6096 = ( n669 & ~n1052 ) | ( n669 & n1461 ) | ( ~n1052 & n1461 ) ;
  assign n6097 = n2104 | n6096 ;
  assign n6098 = n6097 ^ n1958 ^ 1'b0 ;
  assign n6099 = ( ~x79 & x105 ) | ( ~x79 & n6098 ) | ( x105 & n6098 ) ;
  assign n6090 = ( n607 & n2280 ) | ( n607 & n2833 ) | ( n2280 & n2833 ) ;
  assign n6091 = n2891 | n3197 ;
  assign n6092 = n6091 ^ n2296 ^ 1'b0 ;
  assign n6093 = n6092 ^ n1080 ^ x101 ;
  assign n6094 = n6090 | n6093 ;
  assign n6095 = n615 & ~n6094 ;
  assign n6100 = n6099 ^ n6095 ^ 1'b0 ;
  assign n6101 = ( ~n809 & n1108 ) | ( ~n809 & n1442 ) | ( n1108 & n1442 ) ;
  assign n6108 = n1274 | n4771 ;
  assign n6102 = ( n703 & n2707 ) | ( n703 & n5846 ) | ( n2707 & n5846 ) ;
  assign n6103 = n6102 ^ n4431 ^ n1538 ;
  assign n6105 = ( n1610 & ~n2530 ) | ( n1610 & n5343 ) | ( ~n2530 & n5343 ) ;
  assign n6104 = ~n423 & n1721 ;
  assign n6106 = n6105 ^ n6104 ^ 1'b0 ;
  assign n6107 = n6103 & n6106 ;
  assign n6109 = n6108 ^ n6107 ^ 1'b0 ;
  assign n6110 = ~n1183 & n1276 ;
  assign n6111 = n4631 ^ n2530 ^ n2269 ;
  assign n6112 = n5162 & n6111 ;
  assign n6113 = ( n1838 & n2294 ) | ( n1838 & ~n6112 ) | ( n2294 & ~n6112 ) ;
  assign n6114 = ( ~n1212 & n6110 ) | ( ~n1212 & n6113 ) | ( n6110 & n6113 ) ;
  assign n6115 = n6114 ^ n5245 ^ 1'b0 ;
  assign n6116 = n5652 & ~n6115 ;
  assign n6117 = n2581 ^ n1852 ^ x191 ;
  assign n6118 = ( n422 & n3237 ) | ( n422 & ~n6117 ) | ( n3237 & ~n6117 ) ;
  assign n6119 = n6118 ^ n4389 ^ n529 ;
  assign n6126 = n533 | n2633 ;
  assign n6127 = n6126 ^ n1659 ^ n1625 ;
  assign n6128 = n6127 ^ n5586 ^ n4772 ;
  assign n6121 = n735 | n1997 ;
  assign n6122 = n6121 ^ n644 ^ n512 ;
  assign n6123 = n6122 ^ n4134 ^ n658 ;
  assign n6120 = ( n1503 & n1713 ) | ( n1503 & ~n4690 ) | ( n1713 & ~n4690 ) ;
  assign n6124 = n6123 ^ n6120 ^ n2059 ;
  assign n6125 = ( n869 & ~n1048 ) | ( n869 & n6124 ) | ( ~n1048 & n6124 ) ;
  assign n6129 = n6128 ^ n6125 ^ n4245 ;
  assign n6130 = n3743 ^ n1496 ^ 1'b0 ;
  assign n6131 = ( n1081 & n3651 ) | ( n1081 & ~n6130 ) | ( n3651 & ~n6130 ) ;
  assign n6132 = n4608 ^ n2918 ^ x216 ;
  assign n6133 = n2567 & ~n6132 ;
  assign n6134 = n6133 ^ n6113 ^ 1'b0 ;
  assign n6135 = ~n6131 & n6134 ;
  assign n6136 = n6129 & n6135 ;
  assign n6137 = n5560 ^ n1427 ^ x244 ;
  assign n6138 = n1453 ^ n1329 ^ x126 ;
  assign n6139 = n6138 ^ n2096 ^ x44 ;
  assign n6140 = n2542 ^ n1852 ^ n831 ;
  assign n6141 = ( ~n2854 & n4197 ) | ( ~n2854 & n6140 ) | ( n4197 & n6140 ) ;
  assign n6142 = ( ~x221 & n427 ) | ( ~x221 & n6141 ) | ( n427 & n6141 ) ;
  assign n6143 = ( n830 & n6139 ) | ( n830 & ~n6142 ) | ( n6139 & ~n6142 ) ;
  assign n6145 = ( ~n1938 & n2952 ) | ( ~n1938 & n3293 ) | ( n2952 & n3293 ) ;
  assign n6144 = n1605 & ~n4439 ;
  assign n6146 = n6145 ^ n6144 ^ n355 ;
  assign n6147 = n6143 & ~n6146 ;
  assign n6148 = n6147 ^ n4261 ^ 1'b0 ;
  assign n6149 = n3497 & ~n3900 ;
  assign n6150 = n6149 ^ n1459 ^ 1'b0 ;
  assign n6151 = ~n3969 & n6150 ;
  assign n6152 = ( n6137 & ~n6148 ) | ( n6137 & n6151 ) | ( ~n6148 & n6151 ) ;
  assign n6153 = ( n931 & n3867 ) | ( n931 & ~n6152 ) | ( n3867 & ~n6152 ) ;
  assign n6154 = n3609 ^ n1416 ^ 1'b0 ;
  assign n6155 = ( n3612 & ~n4305 ) | ( n3612 & n6154 ) | ( ~n4305 & n6154 ) ;
  assign n6156 = n6155 ^ n3898 ^ x187 ;
  assign n6164 = n2327 ^ n1045 ^ n695 ;
  assign n6165 = ( ~n1223 & n1381 ) | ( ~n1223 & n6164 ) | ( n1381 & n6164 ) ;
  assign n6161 = n3713 ^ n1033 ^ 1'b0 ;
  assign n6162 = ( n1213 & ~n1511 ) | ( n1213 & n6161 ) | ( ~n1511 & n6161 ) ;
  assign n6163 = ~n2511 & n6162 ;
  assign n6166 = n6165 ^ n6163 ^ 1'b0 ;
  assign n6157 = n1187 ^ x59 ^ x56 ;
  assign n6158 = ( n1219 & ~n3014 ) | ( n1219 & n5304 ) | ( ~n3014 & n5304 ) ;
  assign n6159 = n6158 ^ n4597 ^ n518 ;
  assign n6160 = n6157 & n6159 ;
  assign n6167 = n6166 ^ n6160 ^ n569 ;
  assign n6168 = n781 | n2169 ;
  assign n6169 = n6168 ^ n2071 ^ 1'b0 ;
  assign n6170 = n6169 ^ n2245 ^ n736 ;
  assign n6171 = n363 & n3271 ;
  assign n6172 = n6171 ^ n2401 ^ n1588 ;
  assign n6173 = ( n2887 & n4996 ) | ( n2887 & ~n6172 ) | ( n4996 & ~n6172 ) ;
  assign n6174 = ( n1675 & n6170 ) | ( n1675 & n6173 ) | ( n6170 & n6173 ) ;
  assign n6186 = n887 ^ x123 ^ 1'b0 ;
  assign n6187 = n1776 & n6186 ;
  assign n6182 = x110 & ~n1682 ;
  assign n6183 = ( n1609 & ~n1834 ) | ( n1609 & n5843 ) | ( ~n1834 & n5843 ) ;
  assign n6184 = ( n1342 & n6182 ) | ( n1342 & n6183 ) | ( n6182 & n6183 ) ;
  assign n6175 = n4946 ^ n4430 ^ n1999 ;
  assign n6176 = n335 & n1221 ;
  assign n6177 = ~n6175 & n6176 ;
  assign n6178 = n6177 ^ n4973 ^ n729 ;
  assign n6179 = ( n1227 & ~n1834 ) | ( n1227 & n6178 ) | ( ~n1834 & n6178 ) ;
  assign n6180 = n3654 ^ n1007 ^ n310 ;
  assign n6181 = ( n848 & n6179 ) | ( n848 & n6180 ) | ( n6179 & n6180 ) ;
  assign n6185 = n6184 ^ n6181 ^ n5663 ;
  assign n6188 = n6187 ^ n6185 ^ n4021 ;
  assign n6198 = n1944 & n3595 ;
  assign n6199 = n6198 ^ n5296 ^ 1'b0 ;
  assign n6200 = ( n880 & n3300 ) | ( n880 & ~n6199 ) | ( n3300 & ~n6199 ) ;
  assign n6191 = n3206 & ~n3534 ;
  assign n6192 = n622 ^ n468 ^ n345 ;
  assign n6193 = ~n543 & n1398 ;
  assign n6194 = ~n6192 & n6193 ;
  assign n6195 = n6194 ^ n4149 ^ 1'b0 ;
  assign n6196 = n6195 ^ n2221 ^ 1'b0 ;
  assign n6197 = ( n4773 & ~n6191 ) | ( n4773 & n6196 ) | ( ~n6191 & n6196 ) ;
  assign n6201 = n6200 ^ n6197 ^ n2704 ;
  assign n6189 = n4040 ^ n2558 ^ x72 ;
  assign n6190 = ~n5718 & n6189 ;
  assign n6202 = n6201 ^ n6190 ^ n3298 ;
  assign n6203 = n5555 ^ n4842 ^ 1'b0 ;
  assign n6204 = n631 | n2661 ;
  assign n6205 = n6204 ^ n5874 ^ n3298 ;
  assign n6206 = n361 ^ x221 ^ x55 ;
  assign n6207 = n6206 ^ n3819 ^ n1854 ;
  assign n6208 = ( x77 & ~n1428 ) | ( x77 & n2794 ) | ( ~n1428 & n2794 ) ;
  assign n6209 = n2364 & ~n3660 ;
  assign n6210 = ( ~n6207 & n6208 ) | ( ~n6207 & n6209 ) | ( n6208 & n6209 ) ;
  assign n6211 = ~n2164 & n2293 ;
  assign n6212 = n6211 ^ n813 ^ 1'b0 ;
  assign n6213 = ( n839 & n1830 ) | ( n839 & ~n6212 ) | ( n1830 & ~n6212 ) ;
  assign n6214 = n2362 ^ n1935 ^ n469 ;
  assign n6215 = n6214 ^ n4644 ^ n565 ;
  assign n6216 = ( ~n565 & n6213 ) | ( ~n565 & n6215 ) | ( n6213 & n6215 ) ;
  assign n6218 = n1308 | n3669 ;
  assign n6217 = ~n1010 & n4260 ;
  assign n6219 = n6218 ^ n6217 ^ 1'b0 ;
  assign n6220 = n2066 ^ n363 ^ 1'b0 ;
  assign n6221 = n3288 | n6220 ;
  assign n6222 = n1380 ^ n1106 ^ n982 ;
  assign n6223 = ( n1444 & ~n6221 ) | ( n1444 & n6222 ) | ( ~n6221 & n6222 ) ;
  assign n6224 = n4160 ^ n1823 ^ n1700 ;
  assign n6225 = n6224 ^ n1988 ^ 1'b0 ;
  assign n6226 = ~n6223 & n6225 ;
  assign n6227 = ( n1010 & n1617 ) | ( n1010 & n6226 ) | ( n1617 & n6226 ) ;
  assign n6228 = n6227 ^ n2699 ^ n842 ;
  assign n6229 = n6228 ^ n4781 ^ 1'b0 ;
  assign n6230 = n558 & ~n658 ;
  assign n6231 = n6230 ^ n1902 ^ 1'b0 ;
  assign n6232 = n6231 ^ n3450 ^ n1010 ;
  assign n6233 = ~n2818 & n6232 ;
  assign n6234 = n6233 ^ n5494 ^ 1'b0 ;
  assign n6236 = n260 | n651 ;
  assign n6237 = n1241 | n6236 ;
  assign n6235 = n5783 ^ n1904 ^ n590 ;
  assign n6238 = n6237 ^ n6235 ^ n1114 ;
  assign n6240 = n4184 ^ n2487 ^ n848 ;
  assign n6241 = ~n3768 & n6240 ;
  assign n6239 = n2326 & ~n5212 ;
  assign n6242 = n6241 ^ n6239 ^ 1'b0 ;
  assign n6243 = ( n2125 & n6238 ) | ( n2125 & ~n6242 ) | ( n6238 & ~n6242 ) ;
  assign n6244 = n2290 & ~n3297 ;
  assign n6245 = n6244 ^ n3374 ^ 1'b0 ;
  assign n6246 = ~n846 & n6245 ;
  assign n6247 = n3776 & n6246 ;
  assign n6248 = n5367 ^ n3237 ^ 1'b0 ;
  assign n6249 = n6248 ^ n2514 ^ n523 ;
  assign n6250 = n6249 ^ n4844 ^ n4683 ;
  assign n6251 = ~n4878 & n6250 ;
  assign n6252 = n6247 & n6251 ;
  assign n6253 = n457 & ~n6252 ;
  assign n6254 = n1402 ^ n402 ^ 1'b0 ;
  assign n6255 = n876 & n6254 ;
  assign n6256 = n6149 ^ n5836 ^ n3681 ;
  assign n6257 = n3798 ^ n2954 ^ n688 ;
  assign n6258 = n6257 ^ n4618 ^ n302 ;
  assign n6259 = n6258 ^ n4631 ^ 1'b0 ;
  assign n6260 = n6259 ^ n2459 ^ n1658 ;
  assign n6261 = ( n2064 & n3967 ) | ( n2064 & n6260 ) | ( n3967 & n6260 ) ;
  assign n6262 = n2816 ^ n2316 ^ n488 ;
  assign n6266 = n5435 ^ n3326 ^ n2707 ;
  assign n6263 = x191 & ~n2222 ;
  assign n6264 = n6263 ^ n542 ^ 1'b0 ;
  assign n6265 = n6264 ^ n2372 ^ n523 ;
  assign n6267 = n6266 ^ n6265 ^ n863 ;
  assign n6270 = ( n1669 & n2119 ) | ( n1669 & ~n3568 ) | ( n2119 & ~n3568 ) ;
  assign n6268 = n2977 ^ n643 ^ 1'b0 ;
  assign n6269 = ~n2774 & n6268 ;
  assign n6271 = n6270 ^ n6269 ^ 1'b0 ;
  assign n6272 = ~n6267 & n6271 ;
  assign n6273 = n6272 ^ n1964 ^ 1'b0 ;
  assign n6274 = ( ~n2977 & n6262 ) | ( ~n2977 & n6273 ) | ( n6262 & n6273 ) ;
  assign n6275 = n6274 ^ n6248 ^ n3790 ;
  assign n6276 = ~n3577 & n4164 ;
  assign n6277 = n5647 ^ n2162 ^ n1957 ;
  assign n6278 = ( ~n352 & n6276 ) | ( ~n352 & n6277 ) | ( n6276 & n6277 ) ;
  assign n6279 = ( ~n465 & n4718 ) | ( ~n465 & n6278 ) | ( n4718 & n6278 ) ;
  assign n6280 = n6279 ^ n3769 ^ n3291 ;
  assign n6287 = n3568 ^ n3456 ^ n686 ;
  assign n6288 = n6287 ^ n4882 ^ n3130 ;
  assign n6289 = n1657 | n6288 ;
  assign n6290 = n6289 ^ x142 ^ 1'b0 ;
  assign n6291 = n2178 & n6290 ;
  assign n6292 = n6291 ^ n1809 ^ 1'b0 ;
  assign n6286 = n4160 ^ n3875 ^ n2040 ;
  assign n6281 = ~n1448 & n1703 ;
  assign n6282 = ~n2335 & n6281 ;
  assign n6283 = n6282 ^ n5376 ^ x154 ;
  assign n6284 = n3212 & n5466 ;
  assign n6285 = ( n3356 & ~n6283 ) | ( n3356 & n6284 ) | ( ~n6283 & n6284 ) ;
  assign n6293 = n6292 ^ n6286 ^ n6285 ;
  assign n6297 = ( x147 & n439 ) | ( x147 & ~n2557 ) | ( n439 & ~n2557 ) ;
  assign n6294 = n5562 ^ n4061 ^ n877 ;
  assign n6295 = ( n2600 & ~n4896 ) | ( n2600 & n6294 ) | ( ~n4896 & n6294 ) ;
  assign n6296 = n6295 ^ n5751 ^ n1582 ;
  assign n6298 = n6297 ^ n6296 ^ n2031 ;
  assign n6299 = ~n601 & n2020 ;
  assign n6300 = n6299 ^ n2447 ^ 1'b0 ;
  assign n6301 = n3880 ^ n2201 ^ n565 ;
  assign n6302 = n6301 ^ n3969 ^ n2017 ;
  assign n6303 = n4347 ^ n2687 ^ n990 ;
  assign n6304 = ( n1525 & ~n3129 ) | ( n1525 & n5963 ) | ( ~n3129 & n5963 ) ;
  assign n6305 = ~n6303 & n6304 ;
  assign n6306 = ( x157 & ~n6302 ) | ( x157 & n6305 ) | ( ~n6302 & n6305 ) ;
  assign n6307 = n1936 | n3891 ;
  assign n6308 = n6306 | n6307 ;
  assign n6309 = n6308 ^ n3266 ^ n1565 ;
  assign n6310 = n6309 ^ n4039 ^ n3200 ;
  assign n6311 = n6065 ^ n3610 ^ 1'b0 ;
  assign n6312 = n3769 | n6311 ;
  assign n6313 = n992 ^ n544 ^ n392 ;
  assign n6314 = ( x45 & ~n1243 ) | ( x45 & n6313 ) | ( ~n1243 & n6313 ) ;
  assign n6315 = x248 & ~n6314 ;
  assign n6316 = n6315 ^ n2197 ^ 1'b0 ;
  assign n6317 = n1021 | n1770 ;
  assign n6318 = x191 & n711 ;
  assign n6319 = n6318 ^ n5459 ^ 1'b0 ;
  assign n6320 = n890 & n4360 ;
  assign n6321 = n6320 ^ n5128 ^ 1'b0 ;
  assign n6322 = n998 | n6321 ;
  assign n6323 = n6319 & ~n6322 ;
  assign n6324 = ( n6316 & ~n6317 ) | ( n6316 & n6323 ) | ( ~n6317 & n6323 ) ;
  assign n6325 = ( n5003 & n6312 ) | ( n5003 & ~n6324 ) | ( n6312 & ~n6324 ) ;
  assign n6326 = n6292 ^ n3553 ^ n1169 ;
  assign n6327 = n1161 & n6326 ;
  assign n6328 = ( ~x119 & n1606 ) | ( ~x119 & n1617 ) | ( n1606 & n1617 ) ;
  assign n6329 = n6328 ^ n3971 ^ n2894 ;
  assign n6330 = n3650 ^ n2927 ^ n1050 ;
  assign n6331 = ( n5405 & n6329 ) | ( n5405 & ~n6330 ) | ( n6329 & ~n6330 ) ;
  assign n6336 = n3143 ^ n2819 ^ n1778 ;
  assign n6332 = n1879 & ~n1893 ;
  assign n6333 = ~n2410 & n6332 ;
  assign n6334 = n5616 | n6333 ;
  assign n6335 = n6334 ^ n1766 ^ 1'b0 ;
  assign n6337 = n6336 ^ n6335 ^ n5058 ;
  assign n6338 = ~n3763 & n6337 ;
  assign n6339 = n2659 ^ n1715 ^ n319 ;
  assign n6340 = ( n5169 & ~n6338 ) | ( n5169 & n6339 ) | ( ~n6338 & n6339 ) ;
  assign n6341 = n1559 ^ n1352 ^ n1088 ;
  assign n6342 = ( n1103 & n2110 ) | ( n1103 & ~n3743 ) | ( n2110 & ~n3743 ) ;
  assign n6343 = n1731 & ~n6342 ;
  assign n6344 = n6343 ^ n709 ^ 1'b0 ;
  assign n6345 = ( ~n1961 & n6341 ) | ( ~n1961 & n6344 ) | ( n6341 & n6344 ) ;
  assign n6346 = ~n2710 & n6345 ;
  assign n6347 = n6346 ^ n3754 ^ n3648 ;
  assign n6348 = n5043 & ~n6347 ;
  assign n6349 = n6348 ^ n3317 ^ 1'b0 ;
  assign n6350 = ( ~n545 & n1312 ) | ( ~n545 & n2036 ) | ( n1312 & n2036 ) ;
  assign n6351 = n6350 ^ n2285 ^ n688 ;
  assign n6352 = ( n2519 & ~n2659 ) | ( n2519 & n6351 ) | ( ~n2659 & n6351 ) ;
  assign n6353 = n6352 ^ n3893 ^ 1'b0 ;
  assign n6354 = n4577 ^ n662 ^ 1'b0 ;
  assign n6355 = n6354 ^ n2204 ^ n1383 ;
  assign n6356 = n6355 ^ x97 ^ 1'b0 ;
  assign n6357 = n3587 ^ n2283 ^ n1486 ;
  assign n6358 = n6357 ^ n6313 ^ n3416 ;
  assign n6359 = ( n366 & n3259 ) | ( n366 & ~n3744 ) | ( n3259 & ~n3744 ) ;
  assign n6360 = ( x144 & n3208 ) | ( x144 & n3628 ) | ( n3208 & n3628 ) ;
  assign n6361 = ( n1915 & n6359 ) | ( n1915 & ~n6360 ) | ( n6359 & ~n6360 ) ;
  assign n6362 = n6361 ^ n1125 ^ 1'b0 ;
  assign n6363 = n526 & ~n1057 ;
  assign n6364 = n1272 & n6363 ;
  assign n6365 = ( ~n1734 & n2874 ) | ( ~n1734 & n6364 ) | ( n2874 & n6364 ) ;
  assign n6366 = ( n1088 & ~n2848 ) | ( n1088 & n6365 ) | ( ~n2848 & n6365 ) ;
  assign n6367 = x185 & n6366 ;
  assign n6368 = n6367 ^ n1404 ^ 1'b0 ;
  assign n6369 = n6368 ^ n4407 ^ n3573 ;
  assign n6370 = n3754 & n4447 ;
  assign n6371 = n2239 & n6370 ;
  assign n6372 = ( ~n3004 & n4552 ) | ( ~n3004 & n6371 ) | ( n4552 & n6371 ) ;
  assign n6373 = ( n2945 & n3674 ) | ( n2945 & n6372 ) | ( n3674 & n6372 ) ;
  assign n6374 = ( n320 & n1448 ) | ( n320 & ~n1868 ) | ( n1448 & ~n1868 ) ;
  assign n6381 = n4635 ^ n3308 ^ n2146 ;
  assign n6375 = n1135 & ~n1582 ;
  assign n6376 = n6375 ^ n803 ^ 1'b0 ;
  assign n6377 = ~n688 & n2343 ;
  assign n6378 = n1826 & n6377 ;
  assign n6379 = n1255 & ~n6378 ;
  assign n6380 = n6376 & n6379 ;
  assign n6382 = n6381 ^ n6380 ^ x14 ;
  assign n6383 = n6374 & ~n6382 ;
  assign n6384 = ( ~n2060 & n2456 ) | ( ~n2060 & n5454 ) | ( n2456 & n5454 ) ;
  assign n6385 = ( ~n4787 & n6383 ) | ( ~n4787 & n6384 ) | ( n6383 & n6384 ) ;
  assign n6386 = n3668 & n5088 ;
  assign n6387 = ~n2664 & n6386 ;
  assign n6388 = n6387 ^ n5643 ^ n3444 ;
  assign n6389 = n5270 ^ n5094 ^ n4864 ;
  assign n6390 = n480 & n996 ;
  assign n6391 = n6390 ^ n3542 ^ n3014 ;
  assign n6392 = ( x125 & ~n4061 ) | ( x125 & n6391 ) | ( ~n4061 & n6391 ) ;
  assign n6397 = ( x224 & x234 ) | ( x224 & ~n3112 ) | ( x234 & ~n3112 ) ;
  assign n6396 = x99 | n4019 ;
  assign n6393 = n5417 ^ n3026 ^ 1'b0 ;
  assign n6394 = n1547 & ~n2448 ;
  assign n6395 = ( n5734 & n6393 ) | ( n5734 & n6394 ) | ( n6393 & n6394 ) ;
  assign n6398 = n6397 ^ n6396 ^ n6395 ;
  assign n6399 = n3570 ^ n1383 ^ n1107 ;
  assign n6400 = ( ~x170 & n363 ) | ( ~x170 & n2350 ) | ( n363 & n2350 ) ;
  assign n6401 = ( x62 & n840 ) | ( x62 & ~n3144 ) | ( n840 & ~n3144 ) ;
  assign n6402 = ( ~n6399 & n6400 ) | ( ~n6399 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6403 = n6402 ^ n3384 ^ 1'b0 ;
  assign n6415 = ( ~n662 & n2509 ) | ( ~n662 & n3743 ) | ( n2509 & n3743 ) ;
  assign n6413 = n950 & ~n1197 ;
  assign n6408 = n3383 ^ n3191 ^ n2838 ;
  assign n6409 = n6408 ^ n3617 ^ n265 ;
  assign n6410 = n5482 ^ n3614 ^ n2953 ;
  assign n6411 = n4406 ^ n3543 ^ n2018 ;
  assign n6412 = ( ~n6409 & n6410 ) | ( ~n6409 & n6411 ) | ( n6410 & n6411 ) ;
  assign n6404 = n894 & ~n1378 ;
  assign n6414 = n6413 ^ n6412 ^ n6404 ;
  assign n6416 = n6415 ^ n6414 ^ n6023 ;
  assign n6405 = n6404 ^ n4426 ^ n1060 ;
  assign n6406 = n6405 ^ n1504 ^ n571 ;
  assign n6407 = n6406 ^ n5805 ^ n1840 ;
  assign n6417 = n6416 ^ n6407 ^ n1062 ;
  assign n6418 = n6417 ^ n1801 ^ 1'b0 ;
  assign n6419 = n5393 & ~n6418 ;
  assign n6432 = n3260 ^ n892 ^ 1'b0 ;
  assign n6433 = ( n2349 & n3375 ) | ( n2349 & ~n6432 ) | ( n3375 & ~n6432 ) ;
  assign n6420 = n5290 & n5814 ;
  assign n6421 = n6420 ^ n1372 ^ 1'b0 ;
  assign n6422 = ( n897 & n1707 ) | ( n897 & ~n2453 ) | ( n1707 & ~n2453 ) ;
  assign n6423 = n6422 ^ n2262 ^ n2020 ;
  assign n6424 = ( n1667 & n4973 ) | ( n1667 & ~n5310 ) | ( n4973 & ~n5310 ) ;
  assign n6425 = ( ~x215 & n2487 ) | ( ~x215 & n6424 ) | ( n2487 & n6424 ) ;
  assign n6426 = ( n2765 & ~n6423 ) | ( n2765 & n6425 ) | ( ~n6423 & n6425 ) ;
  assign n6427 = n6421 & n6426 ;
  assign n6428 = ~n263 & n3409 ;
  assign n6429 = n6428 ^ n3115 ^ 1'b0 ;
  assign n6430 = n6429 ^ n4364 ^ n2187 ;
  assign n6431 = ( ~n5210 & n6427 ) | ( ~n5210 & n6430 ) | ( n6427 & n6430 ) ;
  assign n6434 = n6433 ^ n6431 ^ n5493 ;
  assign n6435 = n1963 ^ n475 ^ 1'b0 ;
  assign n6436 = n3295 & ~n6031 ;
  assign n6437 = ( ~n3358 & n6435 ) | ( ~n3358 & n6436 ) | ( n6435 & n6436 ) ;
  assign n6438 = n2437 ^ n1049 ^ x174 ;
  assign n6439 = x115 & ~n5477 ;
  assign n6440 = x148 & n6439 ;
  assign n6441 = n848 & n6440 ;
  assign n6445 = n5985 ^ n1219 ^ 1'b0 ;
  assign n6446 = n904 & n6445 ;
  assign n6443 = ( n543 & ~n3148 ) | ( n543 & n3928 ) | ( ~n3148 & n3928 ) ;
  assign n6444 = n6443 ^ n2466 ^ 1'b0 ;
  assign n6442 = n465 & ~n5679 ;
  assign n6447 = n6446 ^ n6444 ^ n6442 ;
  assign n6448 = n6447 ^ n4407 ^ n439 ;
  assign n6449 = ( ~n6438 & n6441 ) | ( ~n6438 & n6448 ) | ( n6441 & n6448 ) ;
  assign n6450 = x29 | n5086 ;
  assign n6451 = ~n867 & n6450 ;
  assign n6452 = n6451 ^ n1486 ^ 1'b0 ;
  assign n6453 = n3913 & n4366 ;
  assign n6454 = ~n6452 & n6453 ;
  assign n6455 = x11 | n6454 ;
  assign n6456 = ( n1200 & ~n2543 ) | ( n1200 & n3375 ) | ( ~n2543 & n3375 ) ;
  assign n6457 = n1208 | n6456 ;
  assign n6458 = n6457 ^ n2659 ^ 1'b0 ;
  assign n6459 = n4120 ^ n3861 ^ n2062 ;
  assign n6460 = n6458 & n6459 ;
  assign n6461 = n6112 ^ n5888 ^ n2716 ;
  assign n6462 = n767 & n5021 ;
  assign n6463 = n1757 & n6462 ;
  assign n6464 = n6463 ^ n4361 ^ n686 ;
  assign n6465 = ( n2145 & ~n3566 ) | ( n2145 & n3752 ) | ( ~n3566 & n3752 ) ;
  assign n6466 = n4904 & ~n6465 ;
  assign n6467 = n6464 & n6466 ;
  assign n6468 = ( ~n633 & n914 ) | ( ~n633 & n4427 ) | ( n914 & n4427 ) ;
  assign n6469 = n2126 & n6468 ;
  assign n6470 = ~n1196 & n6469 ;
  assign n6471 = n3359 ^ n1461 ^ 1'b0 ;
  assign n6472 = n6470 | n6471 ;
  assign n6473 = n1508 | n5976 ;
  assign n6474 = ( n567 & n4992 ) | ( n567 & n6473 ) | ( n4992 & n6473 ) ;
  assign n6475 = x121 & n590 ;
  assign n6476 = n6475 ^ n3315 ^ n3308 ;
  assign n6477 = n6476 ^ n3314 ^ n1197 ;
  assign n6478 = n348 & n1557 ;
  assign n6479 = n6478 ^ n1793 ^ 1'b0 ;
  assign n6484 = ( ~n850 & n1669 ) | ( ~n850 & n2772 ) | ( n1669 & n2772 ) ;
  assign n6480 = n709 & ~n3479 ;
  assign n6481 = ~n2464 & n6480 ;
  assign n6482 = ~n6212 & n6481 ;
  assign n6483 = x81 & ~n6482 ;
  assign n6485 = n6484 ^ n6483 ^ n2602 ;
  assign n6486 = n328 | n545 ;
  assign n6487 = ( ~n6479 & n6485 ) | ( ~n6479 & n6486 ) | ( n6485 & n6486 ) ;
  assign n6488 = n6487 ^ n4694 ^ 1'b0 ;
  assign n6489 = n6477 & n6488 ;
  assign n6492 = n4341 ^ n3376 ^ n1365 ;
  assign n6490 = n4455 ^ n1795 ^ 1'b0 ;
  assign n6491 = x141 & ~n6490 ;
  assign n6493 = n6492 ^ n6491 ^ n1690 ;
  assign n6494 = ( n3633 & n4737 ) | ( n3633 & n6493 ) | ( n4737 & n6493 ) ;
  assign n6495 = n6489 & n6494 ;
  assign n6496 = ( ~n6472 & n6474 ) | ( ~n6472 & n6495 ) | ( n6474 & n6495 ) ;
  assign n6497 = n3007 ^ n1987 ^ n1297 ;
  assign n6498 = n6497 ^ x180 ^ 1'b0 ;
  assign n6499 = x77 & n1453 ;
  assign n6500 = ~x62 & n6499 ;
  assign n6501 = n6500 ^ n2970 ^ n2325 ;
  assign n6502 = n4701 ^ n459 ^ x134 ;
  assign n6503 = ~n6501 & n6502 ;
  assign n6504 = n6503 ^ n5341 ^ n5268 ;
  assign n6505 = ( n4222 & n6498 ) | ( n4222 & n6504 ) | ( n6498 & n6504 ) ;
  assign n6507 = ( x200 & n4091 ) | ( x200 & ~n5154 ) | ( n4091 & ~n5154 ) ;
  assign n6506 = n1747 ^ n1024 ^ x154 ;
  assign n6508 = n6507 ^ n6506 ^ n6374 ;
  assign n6509 = n1335 ^ x38 ^ 1'b0 ;
  assign n6510 = ( n5829 & ~n6178 ) | ( n5829 & n6509 ) | ( ~n6178 & n6509 ) ;
  assign n6517 = ( n2414 & n2428 ) | ( n2414 & n4361 ) | ( n2428 & n4361 ) ;
  assign n6518 = n6517 ^ n6365 ^ 1'b0 ;
  assign n6519 = n2932 & ~n6518 ;
  assign n6516 = ~n4454 & n6480 ;
  assign n6520 = n6519 ^ n6516 ^ n5287 ;
  assign n6511 = n2051 ^ n430 ^ 1'b0 ;
  assign n6512 = n3448 | n6511 ;
  assign n6513 = n1027 & ~n5086 ;
  assign n6514 = n6513 ^ n5335 ^ 1'b0 ;
  assign n6515 = n6512 | n6514 ;
  assign n6521 = n6520 ^ n6515 ^ 1'b0 ;
  assign n6522 = ( n2285 & n4403 ) | ( n2285 & n6521 ) | ( n4403 & n6521 ) ;
  assign n6523 = n6522 ^ n4250 ^ n1676 ;
  assign n6524 = ( ~n1031 & n1787 ) | ( ~n1031 & n5326 ) | ( n1787 & n5326 ) ;
  assign n6525 = n6524 ^ n2211 ^ n1435 ;
  assign n6526 = n2071 & n5368 ;
  assign n6527 = ( n4354 & ~n6415 ) | ( n4354 & n6526 ) | ( ~n6415 & n6526 ) ;
  assign n6528 = n6525 | n6527 ;
  assign n6531 = n2540 ^ n439 ^ 1'b0 ;
  assign n6529 = n3556 ^ n3097 ^ n2797 ;
  assign n6530 = ( ~n3989 & n4833 ) | ( ~n3989 & n6529 ) | ( n4833 & n6529 ) ;
  assign n6532 = n6531 ^ n6530 ^ n3875 ;
  assign n6533 = n6532 ^ n4933 ^ n2022 ;
  assign n6534 = n4187 | n4443 ;
  assign n6540 = n951 | n1862 ;
  assign n6541 = ( n273 & n2120 ) | ( n273 & n6540 ) | ( n2120 & n6540 ) ;
  assign n6542 = ( n760 & ~n1635 ) | ( n760 & n6541 ) | ( ~n1635 & n6541 ) ;
  assign n6543 = n3297 | n6542 ;
  assign n6536 = ( n1083 & n1891 ) | ( n1083 & n5984 ) | ( n1891 & n5984 ) ;
  assign n6537 = ( n1987 & n2950 ) | ( n1987 & n6536 ) | ( n2950 & n6536 ) ;
  assign n6535 = n4353 ^ n2876 ^ n553 ;
  assign n6538 = n6537 ^ n6535 ^ n3543 ;
  assign n6539 = ( n5953 & n6071 ) | ( n5953 & ~n6538 ) | ( n6071 & ~n6538 ) ;
  assign n6544 = n6543 ^ n6539 ^ n3029 ;
  assign n6545 = x253 & ~n5521 ;
  assign n6546 = n6544 & n6545 ;
  assign n6547 = n6534 & ~n6546 ;
  assign n6548 = n660 & n6547 ;
  assign n6549 = n2755 ^ n2110 ^ n1337 ;
  assign n6550 = n6549 ^ n4669 ^ n1052 ;
  assign n6551 = n2929 ^ n1581 ^ 1'b0 ;
  assign n6552 = ~n1863 & n6551 ;
  assign n6553 = n420 | n981 ;
  assign n6554 = ( ~n5361 & n6552 ) | ( ~n5361 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = ( n1496 & n1942 ) | ( n1496 & ~n6554 ) | ( n1942 & ~n6554 ) ;
  assign n6556 = ( n2372 & n3236 ) | ( n2372 & n6555 ) | ( n3236 & n6555 ) ;
  assign n6557 = n378 & ~n6556 ;
  assign n6558 = n6557 ^ n6018 ^ 1'b0 ;
  assign n6564 = n3035 ^ n2136 ^ 1'b0 ;
  assign n6565 = ( n859 & n6301 ) | ( n859 & n6564 ) | ( n6301 & n6564 ) ;
  assign n6559 = ( n976 & ~n1381 ) | ( n976 & n3743 ) | ( ~n1381 & n3743 ) ;
  assign n6560 = n2318 ^ n1190 ^ n1135 ;
  assign n6561 = n6560 ^ n5435 ^ 1'b0 ;
  assign n6562 = n2864 | n6561 ;
  assign n6563 = ( x87 & ~n6559 ) | ( x87 & n6562 ) | ( ~n6559 & n6562 ) ;
  assign n6566 = n6565 ^ n6563 ^ n3978 ;
  assign n6567 = n691 ^ n558 ^ x133 ;
  assign n6568 = n5199 ^ n3204 ^ 1'b0 ;
  assign n6569 = n6567 & n6568 ;
  assign n6570 = n6544 ^ n6256 ^ n3780 ;
  assign n6571 = n1144 | n3849 ;
  assign n6572 = n3394 | n6039 ;
  assign n6573 = ( n2978 & n6571 ) | ( n2978 & ~n6572 ) | ( n6571 & ~n6572 ) ;
  assign n6578 = ( ~x233 & x244 ) | ( ~x233 & n1220 ) | ( x244 & n1220 ) ;
  assign n6576 = ( n619 & ~n2167 ) | ( n619 & n5923 ) | ( ~n2167 & n5923 ) ;
  assign n6577 = n6576 ^ n4454 ^ n2840 ;
  assign n6574 = ( n912 & ~n1858 ) | ( n912 & n1908 ) | ( ~n1858 & n1908 ) ;
  assign n6575 = ( n1462 & ~n1562 ) | ( n1462 & n6574 ) | ( ~n1562 & n6574 ) ;
  assign n6579 = n6578 ^ n6577 ^ n6575 ;
  assign n6580 = n3589 & n6579 ;
  assign n6581 = n6580 ^ n3629 ^ 1'b0 ;
  assign n6582 = n2882 ^ n2426 ^ n2180 ;
  assign n6583 = n6582 ^ n2597 ^ n943 ;
  assign n6584 = n2693 ^ n2054 ^ 1'b0 ;
  assign n6585 = n6584 ^ n1445 ^ 1'b0 ;
  assign n6586 = ( n901 & n6583 ) | ( n901 & ~n6585 ) | ( n6583 & ~n6585 ) ;
  assign n6596 = n589 & n4277 ;
  assign n6597 = n3731 & n6596 ;
  assign n6587 = n4395 ^ n1198 ^ x101 ;
  assign n6588 = n6587 ^ n6076 ^ n4163 ;
  assign n6591 = n5074 ^ n1726 ^ x84 ;
  assign n6592 = ( ~n1342 & n6257 ) | ( ~n1342 & n6591 ) | ( n6257 & n6591 ) ;
  assign n6589 = n2076 ^ n1690 ^ n1609 ;
  assign n6590 = n6589 ^ n6530 ^ n1402 ;
  assign n6593 = n6592 ^ n6590 ^ n2090 ;
  assign n6594 = n6593 ^ n5762 ^ n4234 ;
  assign n6595 = ( x71 & n6588 ) | ( x71 & n6594 ) | ( n6588 & n6594 ) ;
  assign n6598 = n6597 ^ n6595 ^ n6269 ;
  assign n6599 = n6400 ^ n6361 ^ n4935 ;
  assign n6612 = ( n610 & n809 ) | ( n610 & n981 ) | ( n809 & n981 ) ;
  assign n6613 = ( n1202 & n1694 ) | ( n1202 & n1748 ) | ( n1694 & n1748 ) ;
  assign n6614 = n6613 ^ n3324 ^ n2699 ;
  assign n6615 = n6612 & ~n6614 ;
  assign n6616 = n1384 & n6615 ;
  assign n6600 = n2352 ^ n1436 ^ n724 ;
  assign n6601 = n1639 ^ n722 ^ x123 ;
  assign n6602 = ( ~n578 & n1450 ) | ( ~n578 & n2000 ) | ( n1450 & n2000 ) ;
  assign n6603 = n3168 ^ n859 ^ x95 ;
  assign n6604 = ( n813 & n852 ) | ( n813 & n6603 ) | ( n852 & n6603 ) ;
  assign n6605 = n2064 ^ n1509 ^ 1'b0 ;
  assign n6606 = n6604 & n6605 ;
  assign n6607 = n6606 ^ n5379 ^ n1680 ;
  assign n6608 = ~n2327 & n5728 ;
  assign n6609 = ~n6607 & n6608 ;
  assign n6610 = ( n6601 & n6602 ) | ( n6601 & n6609 ) | ( n6602 & n6609 ) ;
  assign n6611 = n6600 | n6610 ;
  assign n6617 = n6616 ^ n6611 ^ 1'b0 ;
  assign n6618 = n1948 ^ n1223 ^ 1'b0 ;
  assign n6619 = ~n1665 & n6618 ;
  assign n6620 = n262 & ~n980 ;
  assign n6621 = n6620 ^ n4603 ^ n2791 ;
  assign n6622 = n4244 ^ n3484 ^ n670 ;
  assign n6623 = ( n1178 & n3744 ) | ( n1178 & ~n6622 ) | ( n3744 & ~n6622 ) ;
  assign n6631 = ( ~x225 & n539 ) | ( ~x225 & n5287 ) | ( n539 & n5287 ) ;
  assign n6629 = n6042 ^ n4631 ^ x147 ;
  assign n6630 = n6629 ^ n6614 ^ x178 ;
  assign n6627 = n989 & ~n1918 ;
  assign n6624 = n1016 ^ x187 ^ 1'b0 ;
  assign n6625 = n6624 ^ n2868 ^ n1685 ;
  assign n6626 = n6625 ^ n2729 ^ n1592 ;
  assign n6628 = n6627 ^ n6626 ^ n1448 ;
  assign n6632 = n6631 ^ n6630 ^ n6628 ;
  assign n6633 = ( n6621 & n6623 ) | ( n6621 & ~n6632 ) | ( n6623 & ~n6632 ) ;
  assign n6644 = ( n3399 & ~n3558 ) | ( n3399 & n4947 ) | ( ~n3558 & n4947 ) ;
  assign n6636 = n4409 ^ n1779 ^ n1031 ;
  assign n6634 = ( n465 & n2917 ) | ( n465 & n5353 ) | ( n2917 & n5353 ) ;
  assign n6635 = n327 & n6634 ;
  assign n6637 = n6636 ^ n6635 ^ 1'b0 ;
  assign n6638 = n587 | n5676 ;
  assign n6639 = n6638 ^ n5290 ^ 1'b0 ;
  assign n6640 = ( n1007 & n1594 ) | ( n1007 & ~n5064 ) | ( n1594 & ~n5064 ) ;
  assign n6641 = n6640 ^ n5114 ^ n3916 ;
  assign n6642 = ( n5463 & n6639 ) | ( n5463 & n6641 ) | ( n6639 & n6641 ) ;
  assign n6643 = ~n6637 & n6642 ;
  assign n6645 = n6644 ^ n6643 ^ 1'b0 ;
  assign n6646 = ~n6633 & n6645 ;
  assign n6647 = ~n6619 & n6646 ;
  assign n6648 = ( ~n3200 & n6617 ) | ( ~n3200 & n6647 ) | ( n6617 & n6647 ) ;
  assign n6649 = n870 | n1961 ;
  assign n6650 = ~n2223 & n4737 ;
  assign n6651 = n4089 & n6650 ;
  assign n6652 = n6649 & n6651 ;
  assign n6653 = n5819 ^ n3398 ^ 1'b0 ;
  assign n6654 = ( x177 & n589 ) | ( x177 & n612 ) | ( n589 & n612 ) ;
  assign n6655 = n6654 ^ n1571 ^ n1399 ;
  assign n6656 = n683 & ~n6655 ;
  assign n6657 = ( ~n2315 & n6653 ) | ( ~n2315 & n6656 ) | ( n6653 & n6656 ) ;
  assign n6658 = ( n972 & ~n2486 ) | ( n972 & n3725 ) | ( ~n2486 & n3725 ) ;
  assign n6659 = ( n2864 & ~n5053 ) | ( n2864 & n6658 ) | ( ~n5053 & n6658 ) ;
  assign n6660 = n3924 ^ n1419 ^ 1'b0 ;
  assign n6661 = n6660 ^ n4565 ^ n2512 ;
  assign n6662 = n1649 ^ n794 ^ n303 ;
  assign n6663 = ( n1656 & ~n2497 ) | ( n1656 & n3087 ) | ( ~n2497 & n3087 ) ;
  assign n6664 = ~n6662 & n6663 ;
  assign n6665 = ~n6661 & n6664 ;
  assign n6666 = n2566 & n6665 ;
  assign n6667 = n3559 & ~n6666 ;
  assign n6668 = n5266 & n6667 ;
  assign n6672 = n5942 ^ n3120 ^ n1897 ;
  assign n6673 = n6672 ^ n2783 ^ n1836 ;
  assign n6669 = n1137 ^ n301 ^ x24 ;
  assign n6670 = n6669 ^ n4403 ^ n884 ;
  assign n6671 = n6670 ^ n3937 ^ n1503 ;
  assign n6674 = n6673 ^ n6671 ^ 1'b0 ;
  assign n6675 = n2746 ^ n2331 ^ n635 ;
  assign n6676 = ( n3873 & ~n4508 ) | ( n3873 & n6675 ) | ( ~n4508 & n6675 ) ;
  assign n6677 = ( n521 & n3187 ) | ( n521 & ~n3997 ) | ( n3187 & ~n3997 ) ;
  assign n6678 = n652 & ~n1821 ;
  assign n6679 = n1656 & n6678 ;
  assign n6680 = ( n378 & ~n427 ) | ( n378 & n6679 ) | ( ~n427 & n6679 ) ;
  assign n6681 = n6680 ^ n2473 ^ n323 ;
  assign n6682 = ( ~n966 & n1689 ) | ( ~n966 & n2427 ) | ( n1689 & n2427 ) ;
  assign n6683 = n2623 & n6682 ;
  assign n6684 = n6681 & n6683 ;
  assign n6685 = n5146 | n6684 ;
  assign n6686 = n4183 ^ n3172 ^ n1888 ;
  assign n6690 = n5159 ^ n3039 ^ 1'b0 ;
  assign n6691 = n5870 ^ n1441 ^ n1297 ;
  assign n6692 = n6690 & n6691 ;
  assign n6693 = n5196 & n6692 ;
  assign n6687 = ( n1703 & ~n3083 ) | ( n1703 & n6108 ) | ( ~n3083 & n6108 ) ;
  assign n6688 = ( n2343 & n4541 ) | ( n2343 & ~n6687 ) | ( n4541 & ~n6687 ) ;
  assign n6689 = n6688 ^ n4933 ^ n2269 ;
  assign n6694 = n6693 ^ n6689 ^ 1'b0 ;
  assign n6695 = ( n6685 & n6686 ) | ( n6685 & ~n6694 ) | ( n6686 & ~n6694 ) ;
  assign n6696 = ( n1069 & n2254 ) | ( n1069 & n5233 ) | ( n2254 & n5233 ) ;
  assign n6697 = n6696 ^ n4386 ^ n562 ;
  assign n6698 = n3998 ^ n3350 ^ n1724 ;
  assign n6699 = ( n4581 & n4900 ) | ( n4581 & ~n6698 ) | ( n4900 & ~n6698 ) ;
  assign n6700 = ( n1135 & n3345 ) | ( n1135 & ~n6699 ) | ( n3345 & ~n6699 ) ;
  assign n6701 = ( n900 & n4037 ) | ( n900 & n6090 ) | ( n4037 & n6090 ) ;
  assign n6702 = ( n575 & ~n6061 ) | ( n575 & n6701 ) | ( ~n6061 & n6701 ) ;
  assign n6703 = n3761 ^ n2606 ^ 1'b0 ;
  assign n6704 = n5102 ^ n1289 ^ n721 ;
  assign n6713 = n284 & ~n2772 ;
  assign n6714 = ~n2305 & n6713 ;
  assign n6712 = ( ~x66 & n898 ) | ( ~x66 & n4166 ) | ( n898 & n4166 ) ;
  assign n6715 = n6714 ^ n6712 ^ n4181 ;
  assign n6708 = n2517 ^ n980 ^ n641 ;
  assign n6709 = n468 & n6708 ;
  assign n6710 = ( n4040 & n6183 ) | ( n4040 & n6709 ) | ( n6183 & n6709 ) ;
  assign n6705 = n2476 ^ n511 ^ 1'b0 ;
  assign n6706 = n1652 | n6705 ;
  assign n6707 = n6706 ^ n5872 ^ x104 ;
  assign n6711 = n6710 ^ n6707 ^ n3721 ;
  assign n6716 = n6715 ^ n6711 ^ n6152 ;
  assign n6718 = ( ~n384 & n1928 ) | ( ~n384 & n2352 ) | ( n1928 & n2352 ) ;
  assign n6717 = n672 | n5894 ;
  assign n6719 = n6718 ^ n6717 ^ 1'b0 ;
  assign n6720 = n2350 ^ n468 ^ n259 ;
  assign n6721 = ( n1340 & ~n2808 ) | ( n1340 & n4457 ) | ( ~n2808 & n4457 ) ;
  assign n6722 = n6721 ^ n989 ^ 1'b0 ;
  assign n6723 = n6720 & ~n6722 ;
  assign n6724 = ( n1898 & n3420 ) | ( n1898 & ~n6723 ) | ( n3420 & ~n6723 ) ;
  assign n6725 = n6724 ^ n2344 ^ 1'b0 ;
  assign n6726 = ~n6719 & n6725 ;
  assign n6727 = n1804 & n5514 ;
  assign n6728 = ~n907 & n6727 ;
  assign n6729 = ( n336 & n4523 ) | ( n336 & ~n6728 ) | ( n4523 & ~n6728 ) ;
  assign n6730 = n3028 & n6729 ;
  assign n6731 = ~n3995 & n6730 ;
  assign n6732 = n6731 ^ n2492 ^ 1'b0 ;
  assign n6733 = ( n593 & n1462 ) | ( n593 & ~n1716 ) | ( n1462 & ~n1716 ) ;
  assign n6734 = ( n1146 & n3192 ) | ( n1146 & ~n6733 ) | ( n3192 & ~n6733 ) ;
  assign n6735 = n3375 & n6734 ;
  assign n6736 = n5971 & n6735 ;
  assign n6737 = ~n2320 & n3088 ;
  assign n6738 = n1228 & ~n2812 ;
  assign n6739 = n6738 ^ n5733 ^ 1'b0 ;
  assign n6740 = ( ~n6366 & n6737 ) | ( ~n6366 & n6739 ) | ( n6737 & n6739 ) ;
  assign n6741 = ( n4858 & n5517 ) | ( n4858 & n6740 ) | ( n5517 & n6740 ) ;
  assign n6745 = ( n739 & n2984 ) | ( n739 & ~n3505 ) | ( n2984 & ~n3505 ) ;
  assign n6743 = ( x221 & n1561 ) | ( x221 & n2863 ) | ( n1561 & n2863 ) ;
  assign n6742 = n393 & n2567 ;
  assign n6744 = n6743 ^ n6742 ^ 1'b0 ;
  assign n6746 = n6745 ^ n6744 ^ n3092 ;
  assign n6747 = ( ~n3746 & n4631 ) | ( ~n3746 & n6746 ) | ( n4631 & n6746 ) ;
  assign n6748 = n6747 ^ n6549 ^ n693 ;
  assign n6752 = n2950 ^ n1719 ^ n1577 ;
  assign n6749 = n3047 ^ n1092 ^ 1'b0 ;
  assign n6750 = ( n884 & n2836 ) | ( n884 & n5067 ) | ( n2836 & n5067 ) ;
  assign n6751 = n6749 & n6750 ;
  assign n6753 = n6752 ^ n6751 ^ n4658 ;
  assign n6754 = n1496 ^ n640 ^ n382 ;
  assign n6755 = ( n1935 & n3152 ) | ( n1935 & ~n6754 ) | ( n3152 & ~n6754 ) ;
  assign n6756 = n2516 ^ n1030 ^ n558 ;
  assign n6757 = n6756 ^ n6696 ^ n6483 ;
  assign n6758 = ~n2058 & n6068 ;
  assign n6759 = n3124 & n6758 ;
  assign n6760 = n6759 ^ n2304 ^ n2244 ;
  assign n6761 = n6586 ^ n2783 ^ 1'b0 ;
  assign n6762 = n2381 & ~n6761 ;
  assign n6772 = ( ~x155 & n1416 ) | ( ~x155 & n1976 ) | ( n1416 & n1976 ) ;
  assign n6773 = n6772 ^ n1724 ^ 1'b0 ;
  assign n6769 = ~n3113 & n6712 ;
  assign n6763 = n5276 ^ n1374 ^ n551 ;
  assign n6764 = n2014 ^ n1804 ^ 1'b0 ;
  assign n6765 = n938 | n6764 ;
  assign n6766 = n2571 | n6765 ;
  assign n6767 = ( n3354 & n5044 ) | ( n3354 & ~n6766 ) | ( n5044 & ~n6766 ) ;
  assign n6768 = ~n6763 & n6767 ;
  assign n6770 = n6769 ^ n6768 ^ 1'b0 ;
  assign n6771 = n6770 ^ n5053 ^ 1'b0 ;
  assign n6774 = n6773 ^ n6771 ^ n4754 ;
  assign n6775 = n1665 ^ n888 ^ 1'b0 ;
  assign n6776 = ~n3679 & n6775 ;
  assign n6777 = ( n4785 & n6336 ) | ( n4785 & ~n6776 ) | ( n6336 & ~n6776 ) ;
  assign n6778 = n6777 ^ n2863 ^ 1'b0 ;
  assign n6779 = ( ~n410 & n3659 ) | ( ~n410 & n4562 ) | ( n3659 & n4562 ) ;
  assign n6780 = ( ~n339 & n908 ) | ( ~n339 & n6779 ) | ( n908 & n6779 ) ;
  assign n6781 = n3776 ^ n1909 ^ 1'b0 ;
  assign n6782 = n6781 ^ n6598 ^ n5551 ;
  assign n6783 = ~x218 & n2858 ;
  assign n6784 = ( ~n1904 & n5343 ) | ( ~n1904 & n6783 ) | ( n5343 & n6783 ) ;
  assign n6785 = n1106 & ~n6784 ;
  assign n6788 = n4557 ^ n1597 ^ 1'b0 ;
  assign n6786 = n3168 ^ n2509 ^ n1492 ;
  assign n6787 = n6786 ^ n6576 ^ n533 ;
  assign n6789 = n6788 ^ n6787 ^ n579 ;
  assign n6790 = n3918 ^ n2231 ^ n744 ;
  assign n6791 = x108 & n3841 ;
  assign n6792 = n6791 ^ n5306 ^ 1'b0 ;
  assign n6793 = n6792 ^ n4563 ^ n286 ;
  assign n6794 = ( ~n6789 & n6790 ) | ( ~n6789 & n6793 ) | ( n6790 & n6793 ) ;
  assign n6795 = n6766 ^ n2811 ^ n1618 ;
  assign n6796 = n6795 ^ n1776 ^ 1'b0 ;
  assign n6797 = ( ~n6785 & n6794 ) | ( ~n6785 & n6796 ) | ( n6794 & n6796 ) ;
  assign n6798 = ~n1961 & n4107 ;
  assign n6799 = n2312 & n6798 ;
  assign n6800 = n5722 & n6799 ;
  assign n6801 = ~n2779 & n4884 ;
  assign n6802 = n1002 ^ n929 ^ n927 ;
  assign n6803 = n6450 ^ n395 ^ 1'b0 ;
  assign n6804 = ( ~n6148 & n6507 ) | ( ~n6148 & n6803 ) | ( n6507 & n6803 ) ;
  assign n6805 = ( n826 & n964 ) | ( n826 & n1334 ) | ( n964 & n1334 ) ;
  assign n6806 = x218 & ~n6805 ;
  assign n6807 = n6806 ^ n4446 ^ 1'b0 ;
  assign n6808 = n6804 & ~n6807 ;
  assign n6809 = ~n6802 & n6808 ;
  assign n6810 = n6809 ^ n5670 ^ 1'b0 ;
  assign n6811 = n4023 ^ n2125 ^ n1707 ;
  assign n6812 = n6811 ^ n2220 ^ 1'b0 ;
  assign n6813 = ~n1075 & n6812 ;
  assign n6814 = ( n1612 & ~n2708 ) | ( n1612 & n6813 ) | ( ~n2708 & n6813 ) ;
  assign n6815 = n1796 ^ n1303 ^ x132 ;
  assign n6816 = n6815 ^ n4932 ^ 1'b0 ;
  assign n6818 = n3027 | n5017 ;
  assign n6819 = n1481 | n6818 ;
  assign n6817 = ~n3212 & n4306 ;
  assign n6820 = n6819 ^ n6817 ^ n373 ;
  assign n6836 = n6493 ^ n5842 ^ n4946 ;
  assign n6826 = n2994 ^ n1983 ^ 1'b0 ;
  assign n6827 = n5195 & n6826 ;
  assign n6828 = n739 ^ n621 ^ n296 ;
  assign n6829 = n6828 ^ n5472 ^ n594 ;
  assign n6830 = n4769 ^ n3743 ^ n2853 ;
  assign n6831 = n6830 ^ n1859 ^ n1345 ;
  assign n6832 = n6831 ^ n3568 ^ n3375 ;
  assign n6833 = n5800 & ~n6832 ;
  assign n6834 = ( ~n6827 & n6829 ) | ( ~n6827 & n6833 ) | ( n6829 & n6833 ) ;
  assign n6835 = n4200 & n6834 ;
  assign n6821 = ( n362 & n367 ) | ( n362 & ~n1967 ) | ( n367 & ~n1967 ) ;
  assign n6822 = ( n1582 & n4688 ) | ( n1582 & ~n6821 ) | ( n4688 & ~n6821 ) ;
  assign n6823 = n6822 ^ n1430 ^ 1'b0 ;
  assign n6824 = n1325 | n6823 ;
  assign n6825 = ( n1455 & n1760 ) | ( n1455 & n6824 ) | ( n1760 & n6824 ) ;
  assign n6837 = n6836 ^ n6835 ^ n6825 ;
  assign n6838 = ( ~n391 & n1132 ) | ( ~n391 & n2441 ) | ( n1132 & n2441 ) ;
  assign n6843 = ( n4109 & n5511 ) | ( n4109 & n6821 ) | ( n5511 & n6821 ) ;
  assign n6844 = n6843 ^ n4371 ^ n3801 ;
  assign n6841 = ( n583 & n694 ) | ( n583 & n1639 ) | ( n694 & n1639 ) ;
  assign n6840 = n4085 & n6776 ;
  assign n6842 = n6841 ^ n6840 ^ 1'b0 ;
  assign n6839 = ( n2838 & ~n3227 ) | ( n2838 & n3715 ) | ( ~n3227 & n3715 ) ;
  assign n6845 = n6844 ^ n6842 ^ n6839 ;
  assign n6846 = n6838 & n6845 ;
  assign n6848 = ( x22 & n418 ) | ( x22 & n1999 ) | ( n418 & n1999 ) ;
  assign n6847 = n2417 & ~n6672 ;
  assign n6849 = n6848 ^ n6847 ^ 1'b0 ;
  assign n6850 = n5187 & ~n6849 ;
  assign n6851 = ( ~n4414 & n5089 ) | ( ~n4414 & n6506 ) | ( n5089 & n6506 ) ;
  assign n6852 = n6553 ^ n5411 ^ n2527 ;
  assign n6853 = n6852 ^ n1994 ^ n1909 ;
  assign n6854 = n3961 ^ n2135 ^ 1'b0 ;
  assign n6855 = n6854 ^ n1467 ^ 1'b0 ;
  assign n6856 = n2783 ^ n380 ^ n330 ;
  assign n6857 = n6856 ^ n909 ^ n629 ;
  assign n6858 = n701 | n1183 ;
  assign n6859 = n6857 & n6858 ;
  assign n6860 = n6859 ^ n6313 ^ 1'b0 ;
  assign n6861 = n6860 ^ n3088 ^ x29 ;
  assign n6862 = n6861 ^ n1067 ^ x87 ;
  assign n6863 = ( n1164 & ~n3127 ) | ( n1164 & n5647 ) | ( ~n3127 & n5647 ) ;
  assign n6864 = n6863 ^ n1987 ^ n686 ;
  assign n6865 = ( n6855 & ~n6862 ) | ( n6855 & n6864 ) | ( ~n6862 & n6864 ) ;
  assign n6866 = n1128 & ~n3629 ;
  assign n6867 = n1134 ^ n860 ^ 1'b0 ;
  assign n6868 = n6866 & n6867 ;
  assign n6871 = x62 & x141 ;
  assign n6872 = n334 & n6871 ;
  assign n6873 = ( n734 & n1026 ) | ( n734 & ~n6872 ) | ( n1026 & ~n6872 ) ;
  assign n6874 = ( ~x202 & n2735 ) | ( ~x202 & n6873 ) | ( n2735 & n6873 ) ;
  assign n6875 = n2002 & ~n6874 ;
  assign n6876 = n6875 ^ n2965 ^ n1454 ;
  assign n6877 = n6876 ^ n1831 ^ 1'b0 ;
  assign n6878 = n3448 | n6877 ;
  assign n6879 = ( ~n1489 & n5641 ) | ( ~n1489 & n6878 ) | ( n5641 & n6878 ) ;
  assign n6880 = n6879 ^ n4684 ^ 1'b0 ;
  assign n6881 = ~n708 & n6880 ;
  assign n6869 = n395 & n1095 ;
  assign n6870 = n6869 ^ n4716 ^ n3163 ;
  assign n6882 = n6881 ^ n6870 ^ n1965 ;
  assign n6889 = n4914 ^ n4600 ^ 1'b0 ;
  assign n6890 = ~n2628 & n6889 ;
  assign n6891 = n6890 ^ n3082 ^ n1082 ;
  assign n6883 = ( n682 & ~n2253 ) | ( n682 & n3679 ) | ( ~n2253 & n3679 ) ;
  assign n6884 = n6883 ^ n5312 ^ n4338 ;
  assign n6885 = ( ~n353 & n6182 ) | ( ~n353 & n6802 ) | ( n6182 & n6802 ) ;
  assign n6886 = n6885 ^ n4610 ^ n2239 ;
  assign n6887 = n1199 & ~n6886 ;
  assign n6888 = ~n6884 & n6887 ;
  assign n6892 = n6891 ^ n6888 ^ n1266 ;
  assign n6893 = n4385 ^ n3448 ^ x134 ;
  assign n6894 = n2336 & ~n6652 ;
  assign n6895 = n6893 & n6894 ;
  assign n6909 = ( n1278 & ~n1818 ) | ( n1278 & n6540 ) | ( ~n1818 & n6540 ) ;
  assign n6910 = ( x199 & n6772 ) | ( x199 & n6909 ) | ( n6772 & n6909 ) ;
  assign n6896 = ( n832 & n966 ) | ( n832 & n3429 ) | ( n966 & n3429 ) ;
  assign n6903 = n4707 ^ n3120 ^ n2485 ;
  assign n6904 = ( ~n852 & n1682 ) | ( ~n852 & n2531 ) | ( n1682 & n2531 ) ;
  assign n6905 = ( n2777 & n6903 ) | ( n2777 & ~n6904 ) | ( n6903 & ~n6904 ) ;
  assign n6906 = ( n922 & ~n1103 ) | ( n922 & n6905 ) | ( ~n1103 & n6905 ) ;
  assign n6898 = n1427 & ~n2291 ;
  assign n6899 = n6898 ^ n3966 ^ n2048 ;
  assign n6900 = ( ~n3906 & n4173 ) | ( ~n3906 & n5619 ) | ( n4173 & n5619 ) ;
  assign n6901 = ( n2877 & n6899 ) | ( n2877 & ~n6900 ) | ( n6899 & ~n6900 ) ;
  assign n6902 = n6901 ^ n2510 ^ n368 ;
  assign n6897 = n5941 ^ n2255 ^ n1551 ;
  assign n6907 = n6906 ^ n6902 ^ n6897 ;
  assign n6908 = n6896 & ~n6907 ;
  assign n6911 = n6910 ^ n6908 ^ 1'b0 ;
  assign n6912 = n6617 ^ n1638 ^ n1627 ;
  assign n6913 = ( ~n3630 & n4294 ) | ( ~n3630 & n4687 ) | ( n4294 & n4687 ) ;
  assign n6914 = n6913 ^ n5539 ^ x22 ;
  assign n6917 = ~n1626 & n3635 ;
  assign n6918 = n1621 & ~n6917 ;
  assign n6919 = ~n4434 & n6918 ;
  assign n6915 = ~n347 & n1160 ;
  assign n6916 = ( ~n2345 & n5966 ) | ( ~n2345 & n6915 ) | ( n5966 & n6915 ) ;
  assign n6920 = n6919 ^ n6916 ^ n2979 ;
  assign n6921 = ~n4325 & n5640 ;
  assign n6922 = n519 & n6921 ;
  assign n6923 = n6922 ^ n1975 ^ n1122 ;
  assign n6924 = ~n3288 & n6923 ;
  assign n6925 = ~n5059 & n6924 ;
  assign n6929 = ~n3870 & n6432 ;
  assign n6926 = n3840 ^ n1073 ^ n623 ;
  assign n6927 = n3412 ^ n1877 ^ 1'b0 ;
  assign n6928 = n6926 & ~n6927 ;
  assign n6930 = n6929 ^ n6928 ^ n1539 ;
  assign n6931 = n6180 ^ n2557 ^ n1242 ;
  assign n6932 = n3807 & n6931 ;
  assign n6933 = ( n5442 & ~n5994 ) | ( n5442 & n6932 ) | ( ~n5994 & n6932 ) ;
  assign n6934 = ( n6741 & ~n6930 ) | ( n6741 & n6933 ) | ( ~n6930 & n6933 ) ;
  assign n6935 = ( ~x146 & n1580 ) | ( ~x146 & n3578 ) | ( n1580 & n3578 ) ;
  assign n6936 = ( ~n1676 & n4882 ) | ( ~n1676 & n6935 ) | ( n4882 & n6935 ) ;
  assign n6937 = n3954 ^ n2137 ^ n1435 ;
  assign n6938 = n6937 ^ n2883 ^ n1467 ;
  assign n6939 = ( n3065 & ~n5000 ) | ( n3065 & n6938 ) | ( ~n5000 & n6938 ) ;
  assign n6940 = n6939 ^ n5836 ^ 1'b0 ;
  assign n6941 = n6940 ^ n5890 ^ x152 ;
  assign n6942 = ( ~n1197 & n6936 ) | ( ~n1197 & n6941 ) | ( n6936 & n6941 ) ;
  assign n6943 = ( ~n692 & n1771 ) | ( ~n692 & n3205 ) | ( n1771 & n3205 ) ;
  assign n6944 = n1999 & ~n3041 ;
  assign n6945 = n3215 ^ n2511 ^ 1'b0 ;
  assign n6946 = ( n6943 & n6944 ) | ( n6943 & ~n6945 ) | ( n6944 & ~n6945 ) ;
  assign n6947 = n6946 ^ n3625 ^ 1'b0 ;
  assign n6949 = x21 & ~n2058 ;
  assign n6950 = n6949 ^ n615 ^ 1'b0 ;
  assign n6948 = ( n623 & n2431 ) | ( n623 & n6792 ) | ( n2431 & n6792 ) ;
  assign n6951 = n6950 ^ n6948 ^ n4774 ;
  assign n6952 = ( n3202 & ~n5438 ) | ( n3202 & n6951 ) | ( ~n5438 & n6951 ) ;
  assign n6953 = n6952 ^ n5365 ^ n3341 ;
  assign n6954 = ( ~n1440 & n6947 ) | ( ~n1440 & n6953 ) | ( n6947 & n6953 ) ;
  assign n6955 = n2112 ^ n883 ^ x158 ;
  assign n6956 = x238 & n6955 ;
  assign n6957 = n3488 & n6956 ;
  assign n6958 = ( ~n1284 & n1983 ) | ( ~n1284 & n2224 ) | ( n1983 & n2224 ) ;
  assign n6959 = ( n3241 & n6021 ) | ( n3241 & ~n6958 ) | ( n6021 & ~n6958 ) ;
  assign n6960 = n926 | n5134 ;
  assign n6961 = n6959 | n6960 ;
  assign n6962 = n700 & ~n1635 ;
  assign n6963 = n6962 ^ n4524 ^ 1'b0 ;
  assign n6969 = ( n343 & ~n2243 ) | ( n343 & n2510 ) | ( ~n2243 & n2510 ) ;
  assign n6967 = n2708 ^ n1734 ^ 1'b0 ;
  assign n6968 = x132 & ~n6967 ;
  assign n6970 = n6969 ^ n6968 ^ n2598 ;
  assign n6971 = n6970 ^ n2016 ^ 1'b0 ;
  assign n6966 = n6208 ^ n1509 ^ x212 ;
  assign n6972 = n6971 ^ n6966 ^ n6178 ;
  assign n6964 = n2984 ^ x239 ^ 1'b0 ;
  assign n6965 = n6964 ^ n3333 ^ n915 ;
  assign n6973 = n6972 ^ n6965 ^ n5427 ;
  assign n6974 = ( n4474 & n6963 ) | ( n4474 & n6973 ) | ( n6963 & n6973 ) ;
  assign n6975 = n2070 ^ n887 ^ n869 ;
  assign n6976 = n3042 & n4580 ;
  assign n6977 = n5502 & n6976 ;
  assign n6978 = n6975 | n6977 ;
  assign n6979 = n645 | n6978 ;
  assign n6980 = ( n4933 & ~n6102 ) | ( n4933 & n6979 ) | ( ~n6102 & n6979 ) ;
  assign n6981 = x112 & ~n3549 ;
  assign n6982 = n6981 ^ n3911 ^ n1120 ;
  assign n6986 = ( x75 & n1850 ) | ( x75 & ~n5593 ) | ( n1850 & ~n5593 ) ;
  assign n6983 = ( n1846 & n2418 ) | ( n1846 & n4612 ) | ( n2418 & n4612 ) ;
  assign n6984 = ( ~n1944 & n2407 ) | ( ~n1944 & n6983 ) | ( n2407 & n6983 ) ;
  assign n6985 = n2799 | n6984 ;
  assign n6987 = n6986 ^ n6985 ^ 1'b0 ;
  assign n6988 = n1953 ^ x147 ^ 1'b0 ;
  assign n6989 = ( n535 & n1356 ) | ( n535 & n4673 ) | ( n1356 & n4673 ) ;
  assign n6990 = n6989 ^ n3097 ^ 1'b0 ;
  assign n6991 = n5276 ^ n1547 ^ n1275 ;
  assign n6992 = n6991 ^ n722 ^ 1'b0 ;
  assign n6993 = n6409 | n6992 ;
  assign n6994 = n6993 ^ n4847 ^ 1'b0 ;
  assign n6995 = n5450 ^ n5088 ^ n3492 ;
  assign n6996 = ( n3480 & ~n6158 ) | ( n3480 & n6995 ) | ( ~n6158 & n6995 ) ;
  assign n6997 = n6994 & n6996 ;
  assign n6998 = ( n6988 & ~n6990 ) | ( n6988 & n6997 ) | ( ~n6990 & n6997 ) ;
  assign n6999 = n2038 ^ n1546 ^ 1'b0 ;
  assign n7000 = ( n3220 & n5394 ) | ( n3220 & n6999 ) | ( n5394 & n6999 ) ;
  assign n7001 = ( n6987 & n6998 ) | ( n6987 & n7000 ) | ( n6998 & n7000 ) ;
  assign n7004 = n1141 ^ n525 ^ 1'b0 ;
  assign n7002 = n4478 | n6765 ;
  assign n7003 = n7002 ^ n6597 ^ n580 ;
  assign n7005 = n7004 ^ n7003 ^ n3044 ;
  assign n7013 = ( n4128 & n4156 ) | ( n4128 & ~n5549 ) | ( n4156 & ~n5549 ) ;
  assign n7014 = ( n1996 & ~n6314 ) | ( n1996 & n7013 ) | ( ~n6314 & n7013 ) ;
  assign n7011 = n4596 ^ n294 ^ x136 ;
  assign n7012 = ( n889 & n6909 ) | ( n889 & n7011 ) | ( n6909 & n7011 ) ;
  assign n7006 = ( n3387 & n4981 ) | ( n3387 & ~n6213 ) | ( n4981 & ~n6213 ) ;
  assign n7007 = ( n1410 & n4659 ) | ( n1410 & n6649 ) | ( n4659 & n6649 ) ;
  assign n7008 = n7007 ^ n3780 ^ 1'b0 ;
  assign n7009 = ( n3007 & ~n7006 ) | ( n3007 & n7008 ) | ( ~n7006 & n7008 ) ;
  assign n7010 = ( n6249 & n6623 ) | ( n6249 & ~n7009 ) | ( n6623 & ~n7009 ) ;
  assign n7015 = n7014 ^ n7012 ^ n7010 ;
  assign n7016 = ( n488 & ~n1063 ) | ( n488 & n3521 ) | ( ~n1063 & n3521 ) ;
  assign n7023 = n2609 ^ n1143 ^ n490 ;
  assign n7022 = n1624 ^ n280 ^ x68 ;
  assign n7017 = ~n2900 & n3558 ;
  assign n7018 = n1893 & n7017 ;
  assign n7019 = n4701 ^ n1923 ^ x159 ;
  assign n7020 = n2090 & n5187 ;
  assign n7021 = ( n7018 & n7019 ) | ( n7018 & n7020 ) | ( n7019 & n7020 ) ;
  assign n7024 = n7023 ^ n7022 ^ n7021 ;
  assign n7025 = n887 ^ n871 ^ n446 ;
  assign n7026 = ( ~n2808 & n5640 ) | ( ~n2808 & n7025 ) | ( n5640 & n7025 ) ;
  assign n7027 = ( ~n3072 & n4738 ) | ( ~n3072 & n7026 ) | ( n4738 & n7026 ) ;
  assign n7028 = n1670 & n5385 ;
  assign n7029 = n1723 & n5281 ;
  assign n7030 = n2966 & ~n7029 ;
  assign n7031 = n272 & n784 ;
  assign n7032 = ~n3645 & n7031 ;
  assign n7033 = n1492 | n3614 ;
  assign n7034 = ( n1125 & n7032 ) | ( n1125 & ~n7033 ) | ( n7032 & ~n7033 ) ;
  assign n7035 = n5981 & n7034 ;
  assign n7036 = n7035 ^ n3459 ^ 1'b0 ;
  assign n7037 = n6552 ^ n682 ^ x152 ;
  assign n7038 = n2979 | n3066 ;
  assign n7039 = n5421 & ~n7038 ;
  assign n7040 = ( n256 & n7037 ) | ( n256 & ~n7039 ) | ( n7037 & ~n7039 ) ;
  assign n7041 = n7040 ^ n1863 ^ 1'b0 ;
  assign n7042 = n4557 ^ n1973 ^ n1303 ;
  assign n7043 = ( x152 & ~n4549 ) | ( x152 & n7042 ) | ( ~n4549 & n7042 ) ;
  assign n7044 = ( n3580 & n5603 ) | ( n3580 & n7043 ) | ( n5603 & n7043 ) ;
  assign n7045 = ( n3088 & n3772 ) | ( n3088 & n6780 ) | ( n3772 & n6780 ) ;
  assign n7047 = n2386 ^ n1682 ^ n1411 ;
  assign n7048 = ( n1609 & n1997 ) | ( n1609 & ~n7047 ) | ( n1997 & ~n7047 ) ;
  assign n7046 = n4618 ^ n3028 ^ n887 ;
  assign n7049 = n7048 ^ n7046 ^ n6706 ;
  assign n7050 = n1138 & ~n6144 ;
  assign n7051 = n7050 ^ n6031 ^ n2827 ;
  assign n7055 = n2292 ^ n1543 ^ 1'b0 ;
  assign n7053 = ( n3282 & n4599 ) | ( n3282 & ~n4771 ) | ( n4599 & ~n4771 ) ;
  assign n7054 = ( n824 & ~n5128 ) | ( n824 & n7053 ) | ( ~n5128 & n7053 ) ;
  assign n7052 = n1437 | n2339 ;
  assign n7056 = n7055 ^ n7054 ^ n7052 ;
  assign n7064 = n3516 ^ n3275 ^ n986 ;
  assign n7065 = n7064 ^ n5981 ^ n861 ;
  assign n7057 = ~n2317 & n6450 ;
  assign n7058 = ~x244 & n7057 ;
  assign n7059 = ~n897 & n1646 ;
  assign n7060 = n7059 ^ n3268 ^ n701 ;
  assign n7061 = ( x43 & ~n836 ) | ( x43 & n7060 ) | ( ~n836 & n7060 ) ;
  assign n7062 = n7061 ^ n4025 ^ n3037 ;
  assign n7063 = ( n4849 & n7058 ) | ( n4849 & n7062 ) | ( n7058 & n7062 ) ;
  assign n7066 = n7065 ^ n7063 ^ n3525 ;
  assign n7067 = n7066 ^ n3422 ^ n1654 ;
  assign n7071 = n5401 ^ n3213 ^ n1865 ;
  assign n7068 = n4087 & n7042 ;
  assign n7069 = n7068 ^ x110 ^ 1'b0 ;
  assign n7070 = n7069 ^ n6252 ^ n1499 ;
  assign n7072 = n7071 ^ n7070 ^ n5717 ;
  assign n7073 = ( ~n7056 & n7067 ) | ( ~n7056 & n7072 ) | ( n7067 & n7072 ) ;
  assign n7074 = ( ~n1715 & n2350 ) | ( ~n1715 & n6718 ) | ( n2350 & n6718 ) ;
  assign n7075 = ( n1781 & n2450 ) | ( n1781 & ~n6266 ) | ( n2450 & ~n6266 ) ;
  assign n7076 = ( x120 & n2554 ) | ( x120 & n2701 ) | ( n2554 & n2701 ) ;
  assign n7077 = n2700 & ~n2841 ;
  assign n7078 = n1751 & n7077 ;
  assign n7079 = ( n1104 & n1919 ) | ( n1104 & ~n3906 ) | ( n1919 & ~n3906 ) ;
  assign n7080 = ( n7076 & n7078 ) | ( n7076 & n7079 ) | ( n7078 & n7079 ) ;
  assign n7081 = ( ~n7074 & n7075 ) | ( ~n7074 & n7080 ) | ( n7075 & n7080 ) ;
  assign n7082 = n3848 ^ n1759 ^ n1499 ;
  assign n7083 = n7082 ^ n4539 ^ n766 ;
  assign n7084 = n1671 & n3638 ;
  assign n7085 = ( n447 & n804 ) | ( n447 & ~n2708 ) | ( n804 & ~n2708 ) ;
  assign n7086 = ( n749 & ~n2014 ) | ( n749 & n7085 ) | ( ~n2014 & n7085 ) ;
  assign n7087 = n1965 & n7086 ;
  assign n7088 = ~n2809 & n7087 ;
  assign n7089 = n7088 ^ n5725 ^ n2371 ;
  assign n7090 = ( n2810 & n7084 ) | ( n2810 & n7089 ) | ( n7084 & n7089 ) ;
  assign n7091 = ~n7083 & n7090 ;
  assign n7092 = n7091 ^ n1402 ^ 1'b0 ;
  assign n7093 = ( x126 & n2454 ) | ( x126 & ~n2752 ) | ( n2454 & ~n2752 ) ;
  assign n7094 = ( n850 & ~n1258 ) | ( n850 & n6493 ) | ( ~n1258 & n6493 ) ;
  assign n7095 = n7011 ^ n4288 ^ n2179 ;
  assign n7096 = ( n7093 & n7094 ) | ( n7093 & ~n7095 ) | ( n7094 & ~n7095 ) ;
  assign n7100 = n402 | n3927 ;
  assign n7101 = ( n431 & n1576 ) | ( n431 & n7100 ) | ( n1576 & n7100 ) ;
  assign n7099 = n2859 ^ x109 ^ 1'b0 ;
  assign n7102 = n7101 ^ n7099 ^ n569 ;
  assign n7098 = n2471 ^ n2459 ^ n539 ;
  assign n7097 = ( x237 & n2338 ) | ( x237 & ~n2945 ) | ( n2338 & ~n2945 ) ;
  assign n7103 = n7102 ^ n7098 ^ n7097 ;
  assign n7104 = ( n2896 & ~n3306 ) | ( n2896 & n4604 ) | ( ~n3306 & n4604 ) ;
  assign n7105 = n7104 ^ n5357 ^ 1'b0 ;
  assign n7106 = ( n2330 & n4119 ) | ( n2330 & ~n7105 ) | ( n4119 & ~n7105 ) ;
  assign n7107 = n2517 ^ n671 ^ n387 ;
  assign n7108 = n7107 ^ n914 ^ n773 ;
  assign n7113 = n2120 & ~n4003 ;
  assign n7114 = ~n2557 & n7113 ;
  assign n7115 = ( n1083 & ~n6282 ) | ( n1083 & n7114 ) | ( ~n6282 & n7114 ) ;
  assign n7109 = n5815 ^ n4761 ^ 1'b0 ;
  assign n7110 = n1174 ^ n413 ^ 1'b0 ;
  assign n7111 = n7110 ^ n6819 ^ n562 ;
  assign n7112 = ( ~n1618 & n7109 ) | ( ~n1618 & n7111 ) | ( n7109 & n7111 ) ;
  assign n7116 = n7115 ^ n7112 ^ n3350 ;
  assign n7117 = n3864 ^ n3445 ^ 1'b0 ;
  assign n7118 = ~n494 & n7117 ;
  assign n7119 = n7118 ^ n5087 ^ x74 ;
  assign n7120 = ( n2842 & ~n6829 ) | ( n2842 & n7119 ) | ( ~n6829 & n7119 ) ;
  assign n7121 = n3296 ^ n1431 ^ 1'b0 ;
  assign n7122 = n2341 ^ n707 ^ x119 ;
  assign n7123 = ~n3689 & n7122 ;
  assign n7124 = n7123 ^ n635 ^ 1'b0 ;
  assign n7125 = n4965 & ~n5101 ;
  assign n7126 = ~n7124 & n7125 ;
  assign n7132 = n5262 ^ n2750 ^ n2698 ;
  assign n7130 = n412 & n5040 ;
  assign n7131 = ( n491 & ~n5112 ) | ( n491 & n7130 ) | ( ~n5112 & n7130 ) ;
  assign n7128 = n2711 & ~n3224 ;
  assign n7127 = ~n522 & n6339 ;
  assign n7129 = n7128 ^ n7127 ^ 1'b0 ;
  assign n7133 = n7132 ^ n7131 ^ n7129 ;
  assign n7134 = n5732 ^ n3437 ^ 1'b0 ;
  assign n7135 = n6856 & n7134 ;
  assign n7145 = n5735 ^ n4721 ^ n502 ;
  assign n7146 = ( n3160 & ~n6446 ) | ( n3160 & n7145 ) | ( ~n6446 & n7145 ) ;
  assign n7136 = n6848 ^ n1493 ^ n535 ;
  assign n7137 = n3732 ^ n856 ^ x248 ;
  assign n7138 = n7137 ^ n1979 ^ 1'b0 ;
  assign n7139 = n543 | n7138 ;
  assign n7140 = n7139 ^ n4798 ^ n476 ;
  assign n7141 = n7140 ^ n4245 ^ n968 ;
  assign n7142 = n1028 & ~n7141 ;
  assign n7143 = n7142 ^ n4142 ^ 1'b0 ;
  assign n7144 = ( n6131 & ~n7136 ) | ( n6131 & n7143 ) | ( ~n7136 & n7143 ) ;
  assign n7147 = n7146 ^ n7144 ^ x130 ;
  assign n7148 = ( n3601 & n3680 ) | ( n3601 & ~n4892 ) | ( n3680 & ~n4892 ) ;
  assign n7159 = n3355 & n5728 ;
  assign n7160 = ~n5689 & n7159 ;
  assign n7161 = n7160 ^ n411 ^ 1'b0 ;
  assign n7155 = n1019 & ~n3490 ;
  assign n7156 = n7155 ^ n1454 ^ 1'b0 ;
  assign n7157 = n3463 ^ n2491 ^ n957 ;
  assign n7158 = ( ~n1864 & n7156 ) | ( ~n1864 & n7157 ) | ( n7156 & n7157 ) ;
  assign n7162 = n7161 ^ n7158 ^ n1726 ;
  assign n7149 = n6232 ^ x248 ^ 1'b0 ;
  assign n7150 = n1886 ^ n476 ^ 1'b0 ;
  assign n7151 = n2230 & n7150 ;
  assign n7152 = n7151 ^ n3390 ^ 1'b0 ;
  assign n7153 = ( n2183 & ~n7149 ) | ( n2183 & n7152 ) | ( ~n7149 & n7152 ) ;
  assign n7154 = n5801 & n7153 ;
  assign n7163 = n7162 ^ n7154 ^ 1'b0 ;
  assign n7166 = n2231 & n3543 ;
  assign n7167 = ( n1271 & n1272 ) | ( n1271 & n2535 ) | ( n1272 & n2535 ) ;
  assign n7168 = ( n5325 & n5831 ) | ( n5325 & n7167 ) | ( n5831 & n7167 ) ;
  assign n7169 = ( n1228 & n1238 ) | ( n1228 & ~n3777 ) | ( n1238 & ~n3777 ) ;
  assign n7170 = ( n2693 & n5529 ) | ( n2693 & n7169 ) | ( n5529 & n7169 ) ;
  assign n7171 = ( n7166 & n7168 ) | ( n7166 & n7170 ) | ( n7168 & n7170 ) ;
  assign n7164 = n5125 ^ n4347 ^ 1'b0 ;
  assign n7165 = n1356 & ~n7164 ;
  assign n7172 = n7171 ^ n7165 ^ n2728 ;
  assign n7173 = ~n6740 & n7172 ;
  assign n7174 = n7173 ^ n3625 ^ 1'b0 ;
  assign n7175 = n4843 ^ n3364 ^ n1207 ;
  assign n7176 = ( n895 & ~n2399 ) | ( n895 & n5088 ) | ( ~n2399 & n5088 ) ;
  assign n7177 = n2162 | n7176 ;
  assign n7178 = n1558 ^ n1191 ^ x240 ;
  assign n7179 = n2680 & n7178 ;
  assign n7180 = ( n7175 & n7177 ) | ( n7175 & ~n7179 ) | ( n7177 & ~n7179 ) ;
  assign n7188 = n432 & n3841 ;
  assign n7189 = n7188 ^ n4707 ^ 1'b0 ;
  assign n7190 = n7189 ^ n6491 ^ n4662 ;
  assign n7181 = n1621 & n2903 ;
  assign n7182 = n304 & n1168 ;
  assign n7183 = ( n2653 & ~n7181 ) | ( n2653 & n7182 ) | ( ~n7181 & n7182 ) ;
  assign n7184 = n4094 ^ n1438 ^ 1'b0 ;
  assign n7185 = n7183 & ~n7184 ;
  assign n7186 = n7185 ^ n1964 ^ 1'b0 ;
  assign n7187 = n2764 & ~n7186 ;
  assign n7191 = n7190 ^ n7187 ^ n846 ;
  assign n7199 = ( n999 & n1208 ) | ( n999 & n2426 ) | ( n1208 & n2426 ) ;
  assign n7194 = n6843 ^ n1266 ^ 1'b0 ;
  assign n7195 = ( n460 & n2257 ) | ( n460 & ~n7194 ) | ( n2257 & ~n7194 ) ;
  assign n7196 = n4212 ^ n3658 ^ n3448 ;
  assign n7197 = ( ~n5329 & n7195 ) | ( ~n5329 & n7196 ) | ( n7195 & n7196 ) ;
  assign n7198 = ~n2213 & n7197 ;
  assign n7192 = n3278 & n5772 ;
  assign n7193 = ( ~n6484 & n6943 ) | ( ~n6484 & n7192 ) | ( n6943 & n7192 ) ;
  assign n7200 = n7199 ^ n7198 ^ n7193 ;
  assign n7217 = n4991 | n5841 ;
  assign n7214 = ~n2192 & n3916 ;
  assign n7215 = n7214 ^ n3335 ^ 1'b0 ;
  assign n7201 = n326 & ~n3272 ;
  assign n7202 = n7201 ^ n1009 ^ 1'b0 ;
  assign n7208 = n1919 ^ n1380 ^ 1'b0 ;
  assign n7209 = n4692 & n7208 ;
  assign n7207 = n2883 ^ n2096 ^ x90 ;
  assign n7203 = ~n1269 & n2008 ;
  assign n7204 = n801 & n7203 ;
  assign n7205 = n7204 ^ n4626 ^ n3661 ;
  assign n7206 = ( n969 & n2493 ) | ( n969 & ~n7205 ) | ( n2493 & ~n7205 ) ;
  assign n7210 = n7209 ^ n7207 ^ n7206 ;
  assign n7211 = ( n5071 & n5424 ) | ( n5071 & ~n7210 ) | ( n5424 & ~n7210 ) ;
  assign n7212 = ( n1675 & n2042 ) | ( n1675 & ~n7211 ) | ( n2042 & ~n7211 ) ;
  assign n7213 = ( n2242 & ~n7202 ) | ( n2242 & n7212 ) | ( ~n7202 & n7212 ) ;
  assign n7216 = n7215 ^ n7213 ^ n3380 ;
  assign n7218 = n7217 ^ n7216 ^ n5845 ;
  assign n7230 = x1 & ~n6625 ;
  assign n7228 = n3733 ^ n2622 ^ 1'b0 ;
  assign n7229 = n2126 & ~n7228 ;
  assign n7227 = n2936 ^ n2103 ^ x217 ;
  assign n7231 = n7230 ^ n7229 ^ n7227 ;
  assign n7232 = n7231 ^ x100 ^ 1'b0 ;
  assign n7223 = x159 & n5754 ;
  assign n7224 = n7223 ^ n2966 ^ 1'b0 ;
  assign n7225 = ( n1787 & ~n6857 ) | ( n1787 & n7224 ) | ( ~n6857 & n7224 ) ;
  assign n7219 = n3576 ^ n1425 ^ 1'b0 ;
  assign n7220 = ~n1550 & n7219 ;
  assign n7221 = n7220 ^ n3794 ^ n1305 ;
  assign n7222 = ( ~n3997 & n5885 ) | ( ~n3997 & n7221 ) | ( n5885 & n7221 ) ;
  assign n7226 = n7225 ^ n7222 ^ n1535 ;
  assign n7233 = n7232 ^ n7226 ^ 1'b0 ;
  assign n7239 = n1363 & n5528 ;
  assign n7240 = ~n2752 & n7239 ;
  assign n7241 = n7240 ^ n6959 ^ n5094 ;
  assign n7234 = n577 & ~n3069 ;
  assign n7235 = n964 & n7234 ;
  assign n7236 = ( ~n3066 & n3394 ) | ( ~n3066 & n7235 ) | ( n3394 & n7235 ) ;
  assign n7237 = ( n1365 & n1864 ) | ( n1365 & ~n4015 ) | ( n1864 & ~n4015 ) ;
  assign n7238 = ( ~n2928 & n7236 ) | ( ~n2928 & n7237 ) | ( n7236 & n7237 ) ;
  assign n7242 = n7241 ^ n7238 ^ n4713 ;
  assign n7251 = n6872 ^ n5380 ^ n2276 ;
  assign n7246 = n2385 ^ n2291 ^ 1'b0 ;
  assign n7247 = n599 & ~n2278 ;
  assign n7248 = n1655 & n7247 ;
  assign n7249 = n7248 ^ x7 ^ 1'b0 ;
  assign n7250 = ( n6739 & ~n7246 ) | ( n6739 & n7249 ) | ( ~n7246 & n7249 ) ;
  assign n7244 = n2827 ^ n1071 ^ 1'b0 ;
  assign n7243 = n3067 & ~n4403 ;
  assign n7245 = n7244 ^ n7243 ^ 1'b0 ;
  assign n7252 = n7251 ^ n7250 ^ n7245 ;
  assign n7253 = n6802 ^ n3769 ^ x38 ;
  assign n7254 = n2196 ^ n1963 ^ 1'b0 ;
  assign n7255 = ~n256 & n7254 ;
  assign n7256 = n5986 & n7255 ;
  assign n7257 = ( n5791 & n7253 ) | ( n5791 & ~n7256 ) | ( n7253 & ~n7256 ) ;
  assign n7259 = ( n1224 & ~n2035 ) | ( n1224 & n2310 ) | ( ~n2035 & n2310 ) ;
  assign n7260 = n7259 ^ n5905 ^ n866 ;
  assign n7261 = n4352 & n7260 ;
  assign n7262 = n5869 & n7261 ;
  assign n7258 = n5166 ^ n1610 ^ x25 ;
  assign n7263 = n7262 ^ n7258 ^ n6765 ;
  assign n7264 = n311 & ~n2412 ;
  assign n7265 = ~n6813 & n7264 ;
  assign n7266 = n4409 ^ n876 ^ n256 ;
  assign n7267 = ~n3075 & n7266 ;
  assign n7268 = n7267 ^ n1328 ^ 1'b0 ;
  assign n7269 = n7268 ^ n4737 ^ n748 ;
  assign n7270 = n3111 & n6068 ;
  assign n7271 = ~n1083 & n7270 ;
  assign n7272 = n7271 ^ n7204 ^ n4311 ;
  assign n7273 = ( n551 & ~n2455 ) | ( n551 & n2782 ) | ( ~n2455 & n2782 ) ;
  assign n7274 = n5849 | n7059 ;
  assign n7275 = ( ~n528 & n7273 ) | ( ~n528 & n7274 ) | ( n7273 & n7274 ) ;
  assign n7276 = ( ~n1627 & n2879 ) | ( ~n1627 & n7275 ) | ( n2879 & n7275 ) ;
  assign n7293 = ( n1041 & ~n3514 ) | ( n1041 & n5843 ) | ( ~n3514 & n5843 ) ;
  assign n7294 = n7293 ^ n3779 ^ n1293 ;
  assign n7288 = x46 & ~n957 ;
  assign n7289 = n7288 ^ n1704 ^ 1'b0 ;
  assign n7290 = ( n623 & n1233 ) | ( n623 & n7289 ) | ( n1233 & n7289 ) ;
  assign n7287 = ( n916 & n3479 ) | ( n916 & ~n6408 ) | ( n3479 & ~n6408 ) ;
  assign n7291 = n7290 ^ n7287 ^ 1'b0 ;
  assign n7292 = ~n2331 & n7291 ;
  assign n7281 = n2157 ^ n1489 ^ 1'b0 ;
  assign n7282 = n2439 ^ n1976 ^ n1882 ;
  assign n7283 = ( ~n1812 & n7281 ) | ( ~n1812 & n7282 ) | ( n7281 & n7282 ) ;
  assign n7284 = ( ~n891 & n5281 ) | ( ~n891 & n7283 ) | ( n5281 & n7283 ) ;
  assign n7285 = n7284 ^ n4088 ^ n3206 ;
  assign n7277 = n410 & n442 ;
  assign n7278 = n949 & ~n7277 ;
  assign n7279 = n7278 ^ n6433 ^ 1'b0 ;
  assign n7280 = ( ~n2557 & n5353 ) | ( ~n2557 & n7279 ) | ( n5353 & n7279 ) ;
  assign n7286 = n7285 ^ n7280 ^ n391 ;
  assign n7295 = n7294 ^ n7292 ^ n7286 ;
  assign n7296 = n2006 | n4531 ;
  assign n7297 = n7296 ^ n2406 ^ 1'b0 ;
  assign n7298 = n2027 ^ n1891 ^ x53 ;
  assign n7299 = n3027 ^ n1889 ^ n839 ;
  assign n7300 = ( n262 & ~n2103 ) | ( n262 & n7299 ) | ( ~n2103 & n7299 ) ;
  assign n7301 = n2115 & n2176 ;
  assign n7302 = ( n4389 & n7300 ) | ( n4389 & ~n7301 ) | ( n7300 & ~n7301 ) ;
  assign n7303 = ( n7297 & n7298 ) | ( n7297 & n7302 ) | ( n7298 & n7302 ) ;
  assign n7304 = ( ~n1568 & n6805 ) | ( ~n1568 & n7303 ) | ( n6805 & n7303 ) ;
  assign n7305 = n7304 ^ x178 ^ 1'b0 ;
  assign n7306 = ~n1834 & n7305 ;
  assign n7307 = n6994 & n7306 ;
  assign n7308 = n7307 ^ n4989 ^ 1'b0 ;
  assign n7309 = n6821 | n7308 ;
  assign n7310 = ( n486 & n2832 ) | ( n486 & ~n7309 ) | ( n2832 & ~n7309 ) ;
  assign n7311 = n7295 & ~n7310 ;
  assign n7312 = ~n2478 & n7311 ;
  assign n7313 = ( ~n413 & n3629 ) | ( ~n413 & n5389 ) | ( n3629 & n5389 ) ;
  assign n7317 = n5662 ^ n2608 ^ n1928 ;
  assign n7314 = n2903 ^ n1530 ^ n972 ;
  assign n7315 = n7314 ^ n3468 ^ 1'b0 ;
  assign n7316 = n7315 ^ n2636 ^ n2511 ;
  assign n7318 = n7317 ^ n7316 ^ 1'b0 ;
  assign n7319 = ~n4191 & n7318 ;
  assign n7320 = n7319 ^ n1042 ^ n413 ;
  assign n7321 = ( n4406 & ~n7313 ) | ( n4406 & n7320 ) | ( ~n7313 & n7320 ) ;
  assign n7325 = ( n1190 & ~n2633 ) | ( n1190 & n2716 ) | ( ~n2633 & n2716 ) ;
  assign n7322 = n5448 ^ n2936 ^ x147 ;
  assign n7323 = ( n4531 & n4679 ) | ( n4531 & n6299 ) | ( n4679 & n6299 ) ;
  assign n7324 = n7322 & n7323 ;
  assign n7326 = n7325 ^ n7324 ^ n3172 ;
  assign n7328 = n2527 ^ x104 ^ 1'b0 ;
  assign n7329 = n2174 & n7328 ;
  assign n7330 = n7329 ^ n579 ^ x191 ;
  assign n7331 = ( n3301 & n3838 ) | ( n3301 & ~n7330 ) | ( n3838 & ~n7330 ) ;
  assign n7327 = n706 & n5462 ;
  assign n7332 = n7331 ^ n7327 ^ n5905 ;
  assign n7333 = n2750 ^ n1984 ^ n1042 ;
  assign n7334 = ( ~n277 & n1296 ) | ( ~n277 & n3605 ) | ( n1296 & n3605 ) ;
  assign n7335 = ( ~n3701 & n4158 ) | ( ~n3701 & n7334 ) | ( n4158 & n7334 ) ;
  assign n7336 = n4049 ^ n3247 ^ 1'b0 ;
  assign n7337 = ~n7335 & n7336 ;
  assign n7338 = ( x34 & n2747 ) | ( x34 & n7337 ) | ( n2747 & n7337 ) ;
  assign n7339 = ( ~n1441 & n7333 ) | ( ~n1441 & n7338 ) | ( n7333 & n7338 ) ;
  assign n7340 = n4768 ^ n1849 ^ x231 ;
  assign n7341 = ( n4446 & n5998 ) | ( n4446 & n7340 ) | ( n5998 & n7340 ) ;
  assign n7342 = n4720 ^ n4603 ^ 1'b0 ;
  assign n7343 = n7342 ^ n7020 ^ n5030 ;
  assign n7344 = ( ~n280 & n7341 ) | ( ~n280 & n7343 ) | ( n7341 & n7343 ) ;
  assign n7345 = ( n3774 & n5147 ) | ( n3774 & n7344 ) | ( n5147 & n7344 ) ;
  assign n7346 = ( n1954 & n2616 ) | ( n1954 & n3311 ) | ( n2616 & n3311 ) ;
  assign n7347 = n7346 ^ n2500 ^ n1212 ;
  assign n7352 = n744 & ~n2081 ;
  assign n7351 = n7169 ^ n3289 ^ n1280 ;
  assign n7353 = n7352 ^ n7351 ^ n4042 ;
  assign n7354 = ( ~n1004 & n5391 ) | ( ~n1004 & n7353 ) | ( n5391 & n7353 ) ;
  assign n7348 = n5076 ^ n5041 ^ n549 ;
  assign n7349 = n4829 ^ n988 ^ 1'b0 ;
  assign n7350 = ( n3018 & ~n7348 ) | ( n3018 & n7349 ) | ( ~n7348 & n7349 ) ;
  assign n7355 = n7354 ^ n7350 ^ n2376 ;
  assign n7356 = n621 | n7355 ;
  assign n7357 = n5157 | n7356 ;
  assign n7359 = ~n1447 & n3887 ;
  assign n7358 = n1431 ^ n1095 ^ x193 ;
  assign n7360 = n7359 ^ n7358 ^ n425 ;
  assign n7361 = ( ~n1700 & n2820 ) | ( ~n1700 & n6684 ) | ( n2820 & n6684 ) ;
  assign n7362 = n7361 ^ n7273 ^ n6786 ;
  assign n7363 = n5526 ^ n1380 ^ n753 ;
  assign n7364 = n1297 & ~n5115 ;
  assign n7365 = ~n7363 & n7364 ;
  assign n7366 = n7362 & n7365 ;
  assign n7369 = ~n760 & n2213 ;
  assign n7370 = n916 & n7369 ;
  assign n7371 = ( n539 & n862 ) | ( n539 & n4509 ) | ( n862 & n4509 ) ;
  assign n7372 = n7371 ^ n2298 ^ 1'b0 ;
  assign n7373 = ~n7370 & n7372 ;
  assign n7367 = ( ~n2046 & n3191 ) | ( ~n2046 & n3407 ) | ( n3191 & n3407 ) ;
  assign n7368 = ( ~n1113 & n3336 ) | ( ~n1113 & n7367 ) | ( n3336 & n7367 ) ;
  assign n7374 = n7373 ^ n7368 ^ 1'b0 ;
  assign n7375 = x166 & x202 ;
  assign n7376 = ~n1573 & n7375 ;
  assign n7377 = ( n1308 & n4049 ) | ( n1308 & ~n6743 ) | ( n4049 & ~n6743 ) ;
  assign n7378 = n5993 ^ n5147 ^ n3123 ;
  assign n7379 = ( ~n1339 & n4310 ) | ( ~n1339 & n7378 ) | ( n4310 & n7378 ) ;
  assign n7380 = ( ~n7376 & n7377 ) | ( ~n7376 & n7379 ) | ( n7377 & n7379 ) ;
  assign n7381 = ( n1598 & ~n4280 ) | ( n1598 & n7380 ) | ( ~n4280 & n7380 ) ;
  assign n7389 = ( n1276 & n2598 ) | ( n1276 & n3397 ) | ( n2598 & n3397 ) ;
  assign n7390 = n7389 ^ n6224 ^ n442 ;
  assign n7387 = n2010 ^ n1215 ^ 1'b0 ;
  assign n7386 = n3194 ^ n1006 ^ n423 ;
  assign n7382 = ( n2188 & n3574 ) | ( n2188 & n7287 ) | ( n3574 & n7287 ) ;
  assign n7383 = n4572 ^ n866 ^ 1'b0 ;
  assign n7384 = n7383 ^ n3211 ^ n2003 ;
  assign n7385 = ( n1646 & n7382 ) | ( n1646 & ~n7384 ) | ( n7382 & ~n7384 ) ;
  assign n7388 = n7387 ^ n7386 ^ n7385 ;
  assign n7391 = n7390 ^ n7388 ^ n4399 ;
  assign n7396 = ( n801 & ~n3625 ) | ( n801 & n4126 ) | ( ~n3625 & n4126 ) ;
  assign n7393 = n3706 ^ n1710 ^ n478 ;
  assign n7392 = ( n1129 & n5264 ) | ( n1129 & ~n6968 ) | ( n5264 & ~n6968 ) ;
  assign n7394 = n7393 ^ n7392 ^ n2871 ;
  assign n7395 = n7394 ^ n2789 ^ n2636 ;
  assign n7397 = n7396 ^ n7395 ^ x28 ;
  assign n7398 = n5217 ^ n2923 ^ x36 ;
  assign n7399 = n5034 ^ n365 ^ x100 ;
  assign n7400 = n5938 & ~n7399 ;
  assign n7401 = n7400 ^ n5900 ^ 1'b0 ;
  assign n7402 = ( x203 & n932 ) | ( x203 & n4005 ) | ( n932 & n4005 ) ;
  assign n7404 = n4101 ^ n1894 ^ n1872 ;
  assign n7405 = n7404 ^ n3455 ^ n2276 ;
  assign n7403 = n6939 ^ n6143 ^ 1'b0 ;
  assign n7406 = n7405 ^ n7403 ^ n2471 ;
  assign n7407 = n7406 ^ n1243 ^ 1'b0 ;
  assign n7408 = ~n7402 & n7407 ;
  assign n7409 = ( n6733 & ~n7401 ) | ( n6733 & n7408 ) | ( ~n7401 & n7408 ) ;
  assign n7410 = ( ~n498 & n1225 ) | ( ~n498 & n1435 ) | ( n1225 & n1435 ) ;
  assign n7411 = n1091 | n5445 ;
  assign n7412 = ( n1340 & ~n1678 ) | ( n1340 & n7411 ) | ( ~n1678 & n7411 ) ;
  assign n7413 = ( n3040 & ~n7410 ) | ( n3040 & n7412 ) | ( ~n7410 & n7412 ) ;
  assign n7414 = n4787 ^ n477 ^ 1'b0 ;
  assign n7415 = n5901 ^ n4882 ^ n576 ;
  assign n7416 = n5204 | n7415 ;
  assign n7417 = n7416 ^ n4538 ^ 1'b0 ;
  assign n7418 = n7417 ^ n3989 ^ n477 ;
  assign n7419 = n7414 & ~n7418 ;
  assign n7420 = ( ~n4159 & n5811 ) | ( ~n4159 & n7419 ) | ( n5811 & n7419 ) ;
  assign n7421 = n1816 & ~n3960 ;
  assign n7422 = n7421 ^ n2585 ^ 1'b0 ;
  assign n7423 = n7422 ^ n5788 ^ n4606 ;
  assign n7424 = n4040 ^ n3570 ^ n3388 ;
  assign n7425 = n7424 ^ n3132 ^ 1'b0 ;
  assign n7426 = n3002 | n7425 ;
  assign n7427 = ( n4280 & n6674 ) | ( n4280 & n7426 ) | ( n6674 & n7426 ) ;
  assign n7428 = n3975 & n7427 ;
  assign n7429 = n5007 & n7428 ;
  assign n7430 = n2342 ^ n1476 ^ x148 ;
  assign n7431 = ( ~n2218 & n3795 ) | ( ~n2218 & n7430 ) | ( n3795 & n7430 ) ;
  assign n7432 = n1924 ^ n764 ^ 1'b0 ;
  assign n7433 = ( n3162 & ~n6543 ) | ( n3162 & n7432 ) | ( ~n6543 & n7432 ) ;
  assign n7434 = n7433 ^ n6391 ^ n2476 ;
  assign n7435 = ( ~n5663 & n7431 ) | ( ~n5663 & n7434 ) | ( n7431 & n7434 ) ;
  assign n7444 = n1149 ^ n934 ^ n442 ;
  assign n7442 = n4924 ^ n1789 ^ x189 ;
  assign n7443 = n7442 ^ n3300 ^ 1'b0 ;
  assign n7445 = n7444 ^ n7443 ^ n2450 ;
  assign n7446 = n7445 ^ n5935 ^ n3320 ;
  assign n7447 = n7446 ^ n5168 ^ 1'b0 ;
  assign n7436 = ( x75 & n2839 ) | ( x75 & n5582 ) | ( n2839 & n5582 ) ;
  assign n7437 = ( n577 & n4644 ) | ( n577 & ~n5676 ) | ( n4644 & ~n5676 ) ;
  assign n7438 = n7437 ^ n6144 ^ n3142 ;
  assign n7439 = ( ~n6675 & n7436 ) | ( ~n6675 & n7438 ) | ( n7436 & n7438 ) ;
  assign n7440 = ( n1405 & n3002 ) | ( n1405 & n7439 ) | ( n3002 & n7439 ) ;
  assign n7441 = n2840 & ~n7440 ;
  assign n7448 = n7447 ^ n7441 ^ 1'b0 ;
  assign n7449 = ( n824 & ~n5748 ) | ( n824 & n7440 ) | ( ~n5748 & n7440 ) ;
  assign n7450 = n779 | n5859 ;
  assign n7451 = ( ~n1804 & n4700 ) | ( ~n1804 & n7450 ) | ( n4700 & n7450 ) ;
  assign n7452 = n7451 ^ n6868 ^ n2111 ;
  assign n7453 = n5425 ^ n1776 ^ n861 ;
  assign n7464 = ( n826 & ~n3836 ) | ( n826 & n4665 ) | ( ~n3836 & n4665 ) ;
  assign n7462 = n744 & ~n5373 ;
  assign n7463 = ( n851 & n4509 ) | ( n851 & n7462 ) | ( n4509 & n7462 ) ;
  assign n7454 = n6612 ^ n5236 ^ 1'b0 ;
  assign n7456 = ( n3029 & n3205 ) | ( n3029 & ~n4603 ) | ( n3205 & ~n4603 ) ;
  assign n7455 = ( n2512 & ~n2600 ) | ( n2512 & n6536 ) | ( ~n2600 & n6536 ) ;
  assign n7457 = n7456 ^ n7455 ^ n6830 ;
  assign n7458 = ( n5537 & n7454 ) | ( n5537 & n7457 ) | ( n7454 & n7457 ) ;
  assign n7459 = n2762 & n2905 ;
  assign n7460 = n472 & ~n7459 ;
  assign n7461 = n7458 & n7460 ;
  assign n7465 = n7464 ^ n7463 ^ n7461 ;
  assign n7466 = n7465 ^ n4183 ^ n2838 ;
  assign n7467 = n2275 ^ n1102 ^ n612 ;
  assign n7468 = n4422 ^ n2372 ^ n760 ;
  assign n7469 = ( n2919 & n4162 ) | ( n2919 & n7468 ) | ( n4162 & n7468 ) ;
  assign n7470 = ( n2732 & n7467 ) | ( n2732 & ~n7469 ) | ( n7467 & ~n7469 ) ;
  assign n7471 = n4298 ^ n1815 ^ 1'b0 ;
  assign n7472 = n7471 ^ n3431 ^ 1'b0 ;
  assign n7473 = n1869 & n7472 ;
  assign n7474 = ( n3037 & n3522 ) | ( n3037 & n7473 ) | ( n3522 & n7473 ) ;
  assign n7478 = n4882 ^ n2272 ^ 1'b0 ;
  assign n7475 = n2766 & ~n4523 ;
  assign n7476 = n7475 ^ n5819 ^ 1'b0 ;
  assign n7477 = ( n2343 & n6017 ) | ( n2343 & ~n7476 ) | ( n6017 & ~n7476 ) ;
  assign n7479 = n7478 ^ n7477 ^ n4982 ;
  assign n7480 = ~n256 & n7479 ;
  assign n7481 = ~n7474 & n7480 ;
  assign n7482 = n4580 ^ n1430 ^ n1030 ;
  assign n7483 = ( n1482 & n1919 ) | ( n1482 & n7482 ) | ( n1919 & n7482 ) ;
  assign n7484 = ( ~n4425 & n4698 ) | ( ~n4425 & n5441 ) | ( n4698 & n5441 ) ;
  assign n7485 = ( n2091 & ~n2289 ) | ( n2091 & n3743 ) | ( ~n2289 & n3743 ) ;
  assign n7486 = n3470 & n7485 ;
  assign n7487 = n7486 ^ n4233 ^ 1'b0 ;
  assign n7488 = ( n6196 & n7484 ) | ( n6196 & n7487 ) | ( n7484 & n7487 ) ;
  assign n7489 = ( n883 & n936 ) | ( n883 & n1806 ) | ( n936 & n1806 ) ;
  assign n7490 = ( ~n715 & n6479 ) | ( ~n715 & n7489 ) | ( n6479 & n7489 ) ;
  assign n7491 = n7490 ^ n7194 ^ n3613 ;
  assign n7492 = n7491 ^ n1355 ^ n1029 ;
  assign n7493 = n7492 ^ n6237 ^ n2844 ;
  assign n7494 = ( n3341 & n7343 ) | ( n3341 & ~n7493 ) | ( n7343 & ~n7493 ) ;
  assign n7495 = ( n973 & n2667 ) | ( n973 & ~n7494 ) | ( n2667 & ~n7494 ) ;
  assign n7496 = ( n7483 & ~n7488 ) | ( n7483 & n7495 ) | ( ~n7488 & n7495 ) ;
  assign n7497 = ( n783 & n2733 ) | ( n783 & n5950 ) | ( n2733 & n5950 ) ;
  assign n7498 = n3689 ^ n1477 ^ 1'b0 ;
  assign n7499 = n3857 | n7498 ;
  assign n7500 = n7499 ^ n2865 ^ 1'b0 ;
  assign n7501 = ~n7497 & n7500 ;
  assign n7502 = ( n2977 & n3464 ) | ( n2977 & n6049 ) | ( n3464 & n6049 ) ;
  assign n7503 = ( ~n1402 & n2555 ) | ( ~n1402 & n4414 ) | ( n2555 & n4414 ) ;
  assign n7504 = n7503 ^ n4156 ^ x74 ;
  assign n7505 = ( n518 & n2091 ) | ( n518 & n3073 ) | ( n2091 & n3073 ) ;
  assign n7506 = ~n2850 & n3086 ;
  assign n7507 = ~n1217 & n7506 ;
  assign n7508 = n2845 ^ x240 ^ 1'b0 ;
  assign n7509 = n7507 | n7508 ;
  assign n7510 = n7505 | n7509 ;
  assign n7511 = n5179 ^ n3168 ^ n1356 ;
  assign n7512 = ( x127 & n778 ) | ( x127 & ~n7511 ) | ( n778 & ~n7511 ) ;
  assign n7513 = n2458 ^ n303 ^ 1'b0 ;
  assign n7514 = ( n2435 & n7512 ) | ( n2435 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7523 = n1819 & ~n5382 ;
  assign n7524 = n5010 & ~n7523 ;
  assign n7525 = ~n6603 & n7524 ;
  assign n7515 = n4537 ^ n3669 ^ n1625 ;
  assign n7516 = ( n509 & ~n5178 ) | ( n509 & n7515 ) | ( ~n5178 & n7515 ) ;
  assign n7517 = ( n503 & n963 ) | ( n503 & ~n2604 ) | ( n963 & ~n2604 ) ;
  assign n7518 = n7517 ^ n4173 ^ n372 ;
  assign n7519 = ( n5184 & ~n7516 ) | ( n5184 & n7518 ) | ( ~n7516 & n7518 ) ;
  assign n7520 = n7519 ^ n430 ^ 1'b0 ;
  assign n7521 = ~n4091 & n7520 ;
  assign n7522 = ( n3028 & n5234 ) | ( n3028 & n7521 ) | ( n5234 & n7521 ) ;
  assign n7526 = n7525 ^ n7522 ^ 1'b0 ;
  assign n7527 = ( n1374 & ~n5338 ) | ( n1374 & n7526 ) | ( ~n5338 & n7526 ) ;
  assign n7528 = n7514 & n7527 ;
  assign n7529 = n7510 & n7528 ;
  assign n7530 = ( n4213 & ~n7504 ) | ( n4213 & n7529 ) | ( ~n7504 & n7529 ) ;
  assign n7531 = ( n3471 & n7502 ) | ( n3471 & n7530 ) | ( n7502 & n7530 ) ;
  assign n7532 = n3996 ^ n1041 ^ x178 ;
  assign n7533 = n923 | n1448 ;
  assign n7534 = n1937 & ~n7533 ;
  assign n7535 = n7534 ^ n3750 ^ 1'b0 ;
  assign n7536 = ( n1475 & ~n7532 ) | ( n1475 & n7535 ) | ( ~n7532 & n7535 ) ;
  assign n7537 = n7536 ^ n6074 ^ n3132 ;
  assign n7540 = n5082 ^ n2524 ^ n1863 ;
  assign n7541 = n5828 ^ n3770 ^ 1'b0 ;
  assign n7542 = n3618 & n7541 ;
  assign n7543 = n855 | n3172 ;
  assign n7544 = n7542 | n7543 ;
  assign n7545 = ( ~n5365 & n6223 ) | ( ~n5365 & n7544 ) | ( n6223 & n7544 ) ;
  assign n7546 = ( ~n3756 & n7540 ) | ( ~n3756 & n7545 ) | ( n7540 & n7545 ) ;
  assign n7538 = n4608 ^ n3606 ^ n1272 ;
  assign n7539 = n7538 ^ n4311 ^ n1638 ;
  assign n7547 = n7546 ^ n7539 ^ n2950 ;
  assign n7548 = n5284 ^ n3929 ^ x90 ;
  assign n7549 = n7548 ^ n7220 ^ n6577 ;
  assign n7550 = ( n3455 & ~n4010 ) | ( n3455 & n7549 ) | ( ~n4010 & n7549 ) ;
  assign n7551 = n7550 ^ n956 ^ x0 ;
  assign n7552 = ~n531 & n3248 ;
  assign n7553 = n7552 ^ n7425 ^ 1'b0 ;
  assign n7554 = n6483 ^ n3210 ^ 1'b0 ;
  assign n7555 = ( x1 & n2841 ) | ( x1 & n4707 ) | ( n2841 & n4707 ) ;
  assign n7556 = ( x0 & n3629 ) | ( x0 & ~n7555 ) | ( n3629 & ~n7555 ) ;
  assign n7557 = n7556 ^ n3799 ^ n2789 ;
  assign n7558 = x209 & ~n7557 ;
  assign n7559 = n7554 & n7558 ;
  assign n7560 = n7559 ^ n1555 ^ x234 ;
  assign n7561 = ( n6593 & ~n7553 ) | ( n6593 & n7560 ) | ( ~n7553 & n7560 ) ;
  assign n7562 = n6380 ^ n2336 ^ n2297 ;
  assign n7563 = ( n2219 & n7023 ) | ( n2219 & ~n7562 ) | ( n7023 & ~n7562 ) ;
  assign n7564 = ( n1765 & ~n5401 ) | ( n1765 & n7563 ) | ( ~n5401 & n7563 ) ;
  assign n7565 = n7564 ^ n3290 ^ 1'b0 ;
  assign n7566 = n1183 & n2473 ;
  assign n7567 = ~n4744 & n7566 ;
  assign n7568 = ( n1955 & n5745 ) | ( n1955 & n7567 ) | ( n5745 & n7567 ) ;
  assign n7569 = n7568 ^ n4195 ^ n1748 ;
  assign n7570 = ( n992 & ~n2692 ) | ( n992 & n4544 ) | ( ~n2692 & n4544 ) ;
  assign n7571 = ( ~n2491 & n6372 ) | ( ~n2491 & n7570 ) | ( n6372 & n7570 ) ;
  assign n7572 = n7171 | n7571 ;
  assign n7573 = n2297 ^ n1758 ^ n538 ;
  assign n7574 = n7573 ^ n2668 ^ n2378 ;
  assign n7575 = x89 & n7574 ;
  assign n7576 = ( n916 & ~n2562 ) | ( n916 & n3429 ) | ( ~n2562 & n3429 ) ;
  assign n7577 = n7576 ^ n3777 ^ n2651 ;
  assign n7578 = ( n589 & ~n4273 ) | ( n589 & n7577 ) | ( ~n4273 & n7577 ) ;
  assign n7579 = n1716 | n3640 ;
  assign n7580 = n7578 | n7579 ;
  assign n7581 = ( n7572 & n7575 ) | ( n7572 & ~n7580 ) | ( n7575 & ~n7580 ) ;
  assign n7589 = ( ~n844 & n1344 ) | ( ~n844 & n3073 ) | ( n1344 & n3073 ) ;
  assign n7582 = n3579 ^ n334 ^ n256 ;
  assign n7583 = ~n5667 & n7582 ;
  assign n7584 = n2130 | n4315 ;
  assign n7585 = ( n2068 & n5278 ) | ( n2068 & n7584 ) | ( n5278 & n7584 ) ;
  assign n7586 = n7101 & n7585 ;
  assign n7587 = n7586 ^ n7353 ^ 1'b0 ;
  assign n7588 = ( ~n3145 & n7583 ) | ( ~n3145 & n7587 ) | ( n7583 & n7587 ) ;
  assign n7590 = n7589 ^ n7588 ^ n2567 ;
  assign n7591 = n6452 ^ n2728 ^ n1808 ;
  assign n7592 = ( n2811 & n6020 ) | ( n2811 & n7591 ) | ( n6020 & n7591 ) ;
  assign n7593 = ( n269 & ~n2625 ) | ( n269 & n6007 ) | ( ~n2625 & n6007 ) ;
  assign n7594 = ~n2608 & n3369 ;
  assign n7603 = ~n362 & n1249 ;
  assign n7604 = ~x57 & n4122 ;
  assign n7605 = n7604 ^ n1766 ^ n1422 ;
  assign n7606 = ( n753 & ~n2078 ) | ( n753 & n7605 ) | ( ~n2078 & n7605 ) ;
  assign n7607 = ( ~n5155 & n7603 ) | ( ~n5155 & n7606 ) | ( n7603 & n7606 ) ;
  assign n7608 = n5445 & n7607 ;
  assign n7609 = n7608 ^ n4859 ^ 1'b0 ;
  assign n7595 = x86 & ~n732 ;
  assign n7596 = ( n2000 & ~n2127 ) | ( n2000 & n3096 ) | ( ~n2127 & n3096 ) ;
  assign n7597 = n7596 ^ n3535 ^ 1'b0 ;
  assign n7598 = n2856 & n7597 ;
  assign n7599 = n7598 ^ n2963 ^ n2880 ;
  assign n7600 = ( ~n4627 & n7595 ) | ( ~n4627 & n7599 ) | ( n7595 & n7599 ) ;
  assign n7601 = ~n2413 & n7600 ;
  assign n7602 = n1271 & n7601 ;
  assign n7610 = n7609 ^ n7602 ^ 1'b0 ;
  assign n7611 = n7594 & n7610 ;
  assign n7612 = ~n3556 & n5564 ;
  assign n7613 = n6303 ^ n4005 ^ n1505 ;
  assign n7614 = ( n999 & n2730 ) | ( n999 & ~n7613 ) | ( n2730 & ~n7613 ) ;
  assign n7615 = ( n3360 & ~n6394 ) | ( n3360 & n7614 ) | ( ~n6394 & n7614 ) ;
  assign n7616 = n7612 & n7615 ;
  assign n7617 = ~n7611 & n7616 ;
  assign n7618 = ( n7592 & n7593 ) | ( n7592 & ~n7617 ) | ( n7593 & ~n7617 ) ;
  assign n7619 = ( n4858 & n6582 ) | ( n4858 & n6815 ) | ( n6582 & n6815 ) ;
  assign n7620 = ( n4014 & ~n4694 ) | ( n4014 & n7619 ) | ( ~n4694 & n7619 ) ;
  assign n7621 = n3870 ^ n2458 ^ 1'b0 ;
  assign n7622 = n6510 & ~n7621 ;
  assign n7623 = ~n1198 & n4978 ;
  assign n7624 = n7623 ^ n5800 ^ 1'b0 ;
  assign n7625 = ( n744 & n6690 ) | ( n744 & ~n7624 ) | ( n6690 & ~n7624 ) ;
  assign n7629 = ( ~n3078 & n4187 ) | ( ~n3078 & n7485 ) | ( n4187 & n7485 ) ;
  assign n7630 = n7629 ^ n4812 ^ n348 ;
  assign n7626 = n4739 ^ n4666 ^ 1'b0 ;
  assign n7627 = n6625 & ~n7626 ;
  assign n7628 = n2626 | n7627 ;
  assign n7631 = n7630 ^ n7628 ^ n1385 ;
  assign n7636 = ( ~n2500 & n4948 ) | ( ~n2500 & n5257 ) | ( n4948 & n5257 ) ;
  assign n7632 = n267 | n1286 ;
  assign n7633 = n3163 | n7109 ;
  assign n7634 = n2052 & ~n7633 ;
  assign n7635 = ( n1585 & n7632 ) | ( n1585 & ~n7634 ) | ( n7632 & ~n7634 ) ;
  assign n7637 = n7636 ^ n7635 ^ n1823 ;
  assign n7639 = ( n3679 & ~n4591 ) | ( n3679 & n6397 ) | ( ~n4591 & n6397 ) ;
  assign n7640 = ( ~n277 & n3258 ) | ( ~n277 & n7639 ) | ( n3258 & n7639 ) ;
  assign n7641 = n7640 ^ n1833 ^ 1'b0 ;
  assign n7638 = n4175 ^ x97 ^ 1'b0 ;
  assign n7642 = n7641 ^ n7638 ^ n2876 ;
  assign n7643 = n6653 ^ n5045 ^ 1'b0 ;
  assign n7644 = n7387 & ~n7643 ;
  assign n7645 = n3753 ^ n3358 ^ n612 ;
  assign n7649 = ( n1393 & ~n3274 ) | ( n1393 & n4802 ) | ( ~n3274 & n4802 ) ;
  assign n7650 = n2322 & n7649 ;
  assign n7651 = n7650 ^ n2920 ^ 1'b0 ;
  assign n7646 = ~n1217 & n1599 ;
  assign n7647 = n7019 | n7646 ;
  assign n7648 = x77 | n7647 ;
  assign n7652 = n7651 ^ n7648 ^ 1'b0 ;
  assign n7653 = n7645 & ~n7652 ;
  assign n7654 = ( n1605 & n4665 ) | ( n1605 & n6314 ) | ( n4665 & n6314 ) ;
  assign n7655 = n7654 ^ n6999 ^ n5382 ;
  assign n7656 = n7213 | n7655 ;
  assign n7657 = n3735 & n7656 ;
  assign n7658 = n3478 ^ n3444 ^ n1021 ;
  assign n7659 = ( n1149 & n6175 ) | ( n1149 & ~n7658 ) | ( n6175 & ~n7658 ) ;
  assign n7660 = ( n608 & n1331 ) | ( n608 & n3015 ) | ( n1331 & n3015 ) ;
  assign n7661 = n4242 & ~n7660 ;
  assign n7662 = n5579 ^ n5154 ^ n748 ;
  assign n7663 = ~n1826 & n3825 ;
  assign n7664 = n3891 & n7663 ;
  assign n7666 = ( n2921 & n3805 ) | ( n2921 & n6195 ) | ( n3805 & n6195 ) ;
  assign n7665 = n469 & ~n2208 ;
  assign n7667 = n7666 ^ n7665 ^ 1'b0 ;
  assign n7668 = ( n7662 & ~n7664 ) | ( n7662 & n7667 ) | ( ~n7664 & n7667 ) ;
  assign n7669 = n2408 ^ n1419 ^ x181 ;
  assign n7670 = ( ~n1491 & n2977 ) | ( ~n1491 & n7669 ) | ( n2977 & n7669 ) ;
  assign n7671 = n5859 ^ n4489 ^ n2895 ;
  assign n7672 = ( ~n893 & n5472 ) | ( ~n893 & n7671 ) | ( n5472 & n7671 ) ;
  assign n7673 = ( n4037 & n7670 ) | ( n4037 & ~n7672 ) | ( n7670 & ~n7672 ) ;
  assign n7674 = n2444 ^ n863 ^ n526 ;
  assign n7675 = n7674 ^ n6425 ^ n4898 ;
  assign n7676 = ( n6800 & n7673 ) | ( n6800 & ~n7675 ) | ( n7673 & ~n7675 ) ;
  assign n7677 = ( x212 & n7668 ) | ( x212 & ~n7676 ) | ( n7668 & ~n7676 ) ;
  assign n7680 = n4115 & ~n7181 ;
  assign n7681 = n7680 ^ n1777 ^ 1'b0 ;
  assign n7678 = n2917 ^ n2269 ^ 1'b0 ;
  assign n7679 = ~n6411 & n7678 ;
  assign n7682 = n7681 ^ n7679 ^ n3633 ;
  assign n7683 = ~n4512 & n7682 ;
  assign n7685 = n6465 ^ n3703 ^ n1829 ;
  assign n7686 = n7685 ^ n6439 ^ n4164 ;
  assign n7684 = n7408 ^ n5007 ^ n3965 ;
  assign n7687 = n7686 ^ n7684 ^ n4780 ;
  assign n7688 = n3154 ^ n2615 ^ 1'b0 ;
  assign n7689 = ( ~x40 & n3606 ) | ( ~x40 & n7688 ) | ( n3606 & n7688 ) ;
  assign n7690 = n724 & ~n2943 ;
  assign n7691 = n7690 ^ n1114 ^ 1'b0 ;
  assign n7692 = ( n1135 & n6720 ) | ( n1135 & ~n7691 ) | ( n6720 & ~n7691 ) ;
  assign n7694 = ~n840 & n862 ;
  assign n7693 = n2809 ^ n2777 ^ n1882 ;
  assign n7695 = n7694 ^ n7693 ^ n663 ;
  assign n7696 = ( n7689 & n7692 ) | ( n7689 & n7695 ) | ( n7692 & n7695 ) ;
  assign n7697 = n4441 ^ n1283 ^ n882 ;
  assign n7698 = ( n994 & n1410 ) | ( n994 & n2784 ) | ( n1410 & n2784 ) ;
  assign n7699 = n7402 & ~n7698 ;
  assign n7700 = ( n1841 & n7119 ) | ( n1841 & n7699 ) | ( n7119 & n7699 ) ;
  assign n7701 = n7700 ^ n901 ^ n893 ;
  assign n7702 = n5889 ^ n4606 ^ 1'b0 ;
  assign n7703 = n6355 | n7702 ;
  assign n7704 = n2343 ^ x201 ^ x130 ;
  assign n7705 = n914 & n6169 ;
  assign n7706 = n7705 ^ n3995 ^ 1'b0 ;
  assign n7707 = n7706 ^ n4599 ^ n4019 ;
  assign n7708 = n7707 ^ n1236 ^ 1'b0 ;
  assign n7709 = ( n488 & n2704 ) | ( n488 & n5454 ) | ( n2704 & n5454 ) ;
  assign n7710 = n7709 ^ n3861 ^ n2522 ;
  assign n7711 = ( ~n7704 & n7708 ) | ( ~n7704 & n7710 ) | ( n7708 & n7710 ) ;
  assign n7712 = n535 & ~n3629 ;
  assign n7713 = n7712 ^ n4708 ^ 1'b0 ;
  assign n7714 = n847 | n1724 ;
  assign n7715 = n7714 ^ n441 ^ 1'b0 ;
  assign n7716 = ( n577 & n5006 ) | ( n577 & n7715 ) | ( n5006 & n7715 ) ;
  assign n7717 = n4109 & n6829 ;
  assign n7718 = ( n364 & ~n7716 ) | ( n364 & n7717 ) | ( ~n7716 & n7717 ) ;
  assign n7719 = ( ~n336 & n776 ) | ( ~n336 & n7718 ) | ( n776 & n7718 ) ;
  assign n7720 = ~n7563 & n7719 ;
  assign n7721 = n7720 ^ n7377 ^ 1'b0 ;
  assign n7722 = n7713 & n7721 ;
  assign n7723 = n782 | n2597 ;
  assign n7724 = n3535 & ~n7723 ;
  assign n7736 = n1599 | n3851 ;
  assign n7733 = ~n482 & n6827 ;
  assign n7734 = n1085 & n7733 ;
  assign n7732 = n3589 | n5283 ;
  assign n7735 = n7734 ^ n7732 ^ n4972 ;
  assign n7727 = n5125 ^ n1957 ^ n353 ;
  assign n7728 = ( n642 & n746 ) | ( n642 & ~n3022 ) | ( n746 & ~n3022 ) ;
  assign n7729 = ( n7317 & ~n7727 ) | ( n7317 & n7728 ) | ( ~n7727 & n7728 ) ;
  assign n7725 = ~n3231 & n5289 ;
  assign n7726 = n7725 ^ n2480 ^ 1'b0 ;
  assign n7730 = n7729 ^ n7726 ^ 1'b0 ;
  assign n7731 = ~n1517 & n7730 ;
  assign n7737 = n7736 ^ n7735 ^ n7731 ;
  assign n7740 = n1073 & n1565 ;
  assign n7741 = n7740 ^ n495 ^ 1'b0 ;
  assign n7742 = n7741 ^ n5524 ^ n1745 ;
  assign n7738 = n1385 ^ n1378 ^ 1'b0 ;
  assign n7739 = ( ~n6066 & n7437 ) | ( ~n6066 & n7738 ) | ( n7437 & n7738 ) ;
  assign n7743 = n7742 ^ n7739 ^ 1'b0 ;
  assign n7744 = n6159 & n7743 ;
  assign n7746 = n6223 ^ n4463 ^ n490 ;
  assign n7747 = n7746 ^ n437 ^ 1'b0 ;
  assign n7745 = n3458 & ~n6860 ;
  assign n7748 = n7747 ^ n7745 ^ n850 ;
  assign n7749 = ( x115 & n410 ) | ( x115 & ~n4821 ) | ( n410 & ~n4821 ) ;
  assign n7750 = n7749 ^ n6917 ^ n1646 ;
  assign n7751 = n1382 | n6117 ;
  assign n7752 = n7750 | n7751 ;
  assign n7753 = n7752 ^ n943 ^ 1'b0 ;
  assign n7754 = n7748 & ~n7753 ;
  assign n7755 = ( n2009 & n3662 ) | ( n2009 & ~n4064 ) | ( n3662 & ~n4064 ) ;
  assign n7756 = ( n5944 & ~n6058 ) | ( n5944 & n7755 ) | ( ~n6058 & n7755 ) ;
  assign n7757 = n6068 ^ n4161 ^ n383 ;
  assign n7758 = ( n399 & n7521 ) | ( n399 & ~n7757 ) | ( n7521 & ~n7757 ) ;
  assign n7777 = n4215 ^ n3911 ^ 1'b0 ;
  assign n7771 = ( ~n1122 & n1856 ) | ( ~n1122 & n2681 ) | ( n1856 & n2681 ) ;
  assign n7772 = n4353 ^ n2307 ^ n2233 ;
  assign n7773 = n3192 & n6524 ;
  assign n7774 = ~n7772 & n7773 ;
  assign n7775 = ( n7410 & n7771 ) | ( n7410 & ~n7774 ) | ( n7771 & ~n7774 ) ;
  assign n7763 = n1474 ^ n1059 ^ x122 ;
  assign n7764 = ( ~x155 & n3376 ) | ( ~x155 & n7763 ) | ( n3376 & n7763 ) ;
  assign n7765 = ( n1618 & n5142 ) | ( n1618 & n5310 ) | ( n5142 & n5310 ) ;
  assign n7766 = ( n1783 & n1842 ) | ( n1783 & ~n7765 ) | ( n1842 & ~n7765 ) ;
  assign n7767 = n6857 ^ n4163 ^ n3598 ;
  assign n7768 = ( ~n482 & n7766 ) | ( ~n482 & n7767 ) | ( n7766 & n7767 ) ;
  assign n7769 = ~n3742 & n7768 ;
  assign n7770 = ~n7764 & n7769 ;
  assign n7776 = n7775 ^ n7770 ^ n5624 ;
  assign n7759 = n1396 ^ n1112 ^ 1'b0 ;
  assign n7760 = n3366 ^ n2819 ^ x94 ;
  assign n7761 = n346 & ~n7760 ;
  assign n7762 = ~n7759 & n7761 ;
  assign n7778 = n7777 ^ n7776 ^ n7762 ;
  assign n7779 = n7778 ^ n532 ^ 1'b0 ;
  assign n7800 = n2881 ^ x165 ^ 1'b0 ;
  assign n7801 = n3913 & ~n7800 ;
  assign n7802 = ~x200 & n7801 ;
  assign n7803 = n7802 ^ n2998 ^ 1'b0 ;
  assign n7804 = n7803 ^ x6 ^ 1'b0 ;
  assign n7790 = n1369 | n3018 ;
  assign n7791 = n7790 ^ n379 ^ 1'b0 ;
  assign n7792 = ( n2976 & n3093 ) | ( n2976 & n6805 ) | ( n3093 & n6805 ) ;
  assign n7793 = n7792 ^ n3266 ^ n2521 ;
  assign n7794 = ( ~n3619 & n7791 ) | ( ~n3619 & n7793 ) | ( n7791 & n7793 ) ;
  assign n7796 = ( n2104 & n2309 ) | ( n2104 & ~n2679 ) | ( n2309 & ~n2679 ) ;
  assign n7795 = n4172 ^ n2389 ^ n868 ;
  assign n7797 = n7796 ^ n7795 ^ n3025 ;
  assign n7798 = ( n853 & n7794 ) | ( n853 & ~n7797 ) | ( n7794 & ~n7797 ) ;
  assign n7785 = n1039 ^ n979 ^ 1'b0 ;
  assign n7786 = n646 | n7785 ;
  assign n7787 = n2772 ^ n2046 ^ 1'b0 ;
  assign n7788 = n7787 ^ n1935 ^ 1'b0 ;
  assign n7789 = ~n7786 & n7788 ;
  assign n7799 = n7798 ^ n7789 ^ n1456 ;
  assign n7783 = n1478 ^ n476 ^ 1'b0 ;
  assign n7780 = n2285 ^ n1374 ^ n1334 ;
  assign n7781 = ( n2315 & n6631 ) | ( n2315 & n7780 ) | ( n6631 & n7780 ) ;
  assign n7782 = n5446 & ~n7781 ;
  assign n7784 = n7783 ^ n7782 ^ 1'b0 ;
  assign n7805 = n7804 ^ n7799 ^ n7784 ;
  assign n7808 = ( ~n594 & n3387 ) | ( ~n594 & n4599 ) | ( n3387 & n4599 ) ;
  assign n7806 = ( n2953 & n5344 ) | ( n2953 & n7707 ) | ( n5344 & n7707 ) ;
  assign n7807 = ( x16 & n5817 ) | ( x16 & ~n7806 ) | ( n5817 & ~n7806 ) ;
  assign n7809 = n7808 ^ n7807 ^ n2852 ;
  assign n7811 = ( n354 & n1305 ) | ( n354 & ~n3795 ) | ( n1305 & ~n3795 ) ;
  assign n7810 = n7431 ^ n696 ^ 1'b0 ;
  assign n7812 = n7811 ^ n7810 ^ 1'b0 ;
  assign n7819 = n6207 ^ n4381 ^ n1361 ;
  assign n7814 = n4693 & ~n7455 ;
  assign n7815 = n954 & n7814 ;
  assign n7816 = n2052 ^ n1972 ^ x57 ;
  assign n7817 = n7816 ^ n2152 ^ 1'b0 ;
  assign n7818 = ( n5189 & n7815 ) | ( n5189 & n7817 ) | ( n7815 & n7817 ) ;
  assign n7820 = n7819 ^ n7818 ^ n7545 ;
  assign n7813 = x22 & ~n2099 ;
  assign n7821 = n7820 ^ n7813 ^ 1'b0 ;
  assign n7822 = n4924 ^ n3078 ^ n2886 ;
  assign n7823 = n405 & ~n6680 ;
  assign n7824 = n7823 ^ n975 ^ 1'b0 ;
  assign n7825 = ( x103 & n868 ) | ( x103 & n3376 ) | ( n868 & n3376 ) ;
  assign n7826 = n1075 | n7825 ;
  assign n7827 = n7826 ^ n1635 ^ 1'b0 ;
  assign n7828 = ( n851 & n2561 ) | ( n851 & ~n5274 ) | ( n2561 & ~n5274 ) ;
  assign n7829 = n7828 ^ n4464 ^ n577 ;
  assign n7830 = n6944 ^ n6140 ^ n3516 ;
  assign n7831 = n3990 | n4478 ;
  assign n7832 = n7830 | n7831 ;
  assign n7833 = n7832 ^ n698 ^ 1'b0 ;
  assign n7834 = ~n7829 & n7833 ;
  assign n7835 = n365 | n2883 ;
  assign n7836 = n7835 ^ n4892 ^ n4396 ;
  assign n7837 = n5136 & n7836 ;
  assign n7838 = ( n1496 & n1647 ) | ( n1496 & ~n4948 ) | ( n1647 & ~n4948 ) ;
  assign n7839 = n7838 ^ n6443 ^ n4017 ;
  assign n7840 = ( ~n3328 & n7837 ) | ( ~n3328 & n7839 ) | ( n7837 & n7839 ) ;
  assign n7841 = ~n569 & n4785 ;
  assign n7842 = ~n2076 & n7841 ;
  assign n7843 = n7842 ^ n4433 ^ 1'b0 ;
  assign n7844 = ( ~n592 & n918 ) | ( ~n592 & n7843 ) | ( n918 & n7843 ) ;
  assign n7845 = n6041 ^ n3327 ^ n2974 ;
  assign n7846 = n7845 ^ n1476 ^ 1'b0 ;
  assign n7847 = ~n2232 & n7846 ;
  assign n7848 = n7847 ^ n4794 ^ n1204 ;
  assign n7849 = ( ~n2979 & n3170 ) | ( ~n2979 & n3925 ) | ( n3170 & n3925 ) ;
  assign n7850 = n5908 & ~n7849 ;
  assign n7851 = n7850 ^ n5632 ^ n2200 ;
  assign n7852 = ( ~x223 & n1517 ) | ( ~x223 & n1900 ) | ( n1517 & n1900 ) ;
  assign n7864 = ( n292 & ~n558 ) | ( n292 & n2295 ) | ( ~n558 & n2295 ) ;
  assign n7865 = ( n501 & ~n2664 ) | ( n501 & n7864 ) | ( ~n2664 & n7864 ) ;
  assign n7866 = n5448 ^ n3889 ^ n2895 ;
  assign n7867 = ( n5379 & ~n7865 ) | ( n5379 & n7866 ) | ( ~n7865 & n7866 ) ;
  assign n7862 = n5769 ^ n2317 ^ n1242 ;
  assign n7853 = n2074 | n5718 ;
  assign n7854 = n7853 ^ n5289 ^ 1'b0 ;
  assign n7855 = ~n525 & n7854 ;
  assign n7856 = n7855 ^ n5627 ^ 1'b0 ;
  assign n7857 = n939 & ~n3655 ;
  assign n7858 = n7857 ^ n5584 ^ 1'b0 ;
  assign n7859 = n278 | n7858 ;
  assign n7860 = n7856 | n7859 ;
  assign n7861 = n4018 & n7860 ;
  assign n7863 = n7862 ^ n7861 ^ 1'b0 ;
  assign n7868 = n7867 ^ n7863 ^ 1'b0 ;
  assign n7869 = ( x216 & n7852 ) | ( x216 & ~n7868 ) | ( n7852 & ~n7868 ) ;
  assign n7871 = ( x39 & n6342 ) | ( x39 & n7454 ) | ( n6342 & n7454 ) ;
  assign n7870 = n6670 ^ n3901 ^ n1363 ;
  assign n7872 = n7871 ^ n7870 ^ n7323 ;
  assign n7873 = n7872 ^ n2938 ^ n870 ;
  assign n7874 = ( x196 & ~n1110 ) | ( x196 & n2818 ) | ( ~n1110 & n2818 ) ;
  assign n7875 = ( ~n839 & n4906 ) | ( ~n839 & n7704 ) | ( n4906 & n7704 ) ;
  assign n7876 = ( n2427 & n7874 ) | ( n2427 & ~n7875 ) | ( n7874 & ~n7875 ) ;
  assign n7877 = ( n3557 & n7008 ) | ( n3557 & n7876 ) | ( n7008 & n7876 ) ;
  assign n7878 = n2773 | n6476 ;
  assign n7879 = ~n3146 & n3616 ;
  assign n7880 = n7878 & n7879 ;
  assign n7881 = ( n2905 & n7715 ) | ( n2905 & n7880 ) | ( n7715 & n7880 ) ;
  assign n7882 = ( n1060 & n4957 ) | ( n1060 & ~n7881 ) | ( n4957 & ~n7881 ) ;
  assign n7883 = n4340 ^ n2072 ^ n531 ;
  assign n7884 = ( n2928 & ~n5856 ) | ( n2928 & n7883 ) | ( ~n5856 & n7883 ) ;
  assign n7886 = n2855 | n6600 ;
  assign n7887 = n7886 ^ n482 ^ 1'b0 ;
  assign n7885 = n6122 ^ n2682 ^ n1885 ;
  assign n7888 = n7887 ^ n7885 ^ n1885 ;
  assign n7889 = n7888 ^ n4879 ^ 1'b0 ;
  assign n7890 = ~n7884 & n7889 ;
  assign n7891 = ( n716 & n840 ) | ( n716 & n2064 ) | ( n840 & n2064 ) ;
  assign n7893 = ( ~n1492 & n1680 ) | ( ~n1492 & n5838 ) | ( n1680 & n5838 ) ;
  assign n7894 = ( ~n2869 & n3044 ) | ( ~n2869 & n7893 ) | ( n3044 & n7893 ) ;
  assign n7892 = ( n596 & n1371 ) | ( n596 & ~n1372 ) | ( n1371 & ~n1372 ) ;
  assign n7895 = n7894 ^ n7892 ^ 1'b0 ;
  assign n7896 = ~n1094 & n7895 ;
  assign n7897 = n7896 ^ n3257 ^ 1'b0 ;
  assign n7898 = ( n5505 & n7891 ) | ( n5505 & ~n7897 ) | ( n7891 & ~n7897 ) ;
  assign n7899 = n716 & n7898 ;
  assign n7900 = n7899 ^ n3655 ^ 1'b0 ;
  assign n7901 = ( ~n2343 & n2583 ) | ( ~n2343 & n4099 ) | ( n2583 & n4099 ) ;
  assign n7902 = ( n1875 & ~n4354 ) | ( n1875 & n7901 ) | ( ~n4354 & n7901 ) ;
  assign n7903 = ( x133 & n6885 ) | ( x133 & n7902 ) | ( n6885 & n7902 ) ;
  assign n7906 = n1596 ^ n1497 ^ x51 ;
  assign n7905 = n7299 ^ n3236 ^ n977 ;
  assign n7904 = n6111 ^ n2182 ^ 1'b0 ;
  assign n7907 = n7906 ^ n7905 ^ n7904 ;
  assign n7908 = n7907 ^ n624 ^ 1'b0 ;
  assign n7915 = n980 ^ n447 ^ x172 ;
  assign n7916 = n7178 & ~n7915 ;
  assign n7917 = n4128 & n7916 ;
  assign n7918 = ( n3405 & ~n3873 ) | ( n3405 & n6680 ) | ( ~n3873 & n6680 ) ;
  assign n7919 = ( n2879 & n7917 ) | ( n2879 & ~n7918 ) | ( n7917 & ~n7918 ) ;
  assign n7909 = n6540 ^ n5223 ^ n333 ;
  assign n7912 = n5997 ^ n604 ^ n317 ;
  assign n7911 = ( n1483 & ~n3754 ) | ( n1483 & n4197 ) | ( ~n3754 & n4197 ) ;
  assign n7910 = n5000 ^ n1962 ^ n447 ;
  assign n7913 = n7912 ^ n7911 ^ n7910 ;
  assign n7914 = ( n4841 & n7909 ) | ( n4841 & ~n7913 ) | ( n7909 & ~n7913 ) ;
  assign n7920 = n7919 ^ n7914 ^ n2344 ;
  assign n7922 = ( n270 & n3458 ) | ( n270 & ~n6317 ) | ( n3458 & ~n6317 ) ;
  assign n7921 = n6647 ^ n1095 ^ 1'b0 ;
  assign n7923 = n7922 ^ n7921 ^ n1059 ;
  assign n7924 = n3316 ^ n1619 ^ 1'b0 ;
  assign n7925 = n554 & ~n7924 ;
  assign n7926 = n7925 ^ n6063 ^ n730 ;
  assign n7927 = n7926 ^ n7403 ^ n1113 ;
  assign n7928 = ( n4427 & n4695 ) | ( n4427 & n5997 ) | ( n4695 & n5997 ) ;
  assign n7929 = ~n875 & n2641 ;
  assign n7930 = n7929 ^ n523 ^ 1'b0 ;
  assign n7931 = n7124 ^ n6148 ^ 1'b0 ;
  assign n7932 = n3561 | n7903 ;
  assign n7933 = n5661 ^ n3707 ^ n469 ;
  assign n7934 = ( n4697 & n6586 ) | ( n4697 & ~n7933 ) | ( n6586 & ~n7933 ) ;
  assign n7935 = x155 & n4635 ;
  assign n7936 = n7935 ^ n1140 ^ 1'b0 ;
  assign n7937 = n339 & ~n697 ;
  assign n7938 = n7937 ^ n929 ^ 1'b0 ;
  assign n7939 = n861 & n2183 ;
  assign n7940 = n740 & n7939 ;
  assign n7941 = ~x205 & n2635 ;
  assign n7942 = ( n7938 & n7940 ) | ( n7938 & ~n7941 ) | ( n7940 & ~n7941 ) ;
  assign n7943 = n7942 ^ n4606 ^ n1410 ;
  assign n7944 = n7943 ^ n2096 ^ n1276 ;
  assign n7945 = n7936 & n7944 ;
  assign n7946 = ~x245 & n2911 ;
  assign n7947 = ( n1493 & n7945 ) | ( n1493 & ~n7946 ) | ( n7945 & ~n7946 ) ;
  assign n7948 = ( n5266 & n5658 ) | ( n5266 & n7947 ) | ( n5658 & n7947 ) ;
  assign n7949 = n7948 ^ n7735 ^ 1'b0 ;
  assign n7950 = ~n5645 & n6197 ;
  assign n7951 = ( n463 & ~n3966 ) | ( n463 & n7950 ) | ( ~n3966 & n7950 ) ;
  assign n7953 = n1642 & n5020 ;
  assign n7952 = n2048 ^ n345 ^ 1'b0 ;
  assign n7954 = n7953 ^ n7952 ^ 1'b0 ;
  assign n7955 = ( x165 & n1469 ) | ( x165 & ~n2464 ) | ( n1469 & ~n2464 ) ;
  assign n7956 = n7955 ^ n3430 ^ n3166 ;
  assign n7957 = n7956 ^ n5716 ^ n4446 ;
  assign n7958 = n7957 ^ n4515 ^ n2597 ;
  assign n7959 = ( ~n4266 & n5522 ) | ( ~n4266 & n7958 ) | ( n5522 & n7958 ) ;
  assign n7960 = n3146 ^ n1019 ^ 1'b0 ;
  assign n7961 = x80 & ~n7960 ;
  assign n7962 = ( n1464 & n1670 ) | ( n1464 & ~n7961 ) | ( n1670 & ~n7961 ) ;
  assign n7963 = n826 | n1586 ;
  assign n7964 = ( n343 & n2093 ) | ( n343 & ~n2464 ) | ( n2093 & ~n2464 ) ;
  assign n7965 = ( ~n2559 & n4011 ) | ( ~n2559 & n4134 ) | ( n4011 & n4134 ) ;
  assign n7966 = n7965 ^ n6616 ^ n1523 ;
  assign n7967 = n7966 ^ n1058 ^ 1'b0 ;
  assign n7968 = n7964 | n7967 ;
  assign n7969 = ( n7962 & n7963 ) | ( n7962 & ~n7968 ) | ( n7963 & ~n7968 ) ;
  assign n7970 = ( n5332 & n5400 ) | ( n5332 & n7919 ) | ( n5400 & n7919 ) ;
  assign n7971 = ( n5640 & ~n5685 ) | ( n5640 & n7970 ) | ( ~n5685 & n7970 ) ;
  assign n7972 = ( n2024 & n5595 ) | ( n2024 & n6419 ) | ( n5595 & n6419 ) ;
  assign n7976 = n5267 ^ n2130 ^ 1'b0 ;
  assign n7975 = n3437 ^ n2072 ^ n1326 ;
  assign n7977 = n7976 ^ n7975 ^ n2970 ;
  assign n7978 = n6359 & ~n7977 ;
  assign n7979 = n1763 & n7978 ;
  assign n7980 = ( ~n4264 & n6516 ) | ( ~n4264 & n7979 ) | ( n6516 & n7979 ) ;
  assign n7973 = ~x228 & n2414 ;
  assign n7974 = n7973 ^ n4450 ^ n3938 ;
  assign n7981 = n7980 ^ n7974 ^ n7322 ;
  assign n7982 = n3349 ^ n2376 ^ 1'b0 ;
  assign n7983 = n911 & n7982 ;
  assign n7984 = ( n2215 & n3750 ) | ( n2215 & n7983 ) | ( n3750 & n7983 ) ;
  assign n7985 = ~n7440 & n7984 ;
  assign n7986 = ~n4849 & n7985 ;
  assign n7987 = n7418 ^ n7285 ^ n5615 ;
  assign n7988 = ( ~n6197 & n7986 ) | ( ~n6197 & n7987 ) | ( n7986 & n7987 ) ;
  assign n7994 = ( n823 & n1901 ) | ( n823 & n3514 ) | ( n1901 & n3514 ) ;
  assign n7995 = ( n592 & n987 ) | ( n592 & n1844 ) | ( n987 & n1844 ) ;
  assign n7996 = n3807 | n7995 ;
  assign n7997 = n2134 & ~n7996 ;
  assign n7998 = ( n3951 & n7994 ) | ( n3951 & ~n7997 ) | ( n7994 & ~n7997 ) ;
  assign n7999 = ( n4017 & n5511 ) | ( n4017 & n7998 ) | ( n5511 & n7998 ) ;
  assign n7989 = n4341 ^ n3178 ^ n957 ;
  assign n7990 = ( ~n318 & n1797 ) | ( ~n318 & n2311 ) | ( n1797 & n2311 ) ;
  assign n7991 = n7990 ^ n3861 ^ n906 ;
  assign n7992 = ( n4663 & n7989 ) | ( n4663 & ~n7991 ) | ( n7989 & ~n7991 ) ;
  assign n7993 = n713 & n7992 ;
  assign n8000 = n7999 ^ n7993 ^ 1'b0 ;
  assign n8027 = n3467 ^ n1412 ^ x37 ;
  assign n8025 = ( n1098 & n4491 ) | ( n1098 & ~n7178 ) | ( n4491 & ~n7178 ) ;
  assign n8026 = n8025 ^ n5056 ^ n2941 ;
  assign n8001 = n4712 ^ n4117 ^ 1'b0 ;
  assign n8002 = ~n1627 & n8001 ;
  assign n8003 = n6969 ^ n4504 ^ n4094 ;
  assign n8004 = n891 ^ n380 ^ x170 ;
  assign n8005 = n8004 ^ n5855 ^ n3794 ;
  assign n8006 = n8003 | n8005 ;
  assign n8007 = ( n4101 & n8002 ) | ( n4101 & n8006 ) | ( n8002 & n8006 ) ;
  assign n8017 = ( x166 & ~n2739 ) | ( x166 & n3246 ) | ( ~n2739 & n3246 ) ;
  assign n8012 = n3792 ^ x19 ^ 1'b0 ;
  assign n8013 = ~n931 & n8012 ;
  assign n8014 = n8013 ^ n5502 ^ n1482 ;
  assign n8010 = n1779 ^ n1671 ^ n1612 ;
  assign n8011 = ( ~n3126 & n4627 ) | ( ~n3126 & n8010 ) | ( n4627 & n8010 ) ;
  assign n8015 = n8014 ^ n8011 ^ 1'b0 ;
  assign n8016 = n649 & ~n8015 ;
  assign n8008 = n1926 ^ n1281 ^ 1'b0 ;
  assign n8009 = n8008 ^ n7523 ^ x46 ;
  assign n8018 = n8017 ^ n8016 ^ n8009 ;
  assign n8019 = n2682 ^ n952 ^ 1'b0 ;
  assign n8020 = n8019 ^ n1666 ^ 1'b0 ;
  assign n8021 = n4992 | n8020 ;
  assign n8022 = n8021 ^ n4243 ^ 1'b0 ;
  assign n8023 = n8018 & ~n8022 ;
  assign n8024 = n8007 & n8023 ;
  assign n8028 = n8027 ^ n8026 ^ n8024 ;
  assign n8029 = n2209 & n8028 ;
  assign n8030 = ( ~x108 & n5179 ) | ( ~x108 & n6483 ) | ( n5179 & n6483 ) ;
  assign n8031 = n6475 ^ n5637 ^ n1180 ;
  assign n8032 = ( ~n5275 & n7023 ) | ( ~n5275 & n8031 ) | ( n7023 & n8031 ) ;
  assign n8033 = ~n8030 & n8032 ;
  assign n8034 = n4409 ^ n3813 ^ n1865 ;
  assign n8035 = n8034 ^ n6336 ^ n3680 ;
  assign n8036 = n8035 ^ n4129 ^ n2052 ;
  assign n8037 = n4148 | n8036 ;
  assign n8038 = n8037 ^ n5257 ^ 1'b0 ;
  assign n8039 = n7727 ^ n1972 ^ n1824 ;
  assign n8040 = ( n6890 & n8038 ) | ( n6890 & ~n8039 ) | ( n8038 & ~n8039 ) ;
  assign n8041 = ( n7255 & n8033 ) | ( n7255 & n8040 ) | ( n8033 & n8040 ) ;
  assign n8042 = ~n926 & n2336 ;
  assign n8043 = ( n1775 & n5064 ) | ( n1775 & n8042 ) | ( n5064 & n8042 ) ;
  assign n8044 = n8043 ^ n1204 ^ 1'b0 ;
  assign n8045 = n7266 ^ n3435 ^ n2191 ;
  assign n8046 = n6412 | n6482 ;
  assign n8047 = ( n5310 & n8045 ) | ( n5310 & n8046 ) | ( n8045 & n8046 ) ;
  assign n8048 = ~n761 & n3910 ;
  assign n8049 = n8048 ^ n3136 ^ 1'b0 ;
  assign n8050 = n2592 & ~n8049 ;
  assign n8051 = ( n447 & ~n898 ) | ( n447 & n1834 ) | ( ~n898 & n1834 ) ;
  assign n8052 = ( n2495 & n4978 ) | ( n2495 & n8051 ) | ( n4978 & n8051 ) ;
  assign n8053 = ( n4609 & n6269 ) | ( n4609 & ~n8052 ) | ( n6269 & ~n8052 ) ;
  assign n8054 = ~n4992 & n5128 ;
  assign n8055 = ( n2916 & n3774 ) | ( n2916 & n4375 ) | ( n3774 & n4375 ) ;
  assign n8056 = n6287 ^ n4698 ^ n2773 ;
  assign n8057 = n8056 ^ n7217 ^ x167 ;
  assign n8058 = ( ~x218 & n8055 ) | ( ~x218 & n8057 ) | ( n8055 & n8057 ) ;
  assign n8059 = n6910 ^ n5693 ^ n5056 ;
  assign n8060 = n7039 ^ n1860 ^ 1'b0 ;
  assign n8061 = ( n7697 & n8059 ) | ( n7697 & n8060 ) | ( n8059 & n8060 ) ;
  assign n8062 = ( ~x105 & n4160 ) | ( ~x105 & n6160 ) | ( n4160 & n6160 ) ;
  assign n8063 = ( n262 & n6756 ) | ( n262 & ~n7794 ) | ( n6756 & ~n7794 ) ;
  assign n8064 = ( n3250 & n4497 ) | ( n3250 & ~n6750 ) | ( n4497 & ~n6750 ) ;
  assign n8065 = ( ~n846 & n1021 ) | ( ~n846 & n2591 ) | ( n1021 & n2591 ) ;
  assign n8066 = n778 & n3410 ;
  assign n8067 = n8066 ^ n828 ^ 1'b0 ;
  assign n8068 = n8065 & n8067 ;
  assign n8069 = n8068 ^ n3318 ^ 1'b0 ;
  assign n8070 = n4553 ^ n4368 ^ n1182 ;
  assign n8071 = ( n1443 & n6805 ) | ( n1443 & ~n7904 ) | ( n6805 & ~n7904 ) ;
  assign n8072 = ( n2698 & ~n2731 ) | ( n2698 & n8071 ) | ( ~n2731 & n8071 ) ;
  assign n8073 = ~n981 & n2728 ;
  assign n8074 = n8073 ^ n2774 ^ 1'b0 ;
  assign n8075 = n7327 & ~n8074 ;
  assign n8076 = n580 & ~n7495 ;
  assign n8077 = ( ~n5161 & n5164 ) | ( ~n5161 & n7925 ) | ( n5164 & n7925 ) ;
  assign n8078 = ( ~n3652 & n5173 ) | ( ~n3652 & n5795 ) | ( n5173 & n5795 ) ;
  assign n8081 = n6669 ^ n3102 ^ x94 ;
  assign n8079 = n5950 ^ n5940 ^ 1'b0 ;
  assign n8080 = ~n7995 & n8079 ;
  assign n8082 = n8081 ^ n8080 ^ n589 ;
  assign n8083 = ( ~n7483 & n8078 ) | ( ~n7483 & n8082 ) | ( n8078 & n8082 ) ;
  assign n8084 = n8083 ^ n4631 ^ n3096 ;
  assign n8085 = n8077 & ~n8084 ;
  assign n8086 = ~n8076 & n8085 ;
  assign n8087 = n4357 ^ n943 ^ 1'b0 ;
  assign n8088 = ( n1430 & ~n2132 ) | ( n1430 & n3105 ) | ( ~n2132 & n3105 ) ;
  assign n8091 = n5188 ^ n1221 ^ x242 ;
  assign n8089 = n4647 ^ n4473 ^ 1'b0 ;
  assign n8090 = n1008 & n8089 ;
  assign n8092 = n8091 ^ n8090 ^ x236 ;
  assign n8093 = n1875 & ~n8092 ;
  assign n8094 = ( n8087 & n8088 ) | ( n8087 & n8093 ) | ( n8088 & n8093 ) ;
  assign n8095 = n4023 ^ n2238 ^ x228 ;
  assign n8096 = ( x22 & n2829 ) | ( x22 & ~n7801 ) | ( n2829 & ~n7801 ) ;
  assign n8097 = ( n3680 & n4957 ) | ( n3680 & n8096 ) | ( n4957 & n8096 ) ;
  assign n8098 = n8095 & ~n8097 ;
  assign n8099 = n8098 ^ n5190 ^ 1'b0 ;
  assign n8104 = n3139 ^ n1447 ^ n384 ;
  assign n8102 = n471 ^ n363 ^ x53 ;
  assign n8103 = n8102 ^ n6752 ^ n463 ;
  assign n8100 = ( n2671 & ~n3395 ) | ( n2671 & n5365 ) | ( ~n3395 & n5365 ) ;
  assign n8101 = n8100 ^ n6071 ^ n3634 ;
  assign n8105 = n8104 ^ n8103 ^ n8101 ;
  assign n8106 = ( ~n8094 & n8099 ) | ( ~n8094 & n8105 ) | ( n8099 & n8105 ) ;
  assign n8107 = n2273 & n3214 ;
  assign n8108 = n8107 ^ n7325 ^ 1'b0 ;
  assign n8109 = n4215 & ~n8108 ;
  assign n8110 = n8109 ^ n7359 ^ 1'b0 ;
  assign n8111 = ( n1839 & n3218 ) | ( n1839 & n8110 ) | ( n3218 & n8110 ) ;
  assign n8112 = ( ~n690 & n3119 ) | ( ~n690 & n7941 ) | ( n3119 & n7941 ) ;
  assign n8113 = n8112 ^ x116 ^ 1'b0 ;
  assign n8119 = ~n2223 & n8096 ;
  assign n8120 = n8119 ^ n3209 ^ 1'b0 ;
  assign n8116 = ( n578 & n3932 ) | ( n578 & n5806 ) | ( n3932 & n5806 ) ;
  assign n8114 = n928 & n2739 ;
  assign n8115 = ~n6943 & n8114 ;
  assign n8117 = n8116 ^ n8115 ^ n5482 ;
  assign n8118 = ( n1575 & n3010 ) | ( n1575 & n8117 ) | ( n3010 & n8117 ) ;
  assign n8121 = n8120 ^ n8118 ^ n4217 ;
  assign n8122 = n3268 & ~n8121 ;
  assign n8123 = n8113 & n8122 ;
  assign n8124 = n7972 ^ n1988 ^ x43 ;
  assign n8125 = n2216 | n8124 ;
  assign n8127 = ( n2651 & ~n3750 ) | ( n2651 & n4075 ) | ( ~n3750 & n4075 ) ;
  assign n8128 = n2674 | n8127 ;
  assign n8129 = n8128 ^ n6625 ^ 1'b0 ;
  assign n8126 = ~n2187 & n3780 ;
  assign n8130 = n8129 ^ n8126 ^ n2048 ;
  assign n8131 = ( n2320 & n2912 ) | ( n2320 & ~n8130 ) | ( n2912 & ~n8130 ) ;
  assign n8132 = n1406 | n6282 ;
  assign n8133 = n8132 ^ n3629 ^ 1'b0 ;
  assign n8134 = n8131 | n8133 ;
  assign n8136 = n4785 & n5459 ;
  assign n8137 = ~n2857 & n8136 ;
  assign n8135 = ( n1142 & n1679 ) | ( n1142 & ~n4604 ) | ( n1679 & ~n4604 ) ;
  assign n8138 = n8137 ^ n8135 ^ n5907 ;
  assign n8139 = ~n3752 & n8138 ;
  assign n8140 = n7964 ^ n1025 ^ x253 ;
  assign n8141 = n2637 & n8140 ;
  assign n8142 = n8141 ^ n594 ^ 1'b0 ;
  assign n8143 = n8142 ^ n7771 ^ 1'b0 ;
  assign n8145 = n2232 | n3479 ;
  assign n8146 = ( n1164 & n1310 ) | ( n1164 & n6787 ) | ( n1310 & n6787 ) ;
  assign n8147 = ( ~n496 & n8145 ) | ( ~n496 & n8146 ) | ( n8145 & n8146 ) ;
  assign n8154 = n817 & n2528 ;
  assign n8155 = n4045 & n8154 ;
  assign n8148 = ~n410 & n2971 ;
  assign n8149 = ( ~n1831 & n2510 ) | ( ~n1831 & n4307 ) | ( n2510 & n4307 ) ;
  assign n8150 = n8149 ^ n5560 ^ n4788 ;
  assign n8151 = ~n7727 & n8150 ;
  assign n8152 = n8148 & ~n8151 ;
  assign n8153 = n8152 ^ n7281 ^ 1'b0 ;
  assign n8156 = n8155 ^ n8153 ^ n5249 ;
  assign n8157 = ( n2421 & n8147 ) | ( n2421 & n8156 ) | ( n8147 & n8156 ) ;
  assign n8144 = n3582 | n3639 ;
  assign n8158 = n8157 ^ n8144 ^ 1'b0 ;
  assign n8163 = ( n1434 & ~n3166 ) | ( n1434 & n7511 ) | ( ~n3166 & n7511 ) ;
  assign n8161 = n3750 ^ n1889 ^ n496 ;
  assign n8162 = n2024 | n8161 ;
  assign n8159 = n6552 ^ n5212 ^ 1'b0 ;
  assign n8160 = n328 & ~n8159 ;
  assign n8164 = n8163 ^ n8162 ^ n8160 ;
  assign n8165 = ( n468 & n6723 ) | ( n468 & n8164 ) | ( n6723 & n8164 ) ;
  assign n8166 = n1945 | n5628 ;
  assign n8167 = n3306 & ~n3879 ;
  assign n8168 = ( n485 & n4571 ) | ( n485 & n8167 ) | ( n4571 & n8167 ) ;
  assign n8169 = n7709 ^ n5374 ^ n4063 ;
  assign n8170 = ( ~n6644 & n8168 ) | ( ~n6644 & n8169 ) | ( n8168 & n8169 ) ;
  assign n8171 = n8170 ^ n1483 ^ 1'b0 ;
  assign n8172 = n1719 ^ n1098 ^ 1'b0 ;
  assign n8173 = n8172 ^ n7112 ^ 1'b0 ;
  assign n8182 = n3981 ^ x185 ^ 1'b0 ;
  assign n8178 = ( n938 & ~n1491 ) | ( n938 & n4720 ) | ( ~n1491 & n4720 ) ;
  assign n8179 = n8178 ^ n4600 ^ n2712 ;
  assign n8174 = x11 & n1263 ;
  assign n8175 = n8174 ^ n4180 ^ 1'b0 ;
  assign n8176 = n8175 ^ n2404 ^ x89 ;
  assign n8177 = ( ~n933 & n996 ) | ( ~n933 & n8176 ) | ( n996 & n8176 ) ;
  assign n8180 = n8179 ^ n8177 ^ n3177 ;
  assign n8181 = ( ~n3399 & n7837 ) | ( ~n3399 & n8180 ) | ( n7837 & n8180 ) ;
  assign n8183 = n8182 ^ n8181 ^ n4378 ;
  assign n8184 = ( n828 & ~n1110 ) | ( n828 & n1431 ) | ( ~n1110 & n1431 ) ;
  assign n8185 = n8184 ^ n3598 ^ 1'b0 ;
  assign n8186 = ~n1991 & n8185 ;
  assign n8187 = n3893 & n4822 ;
  assign n8188 = ~n8186 & n8187 ;
  assign n8189 = ( ~n1434 & n6866 ) | ( ~n1434 & n8188 ) | ( n6866 & n8188 ) ;
  assign n8190 = n7746 ^ n4612 ^ n1637 ;
  assign n8191 = n3784 ^ n2418 ^ n418 ;
  assign n8192 = ~n536 & n8191 ;
  assign n8193 = n8192 ^ x131 ^ 1'b0 ;
  assign n8194 = n1161 | n8193 ;
  assign n8195 = n1445 & n8194 ;
  assign n8196 = n5083 & n8195 ;
  assign n8204 = n1255 ^ n859 ^ n348 ;
  assign n8205 = ~n3133 & n8204 ;
  assign n8200 = n622 & ~n6266 ;
  assign n8201 = ~n2316 & n8200 ;
  assign n8202 = n8201 ^ n6827 ^ n869 ;
  assign n8203 = ( n877 & n993 ) | ( n877 & n8202 ) | ( n993 & n8202 ) ;
  assign n8199 = n6763 ^ n6062 ^ n1301 ;
  assign n8206 = n8205 ^ n8203 ^ n8199 ;
  assign n8197 = ( ~n1481 & n2516 ) | ( ~n1481 & n7994 ) | ( n2516 & n7994 ) ;
  assign n8198 = n784 & ~n8197 ;
  assign n8207 = n8206 ^ n8198 ^ 1'b0 ;
  assign n8210 = n4105 ^ n1511 ^ 1'b0 ;
  assign n8211 = n8210 ^ n5169 ^ 1'b0 ;
  assign n8208 = n1907 | n5736 ;
  assign n8209 = n8208 ^ n4026 ^ 1'b0 ;
  assign n8212 = n8211 ^ n8209 ^ n2646 ;
  assign n8222 = n5146 ^ n2859 ^ n518 ;
  assign n8213 = ( n2192 & ~n2196 ) | ( n2192 & n2483 ) | ( ~n2196 & n2483 ) ;
  assign n8214 = ( n1840 & n2912 ) | ( n1840 & n8213 ) | ( n2912 & n8213 ) ;
  assign n8215 = n8214 ^ n818 ^ n548 ;
  assign n8216 = ( ~n680 & n4573 ) | ( ~n680 & n8215 ) | ( n4573 & n8215 ) ;
  assign n8217 = ~n2179 & n6613 ;
  assign n8218 = n8217 ^ n6103 ^ 1'b0 ;
  assign n8219 = ( n974 & n1800 ) | ( n974 & n7556 ) | ( n1800 & n7556 ) ;
  assign n8220 = n8219 ^ n6072 ^ n1822 ;
  assign n8221 = ( ~n8216 & n8218 ) | ( ~n8216 & n8220 ) | ( n8218 & n8220 ) ;
  assign n8223 = n8222 ^ n8221 ^ n518 ;
  assign n8224 = n5000 ^ x136 ^ 1'b0 ;
  assign n8231 = n670 & n4785 ;
  assign n8232 = n2973 & n8231 ;
  assign n8233 = ( x250 & ~n3798 ) | ( x250 & n8232 ) | ( ~n3798 & n8232 ) ;
  assign n8225 = n2117 ^ n1428 ^ n299 ;
  assign n8226 = n2027 & n4476 ;
  assign n8227 = ( ~n2194 & n2350 ) | ( ~n2194 & n8226 ) | ( n2350 & n8226 ) ;
  assign n8228 = ( n2348 & n8225 ) | ( n2348 & n8227 ) | ( n8225 & n8227 ) ;
  assign n8229 = n8228 ^ n2848 ^ n1552 ;
  assign n8230 = ( ~n1707 & n3554 ) | ( ~n1707 & n8229 ) | ( n3554 & n8229 ) ;
  assign n8234 = n8233 ^ n8230 ^ n5393 ;
  assign n8235 = ~n6958 & n8234 ;
  assign n8236 = n8235 ^ n4679 ^ 1'b0 ;
  assign n8242 = n962 & n3153 ;
  assign n8243 = n8242 ^ n2671 ^ x24 ;
  assign n8239 = n3545 ^ n1074 ^ x1 ;
  assign n8240 = n8239 ^ n1533 ^ 1'b0 ;
  assign n8241 = n8240 ^ n2294 ^ x14 ;
  assign n8244 = n8243 ^ n8241 ^ n3142 ;
  assign n8237 = ( x109 & ~n2374 ) | ( x109 & n2546 ) | ( ~n2374 & n2546 ) ;
  assign n8238 = n6837 & ~n8237 ;
  assign n8245 = n8244 ^ n8238 ^ n1325 ;
  assign n8246 = n8245 ^ n4574 ^ n4070 ;
  assign n8247 = n7781 ^ n3057 ^ n1153 ;
  assign n8249 = n1904 ^ n1785 ^ x184 ;
  assign n8248 = n1858 & n7101 ;
  assign n8250 = n8249 ^ n8248 ^ 1'b0 ;
  assign n8251 = n8247 | n8250 ;
  assign n8252 = ( x237 & ~n4318 ) | ( x237 & n8179 ) | ( ~n4318 & n8179 ) ;
  assign n8253 = n1610 ^ x43 ^ 1'b0 ;
  assign n8254 = n8252 & n8253 ;
  assign n8255 = ( n581 & ~n1483 ) | ( n581 & n8254 ) | ( ~n1483 & n8254 ) ;
  assign n8258 = n2090 & ~n4502 ;
  assign n8259 = ( n3137 & n4731 ) | ( n3137 & ~n8258 ) | ( n4731 & ~n8258 ) ;
  assign n8256 = n6948 ^ n4504 ^ n1473 ;
  assign n8257 = n1143 | n8256 ;
  assign n8260 = n8259 ^ n8257 ^ 1'b0 ;
  assign n8261 = ( n8251 & n8255 ) | ( n8251 & ~n8260 ) | ( n8255 & ~n8260 ) ;
  assign n8262 = n4900 ^ n4371 ^ 1'b0 ;
  assign n8263 = n2860 ^ n1951 ^ x110 ;
  assign n8264 = n8263 ^ n2677 ^ 1'b0 ;
  assign n8265 = n8264 ^ n4378 ^ 1'b0 ;
  assign n8266 = n8262 & ~n8265 ;
  assign n8270 = n420 & ~n5255 ;
  assign n8267 = n720 ^ n604 ^ 1'b0 ;
  assign n8268 = n8267 ^ n6108 ^ n3034 ;
  assign n8269 = n8268 ^ n7248 ^ n3994 ;
  assign n8271 = n8270 ^ n8269 ^ n2307 ;
  assign n8272 = ( n906 & n4509 ) | ( n906 & ~n6121 ) | ( n4509 & ~n6121 ) ;
  assign n8273 = n8272 ^ n2348 ^ 1'b0 ;
  assign n8274 = n8025 & ~n8273 ;
  assign n8275 = ~n2816 & n8274 ;
  assign n8276 = ~n8271 & n8275 ;
  assign n8278 = ( n778 & n4135 ) | ( n778 & n7713 ) | ( n4135 & n7713 ) ;
  assign n8279 = n8278 ^ n3657 ^ n1935 ;
  assign n8280 = ~n588 & n1293 ;
  assign n8281 = n8280 ^ n982 ^ 1'b0 ;
  assign n8282 = ( ~n2723 & n6943 ) | ( ~n2723 & n8281 ) | ( n6943 & n8281 ) ;
  assign n8283 = ( ~x131 & n8279 ) | ( ~x131 & n8282 ) | ( n8279 & n8282 ) ;
  assign n8277 = n875 & n5043 ;
  assign n8284 = n8283 ^ n8277 ^ 1'b0 ;
  assign n8287 = n1890 & n4977 ;
  assign n8288 = n3277 & n8287 ;
  assign n8289 = n8288 ^ n1422 ^ x113 ;
  assign n8285 = ( ~n2528 & n3060 ) | ( ~n2528 & n5472 ) | ( n3060 & n5472 ) ;
  assign n8286 = n8285 ^ n5048 ^ n4752 ;
  assign n8290 = n8289 ^ n8286 ^ n7571 ;
  assign n8291 = n8290 ^ n7294 ^ 1'b0 ;
  assign n8292 = x141 & n5284 ;
  assign n8293 = n4163 ^ x119 ^ x111 ;
  assign n8294 = ( x122 & n579 ) | ( x122 & ~n8293 ) | ( n579 & ~n8293 ) ;
  assign n8295 = ( ~n1123 & n1278 ) | ( ~n1123 & n8294 ) | ( n1278 & n8294 ) ;
  assign n8296 = n8295 ^ n4647 ^ 1'b0 ;
  assign n8297 = ( ~n3771 & n5676 ) | ( ~n3771 & n8296 ) | ( n5676 & n8296 ) ;
  assign n8298 = ( ~n1451 & n5648 ) | ( ~n1451 & n8297 ) | ( n5648 & n8297 ) ;
  assign n8299 = ( n1435 & n3779 ) | ( n1435 & n6303 ) | ( n3779 & n6303 ) ;
  assign n8300 = n567 ^ n348 ^ 1'b0 ;
  assign n8301 = n8299 | n8300 ;
  assign n8302 = n8301 ^ n5793 ^ 1'b0 ;
  assign n8303 = n8302 ^ n2023 ^ n564 ;
  assign n8304 = ~n5678 & n8303 ;
  assign n8305 = n5201 ^ n2841 ^ 1'b0 ;
  assign n8306 = n8204 ^ n2478 ^ 1'b0 ;
  assign n8307 = n8305 | n8306 ;
  assign n8308 = ( n2765 & ~n3370 ) | ( n2765 & n6376 ) | ( ~n3370 & n6376 ) ;
  assign n8309 = ( ~n2271 & n4434 ) | ( ~n2271 & n6779 ) | ( n4434 & n6779 ) ;
  assign n8310 = ( ~n3061 & n4443 ) | ( ~n3061 & n8309 ) | ( n4443 & n8309 ) ;
  assign n8311 = ~n3504 & n8310 ;
  assign n8312 = n707 & n8311 ;
  assign n8313 = n8308 & ~n8312 ;
  assign n8314 = n7180 ^ n1476 ^ 1'b0 ;
  assign n8319 = ( n797 & n5770 ) | ( n797 & n6390 ) | ( n5770 & n6390 ) ;
  assign n8315 = n4783 ^ n2396 ^ n282 ;
  assign n8316 = n8315 ^ n2399 ^ n384 ;
  assign n8317 = n8316 ^ x166 ^ 1'b0 ;
  assign n8318 = ( n2921 & n6856 ) | ( n2921 & n8317 ) | ( n6856 & n8317 ) ;
  assign n8320 = n8319 ^ n8318 ^ n6439 ;
  assign n8321 = n3316 & ~n5012 ;
  assign n8322 = ~n2335 & n8321 ;
  assign n8323 = ( ~n667 & n8320 ) | ( ~n667 & n8322 ) | ( n8320 & n8322 ) ;
  assign n8325 = n7058 ^ n5797 ^ n2887 ;
  assign n8326 = ( n2096 & ~n2159 ) | ( n2096 & n6763 ) | ( ~n2159 & n6763 ) ;
  assign n8327 = n7220 & n8326 ;
  assign n8328 = ~n8325 & n8327 ;
  assign n8324 = n1359 | n6237 ;
  assign n8329 = n8328 ^ n8324 ^ n2026 ;
  assign n8335 = n979 ^ n373 ^ 1'b0 ;
  assign n8336 = x19 & n8335 ;
  assign n8330 = n6212 ^ n3324 ^ n486 ;
  assign n8331 = n8330 ^ n1207 ^ 1'b0 ;
  assign n8332 = n7260 & ~n8331 ;
  assign n8333 = n4798 ^ n3363 ^ n739 ;
  assign n8334 = ( n6979 & ~n8332 ) | ( n6979 & n8333 ) | ( ~n8332 & n8333 ) ;
  assign n8337 = n8336 ^ n8334 ^ n5962 ;
  assign n8344 = ( ~n1356 & n2528 ) | ( ~n1356 & n4176 ) | ( n2528 & n4176 ) ;
  assign n8341 = n7352 ^ n3945 ^ n3753 ;
  assign n8338 = n6506 ^ n2107 ^ n1894 ;
  assign n8339 = ( ~n3681 & n3939 ) | ( ~n3681 & n4090 ) | ( n3939 & n4090 ) ;
  assign n8340 = ( n3495 & ~n8338 ) | ( n3495 & n8339 ) | ( ~n8338 & n8339 ) ;
  assign n8342 = n8341 ^ n8340 ^ n5394 ;
  assign n8343 = n8342 ^ n8252 ^ n2048 ;
  assign n8345 = n8344 ^ n8343 ^ n1056 ;
  assign n8347 = x26 & x36 ;
  assign n8348 = ~n904 & n8347 ;
  assign n8349 = n3255 ^ n1697 ^ 1'b0 ;
  assign n8350 = n8348 | n8349 ;
  assign n8351 = n8350 ^ n396 ^ 1'b0 ;
  assign n8352 = n1411 & n8351 ;
  assign n8346 = ( n271 & ~n959 ) | ( n271 & n7137 ) | ( ~n959 & n7137 ) ;
  assign n8353 = n8352 ^ n8346 ^ 1'b0 ;
  assign n8354 = ( ~n1739 & n2206 ) | ( ~n1739 & n6540 ) | ( n2206 & n6540 ) ;
  assign n8355 = n3361 ^ n2527 ^ n1532 ;
  assign n8356 = n8035 ^ n5472 ^ n4572 ;
  assign n8357 = n8356 ^ n3376 ^ n1790 ;
  assign n8358 = n8087 ^ n3367 ^ n2117 ;
  assign n8359 = ( n1177 & ~n5834 ) | ( n1177 & n8358 ) | ( ~n5834 & n8358 ) ;
  assign n8360 = ( ~n8355 & n8357 ) | ( ~n8355 & n8359 ) | ( n8357 & n8359 ) ;
  assign n8363 = x24 & n2899 ;
  assign n8364 = n707 & n8363 ;
  assign n8365 = n2425 ^ n2103 ^ x60 ;
  assign n8366 = ( n7139 & ~n8364 ) | ( n7139 & n8365 ) | ( ~n8364 & n8365 ) ;
  assign n8361 = n3105 & ~n3473 ;
  assign n8362 = n2091 & n8361 ;
  assign n8367 = n8366 ^ n8362 ^ n6223 ;
  assign n8369 = ( n975 & n2133 ) | ( n975 & n2647 ) | ( n2133 & n2647 ) ;
  assign n8368 = n7918 ^ n4619 ^ n1136 ;
  assign n8370 = n8369 ^ n8368 ^ n6642 ;
  assign n8374 = ( n3361 & n7118 ) | ( n3361 & n8115 ) | ( n7118 & n8115 ) ;
  assign n8371 = n1960 | n7909 ;
  assign n8372 = n8371 ^ n6294 ^ 1'b0 ;
  assign n8373 = n6814 | n8372 ;
  assign n8375 = n8374 ^ n8373 ^ 1'b0 ;
  assign n8376 = n2956 | n3154 ;
  assign n8377 = ( n288 & ~n6002 ) | ( n288 & n8376 ) | ( ~n6002 & n8376 ) ;
  assign n8378 = n1730 ^ n1700 ^ 1'b0 ;
  assign n8379 = n5151 ^ n2714 ^ 1'b0 ;
  assign n8380 = ( n2339 & ~n8378 ) | ( n2339 & n8379 ) | ( ~n8378 & n8379 ) ;
  assign n8381 = ( n1395 & n1924 ) | ( n1395 & ~n7905 ) | ( n1924 & ~n7905 ) ;
  assign n8382 = ~n2191 & n5149 ;
  assign n8383 = n8381 | n8382 ;
  assign n8384 = ( x167 & n2180 ) | ( x167 & n7933 ) | ( n2180 & n7933 ) ;
  assign n8385 = n8384 ^ n7118 ^ 1'b0 ;
  assign n8386 = n4693 & n8385 ;
  assign n8387 = n4531 ^ n2627 ^ n716 ;
  assign n8388 = n2535 & n8387 ;
  assign n8389 = ( n5644 & ~n7122 ) | ( n5644 & n8388 ) | ( ~n7122 & n8388 ) ;
  assign n8390 = ( n8383 & ~n8386 ) | ( n8383 & n8389 ) | ( ~n8386 & n8389 ) ;
  assign n8393 = ( ~n993 & n1568 ) | ( ~n993 & n2864 ) | ( n1568 & n2864 ) ;
  assign n8394 = n8393 ^ n5719 ^ n258 ;
  assign n8395 = ( n1928 & n2082 ) | ( n1928 & n3353 ) | ( n2082 & n3353 ) ;
  assign n8396 = ( n654 & n5961 ) | ( n654 & n8395 ) | ( n5961 & n8395 ) ;
  assign n8397 = ( ~n5187 & n8394 ) | ( ~n5187 & n8396 ) | ( n8394 & n8396 ) ;
  assign n8391 = ( n2824 & n3797 ) | ( n2824 & n3856 ) | ( n3797 & n3856 ) ;
  assign n8392 = n3402 & n8391 ;
  assign n8398 = n8397 ^ n8392 ^ 1'b0 ;
  assign n8404 = ( n1749 & ~n3963 ) | ( n1749 & n5446 ) | ( ~n3963 & n5446 ) ;
  assign n8403 = n5355 & ~n6775 ;
  assign n8405 = n8404 ^ n8403 ^ 1'b0 ;
  assign n8399 = n5034 ^ n3146 ^ n1696 ;
  assign n8400 = n1446 & ~n8399 ;
  assign n8401 = n4662 ^ n3860 ^ 1'b0 ;
  assign n8402 = ( ~n1780 & n8400 ) | ( ~n1780 & n8401 ) | ( n8400 & n8401 ) ;
  assign n8406 = n8405 ^ n8402 ^ n5593 ;
  assign n8407 = n6196 ^ n5794 ^ 1'b0 ;
  assign n8408 = ( n2414 & n5997 ) | ( n2414 & n7433 ) | ( n5997 & n7433 ) ;
  assign n8409 = n1656 & n2113 ;
  assign n8410 = ( n1253 & n3599 ) | ( n1253 & ~n6991 ) | ( n3599 & ~n6991 ) ;
  assign n8411 = ( n669 & ~n7052 ) | ( n669 & n8410 ) | ( ~n7052 & n8410 ) ;
  assign n8412 = n6500 ^ n5082 ^ n1896 ;
  assign n8413 = ( n328 & n4954 ) | ( n328 & n5367 ) | ( n4954 & n5367 ) ;
  assign n8414 = n8093 ^ n6435 ^ 1'b0 ;
  assign n8415 = ( n8412 & ~n8413 ) | ( n8412 & n8414 ) | ( ~n8413 & n8414 ) ;
  assign n8416 = n5471 ^ n4312 ^ 1'b0 ;
  assign n8417 = n1108 | n8416 ;
  assign n8418 = n8417 ^ n995 ^ 1'b0 ;
  assign n8419 = n4327 ^ n1008 ^ n870 ;
  assign n8420 = n4540 & n8419 ;
  assign n8421 = ~n1416 & n8420 ;
  assign n8422 = n6157 ^ n3400 ^ 1'b0 ;
  assign n8423 = n8422 ^ n8169 ^ n4725 ;
  assign n8424 = n2938 ^ n2755 ^ 1'b0 ;
  assign n8425 = n3543 & n8424 ;
  assign n8426 = n8425 ^ n5983 ^ n1989 ;
  assign n8427 = n846 ^ n406 ^ n375 ;
  assign n8428 = n636 & n4889 ;
  assign n8429 = n8428 ^ n3176 ^ n553 ;
  assign n8430 = ( n8426 & n8427 ) | ( n8426 & ~n8429 ) | ( n8427 & ~n8429 ) ;
  assign n8434 = ( x135 & ~n1056 ) | ( x135 & n3927 ) | ( ~n1056 & n3927 ) ;
  assign n8435 = n6290 & ~n6530 ;
  assign n8436 = n8435 ^ n2403 ^ 1'b0 ;
  assign n8439 = n3495 ^ n1474 ^ n631 ;
  assign n8440 = n8439 ^ n1831 ^ n642 ;
  assign n8437 = n2910 ^ n2676 ^ 1'b0 ;
  assign n8438 = ~n1414 & n8437 ;
  assign n8441 = n8440 ^ n8438 ^ 1'b0 ;
  assign n8442 = ( ~n3177 & n8436 ) | ( ~n3177 & n8441 ) | ( n8436 & n8441 ) ;
  assign n8443 = n8442 ^ n1811 ^ 1'b0 ;
  assign n8444 = ~n8434 & n8443 ;
  assign n8431 = x236 & ~n399 ;
  assign n8432 = n8431 ^ n4238 ^ n3281 ;
  assign n8433 = ( n4406 & n5587 ) | ( n4406 & ~n8432 ) | ( n5587 & ~n8432 ) ;
  assign n8445 = n8444 ^ n8433 ^ n4310 ;
  assign n8446 = ~n1205 & n4352 ;
  assign n8447 = ~n523 & n8446 ;
  assign n8448 = ( x175 & ~n4142 ) | ( x175 & n8447 ) | ( ~n4142 & n8447 ) ;
  assign n8449 = ( ~n8430 & n8445 ) | ( ~n8430 & n8448 ) | ( n8445 & n8448 ) ;
  assign n8451 = n5822 ^ n2384 ^ n871 ;
  assign n8450 = n4526 ^ n477 ^ 1'b0 ;
  assign n8452 = n8451 ^ n8450 ^ n1159 ;
  assign n8453 = ( ~n328 & n4366 ) | ( ~n328 & n8452 ) | ( n4366 & n8452 ) ;
  assign n8454 = ( n2097 & ~n2240 ) | ( n2097 & n4653 ) | ( ~n2240 & n4653 ) ;
  assign n8459 = n545 | n1290 ;
  assign n8457 = n4948 ^ n870 ^ n678 ;
  assign n8458 = n8457 ^ n2035 ^ x83 ;
  assign n8455 = n7887 ^ n5950 ^ n797 ;
  assign n8456 = n1525 & ~n8455 ;
  assign n8460 = n8459 ^ n8458 ^ n8456 ;
  assign n8470 = ( ~n387 & n3422 ) | ( ~n387 & n5706 ) | ( n3422 & n5706 ) ;
  assign n8471 = ( x207 & n3852 ) | ( x207 & ~n8002 ) | ( n3852 & ~n8002 ) ;
  assign n8472 = ( ~n1294 & n8470 ) | ( ~n1294 & n8471 ) | ( n8470 & n8471 ) ;
  assign n8469 = n5142 & n5938 ;
  assign n8473 = n8472 ^ n8469 ^ 1'b0 ;
  assign n8474 = ~n1577 & n8473 ;
  assign n8475 = n660 & n8474 ;
  assign n8461 = n7654 ^ n4763 ^ n4692 ;
  assign n8462 = n5887 ^ n2034 ^ x169 ;
  assign n8463 = ( n901 & n8461 ) | ( n901 & ~n8462 ) | ( n8461 & ~n8462 ) ;
  assign n8464 = ( n2049 & n2993 ) | ( n2049 & ~n5849 ) | ( n2993 & ~n5849 ) ;
  assign n8465 = n6090 & n8464 ;
  assign n8466 = n8465 ^ n2863 ^ 1'b0 ;
  assign n8467 = n8466 ^ n1970 ^ 1'b0 ;
  assign n8468 = ( n2038 & ~n8463 ) | ( n2038 & n8467 ) | ( ~n8463 & n8467 ) ;
  assign n8476 = n8475 ^ n8468 ^ n5898 ;
  assign n8477 = n5583 ^ n2983 ^ n2378 ;
  assign n8478 = ( x208 & n6285 ) | ( x208 & n8477 ) | ( n6285 & n8477 ) ;
  assign n8479 = ( ~n3639 & n3768 ) | ( ~n3639 & n6811 ) | ( n3768 & n6811 ) ;
  assign n8480 = n8323 ^ n7940 ^ 1'b0 ;
  assign n8481 = n8479 | n8480 ;
  assign n8487 = n8081 ^ n5304 ^ 1'b0 ;
  assign n8488 = n8383 ^ n7330 ^ 1'b0 ;
  assign n8489 = ~n8487 & n8488 ;
  assign n8484 = n6052 ^ n2601 ^ n1991 ;
  assign n8483 = n2604 ^ n1715 ^ 1'b0 ;
  assign n8485 = n8484 ^ n8483 ^ n1675 ;
  assign n8482 = ( ~n1952 & n2459 ) | ( ~n1952 & n6830 ) | ( n2459 & n6830 ) ;
  assign n8486 = n8485 ^ n8482 ^ n3365 ;
  assign n8490 = n8489 ^ n8486 ^ n1629 ;
  assign n8491 = n7095 ^ n3401 ^ n3116 ;
  assign n8492 = n6042 ^ n812 ^ n471 ;
  assign n8493 = n642 | n8492 ;
  assign n8494 = n8493 ^ n2664 ^ n1595 ;
  assign n8495 = ~n4783 & n8494 ;
  assign n8496 = n8491 & n8495 ;
  assign n8497 = ( ~n547 & n938 ) | ( ~n547 & n1428 ) | ( n938 & n1428 ) ;
  assign n8498 = n8497 ^ n6654 ^ 1'b0 ;
  assign n8499 = ( n2965 & ~n4357 ) | ( n2965 & n4806 ) | ( ~n4357 & n4806 ) ;
  assign n8500 = n8389 ^ n4010 ^ 1'b0 ;
  assign n8508 = n938 | n1963 ;
  assign n8509 = n8508 ^ x58 ^ 1'b0 ;
  assign n8503 = n3929 ^ n287 ^ 1'b0 ;
  assign n8501 = ( n1404 & n2858 ) | ( n1404 & ~n5285 ) | ( n2858 & ~n5285 ) ;
  assign n8502 = ( n3272 & n7842 ) | ( n3272 & n8501 ) | ( n7842 & n8501 ) ;
  assign n8504 = n8503 ^ n8502 ^ 1'b0 ;
  assign n8505 = ( n3972 & ~n6165 ) | ( n3972 & n7304 ) | ( ~n6165 & n7304 ) ;
  assign n8506 = n3434 & n4437 ;
  assign n8507 = ( n8504 & n8505 ) | ( n8504 & n8506 ) | ( n8505 & n8506 ) ;
  assign n8510 = n8509 ^ n8507 ^ 1'b0 ;
  assign n8511 = n6412 ^ n5216 ^ n2660 ;
  assign n8512 = n5316 ^ x10 ^ 1'b0 ;
  assign n8513 = ( n8325 & ~n8511 ) | ( n8325 & n8512 ) | ( ~n8511 & n8512 ) ;
  assign n8514 = ~n316 & n7542 ;
  assign n8515 = n3791 & n8514 ;
  assign n8516 = n5152 ^ n5013 ^ n544 ;
  assign n8517 = ( n535 & ~n3106 ) | ( n535 & n7165 ) | ( ~n3106 & n7165 ) ;
  assign n8518 = ~n8516 & n8517 ;
  assign n8519 = ~n7294 & n8518 ;
  assign n8520 = n1871 & ~n8519 ;
  assign n8521 = ~n3294 & n8520 ;
  assign n8522 = n8521 ^ n3096 ^ n623 ;
  assign n8523 = n5103 ^ n4651 ^ 1'b0 ;
  assign n8524 = n3741 & ~n8523 ;
  assign n8525 = n7324 & n8524 ;
  assign n8530 = ~n1782 & n3418 ;
  assign n8526 = ( n3422 & n4434 ) | ( n3422 & n7385 ) | ( n4434 & n7385 ) ;
  assign n8527 = n7418 ^ n5367 ^ n998 ;
  assign n8528 = ( ~n3971 & n4809 ) | ( ~n3971 & n8527 ) | ( n4809 & n8527 ) ;
  assign n8529 = ( ~n839 & n8526 ) | ( ~n839 & n8528 ) | ( n8526 & n8528 ) ;
  assign n8531 = n8530 ^ n8529 ^ n7457 ;
  assign n8532 = n6154 ^ n801 ^ 1'b0 ;
  assign n8533 = n3950 & n8532 ;
  assign n8534 = n8533 ^ n6610 ^ n4901 ;
  assign n8535 = n8534 ^ n2165 ^ 1'b0 ;
  assign n8536 = n1405 & n8535 ;
  assign n8537 = n5306 ^ n2457 ^ n1264 ;
  assign n8538 = ( ~n1112 & n6831 ) | ( ~n1112 & n8537 ) | ( n6831 & n8537 ) ;
  assign n8539 = n8538 ^ n6766 ^ n818 ;
  assign n8545 = n3633 ^ n2623 ^ n1393 ;
  assign n8540 = ~n1379 & n1842 ;
  assign n8541 = n2303 & n8540 ;
  assign n8542 = n4714 ^ n3275 ^ n623 ;
  assign n8543 = ( n2415 & ~n3855 ) | ( n2415 & n8542 ) | ( ~n3855 & n8542 ) ;
  assign n8544 = ~n8541 & n8543 ;
  assign n8546 = n8545 ^ n8544 ^ 1'b0 ;
  assign n8547 = n8546 ^ n7638 ^ n3664 ;
  assign n8548 = ( n3365 & ~n7843 ) | ( n3365 & n7910 ) | ( ~n7843 & n7910 ) ;
  assign n8549 = ( n3097 & n7884 ) | ( n3097 & n7923 ) | ( n7884 & n7923 ) ;
  assign n8550 = ( n838 & n1166 ) | ( n838 & ~n2902 ) | ( n1166 & ~n2902 ) ;
  assign n8551 = n8550 ^ n7182 ^ n1429 ;
  assign n8552 = n8551 ^ x174 ^ 1'b0 ;
  assign n8553 = n5852 & ~n8552 ;
  assign n8554 = ( x86 & n1056 ) | ( x86 & ~n8553 ) | ( n1056 & ~n8553 ) ;
  assign n8555 = ( n1641 & ~n3354 ) | ( n1641 & n4714 ) | ( ~n3354 & n4714 ) ;
  assign n8556 = n8555 ^ n1198 ^ 1'b0 ;
  assign n8557 = n8554 & n8556 ;
  assign n8558 = ( n6781 & n6816 ) | ( n6781 & ~n8557 ) | ( n6816 & ~n8557 ) ;
  assign n8559 = n3866 ^ n2860 ^ n1629 ;
  assign n8560 = n7787 ^ n4823 ^ 1'b0 ;
  assign n8561 = n8559 & n8560 ;
  assign n8562 = n8561 ^ n7102 ^ n459 ;
  assign n8563 = ( n312 & ~n518 ) | ( n312 & n746 ) | ( ~n518 & n746 ) ;
  assign n8564 = n3213 ^ n1544 ^ n987 ;
  assign n8565 = n5603 ^ n3860 ^ n533 ;
  assign n8566 = ( ~n3277 & n8564 ) | ( ~n3277 & n8565 ) | ( n8564 & n8565 ) ;
  assign n8567 = ( ~n566 & n8563 ) | ( ~n566 & n8566 ) | ( n8563 & n8566 ) ;
  assign n8568 = x91 & x104 ;
  assign n8569 = ~x199 & n8568 ;
  assign n8570 = n8569 ^ n3177 ^ 1'b0 ;
  assign n8571 = ( n2459 & n4002 ) | ( n2459 & n4694 ) | ( n4002 & n4694 ) ;
  assign n8572 = n1387 & ~n4222 ;
  assign n8573 = n8571 & n8572 ;
  assign n8574 = ~n7994 & n8573 ;
  assign n8575 = ( ~n891 & n1973 ) | ( ~n891 & n4915 ) | ( n1973 & n4915 ) ;
  assign n8576 = n8081 ^ n7803 ^ 1'b0 ;
  assign n8577 = ~n2080 & n8576 ;
  assign n8578 = ( n6033 & n8575 ) | ( n6033 & n8577 ) | ( n8575 & n8577 ) ;
  assign n8579 = n6660 ^ n4131 ^ n2462 ;
  assign n8580 = ( n1646 & n2040 ) | ( n1646 & n6937 ) | ( n2040 & n6937 ) ;
  assign n8581 = ( n336 & ~n426 ) | ( n336 & n5463 ) | ( ~n426 & n5463 ) ;
  assign n8582 = ( n3453 & n7503 ) | ( n3453 & n8581 ) | ( n7503 & n8581 ) ;
  assign n8583 = n8582 ^ n5238 ^ 1'b0 ;
  assign n8584 = ~n8580 & n8583 ;
  assign n8585 = n8137 ^ n5902 ^ n1399 ;
  assign n8586 = n4563 ^ n3731 ^ n1956 ;
  assign n8587 = n8585 & n8586 ;
  assign n8588 = n8587 ^ n3814 ^ 1'b0 ;
  assign n8589 = ( ~n3315 & n8025 ) | ( ~n3315 & n8588 ) | ( n8025 & n8588 ) ;
  assign n8590 = ( n2523 & n2718 ) | ( n2523 & ~n3376 ) | ( n2718 & ~n3376 ) ;
  assign n8591 = ( x181 & ~n2295 ) | ( x181 & n8590 ) | ( ~n2295 & n8590 ) ;
  assign n8592 = n1233 & n8591 ;
  assign n8593 = n2555 & n8592 ;
  assign n8594 = n8593 ^ n5740 ^ n629 ;
  assign n8595 = n6287 ^ n2658 ^ 1'b0 ;
  assign n8596 = ( n5160 & n8149 ) | ( n5160 & ~n8595 ) | ( n8149 & ~n8595 ) ;
  assign n8597 = ( n3242 & n8584 ) | ( n3242 & ~n8596 ) | ( n8584 & ~n8596 ) ;
  assign n8598 = n6473 | n7780 ;
  assign n8599 = n2970 ^ n2180 ^ 1'b0 ;
  assign n8600 = n8599 ^ n4633 ^ 1'b0 ;
  assign n8601 = ( n2406 & n7016 ) | ( n2406 & n8600 ) | ( n7016 & n8600 ) ;
  assign n8615 = ( n995 & ~n2326 ) | ( n995 & n4020 ) | ( ~n2326 & n4020 ) ;
  assign n8602 = n437 & ~n1042 ;
  assign n8603 = n7715 & n8602 ;
  assign n8604 = ( n4941 & n5822 ) | ( n4941 & ~n8603 ) | ( n5822 & ~n8603 ) ;
  assign n8605 = n4062 ^ n661 ^ x225 ;
  assign n8606 = ~n3563 & n8605 ;
  assign n8607 = n7456 ^ n3060 ^ n305 ;
  assign n8608 = ( n4988 & n8606 ) | ( n4988 & n8607 ) | ( n8606 & n8607 ) ;
  assign n8609 = ( n5398 & n8604 ) | ( n5398 & n8608 ) | ( n8604 & n8608 ) ;
  assign n8610 = ( n1529 & n7130 ) | ( n1529 & n8609 ) | ( n7130 & n8609 ) ;
  assign n8611 = n3026 ^ n2957 ^ n2679 ;
  assign n8612 = n7053 ^ n4424 ^ 1'b0 ;
  assign n8613 = ( n678 & n8611 ) | ( n678 & ~n8612 ) | ( n8611 & ~n8612 ) ;
  assign n8614 = n8610 | n8613 ;
  assign n8616 = n8615 ^ n8614 ^ 1'b0 ;
  assign n8617 = n1511 ^ n1116 ^ n665 ;
  assign n8618 = ( ~n3182 & n5253 ) | ( ~n3182 & n8617 ) | ( n5253 & n8617 ) ;
  assign n8619 = n8618 ^ n4051 ^ n639 ;
  assign n8620 = ( n2200 & n2723 ) | ( n2200 & ~n4625 ) | ( n2723 & ~n4625 ) ;
  assign n8621 = n2389 | n8620 ;
  assign n8622 = n8619 | n8621 ;
  assign n8626 = n4585 ^ n2787 ^ n1015 ;
  assign n8623 = n2135 | n2391 ;
  assign n8624 = n6833 | n8623 ;
  assign n8625 = ~n7059 & n8624 ;
  assign n8627 = n8626 ^ n8625 ^ 1'b0 ;
  assign n8628 = ( ~n1044 & n2122 ) | ( ~n1044 & n2583 ) | ( n2122 & n2583 ) ;
  assign n8629 = ( n4299 & n5344 ) | ( n4299 & n7282 ) | ( n5344 & n7282 ) ;
  assign n8630 = x61 & ~n8629 ;
  assign n8631 = n8630 ^ n2784 ^ 1'b0 ;
  assign n8632 = ( n5191 & n8628 ) | ( n5191 & ~n8631 ) | ( n8628 & ~n8631 ) ;
  assign n8633 = n4833 ^ n3492 ^ n3088 ;
  assign n8634 = n4375 ^ n1389 ^ 1'b0 ;
  assign n8635 = ( n2405 & n8633 ) | ( n2405 & ~n8634 ) | ( n8633 & ~n8634 ) ;
  assign n8636 = ( n1583 & ~n4978 ) | ( n1583 & n5417 ) | ( ~n4978 & n5417 ) ;
  assign n8637 = ( n1713 & n6297 ) | ( n1713 & ~n8636 ) | ( n6297 & ~n8636 ) ;
  assign n8638 = ( n3844 & n5432 ) | ( n3844 & n8637 ) | ( n5432 & n8637 ) ;
  assign n8639 = ( n4764 & n8635 ) | ( n4764 & n8638 ) | ( n8635 & n8638 ) ;
  assign n8640 = n389 | n3088 ;
  assign n8641 = n2618 | n8640 ;
  assign n8642 = n1662 & ~n8641 ;
  assign n8643 = n4282 ^ x251 ^ 1'b0 ;
  assign n8644 = n8642 | n8643 ;
  assign n8647 = ( n3073 & n3225 ) | ( n3073 & ~n4742 ) | ( n3225 & ~n4742 ) ;
  assign n8645 = n3869 & ~n6721 ;
  assign n8646 = n7557 & n8645 ;
  assign n8648 = n8647 ^ n8646 ^ n606 ;
  assign n8649 = n8648 ^ n2258 ^ 1'b0 ;
  assign n8650 = ~x143 & n8649 ;
  assign n8654 = n3350 ^ n1475 ^ 1'b0 ;
  assign n8655 = n2322 & n8654 ;
  assign n8651 = ( n654 & ~n7915 ) | ( n654 & n8293 ) | ( ~n7915 & n8293 ) ;
  assign n8652 = n8651 ^ n1942 ^ n1836 ;
  assign n8653 = n8652 ^ n3019 ^ n1043 ;
  assign n8656 = n8655 ^ n8653 ^ n2191 ;
  assign n8657 = n6559 ^ x165 ^ 1'b0 ;
  assign n8658 = n8657 ^ n7950 ^ n2662 ;
  assign n8659 = n6668 | n7945 ;
  assign n8660 = n1166 & ~n8659 ;
  assign n8661 = ( n6190 & ~n6204 ) | ( n6190 & n8660 ) | ( ~n6204 & n8660 ) ;
  assign n8662 = n8233 ^ n6626 ^ 1'b0 ;
  assign n8663 = n8662 ^ n2962 ^ 1'b0 ;
  assign n8667 = ( n3652 & n4596 ) | ( n3652 & n5148 ) | ( n4596 & n5148 ) ;
  assign n8664 = n6110 ^ n1068 ^ 1'b0 ;
  assign n8665 = n2950 & n8664 ;
  assign n8666 = n8665 ^ n6984 ^ n889 ;
  assign n8668 = n8667 ^ n8666 ^ n2690 ;
  assign n8669 = n669 & n4247 ;
  assign n8670 = ~n8668 & n8669 ;
  assign n8671 = ( n2509 & ~n8229 ) | ( n2509 & n8241 ) | ( ~n8229 & n8241 ) ;
  assign n8672 = ( ~n576 & n6162 ) | ( ~n576 & n6448 ) | ( n6162 & n6448 ) ;
  assign n8673 = n7073 ^ n4509 ^ 1'b0 ;
  assign n8674 = n4768 ^ n4581 ^ 1'b0 ;
  assign n8675 = n8674 ^ n3618 ^ n1739 ;
  assign n8676 = ( ~n324 & n2698 ) | ( ~n324 & n2885 ) | ( n2698 & n2885 ) ;
  assign n8677 = n2937 ^ n1738 ^ 1'b0 ;
  assign n8678 = ( n6207 & n8676 ) | ( n6207 & ~n8677 ) | ( n8676 & ~n8677 ) ;
  assign n8679 = ( n1319 & n3494 ) | ( n1319 & n8678 ) | ( n3494 & n8678 ) ;
  assign n8680 = n8679 ^ n3887 ^ 1'b0 ;
  assign n8681 = n5946 | n8680 ;
  assign n8684 = ( ~n331 & n1961 ) | ( ~n331 & n6939 ) | ( n1961 & n6939 ) ;
  assign n8682 = ( ~n582 & n1064 ) | ( ~n582 & n3012 ) | ( n1064 & n3012 ) ;
  assign n8683 = n8682 ^ n4937 ^ n3078 ;
  assign n8685 = n8684 ^ n8683 ^ n1477 ;
  assign n8699 = n5391 ^ n4699 ^ n2824 ;
  assign n8698 = n3360 ^ n1696 ^ n1406 ;
  assign n8700 = n8699 ^ n8698 ^ n1289 ;
  assign n8686 = ( x4 & ~n1608 ) | ( x4 & n3296 ) | ( ~n1608 & n3296 ) ;
  assign n8687 = n3579 ^ n3136 ^ x88 ;
  assign n8688 = ( n6395 & n8686 ) | ( n6395 & ~n8687 ) | ( n8686 & ~n8687 ) ;
  assign n8689 = n5664 ^ n3655 ^ n844 ;
  assign n8690 = n2698 ^ n2458 ^ n918 ;
  assign n8691 = n8690 ^ n2216 ^ n2131 ;
  assign n8692 = n3254 ^ n661 ^ 1'b0 ;
  assign n8693 = n2452 | n7431 ;
  assign n8694 = n8692 & ~n8693 ;
  assign n8695 = ( n8689 & ~n8691 ) | ( n8689 & n8694 ) | ( ~n8691 & n8694 ) ;
  assign n8696 = n7006 & ~n8695 ;
  assign n8697 = n8688 & n8696 ;
  assign n8701 = n8700 ^ n8697 ^ n6501 ;
  assign n8702 = n8701 ^ n2474 ^ n1346 ;
  assign n8703 = ( ~x62 & n941 ) | ( ~x62 & n8702 ) | ( n941 & n8702 ) ;
  assign n8704 = n8703 ^ n8094 ^ n1951 ;
  assign n8705 = ( n2690 & n7592 ) | ( n2690 & ~n8050 ) | ( n7592 & ~n8050 ) ;
  assign n8706 = n1324 & ~n5466 ;
  assign n8707 = n8706 ^ n8426 ^ n3292 ;
  assign n8711 = n4215 ^ n3641 ^ 1'b0 ;
  assign n8708 = n3269 ^ n1420 ^ 1'b0 ;
  assign n8709 = ( ~n3014 & n4627 ) | ( ~n3014 & n7792 ) | ( n4627 & n7792 ) ;
  assign n8710 = ( n3245 & ~n8708 ) | ( n3245 & n8709 ) | ( ~n8708 & n8709 ) ;
  assign n8712 = n8711 ^ n8710 ^ n8511 ;
  assign n8713 = n4934 ^ n425 ^ n258 ;
  assign n8714 = ( n6121 & ~n6604 ) | ( n6121 & n8713 ) | ( ~n6604 & n8713 ) ;
  assign n8715 = n8714 ^ n3072 ^ n1125 ;
  assign n8716 = n7715 ^ x128 ^ 1'b0 ;
  assign n8719 = ( n415 & n2164 ) | ( n415 & n4683 ) | ( n2164 & n4683 ) ;
  assign n8720 = ( ~x146 & n1161 ) | ( ~x146 & n8719 ) | ( n1161 & n8719 ) ;
  assign n8717 = n6282 | n6472 ;
  assign n8718 = n3755 | n8717 ;
  assign n8721 = n8720 ^ n8718 ^ 1'b0 ;
  assign n8722 = ( n6676 & ~n8716 ) | ( n6676 & n8721 ) | ( ~n8716 & n8721 ) ;
  assign n8723 = ( n5199 & n5885 ) | ( n5199 & n6346 ) | ( n5885 & n6346 ) ;
  assign n8728 = ( n2592 & n3040 ) | ( n2592 & ~n6578 ) | ( n3040 & ~n6578 ) ;
  assign n8729 = n8728 ^ n3728 ^ n2099 ;
  assign n8725 = n1143 ^ n1108 ^ n871 ;
  assign n8724 = n5439 ^ n3597 ^ n2571 ;
  assign n8726 = n8725 ^ n8724 ^ 1'b0 ;
  assign n8727 = n324 & ~n8726 ;
  assign n8730 = n8729 ^ n8727 ^ n2317 ;
  assign n8733 = n1464 & ~n1678 ;
  assign n8734 = n2863 & n8733 ;
  assign n8731 = ( n409 & ~n1139 ) | ( n409 & n1902 ) | ( ~n1139 & n1902 ) ;
  assign n8732 = n8731 ^ n3729 ^ n1001 ;
  assign n8735 = n8734 ^ n8732 ^ n1432 ;
  assign n8736 = n3579 ^ n2627 ^ n950 ;
  assign n8737 = n4707 ^ n4308 ^ n2907 ;
  assign n8738 = ( n1795 & ~n2636 ) | ( n1795 & n8737 ) | ( ~n2636 & n8737 ) ;
  assign n8739 = n2022 ^ n1264 ^ 1'b0 ;
  assign n8740 = n8738 & ~n8739 ;
  assign n8741 = ~n1342 & n8740 ;
  assign n8742 = n8741 ^ n2469 ^ 1'b0 ;
  assign n8743 = ( x76 & ~n8736 ) | ( x76 & n8742 ) | ( ~n8736 & n8742 ) ;
  assign n8744 = ( ~n2976 & n8735 ) | ( ~n2976 & n8743 ) | ( n8735 & n8743 ) ;
  assign n8745 = n5077 & n8744 ;
  assign n8746 = ( ~n5732 & n6329 ) | ( ~n5732 & n8031 ) | ( n6329 & n8031 ) ;
  assign n8747 = n1129 ^ x235 ^ x93 ;
  assign n8748 = n8747 ^ n5289 ^ n3594 ;
  assign n8749 = n363 & n8748 ;
  assign n8750 = ~n8746 & n8749 ;
  assign n8751 = ( ~n728 & n8745 ) | ( ~n728 & n8750 ) | ( n8745 & n8750 ) ;
  assign n8752 = n3835 ^ n3165 ^ 1'b0 ;
  assign n8753 = ( ~n4566 & n8247 ) | ( ~n4566 & n8440 ) | ( n8247 & n8440 ) ;
  assign n8754 = n5043 & n6479 ;
  assign n8755 = n8754 ^ n7455 ^ 1'b0 ;
  assign n8756 = n8755 ^ n2790 ^ 1'b0 ;
  assign n8757 = ( n2386 & n3985 ) | ( n2386 & n4204 ) | ( n3985 & n4204 ) ;
  assign n8759 = n948 & n1447 ;
  assign n8760 = n8759 ^ x68 ^ 1'b0 ;
  assign n8758 = n7325 ^ n6423 ^ n1744 ;
  assign n8761 = n8760 ^ n8758 ^ n3434 ;
  assign n8762 = ( n1308 & ~n1441 ) | ( n1308 & n5357 ) | ( ~n1441 & n5357 ) ;
  assign n8767 = ( n2457 & n6537 ) | ( n2457 & n7376 ) | ( n6537 & n7376 ) ;
  assign n8768 = n3614 | n8767 ;
  assign n8763 = n310 | n496 ;
  assign n8764 = n8763 ^ n4003 ^ 1'b0 ;
  assign n8765 = n8431 ^ n4457 ^ n3608 ;
  assign n8766 = ( n3889 & n8764 ) | ( n3889 & n8765 ) | ( n8764 & n8765 ) ;
  assign n8769 = n8768 ^ n8766 ^ n4159 ;
  assign n8770 = ( n8299 & n8762 ) | ( n8299 & ~n8769 ) | ( n8762 & ~n8769 ) ;
  assign n8771 = ( n8757 & n8761 ) | ( n8757 & ~n8770 ) | ( n8761 & ~n8770 ) ;
  assign n8772 = ( n2152 & ~n3213 ) | ( n2152 & n6597 ) | ( ~n3213 & n6597 ) ;
  assign n8773 = ( n1782 & n6815 ) | ( n1782 & ~n7018 ) | ( n6815 & ~n7018 ) ;
  assign n8774 = n8773 ^ n2669 ^ 1'b0 ;
  assign n8775 = n6297 & ~n8774 ;
  assign n8776 = ( n3020 & n8772 ) | ( n3020 & n8775 ) | ( n8772 & n8775 ) ;
  assign n8777 = ( ~n4506 & n7246 ) | ( ~n4506 & n8395 ) | ( n7246 & n8395 ) ;
  assign n8778 = n8777 ^ n4403 ^ 1'b0 ;
  assign n8779 = n7713 & n8778 ;
  assign n8784 = ( n459 & n2732 ) | ( n459 & ~n2885 ) | ( n2732 & ~n2885 ) ;
  assign n8785 = n3154 ^ n948 ^ 1'b0 ;
  assign n8786 = n8785 ^ n5021 ^ n569 ;
  assign n8787 = n7562 ^ n7340 ^ n4436 ;
  assign n8788 = n1140 & n5179 ;
  assign n8789 = ~n8787 & n8788 ;
  assign n8790 = n8789 ^ n1162 ^ 1'b0 ;
  assign n8791 = n2498 & n8790 ;
  assign n8792 = ( n8784 & n8786 ) | ( n8784 & n8791 ) | ( n8786 & n8791 ) ;
  assign n8783 = n6293 ^ n6124 ^ 1'b0 ;
  assign n8780 = ~n4761 & n6480 ;
  assign n8781 = n2230 & ~n8780 ;
  assign n8782 = ~n6876 & n8781 ;
  assign n8793 = n8792 ^ n8783 ^ n8782 ;
  assign n8794 = n1889 & n7221 ;
  assign n8795 = ( n1888 & n7946 ) | ( n1888 & ~n8794 ) | ( n7946 & ~n8794 ) ;
  assign n8796 = n8795 ^ n2912 ^ 1'b0 ;
  assign n8797 = n3601 ^ n3075 ^ n2723 ;
  assign n8798 = n6564 ^ n4426 ^ 1'b0 ;
  assign n8799 = n8797 | n8798 ;
  assign n8800 = n8799 ^ n7055 ^ 1'b0 ;
  assign n8801 = n8800 ^ n3399 ^ 1'b0 ;
  assign n8804 = n4891 ^ n3616 ^ n1256 ;
  assign n8802 = ( n256 & n2684 ) | ( n256 & n4447 ) | ( n2684 & n4447 ) ;
  assign n8803 = n8802 ^ n5029 ^ n4403 ;
  assign n8805 = n8804 ^ n8803 ^ n5524 ;
  assign n8809 = n4748 ^ n4701 ^ 1'b0 ;
  assign n8810 = n631 | n8809 ;
  assign n8806 = n6737 ^ n773 ^ x18 ;
  assign n8807 = n4039 & ~n8806 ;
  assign n8808 = n8807 ^ n3923 ^ n1997 ;
  assign n8811 = n8810 ^ n8808 ^ n1455 ;
  assign n8812 = n2843 & n6422 ;
  assign n8813 = n8812 ^ n1001 ^ 1'b0 ;
  assign n8814 = n6991 ^ n4143 ^ 1'b0 ;
  assign n8815 = n8813 & ~n8814 ;
  assign n8816 = n6293 & ~n8815 ;
  assign n8817 = ( n1097 & n4378 ) | ( n1097 & ~n8816 ) | ( n4378 & ~n8816 ) ;
  assign n8818 = ( n626 & n1822 ) | ( n626 & n3261 ) | ( n1822 & n3261 ) ;
  assign n8819 = ( n1852 & ~n3476 ) | ( n1852 & n8818 ) | ( ~n3476 & n8818 ) ;
  assign n8820 = n4349 ^ n4216 ^ n1058 ;
  assign n8821 = ( n1742 & n8819 ) | ( n1742 & ~n8820 ) | ( n8819 & ~n8820 ) ;
  assign n8830 = n4468 ^ n3644 ^ n770 ;
  assign n8826 = n7694 ^ n3079 ^ n565 ;
  assign n8827 = n7808 ^ n2350 ^ n321 ;
  assign n8828 = ( n4073 & n8826 ) | ( n4073 & ~n8827 ) | ( n8826 & ~n8827 ) ;
  assign n8825 = ~n1082 & n7250 ;
  assign n8829 = n8828 ^ n8825 ^ n3721 ;
  assign n8831 = n8830 ^ n8829 ^ 1'b0 ;
  assign n8822 = n581 & n3132 ;
  assign n8823 = x197 | n8822 ;
  assign n8824 = n1541 & n8823 ;
  assign n8832 = n8831 ^ n8824 ^ 1'b0 ;
  assign n8833 = n3915 ^ n3703 ^ n2721 ;
  assign n8834 = n4192 ^ n3750 ^ n2077 ;
  assign n8835 = ( n2925 & n3534 ) | ( n2925 & ~n8834 ) | ( n3534 & ~n8834 ) ;
  assign n8837 = ( ~n3315 & n4108 ) | ( ~n3315 & n5637 ) | ( n4108 & n5637 ) ;
  assign n8838 = n8837 ^ n5470 ^ 1'b0 ;
  assign n8839 = n1477 & ~n8838 ;
  assign n8836 = n5022 ^ n3562 ^ n2853 ;
  assign n8840 = n8839 ^ n8836 ^ n4133 ;
  assign n8841 = n1914 & ~n8840 ;
  assign n8842 = ( n311 & ~n8835 ) | ( n311 & n8841 ) | ( ~n8835 & n8841 ) ;
  assign n8843 = n8833 & ~n8842 ;
  assign n8847 = n696 & ~n3387 ;
  assign n8848 = ~n1608 & n8847 ;
  assign n8849 = ( ~n1646 & n3435 ) | ( ~n1646 & n8848 ) | ( n3435 & n8848 ) ;
  assign n8844 = ( n1821 & n2028 ) | ( n1821 & n3930 ) | ( n2028 & n3930 ) ;
  assign n8845 = n7555 ^ n5215 ^ n1352 ;
  assign n8846 = ( n6497 & ~n8844 ) | ( n6497 & n8845 ) | ( ~n8844 & n8845 ) ;
  assign n8850 = n8849 ^ n8846 ^ n2010 ;
  assign n8859 = n3355 & n3550 ;
  assign n8860 = ~n1455 & n8859 ;
  assign n8861 = n7858 ^ n4481 ^ 1'b0 ;
  assign n8862 = ~n8860 & n8861 ;
  assign n8851 = n1748 ^ n749 ^ 1'b0 ;
  assign n8852 = ( n1407 & n3451 ) | ( n1407 & ~n8851 ) | ( n3451 & ~n8851 ) ;
  assign n8853 = n4754 & ~n6264 ;
  assign n8854 = n8853 ^ n6215 ^ 1'b0 ;
  assign n8855 = n2495 | n8854 ;
  assign n8856 = n8855 ^ n1686 ^ 1'b0 ;
  assign n8857 = ~n8852 & n8856 ;
  assign n8858 = n8857 ^ n6137 ^ 1'b0 ;
  assign n8863 = n8862 ^ n8858 ^ 1'b0 ;
  assign n8864 = n7778 & n8863 ;
  assign n8871 = n5778 ^ n3245 ^ n1322 ;
  assign n8870 = ~n1321 & n3564 ;
  assign n8872 = n8871 ^ n8870 ^ 1'b0 ;
  assign n8873 = n8872 ^ n1793 ^ n1761 ;
  assign n8866 = ~n341 & n476 ;
  assign n8867 = ~n6524 & n8866 ;
  assign n8868 = n8867 ^ n4021 ^ 1'b0 ;
  assign n8865 = ( n434 & n5748 ) | ( n434 & n7443 ) | ( n5748 & n7443 ) ;
  assign n8869 = n8868 ^ n8865 ^ n5153 ;
  assign n8874 = n8873 ^ n8869 ^ x89 ;
  assign n8875 = ( n5762 & n8263 ) | ( n5762 & n8874 ) | ( n8263 & n8874 ) ;
  assign n8876 = ( n3021 & ~n5396 ) | ( n3021 & n8761 ) | ( ~n5396 & n8761 ) ;
  assign n8877 = n809 & ~n1296 ;
  assign n8878 = ~x2 & n8877 ;
  assign n8879 = ( n7053 & ~n8876 ) | ( n7053 & n8878 ) | ( ~n8876 & n8878 ) ;
  assign n8880 = n8879 ^ n2926 ^ n1609 ;
  assign n8881 = ~n2491 & n6391 ;
  assign n8882 = n8881 ^ n5161 ^ n2647 ;
  assign n8883 = n8882 ^ n1557 ^ n321 ;
  assign n8884 = n5808 ^ n1320 ^ x125 ;
  assign n8885 = n1063 | n5815 ;
  assign n8886 = ( n1916 & n4359 ) | ( n1916 & n6883 ) | ( n4359 & n6883 ) ;
  assign n8887 = n8886 ^ n6600 ^ n1022 ;
  assign n8888 = ~n8687 & n8887 ;
  assign n8889 = n8888 ^ x152 ^ 1'b0 ;
  assign n8890 = ~n8885 & n8889 ;
  assign n8891 = ( n7686 & n8884 ) | ( n7686 & ~n8890 ) | ( n8884 & ~n8890 ) ;
  assign n8892 = n5040 ^ n1757 ^ 1'b0 ;
  assign n8893 = n2271 | n8892 ;
  assign n8894 = n8760 | n8893 ;
  assign n8895 = n8894 ^ n1638 ^ 1'b0 ;
  assign n8896 = n3132 ^ n391 ^ x137 ;
  assign n8897 = n8896 ^ n4595 ^ n448 ;
  assign n8898 = ( n1069 & n7857 ) | ( n1069 & n8897 ) | ( n7857 & n8897 ) ;
  assign n8899 = ( n286 & ~n4314 ) | ( n286 & n6987 ) | ( ~n4314 & n6987 ) ;
  assign n8900 = ( n308 & ~n1986 ) | ( n308 & n5560 ) | ( ~n1986 & n5560 ) ;
  assign n8901 = n5268 ^ n3019 ^ n1768 ;
  assign n8902 = ( ~n4806 & n8900 ) | ( ~n4806 & n8901 ) | ( n8900 & n8901 ) ;
  assign n8903 = n8358 | n8902 ;
  assign n8904 = ( n8472 & ~n8899 ) | ( n8472 & n8903 ) | ( ~n8899 & n8903 ) ;
  assign n8908 = n4636 ^ n4315 ^ n2895 ;
  assign n8909 = n8908 ^ n506 ^ n424 ;
  assign n8905 = n5148 ^ n1757 ^ n1101 ;
  assign n8906 = n8905 ^ n6507 ^ n912 ;
  assign n8907 = n8906 ^ n8505 ^ n7032 ;
  assign n8910 = n8909 ^ n8907 ^ n4556 ;
  assign n8911 = n5403 ^ x151 ^ 1'b0 ;
  assign n8912 = n8910 & n8911 ;
  assign n8913 = ( n1117 & n8904 ) | ( n1117 & n8912 ) | ( n8904 & n8912 ) ;
  assign n8916 = n4752 ^ n1677 ^ 1'b0 ;
  assign n8917 = n5065 & n8916 ;
  assign n8914 = n2919 ^ n2253 ^ n1367 ;
  assign n8915 = n8914 ^ n7420 ^ n4427 ;
  assign n8918 = n8917 ^ n8915 ^ n3994 ;
  assign n8922 = n6025 ^ n4961 ^ n1462 ;
  assign n8919 = ( n1738 & n2178 ) | ( n1738 & ~n3018 ) | ( n2178 & ~n3018 ) ;
  assign n8920 = n8919 ^ n6456 ^ n6187 ;
  assign n8921 = ~n3831 & n8920 ;
  assign n8923 = n8922 ^ n8921 ^ 1'b0 ;
  assign n8924 = n8509 ^ n7143 ^ n5179 ;
  assign n8925 = n8924 ^ n5110 ^ n3297 ;
  assign n8933 = ( n341 & n1304 ) | ( n341 & n1778 ) | ( n1304 & n1778 ) ;
  assign n8934 = n8933 ^ n1678 ^ n1479 ;
  assign n8935 = n8934 ^ n6662 ^ n5800 ;
  assign n8926 = n6154 ^ n4947 ^ n4892 ;
  assign n8928 = n3913 ^ n2304 ^ x200 ;
  assign n8929 = n8928 ^ n3118 ^ 1'b0 ;
  assign n8930 = n6077 | n8929 ;
  assign n8927 = ( ~n487 & n3058 ) | ( ~n487 & n4575 ) | ( n3058 & n4575 ) ;
  assign n8931 = n8930 ^ n8927 ^ 1'b0 ;
  assign n8932 = n8926 & ~n8931 ;
  assign n8936 = n8935 ^ n8932 ^ n5448 ;
  assign n8937 = n7828 ^ n2696 ^ n1349 ;
  assign n8938 = n3922 | n7651 ;
  assign n8939 = n8938 ^ n3191 ^ n658 ;
  assign n8945 = ( ~n1430 & n1803 ) | ( ~n1430 & n8652 ) | ( n1803 & n8652 ) ;
  assign n8946 = ( n944 & ~n8205 ) | ( n944 & n8945 ) | ( ~n8205 & n8945 ) ;
  assign n8940 = n1270 | n3898 ;
  assign n8941 = n8940 ^ n5255 ^ 1'b0 ;
  assign n8942 = ( ~n439 & n6938 ) | ( ~n439 & n8941 ) | ( n6938 & n8941 ) ;
  assign n8943 = ( n1782 & ~n2414 ) | ( n1782 & n6630 ) | ( ~n2414 & n6630 ) ;
  assign n8944 = n8942 & ~n8943 ;
  assign n8947 = n8946 ^ n8944 ^ 1'b0 ;
  assign n8948 = ( n3014 & ~n3090 ) | ( n3014 & n8947 ) | ( ~n3090 & n8947 ) ;
  assign n8950 = n8002 ^ n6787 ^ n2151 ;
  assign n8951 = n8950 ^ n4344 ^ n753 ;
  assign n8952 = ~n2278 & n5804 ;
  assign n8953 = n8952 ^ n3210 ^ 1'b0 ;
  assign n8954 = n8953 ^ n909 ^ 1'b0 ;
  assign n8955 = n8951 | n8954 ;
  assign n8949 = ( n1814 & ~n2145 ) | ( n1814 & n8279 ) | ( ~n2145 & n8279 ) ;
  assign n8956 = n8955 ^ n8949 ^ n7962 ;
  assign n8962 = n3257 ^ n2325 ^ x216 ;
  assign n8960 = ( n479 & n4256 ) | ( n479 & ~n7534 ) | ( n4256 & ~n7534 ) ;
  assign n8961 = n8960 ^ n5751 ^ 1'b0 ;
  assign n8957 = ( ~n968 & n1282 ) | ( ~n968 & n3705 ) | ( n1282 & n3705 ) ;
  assign n8958 = n8957 ^ n882 ^ 1'b0 ;
  assign n8959 = n8958 ^ n8700 ^ n7107 ;
  assign n8963 = n8962 ^ n8961 ^ n8959 ;
  assign n8967 = n4993 ^ n2530 ^ n688 ;
  assign n8966 = n6844 & ~n7503 ;
  assign n8968 = n8967 ^ n8966 ^ 1'b0 ;
  assign n8969 = n8968 ^ n7141 ^ n1634 ;
  assign n8964 = n3786 ^ n1903 ^ n1784 ;
  assign n8965 = ( ~n1590 & n1866 ) | ( ~n1590 & n8964 ) | ( n1866 & n8964 ) ;
  assign n8970 = n8969 ^ n8965 ^ n8933 ;
  assign n8971 = n4474 & ~n5115 ;
  assign n8972 = ~n1023 & n1977 ;
  assign n8973 = n8972 ^ n2682 ^ x77 ;
  assign n8974 = n803 & n6169 ;
  assign n8975 = n8974 ^ x169 ^ 1'b0 ;
  assign n8976 = n8975 ^ n6145 ^ n2597 ;
  assign n8977 = n8976 ^ n8504 ^ n4904 ;
  assign n8978 = n8973 | n8977 ;
  assign n8979 = n8971 | n8978 ;
  assign n8981 = ( x87 & x195 ) | ( x87 & n1257 ) | ( x195 & n1257 ) ;
  assign n8982 = ( ~n1081 & n7781 ) | ( ~n1081 & n8981 ) | ( n7781 & n8981 ) ;
  assign n8983 = ( n1793 & n4801 ) | ( n1793 & ~n5881 ) | ( n4801 & ~n5881 ) ;
  assign n8984 = n5104 ^ n4173 ^ 1'b0 ;
  assign n8985 = n8984 ^ n3835 ^ x114 ;
  assign n8986 = ( n8982 & ~n8983 ) | ( n8982 & n8985 ) | ( ~n8983 & n8985 ) ;
  assign n8980 = n8008 ^ n1125 ^ x217 ;
  assign n8987 = n8986 ^ n8980 ^ 1'b0 ;
  assign n8988 = ~n1791 & n3093 ;
  assign n8989 = n8988 ^ n1256 ^ 1'b0 ;
  assign n8990 = n8989 ^ n824 ^ n316 ;
  assign n8991 = ( x172 & ~n1060 ) | ( x172 & n8990 ) | ( ~n1060 & n8990 ) ;
  assign n8992 = n8991 ^ n7394 ^ n6222 ;
  assign n8993 = ~n7793 & n8992 ;
  assign n8994 = n8993 ^ n4618 ^ 1'b0 ;
  assign n8995 = n4064 ^ n926 ^ 1'b0 ;
  assign n8996 = n906 & n8995 ;
  assign n8997 = n1620 | n8996 ;
  assign n8998 = ( ~n4991 & n7615 ) | ( ~n4991 & n8997 ) | ( n7615 & n8997 ) ;
  assign n8999 = n3235 & ~n8998 ;
  assign n9000 = n8999 ^ n8609 ^ 1'b0 ;
  assign n9001 = n2096 | n9000 ;
  assign n9002 = n7768 & n9001 ;
  assign n9003 = ~n8994 & n9002 ;
  assign n9012 = ( n702 & n891 ) | ( n702 & n7573 ) | ( n891 & n7573 ) ;
  assign n9010 = ( n5299 & n7118 ) | ( n5299 & n8341 ) | ( n7118 & n8341 ) ;
  assign n9008 = n2511 | n8647 ;
  assign n9009 = n9008 ^ n2262 ^ 1'b0 ;
  assign n9011 = n9010 ^ n9009 ^ n2006 ;
  assign n9013 = n9012 ^ n9011 ^ n6128 ;
  assign n9004 = n5278 ^ n4063 ^ 1'b0 ;
  assign n9005 = n4088 & n9004 ;
  assign n9006 = n2302 | n5155 ;
  assign n9007 = n9005 & ~n9006 ;
  assign n9014 = n9013 ^ n9007 ^ 1'b0 ;
  assign n9015 = n9014 ^ n7468 ^ x9 ;
  assign n9016 = n426 | n8048 ;
  assign n9017 = n9016 ^ n2240 ^ n308 ;
  assign n9018 = n4783 ^ n1738 ^ 1'b0 ;
  assign n9019 = ( n3108 & n9017 ) | ( n3108 & n9018 ) | ( n9017 & n9018 ) ;
  assign n9026 = n3617 ^ n2971 ^ n2604 ;
  assign n9022 = n4043 ^ n1795 ^ n1179 ;
  assign n9023 = n2880 & n9022 ;
  assign n9024 = n1658 & n9023 ;
  assign n9025 = ~n888 & n9024 ;
  assign n9027 = n9026 ^ n9025 ^ n6094 ;
  assign n9020 = ( n1582 & ~n6883 ) | ( n1582 & n8172 ) | ( ~n6883 & n8172 ) ;
  assign n9021 = ~n7600 & n9020 ;
  assign n9028 = n9027 ^ n9021 ^ 1'b0 ;
  assign n9029 = n3778 ^ n1149 ^ 1'b0 ;
  assign n9030 = n9029 ^ n4096 ^ n3603 ;
  assign n9031 = n8317 & n9030 ;
  assign n9032 = n8288 & n9031 ;
  assign n9033 = n6020 ^ n3277 ^ n1041 ;
  assign n9034 = n3635 & ~n4151 ;
  assign n9035 = ( n2347 & n5603 ) | ( n2347 & ~n9034 ) | ( n5603 & ~n9034 ) ;
  assign n9036 = ( n6591 & ~n9033 ) | ( n6591 & n9035 ) | ( ~n9033 & n9035 ) ;
  assign n9037 = ( n3660 & n8118 ) | ( n3660 & n9036 ) | ( n8118 & n9036 ) ;
  assign n9040 = ( n335 & ~n3173 ) | ( n335 & n7085 ) | ( ~n3173 & n7085 ) ;
  assign n9041 = n9040 ^ n2933 ^ 1'b0 ;
  assign n9043 = n2459 ^ x23 ^ 1'b0 ;
  assign n9044 = n2402 & n9043 ;
  assign n9045 = ~n5049 & n9044 ;
  assign n9046 = ~n2752 & n9045 ;
  assign n9042 = ( ~n682 & n986 ) | ( ~n682 & n2034 ) | ( n986 & n2034 ) ;
  assign n9047 = n9046 ^ n9042 ^ 1'b0 ;
  assign n9048 = n9041 & ~n9047 ;
  assign n9038 = n8483 ^ n4258 ^ n1255 ;
  assign n9039 = n8505 & ~n9038 ;
  assign n9049 = n9048 ^ n9039 ^ 1'b0 ;
  assign n9050 = n3765 ^ n1822 ^ 1'b0 ;
  assign n9051 = ( ~x48 & n4133 ) | ( ~x48 & n4504 ) | ( n4133 & n4504 ) ;
  assign n9052 = ( n4899 & n8225 ) | ( n4899 & n8564 ) | ( n8225 & n8564 ) ;
  assign n9053 = ( n1114 & n2162 ) | ( n1114 & ~n5253 ) | ( n2162 & ~n5253 ) ;
  assign n9054 = n9053 ^ n2429 ^ n1117 ;
  assign n9055 = ( ~n9051 & n9052 ) | ( ~n9051 & n9054 ) | ( n9052 & n9054 ) ;
  assign n9056 = ( x97 & n3391 ) | ( x97 & ~n9055 ) | ( n3391 & ~n9055 ) ;
  assign n9085 = n7394 ^ n5873 ^ n4164 ;
  assign n9081 = n6083 ^ n387 ^ x114 ;
  assign n9082 = n7874 ^ n1885 ^ n1404 ;
  assign n9083 = n9082 ^ n4151 ^ n1113 ;
  assign n9084 = n9081 & n9083 ;
  assign n9086 = n9085 ^ n9084 ^ 1'b0 ;
  assign n9057 = n2232 | n4890 ;
  assign n9065 = n1703 ^ n1225 ^ 1'b0 ;
  assign n9066 = n7796 & n9065 ;
  assign n9067 = n9066 ^ n6541 ^ n480 ;
  assign n9068 = ( n330 & ~n3377 ) | ( n330 & n9067 ) | ( ~n3377 & n9067 ) ;
  assign n9058 = n6682 ^ n2137 ^ n1968 ;
  assign n9059 = n1130 ^ n1107 ^ n582 ;
  assign n9060 = n7316 ^ n5168 ^ 1'b0 ;
  assign n9061 = ( n2094 & n9059 ) | ( n2094 & ~n9060 ) | ( n9059 & ~n9060 ) ;
  assign n9062 = ( n425 & ~n9058 ) | ( n425 & n9061 ) | ( ~n9058 & n9061 ) ;
  assign n9063 = n9062 ^ n2909 ^ 1'b0 ;
  assign n9064 = n6006 & ~n9063 ;
  assign n9069 = n9068 ^ n9064 ^ n4868 ;
  assign n9070 = ( n4847 & n9057 ) | ( n4847 & n9069 ) | ( n9057 & n9069 ) ;
  assign n9073 = n5648 ^ n3770 ^ 1'b0 ;
  assign n9074 = n1329 & n9073 ;
  assign n9071 = n1060 & n3604 ;
  assign n9072 = n9071 ^ n2349 ^ 1'b0 ;
  assign n9075 = n9074 ^ n9072 ^ x219 ;
  assign n9076 = ( ~n4948 & n7099 ) | ( ~n4948 & n9075 ) | ( n7099 & n9075 ) ;
  assign n9077 = n1069 | n9076 ;
  assign n9078 = ~n8983 & n9077 ;
  assign n9079 = ~n9070 & n9078 ;
  assign n9080 = n5901 | n9079 ;
  assign n9087 = n9086 ^ n9080 ^ 1'b0 ;
  assign n9088 = n7332 ^ n7319 ^ n4267 ;
  assign n9089 = x17 & n626 ;
  assign n9090 = ~n1714 & n9089 ;
  assign n9091 = n8191 ^ n334 ^ 1'b0 ;
  assign n9092 = ( n1233 & ~n9090 ) | ( n1233 & n9091 ) | ( ~n9090 & n9091 ) ;
  assign n9093 = ( n708 & n1465 ) | ( n708 & ~n1955 ) | ( n1465 & ~n1955 ) ;
  assign n9094 = n5284 & ~n9093 ;
  assign n9095 = ( n4506 & n9092 ) | ( n4506 & n9094 ) | ( n9092 & n9094 ) ;
  assign n9096 = n7209 ^ n2395 ^ n1069 ;
  assign n9097 = n5176 ^ n2940 ^ n1994 ;
  assign n9098 = n4335 & n9097 ;
  assign n9099 = ~n9096 & n9098 ;
  assign n9100 = ( n5871 & n6112 ) | ( n5871 & n7490 ) | ( n6112 & n7490 ) ;
  assign n9101 = n9100 ^ n3236 ^ 1'b0 ;
  assign n9102 = n6455 ^ n1517 ^ 1'b0 ;
  assign n9103 = n1545 ^ x137 ^ 1'b0 ;
  assign n9104 = n5388 | n9103 ;
  assign n9105 = ~n1061 & n1554 ;
  assign n9106 = n9105 ^ n2515 ^ 1'b0 ;
  assign n9107 = n805 ^ n576 ^ x240 ;
  assign n9108 = n9106 & ~n9107 ;
  assign n9109 = ( ~n8009 & n9104 ) | ( ~n8009 & n9108 ) | ( n9104 & n9108 ) ;
  assign n9110 = ~n2524 & n6240 ;
  assign n9111 = n9110 ^ n2465 ^ 1'b0 ;
  assign n9112 = n1592 | n9111 ;
  assign n9113 = ~n909 & n3149 ;
  assign n9114 = ~n2504 & n9113 ;
  assign n9115 = n9114 ^ n7571 ^ 1'b0 ;
  assign n9116 = n833 & n9115 ;
  assign n9117 = ( n3702 & n5822 ) | ( n3702 & ~n9116 ) | ( n5822 & ~n9116 ) ;
  assign n9118 = ( n4208 & n6993 ) | ( n4208 & n8601 ) | ( n6993 & n8601 ) ;
  assign n9126 = n6316 ^ n3486 ^ n277 ;
  assign n9122 = n6720 ^ n6507 ^ 1'b0 ;
  assign n9123 = n958 & n9122 ;
  assign n9124 = ~n406 & n9123 ;
  assign n9125 = ~n797 & n9124 ;
  assign n9119 = n1275 ^ n904 ^ 1'b0 ;
  assign n9120 = n1724 & ~n9119 ;
  assign n9121 = n9120 ^ n5764 ^ n3230 ;
  assign n9127 = n9126 ^ n9125 ^ n9121 ;
  assign n9129 = x166 & ~n2920 ;
  assign n9130 = ~n3875 & n9129 ;
  assign n9131 = ~n6578 & n9130 ;
  assign n9132 = ( n1887 & n3295 ) | ( n1887 & ~n9131 ) | ( n3295 & ~n9131 ) ;
  assign n9128 = n4647 ^ n4465 ^ 1'b0 ;
  assign n9133 = n9132 ^ n9128 ^ 1'b0 ;
  assign n9139 = n1751 ^ n1123 ^ 1'b0 ;
  assign n9140 = n2786 | n9139 ;
  assign n9141 = n5424 | n9140 ;
  assign n9134 = ~n1174 & n5070 ;
  assign n9135 = n1840 & n9134 ;
  assign n9136 = n2789 | n9135 ;
  assign n9137 = n9136 ^ n1180 ^ 1'b0 ;
  assign n9138 = n1268 & ~n9137 ;
  assign n9142 = n9141 ^ n9138 ^ 1'b0 ;
  assign n9143 = n3962 ^ n3855 ^ n2732 ;
  assign n9144 = ( n2718 & ~n7436 ) | ( n2718 & n9143 ) | ( ~n7436 & n9143 ) ;
  assign n9145 = ( ~n5237 & n5670 ) | ( ~n5237 & n9144 ) | ( n5670 & n9144 ) ;
  assign n9146 = ( n1064 & n2996 ) | ( n1064 & n9145 ) | ( n2996 & n9145 ) ;
  assign n9147 = n3682 & n8017 ;
  assign n9155 = ( n3128 & n4244 ) | ( n3128 & n8582 ) | ( n4244 & n8582 ) ;
  assign n9156 = n9155 ^ n761 ^ 1'b0 ;
  assign n9148 = n3153 & n4743 ;
  assign n9149 = n8731 ^ n4509 ^ x86 ;
  assign n9150 = n9149 ^ n1103 ^ 1'b0 ;
  assign n9151 = ~n9148 & n9150 ;
  assign n9152 = n9151 ^ n7019 ^ n4862 ;
  assign n9153 = n2425 ^ n517 ^ 1'b0 ;
  assign n9154 = ~n9152 & n9153 ;
  assign n9157 = n9156 ^ n9154 ^ 1'b0 ;
  assign n9158 = n1537 | n9157 ;
  assign n9159 = n9147 & ~n9158 ;
  assign n9160 = n3653 ^ n2994 ^ n1845 ;
  assign n9161 = n9160 ^ n7081 ^ n1040 ;
  assign n9162 = n5640 ^ n5479 ^ n5212 ;
  assign n9163 = ~n3671 & n3928 ;
  assign n9164 = n9162 & n9163 ;
  assign n9165 = ( n894 & n3420 ) | ( n894 & n9164 ) | ( n3420 & n9164 ) ;
  assign n9173 = ( n2059 & n4712 ) | ( n2059 & n6928 ) | ( n4712 & n6928 ) ;
  assign n9166 = ( n468 & n1795 ) | ( n468 & n5330 ) | ( n1795 & n5330 ) ;
  assign n9167 = n359 & ~n6903 ;
  assign n9168 = n9167 ^ n6813 ^ 1'b0 ;
  assign n9169 = n926 | n7940 ;
  assign n9170 = n9168 & ~n9169 ;
  assign n9171 = n5986 & ~n9170 ;
  assign n9172 = ~n9166 & n9171 ;
  assign n9174 = n9173 ^ n9172 ^ n6916 ;
  assign n9175 = n9174 ^ n8923 ^ n8405 ;
  assign n9177 = n482 | n7795 ;
  assign n9176 = ( ~x181 & n6830 ) | ( ~x181 & n8425 ) | ( n6830 & n8425 ) ;
  assign n9178 = n9177 ^ n9176 ^ n9140 ;
  assign n9179 = ( ~n5916 & n6014 ) | ( ~n5916 & n9178 ) | ( n6014 & n9178 ) ;
  assign n9180 = ( ~n1266 & n1692 ) | ( ~n1266 & n9131 ) | ( n1692 & n9131 ) ;
  assign n9181 = n1529 | n4820 ;
  assign n9182 = n947 | n9181 ;
  assign n9183 = ( n8440 & n8888 ) | ( n8440 & n9182 ) | ( n8888 & n9182 ) ;
  assign n9184 = ( n8395 & n9180 ) | ( n8395 & n9183 ) | ( n9180 & n9183 ) ;
  assign n9185 = n1079 ^ x216 ^ 1'b0 ;
  assign n9186 = n9185 ^ n8307 ^ n319 ;
  assign n9198 = n824 | n1164 ;
  assign n9199 = n3224 & n9198 ;
  assign n9187 = n4254 ^ n2046 ^ 1'b0 ;
  assign n9188 = ~n1450 & n9187 ;
  assign n9189 = ~n2385 & n3889 ;
  assign n9190 = n2610 & ~n9189 ;
  assign n9191 = ~n375 & n9190 ;
  assign n9192 = n5565 ^ n2094 ^ n1591 ;
  assign n9193 = n6836 ^ n5215 ^ n1372 ;
  assign n9194 = ( n1443 & n9192 ) | ( n1443 & n9193 ) | ( n9192 & n9193 ) ;
  assign n9195 = n9191 | n9194 ;
  assign n9196 = n9188 & n9195 ;
  assign n9197 = ~n6598 & n9196 ;
  assign n9200 = n9199 ^ n9197 ^ n6188 ;
  assign n9204 = n7006 ^ n4189 ^ n743 ;
  assign n9201 = ~n5698 & n8168 ;
  assign n9202 = n1595 & n9201 ;
  assign n9203 = ( n6100 & n6292 ) | ( n6100 & n9202 ) | ( n6292 & n9202 ) ;
  assign n9205 = n9204 ^ n9203 ^ n2966 ;
  assign n9206 = n4237 ^ n4150 ^ 1'b0 ;
  assign n9207 = n8886 ^ n4094 ^ n372 ;
  assign n9208 = n415 & n9207 ;
  assign n9209 = ~n9206 & n9208 ;
  assign n9210 = n9209 ^ n1991 ^ 1'b0 ;
  assign n9211 = n1325 & n9210 ;
  assign n9212 = n805 & ~n3329 ;
  assign n9214 = n5875 ^ n869 ^ n348 ;
  assign n9213 = ( ~n4375 & n7546 ) | ( ~n4375 & n7687 ) | ( n7546 & n7687 ) ;
  assign n9215 = n9214 ^ n9213 ^ n8683 ;
  assign n9224 = n8802 ^ n7746 ^ n2371 ;
  assign n9222 = n1440 | n2770 ;
  assign n9218 = n2080 ^ n1641 ^ n432 ;
  assign n9219 = x28 & ~n9218 ;
  assign n9220 = n2694 & n9219 ;
  assign n9221 = ( n2272 & ~n2519 ) | ( n2272 & n9220 ) | ( ~n2519 & n9220 ) ;
  assign n9216 = n5550 ^ n839 ^ n772 ;
  assign n9217 = ( n2703 & n7578 ) | ( n2703 & n9216 ) | ( n7578 & n9216 ) ;
  assign n9223 = n9222 ^ n9221 ^ n9217 ;
  assign n9225 = n9224 ^ n9223 ^ n3713 ;
  assign n9227 = n2623 ^ n654 ^ 1'b0 ;
  assign n9228 = n9227 ^ n1561 ^ 1'b0 ;
  assign n9229 = n3786 | n9228 ;
  assign n9226 = ( x19 & ~n532 ) | ( x19 & n2027 ) | ( ~n532 & n2027 ) ;
  assign n9230 = n9229 ^ n9226 ^ n3927 ;
  assign n9231 = n3463 ^ n385 ^ 1'b0 ;
  assign n9232 = ( n1492 & ~n5497 ) | ( n1492 & n9231 ) | ( ~n5497 & n9231 ) ;
  assign n9233 = n7039 | n9232 ;
  assign n9234 = n9233 ^ n3192 ^ 1'b0 ;
  assign n9235 = ( x72 & ~n511 ) | ( x72 & n6909 ) | ( ~n511 & n6909 ) ;
  assign n9236 = n9235 ^ n6365 ^ n3747 ;
  assign n9237 = ( n3735 & ~n9176 ) | ( n3735 & n9236 ) | ( ~n9176 & n9236 ) ;
  assign n9238 = n1840 | n2242 ;
  assign n9239 = n9238 ^ n745 ^ 1'b0 ;
  assign n9240 = n9239 ^ n6025 ^ n5852 ;
  assign n9241 = ( n8835 & ~n9237 ) | ( n8835 & n9240 ) | ( ~n9237 & n9240 ) ;
  assign n9242 = n2510 & ~n6093 ;
  assign n9244 = n5736 ^ n3020 ^ n1893 ;
  assign n9245 = n9244 ^ n2804 ^ 1'b0 ;
  assign n9246 = n8213 & ~n9245 ;
  assign n9247 = n7393 ^ n862 ^ 1'b0 ;
  assign n9248 = n9246 & n9247 ;
  assign n9243 = ( n817 & n3412 ) | ( n817 & ~n7235 ) | ( n3412 & ~n7235 ) ;
  assign n9249 = n9248 ^ n9243 ^ n3645 ;
  assign n9250 = n8056 ^ n6113 ^ n1326 ;
  assign n9251 = ( ~n1337 & n9249 ) | ( ~n1337 & n9250 ) | ( n9249 & n9250 ) ;
  assign n9252 = n5134 ^ n1233 ^ 1'b0 ;
  assign n9253 = ~n387 & n3689 ;
  assign n9254 = ( ~n1172 & n8487 ) | ( ~n1172 & n9253 ) | ( n8487 & n9253 ) ;
  assign n9255 = ( n577 & n9252 ) | ( n577 & ~n9254 ) | ( n9252 & ~n9254 ) ;
  assign n9256 = n5341 ^ n1552 ^ 1'b0 ;
  assign n9257 = n6666 ^ n6549 ^ n5894 ;
  assign n9258 = n9257 ^ n6863 ^ n6827 ;
  assign n9259 = ( n4344 & n9256 ) | ( n4344 & n9258 ) | ( n9256 & n9258 ) ;
  assign n9260 = ( ~n1673 & n3843 ) | ( ~n1673 & n9259 ) | ( n3843 & n9259 ) ;
  assign n9261 = n1568 ^ n1258 ^ n948 ;
  assign n9262 = n9261 ^ n7130 ^ n1555 ;
  assign n9263 = n9262 ^ n5698 ^ x6 ;
  assign n9272 = n2839 ^ n1690 ^ x149 ;
  assign n9269 = n1315 ^ n1045 ^ n880 ;
  assign n9270 = ( ~n1473 & n1585 ) | ( ~n1473 & n9269 ) | ( n1585 & n9269 ) ;
  assign n9271 = n9270 ^ n1973 ^ n514 ;
  assign n9273 = n9272 ^ n9271 ^ n3433 ;
  assign n9266 = ( x164 & n3700 ) | ( x164 & ~n7749 ) | ( n3700 & ~n7749 ) ;
  assign n9267 = ( n1203 & n7573 ) | ( n1203 & n9266 ) | ( n7573 & n9266 ) ;
  assign n9268 = ~n4876 & n9267 ;
  assign n9274 = n9273 ^ n9268 ^ n3583 ;
  assign n9264 = n6874 ^ n6344 ^ n4925 ;
  assign n9265 = ( n2804 & n3538 ) | ( n2804 & ~n9264 ) | ( n3538 & ~n9264 ) ;
  assign n9275 = n9274 ^ n9265 ^ n2612 ;
  assign n9276 = ~n2428 & n6143 ;
  assign n9277 = ( ~x52 & n5625 ) | ( ~x52 & n9276 ) | ( n5625 & n9276 ) ;
  assign n9278 = n4230 ^ n1918 ^ 1'b0 ;
  assign n9279 = n9278 ^ n8036 ^ n6352 ;
  assign n9280 = n4256 & n9279 ;
  assign n9281 = ( ~n2394 & n4806 ) | ( ~n2394 & n5505 ) | ( n4806 & n5505 ) ;
  assign n9282 = x16 & ~n1566 ;
  assign n9283 = n9282 ^ n3778 ^ 1'b0 ;
  assign n9284 = ( n1753 & ~n7519 ) | ( n1753 & n9283 ) | ( ~n7519 & n9283 ) ;
  assign n9285 = n9281 | n9284 ;
  assign n9286 = n9285 ^ n1841 ^ 1'b0 ;
  assign n9287 = n8720 & ~n9286 ;
  assign n9288 = n9287 ^ n1102 ^ 1'b0 ;
  assign n9289 = ( n697 & n9280 ) | ( n697 & n9288 ) | ( n9280 & n9288 ) ;
  assign n9290 = n4832 ^ n4549 ^ 1'b0 ;
  assign n9291 = ~n318 & n9290 ;
  assign n9292 = n673 & n962 ;
  assign n9293 = ( n766 & n1505 ) | ( n766 & n9292 ) | ( n1505 & n9292 ) ;
  assign n9294 = ( n770 & n1296 ) | ( n770 & n1344 ) | ( n1296 & n1344 ) ;
  assign n9295 = ( n1098 & n1430 ) | ( n1098 & n9294 ) | ( n1430 & n9294 ) ;
  assign n9296 = n5745 ^ n1374 ^ n536 ;
  assign n9297 = n5661 ^ n1195 ^ n414 ;
  assign n9298 = n9297 ^ n4994 ^ 1'b0 ;
  assign n9299 = n8618 & n9298 ;
  assign n9300 = n9299 ^ n387 ^ 1'b0 ;
  assign n9301 = n9296 & ~n9300 ;
  assign n9302 = ( n4145 & n6422 ) | ( n4145 & n9301 ) | ( n6422 & n9301 ) ;
  assign n9303 = n4035 ^ n3918 ^ n1002 ;
  assign n9304 = ( n9295 & ~n9302 ) | ( n9295 & n9303 ) | ( ~n9302 & n9303 ) ;
  assign n9314 = n2583 ^ n473 ^ x254 ;
  assign n9308 = ~n655 & n5846 ;
  assign n9309 = ( ~n427 & n3745 ) | ( ~n427 & n9308 ) | ( n3745 & n9308 ) ;
  assign n9310 = n9309 ^ n8706 ^ n1868 ;
  assign n9311 = ( x165 & n6027 ) | ( x165 & n9310 ) | ( n6027 & n9310 ) ;
  assign n9312 = n7378 ^ n5290 ^ n1964 ;
  assign n9313 = n9311 & n9312 ;
  assign n9315 = n9314 ^ n9313 ^ 1'b0 ;
  assign n9305 = ( n2909 & ~n5015 ) | ( n2909 & n5783 ) | ( ~n5015 & n5783 ) ;
  assign n9306 = ( ~n1826 & n2835 ) | ( ~n1826 & n9305 ) | ( n2835 & n9305 ) ;
  assign n9307 = n9306 ^ n5573 ^ 1'b0 ;
  assign n9316 = n9315 ^ n9307 ^ n1405 ;
  assign n9317 = ( n5505 & ~n9304 ) | ( n5505 & n9316 ) | ( ~n9304 & n9316 ) ;
  assign n9318 = ~n3747 & n8316 ;
  assign n9319 = ( n1990 & ~n7367 ) | ( n1990 & n9318 ) | ( ~n7367 & n9318 ) ;
  assign n9320 = ( ~n465 & n2361 ) | ( ~n465 & n2516 ) | ( n2361 & n2516 ) ;
  assign n9321 = n9319 | n9320 ;
  assign n9322 = n9321 ^ n3541 ^ 1'b0 ;
  assign n9323 = ( n1180 & n3841 ) | ( n1180 & ~n6708 ) | ( n3841 & ~n6708 ) ;
  assign n9330 = ( x53 & n568 ) | ( x53 & ~n1963 ) | ( n568 & ~n1963 ) ;
  assign n9324 = n2631 ^ n2248 ^ 1'b0 ;
  assign n9325 = ~n1717 & n9324 ;
  assign n9326 = n9325 ^ n2828 ^ n559 ;
  assign n9327 = ( ~n3347 & n8034 ) | ( ~n3347 & n9326 ) | ( n8034 & n9326 ) ;
  assign n9328 = n9327 ^ n815 ^ 1'b0 ;
  assign n9329 = ( ~n914 & n1326 ) | ( ~n914 & n9328 ) | ( n1326 & n9328 ) ;
  assign n9331 = n9330 ^ n9329 ^ 1'b0 ;
  assign n9332 = ( n2747 & ~n5975 ) | ( n2747 & n9331 ) | ( ~n5975 & n9331 ) ;
  assign n9333 = n9332 ^ n3084 ^ n1482 ;
  assign n9334 = n9333 ^ n8732 ^ 1'b0 ;
  assign n9335 = n9323 | n9334 ;
  assign n9336 = n8425 ^ n6816 ^ n6679 ;
  assign n9344 = n7274 ^ x65 ^ 1'b0 ;
  assign n9345 = n5135 & ~n9344 ;
  assign n9340 = ~n1296 & n1646 ;
  assign n9341 = n9340 ^ x233 ^ 1'b0 ;
  assign n9339 = n7624 ^ n7074 ^ n4883 ;
  assign n9342 = n9341 ^ n9339 ^ n7199 ;
  assign n9337 = n4227 ^ n853 ^ n702 ;
  assign n9338 = n7112 | n9337 ;
  assign n9343 = n9342 ^ n9338 ^ 1'b0 ;
  assign n9346 = n9345 ^ n9343 ^ n494 ;
  assign n9347 = ( n3383 & ~n4860 ) | ( n3383 & n5020 ) | ( ~n4860 & n5020 ) ;
  assign n9349 = ( ~n1848 & n2538 ) | ( ~n1848 & n3786 ) | ( n2538 & n3786 ) ;
  assign n9348 = ( n2894 & n3663 ) | ( n2894 & ~n5829 ) | ( n3663 & ~n5829 ) ;
  assign n9350 = n9349 ^ n9348 ^ n8922 ;
  assign n9351 = ( ~n8032 & n9347 ) | ( ~n8032 & n9350 ) | ( n9347 & n9350 ) ;
  assign n9353 = n3703 ^ n3209 ^ n2024 ;
  assign n9352 = n5735 ^ n4295 ^ n1065 ;
  assign n9354 = n9353 ^ n9352 ^ n5059 ;
  assign n9355 = ( x253 & n3308 ) | ( x253 & ~n9354 ) | ( n3308 & ~n9354 ) ;
  assign n9356 = n2677 ^ n2587 ^ 1'b0 ;
  assign n9357 = n5026 | n9356 ;
  assign n9358 = n9357 ^ n3196 ^ 1'b0 ;
  assign n9360 = n6822 ^ n6139 ^ n2003 ;
  assign n9359 = ~n2342 & n3824 ;
  assign n9361 = n9360 ^ n9359 ^ n8278 ;
  assign n9362 = n4764 ^ n2864 ^ 1'b0 ;
  assign n9363 = n9361 | n9362 ;
  assign n9364 = ( n4318 & n6109 ) | ( n4318 & n9363 ) | ( n6109 & n9363 ) ;
  assign n9365 = n9358 & ~n9364 ;
  assign n9366 = ~n1773 & n9365 ;
  assign n9367 = n9366 ^ n5222 ^ n2949 ;
  assign n9368 = n8471 ^ n4997 ^ n663 ;
  assign n9369 = n9368 ^ n3353 ^ n1410 ;
  assign n9370 = n9369 ^ n8209 ^ 1'b0 ;
  assign n9371 = ( ~n3388 & n3880 ) | ( ~n3388 & n7076 ) | ( n3880 & n7076 ) ;
  assign n9372 = ( ~n1047 & n1726 ) | ( ~n1047 & n1766 ) | ( n1726 & n1766 ) ;
  assign n9373 = ( ~n2046 & n5209 ) | ( ~n2046 & n9372 ) | ( n5209 & n9372 ) ;
  assign n9374 = ( n3767 & ~n8067 ) | ( n3767 & n8748 ) | ( ~n8067 & n8748 ) ;
  assign n9380 = n3250 ^ n525 ^ 1'b0 ;
  assign n9381 = n9380 ^ n3985 ^ 1'b0 ;
  assign n9379 = n5982 ^ n3505 ^ 1'b0 ;
  assign n9382 = n9381 ^ n9379 ^ n1630 ;
  assign n9375 = ( ~x65 & n2790 ) | ( ~x65 & n8004 ) | ( n2790 & n8004 ) ;
  assign n9376 = n9375 ^ n7707 ^ 1'b0 ;
  assign n9377 = ~n7211 & n9376 ;
  assign n9378 = n2981 & n9377 ;
  assign n9383 = n9382 ^ n9378 ^ n2856 ;
  assign n9384 = n6475 ^ n6316 ^ n4757 ;
  assign n9385 = ( n2768 & n8687 ) | ( n2768 & ~n9384 ) | ( n8687 & ~n9384 ) ;
  assign n9386 = n4822 & n9385 ;
  assign n9387 = ~n284 & n9386 ;
  assign n9388 = n6261 & ~n8631 ;
  assign n9389 = n9387 & n9388 ;
  assign n9390 = ~n7499 & n9389 ;
  assign n9391 = n5439 ^ n3927 ^ 1'b0 ;
  assign n9392 = n8167 ^ n2626 ^ n561 ;
  assign n9393 = ( n1753 & ~n9391 ) | ( n1753 & n9392 ) | ( ~n9391 & n9392 ) ;
  assign n9394 = n4854 ^ n2313 ^ 1'b0 ;
  assign n9395 = ~n8286 & n9394 ;
  assign n9396 = n5330 ^ n4783 ^ x234 ;
  assign n9397 = n9396 ^ n7640 ^ n7549 ;
  assign n9398 = ( n3789 & ~n9395 ) | ( n3789 & n9397 ) | ( ~n9395 & n9397 ) ;
  assign n9399 = n5875 ^ n3910 ^ n416 ;
  assign n9400 = n8160 ^ n2032 ^ 1'b0 ;
  assign n9401 = ~n1325 & n9400 ;
  assign n9402 = ( n805 & n9399 ) | ( n805 & n9401 ) | ( n9399 & n9401 ) ;
  assign n9403 = n3752 ^ n790 ^ 1'b0 ;
  assign n9404 = ( ~n790 & n9262 ) | ( ~n790 & n9403 ) | ( n9262 & n9403 ) ;
  assign n9405 = ( n2786 & n9402 ) | ( n2786 & n9404 ) | ( n9402 & n9404 ) ;
  assign n9406 = n2600 ^ x101 ^ 1'b0 ;
  assign n9407 = ~n1074 & n9406 ;
  assign n9408 = n9407 ^ n8425 ^ 1'b0 ;
  assign n9409 = ~n4504 & n9408 ;
  assign n9410 = ( n2787 & ~n5000 ) | ( n2787 & n6577 ) | ( ~n5000 & n6577 ) ;
  assign n9411 = ~n699 & n1844 ;
  assign n9412 = n9411 ^ n8154 ^ x97 ;
  assign n9413 = ( n9409 & n9410 ) | ( n9409 & ~n9412 ) | ( n9410 & ~n9412 ) ;
  assign n9416 = n1606 ^ n1525 ^ x49 ;
  assign n9414 = n4036 ^ n4017 ^ n2439 ;
  assign n9415 = n9414 ^ n2140 ^ n1659 ;
  assign n9417 = n9416 ^ n9415 ^ n1864 ;
  assign n9418 = ( n1489 & ~n4747 ) | ( n1489 & n7489 ) | ( ~n4747 & n7489 ) ;
  assign n9419 = ~n624 & n6603 ;
  assign n9420 = ( n4854 & n9418 ) | ( n4854 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9421 = n2245 ^ n1256 ^ x59 ;
  assign n9422 = ( n7137 & n7540 ) | ( n7137 & ~n9421 ) | ( n7540 & ~n9421 ) ;
  assign n9423 = n9422 ^ n4959 ^ 1'b0 ;
  assign n9429 = ( n1465 & ~n2510 ) | ( n1465 & n4647 ) | ( ~n2510 & n4647 ) ;
  assign n9430 = ( n3522 & ~n7225 ) | ( n3522 & n9429 ) | ( ~n7225 & n9429 ) ;
  assign n9428 = n3888 ^ n1872 ^ n393 ;
  assign n9431 = n9430 ^ n9428 ^ n5117 ;
  assign n9432 = n9431 ^ n2097 ^ n601 ;
  assign n9424 = ( n545 & ~n4502 ) | ( n545 & n4714 ) | ( ~n4502 & n4714 ) ;
  assign n9425 = n9424 ^ n4822 ^ n3872 ;
  assign n9426 = n9425 ^ n4042 ^ n2014 ;
  assign n9427 = n9426 ^ n7445 ^ n3010 ;
  assign n9433 = n9432 ^ n9427 ^ x8 ;
  assign n9441 = n6972 ^ n1162 ^ 1'b0 ;
  assign n9434 = n4158 & ~n5080 ;
  assign n9435 = ~n5446 & n9434 ;
  assign n9438 = ( ~x139 & n5832 ) | ( ~x139 & n6590 ) | ( n5832 & n6590 ) ;
  assign n9436 = n7614 ^ n6917 ^ 1'b0 ;
  assign n9437 = ~n8785 & n9436 ;
  assign n9439 = n9438 ^ n9437 ^ 1'b0 ;
  assign n9440 = n9435 | n9439 ;
  assign n9442 = n9441 ^ n9440 ^ n6179 ;
  assign n9443 = ( n1695 & n2797 ) | ( n1695 & ~n6292 ) | ( n2797 & ~n6292 ) ;
  assign n9444 = ( n1741 & n2084 ) | ( n1741 & n9443 ) | ( n2084 & n9443 ) ;
  assign n9451 = ( ~n811 & n6000 ) | ( ~n811 & n8436 ) | ( n6000 & n8436 ) ;
  assign n9446 = n364 & ~n3195 ;
  assign n9447 = ~n6739 & n9446 ;
  assign n9448 = ( ~n5472 & n7255 ) | ( ~n5472 & n9447 ) | ( n7255 & n9447 ) ;
  assign n9449 = n6329 & ~n9448 ;
  assign n9450 = ~n9297 & n9449 ;
  assign n9445 = n6669 ^ n6276 ^ n4223 ;
  assign n9452 = n9451 ^ n9450 ^ n9445 ;
  assign n9453 = n9452 ^ n6485 ^ 1'b0 ;
  assign n9454 = n7393 ^ n3594 ^ n1543 ;
  assign n9455 = ( n725 & n2331 ) | ( n725 & ~n9454 ) | ( n2331 & ~n9454 ) ;
  assign n9456 = n9455 ^ n8483 ^ n7198 ;
  assign n9457 = ( n1211 & ~n8684 ) | ( n1211 & n9456 ) | ( ~n8684 & n9456 ) ;
  assign n9458 = n9457 ^ n7534 ^ 1'b0 ;
  assign n9459 = ~n8502 & n9458 ;
  assign n9461 = ( ~x103 & n2721 ) | ( ~x103 & n7392 ) | ( n2721 & n7392 ) ;
  assign n9460 = n3090 ^ n2456 ^ n2345 ;
  assign n9462 = n9461 ^ n9460 ^ n4991 ;
  assign n9463 = n9462 ^ n7890 ^ n3794 ;
  assign n9464 = ( n782 & ~n1823 ) | ( n782 & n4673 ) | ( ~n1823 & n4673 ) ;
  assign n9466 = n2752 ^ n2724 ^ 1'b0 ;
  assign n9467 = n9466 ^ n7535 ^ n1964 ;
  assign n9465 = n1155 & ~n1363 ;
  assign n9468 = n9467 ^ n9465 ^ 1'b0 ;
  assign n9469 = n9464 | n9468 ;
  assign n9470 = n9469 ^ n666 ^ 1'b0 ;
  assign n9471 = n8559 & ~n9470 ;
  assign n9472 = n8687 ^ n6714 ^ n1759 ;
  assign n9473 = n9399 ^ n7807 ^ n6122 ;
  assign n9474 = ( n4816 & n9472 ) | ( n4816 & n9473 ) | ( n9472 & n9473 ) ;
  assign n9481 = n8740 ^ n1776 ^ n462 ;
  assign n9477 = n3271 ^ n1284 ^ 1'b0 ;
  assign n9478 = n1522 & ~n9477 ;
  assign n9475 = x200 | n2484 ;
  assign n9476 = n9475 ^ n2511 ^ n806 ;
  assign n9479 = n9478 ^ n9476 ^ n1598 ;
  assign n9480 = n6286 & n9479 ;
  assign n9482 = n9481 ^ n9480 ^ n2601 ;
  assign n9483 = n9482 ^ n1279 ^ n778 ;
  assign n9484 = n810 & ~n2430 ;
  assign n9485 = n9484 ^ n4959 ^ n2733 ;
  assign n9486 = n4914 ^ n3088 ^ n1345 ;
  assign n9487 = n9485 | n9486 ;
  assign n9497 = n6959 ^ n1374 ^ x130 ;
  assign n9489 = n6576 ^ n4747 ^ n2299 ;
  assign n9488 = n4341 ^ n1587 ^ 1'b0 ;
  assign n9490 = n9489 ^ n9488 ^ n7064 ;
  assign n9491 = n9490 ^ n6479 ^ n1402 ;
  assign n9492 = n2776 ^ n1739 ^ n804 ;
  assign n9493 = n9492 ^ n2956 ^ 1'b0 ;
  assign n9494 = ( x180 & n1299 ) | ( x180 & n6262 ) | ( n1299 & n6262 ) ;
  assign n9495 = ( n1371 & ~n8493 ) | ( n1371 & n9494 ) | ( ~n8493 & n9494 ) ;
  assign n9496 = ( n9491 & n9493 ) | ( n9491 & ~n9495 ) | ( n9493 & ~n9495 ) ;
  assign n9498 = n9497 ^ n9496 ^ n8667 ;
  assign n9501 = n2646 ^ n2237 ^ n2084 ;
  assign n9499 = n700 & n2063 ;
  assign n9500 = ( n7999 & ~n8399 ) | ( n7999 & n9499 ) | ( ~n8399 & n9499 ) ;
  assign n9502 = n9501 ^ n9500 ^ 1'b0 ;
  assign n9503 = n9498 & n9502 ;
  assign n9504 = n5195 ^ n1362 ^ n1286 ;
  assign n9505 = n6112 & n9504 ;
  assign n9506 = n969 | n9505 ;
  assign n9507 = n4948 | n9506 ;
  assign n9508 = ( n303 & n3882 ) | ( n303 & ~n9507 ) | ( n3882 & ~n9507 ) ;
  assign n9511 = n4161 & ~n8928 ;
  assign n9512 = n3580 & n9511 ;
  assign n9510 = n3982 ^ n1396 ^ n431 ;
  assign n9509 = n5805 ^ n350 ^ 1'b0 ;
  assign n9513 = n9512 ^ n9510 ^ n9509 ;
  assign n9517 = n7589 ^ n5485 ^ 1'b0 ;
  assign n9514 = n2455 ^ n1923 ^ 1'b0 ;
  assign n9515 = ( n1357 & ~n1500 ) | ( n1357 & n5255 ) | ( ~n1500 & n5255 ) ;
  assign n9516 = ( n1867 & ~n9514 ) | ( n1867 & n9515 ) | ( ~n9514 & n9515 ) ;
  assign n9518 = n9517 ^ n9516 ^ n2993 ;
  assign n9519 = ~n2009 & n9518 ;
  assign n9523 = n3372 ^ n2987 ^ n2383 ;
  assign n9520 = ( n2800 & ~n3336 ) | ( n2800 & n5982 ) | ( ~n3336 & n5982 ) ;
  assign n9521 = n2730 ^ x55 ^ 1'b0 ;
  assign n9522 = ~n9520 & n9521 ;
  assign n9524 = n9523 ^ n9522 ^ 1'b0 ;
  assign n9525 = ( ~n1840 & n8825 ) | ( ~n1840 & n9524 ) | ( n8825 & n9524 ) ;
  assign n9526 = n7787 ^ n4180 ^ 1'b0 ;
  assign n9527 = n7655 & n9526 ;
  assign n9528 = ( n2501 & n4206 ) | ( n2501 & n9527 ) | ( n4206 & n9527 ) ;
  assign n9529 = n6905 ^ n3337 ^ n699 ;
  assign n9530 = n4530 ^ n542 ^ x201 ;
  assign n9531 = ( n8908 & ~n9529 ) | ( n8908 & n9530 ) | ( ~n9529 & n9530 ) ;
  assign n9532 = ~n5258 & n7810 ;
  assign n9533 = n9532 ^ n6714 ^ n3118 ;
  assign n9534 = n2735 & n9120 ;
  assign n9535 = n9534 ^ n2138 ^ 1'b0 ;
  assign n9536 = ~n1511 & n3951 ;
  assign n9537 = n9535 & n9536 ;
  assign n9538 = n7742 & ~n9537 ;
  assign n9539 = n9538 ^ n8961 ^ 1'b0 ;
  assign n9540 = n2877 ^ n364 ^ x117 ;
  assign n9541 = n9540 ^ n2005 ^ 1'b0 ;
  assign n9542 = ~n3635 & n9541 ;
  assign n9543 = ( n5956 & n9411 ) | ( n5956 & ~n9542 ) | ( n9411 & ~n9542 ) ;
  assign n9544 = n270 & n1152 ;
  assign n9545 = n396 & n9544 ;
  assign n9546 = n9545 ^ n5160 ^ n2152 ;
  assign n9547 = n6266 | n9012 ;
  assign n9548 = n6286 | n9547 ;
  assign n9549 = n8690 ^ n2017 ^ n1261 ;
  assign n9550 = n7455 ^ n1036 ^ n1023 ;
  assign n9551 = ( n3528 & ~n5013 ) | ( n3528 & n9550 ) | ( ~n5013 & n9550 ) ;
  assign n9552 = n956 | n9551 ;
  assign n9553 = n5638 | n9552 ;
  assign n9554 = ( n9548 & n9549 ) | ( n9548 & ~n9553 ) | ( n9549 & ~n9553 ) ;
  assign n9555 = n6874 ^ n5374 ^ n5022 ;
  assign n9556 = ~n1428 & n3154 ;
  assign n9557 = ( n6830 & n9555 ) | ( n6830 & ~n9556 ) | ( n9555 & ~n9556 ) ;
  assign n9558 = n4667 & ~n9557 ;
  assign n9559 = ~n4688 & n9558 ;
  assign n9560 = n8127 ^ n7538 ^ n5221 ;
  assign n9561 = ( x149 & n9559 ) | ( x149 & ~n9560 ) | ( n9559 & ~n9560 ) ;
  assign n9562 = n3270 & ~n9107 ;
  assign n9563 = n9562 ^ n2789 ^ 1'b0 ;
  assign n9564 = n9563 ^ n4305 ^ 1'b0 ;
  assign n9565 = n9564 ^ n6657 ^ n537 ;
  assign n9566 = n1698 ^ n1336 ^ n271 ;
  assign n9567 = ( ~n672 & n1183 ) | ( ~n672 & n1623 ) | ( n1183 & n1623 ) ;
  assign n9568 = n9567 ^ n2566 ^ 1'b0 ;
  assign n9569 = ( n2130 & n9566 ) | ( n2130 & ~n9568 ) | ( n9566 & ~n9568 ) ;
  assign n9575 = n690 | n2041 ;
  assign n9574 = ( x86 & ~n1636 ) | ( x86 & n6304 ) | ( ~n1636 & n6304 ) ;
  assign n9570 = ~n2221 & n7468 ;
  assign n9571 = ~n8118 & n9570 ;
  assign n9572 = n9571 ^ n2090 ^ n462 ;
  assign n9573 = ( n595 & n3369 ) | ( n595 & n9572 ) | ( n3369 & n9572 ) ;
  assign n9576 = n9575 ^ n9574 ^ n9573 ;
  assign n9577 = ( ~n8528 & n9569 ) | ( ~n8528 & n9576 ) | ( n9569 & n9576 ) ;
  assign n9599 = n540 ^ x205 ^ 1'b0 ;
  assign n9600 = n1685 & n9599 ;
  assign n9601 = n9600 ^ n704 ^ 1'b0 ;
  assign n9602 = n2519 & n4721 ;
  assign n9603 = n1860 | n3110 ;
  assign n9604 = n9603 ^ n3427 ^ 1'b0 ;
  assign n9605 = ~x93 & n9604 ;
  assign n9613 = n6955 ^ n2458 ^ n1899 ;
  assign n9610 = n631 & n7645 ;
  assign n9606 = ( n2356 & n3764 ) | ( n2356 & n5331 ) | ( n3764 & n5331 ) ;
  assign n9607 = n742 & ~n2100 ;
  assign n9608 = n9607 ^ n864 ^ 1'b0 ;
  assign n9609 = ( ~n4219 & n9606 ) | ( ~n4219 & n9608 ) | ( n9606 & n9608 ) ;
  assign n9611 = n9610 ^ n9609 ^ n3020 ;
  assign n9612 = ( ~n2191 & n2821 ) | ( ~n2191 & n9611 ) | ( n2821 & n9611 ) ;
  assign n9614 = n9613 ^ n9612 ^ n6813 ;
  assign n9615 = ( n9602 & ~n9605 ) | ( n9602 & n9614 ) | ( ~n9605 & n9614 ) ;
  assign n9616 = ( n2348 & n9601 ) | ( n2348 & ~n9615 ) | ( n9601 & ~n9615 ) ;
  assign n9594 = ( n1418 & n1904 ) | ( n1418 & ~n6813 ) | ( n1904 & ~n6813 ) ;
  assign n9595 = ( n974 & ~n1425 ) | ( n974 & n1776 ) | ( ~n1425 & n1776 ) ;
  assign n9596 = n4721 ^ n3018 ^ n2436 ;
  assign n9597 = n9596 ^ n874 ^ x195 ;
  assign n9598 = ( n9594 & n9595 ) | ( n9594 & n9597 ) | ( n9595 & n9597 ) ;
  assign n9581 = n1580 & ~n3561 ;
  assign n9582 = n2322 & n9581 ;
  assign n9583 = n9582 ^ n2563 ^ 1'b0 ;
  assign n9578 = ( n269 & n2493 ) | ( n269 & ~n5128 ) | ( n2493 & ~n5128 ) ;
  assign n9579 = ( n1193 & n3345 ) | ( n1193 & n9578 ) | ( n3345 & n9578 ) ;
  assign n9580 = n5041 & n9579 ;
  assign n9584 = n9583 ^ n9580 ^ 1'b0 ;
  assign n9585 = ( n2195 & n3474 ) | ( n2195 & ~n9584 ) | ( n3474 & ~n9584 ) ;
  assign n9586 = n9585 ^ n4973 ^ 1'b0 ;
  assign n9587 = ( n613 & ~n2399 ) | ( n613 & n3619 ) | ( ~n2399 & n3619 ) ;
  assign n9588 = ( n525 & ~n6228 ) | ( n525 & n9587 ) | ( ~n6228 & n9587 ) ;
  assign n9589 = n6199 ^ n2231 ^ x181 ;
  assign n9590 = n2628 ^ n658 ^ 1'b0 ;
  assign n9591 = ~n9589 & n9590 ;
  assign n9592 = n9588 & n9591 ;
  assign n9593 = ~n9586 & n9592 ;
  assign n9617 = n9616 ^ n9598 ^ n9593 ;
  assign n9619 = ( ~n2444 & n3592 ) | ( ~n2444 & n8699 ) | ( n3592 & n8699 ) ;
  assign n9620 = n9619 ^ n2200 ^ n2032 ;
  assign n9618 = n4966 | n8682 ;
  assign n9621 = n9620 ^ n9618 ^ 1'b0 ;
  assign n9622 = ~n3029 & n8957 ;
  assign n9623 = n9622 ^ n3616 ^ 1'b0 ;
  assign n9624 = n6114 ^ n4341 ^ n3326 ;
  assign n9625 = n9624 ^ n4546 ^ n4513 ;
  assign n9626 = ~n9623 & n9625 ;
  assign n9627 = n9626 ^ n2027 ^ 1'b0 ;
  assign n9628 = ( n1766 & ~n7170 ) | ( n1766 & n8245 ) | ( ~n7170 & n8245 ) ;
  assign n9632 = n4685 ^ n2173 ^ n2003 ;
  assign n9629 = n8228 ^ n3023 ^ n2862 ;
  assign n9630 = ( n1113 & ~n1623 ) | ( n1113 & n7394 ) | ( ~n1623 & n7394 ) ;
  assign n9631 = ( n6022 & n9629 ) | ( n6022 & n9630 ) | ( n9629 & n9630 ) ;
  assign n9633 = n9632 ^ n9631 ^ n5742 ;
  assign n9634 = ( n9627 & n9628 ) | ( n9627 & n9633 ) | ( n9628 & n9633 ) ;
  assign n9635 = x66 & ~x227 ;
  assign n9636 = n635 | n9635 ;
  assign n9637 = n1410 & n7483 ;
  assign n9638 = x192 & n9637 ;
  assign n9639 = ~n8837 & n9638 ;
  assign n9640 = n3275 ^ n2451 ^ n905 ;
  assign n9641 = n1026 ^ n658 ^ 1'b0 ;
  assign n9642 = ( n2991 & ~n9640 ) | ( n2991 & n9641 ) | ( ~n9640 & n9641 ) ;
  assign n9643 = n9642 ^ n8481 ^ 1'b0 ;
  assign n9644 = n9639 | n9643 ;
  assign n9645 = ~n3501 & n7808 ;
  assign n9646 = n8885 ^ n3844 ^ n1242 ;
  assign n9647 = ( ~n3501 & n3505 ) | ( ~n3501 & n9646 ) | ( n3505 & n9646 ) ;
  assign n9648 = n9226 ^ n2815 ^ n883 ;
  assign n9649 = n9648 ^ n8501 ^ n5884 ;
  assign n9650 = n9649 ^ n1046 ^ 1'b0 ;
  assign n9651 = ~n2966 & n9650 ;
  assign n9652 = n6936 ^ n4684 ^ n1020 ;
  assign n9653 = ( n1690 & ~n3924 ) | ( n1690 & n7334 ) | ( ~n3924 & n7334 ) ;
  assign n9654 = n2880 & ~n5903 ;
  assign n9655 = ( x246 & ~n8103 ) | ( x246 & n9654 ) | ( ~n8103 & n9654 ) ;
  assign n9656 = ~n2457 & n9655 ;
  assign n9657 = n9656 ^ n2977 ^ 1'b0 ;
  assign n9658 = n9657 ^ n6870 ^ n2787 ;
  assign n9659 = ( n1900 & n9653 ) | ( n1900 & ~n9658 ) | ( n9653 & ~n9658 ) ;
  assign n9660 = n2929 ^ n2506 ^ n1957 ;
  assign n9661 = ( ~n387 & n1908 ) | ( ~n387 & n9660 ) | ( n1908 & n9660 ) ;
  assign n9662 = ( n579 & ~n5035 ) | ( n579 & n9661 ) | ( ~n5035 & n9661 ) ;
  assign n9663 = ( n1991 & n6531 ) | ( n1991 & ~n9662 ) | ( n6531 & ~n9662 ) ;
  assign n9666 = n1322 ^ n1159 ^ x76 ;
  assign n9667 = n6629 ^ n1282 ^ 1'b0 ;
  assign n9668 = n9666 & n9667 ;
  assign n9665 = ( n3946 & ~n8977 ) | ( n3946 & n9660 ) | ( ~n8977 & n9660 ) ;
  assign n9664 = n7513 ^ n5275 ^ 1'b0 ;
  assign n9669 = n9668 ^ n9665 ^ n9664 ;
  assign n9670 = ( ~x188 & n1714 ) | ( ~x188 & n5549 ) | ( n1714 & n5549 ) ;
  assign n9671 = n9670 ^ n8691 ^ x125 ;
  assign n9672 = ( n3683 & n5144 ) | ( n3683 & ~n8297 ) | ( n5144 & ~n8297 ) ;
  assign n9673 = n4622 ^ n3888 ^ n705 ;
  assign n9674 = n9673 ^ n6881 ^ n4296 ;
  assign n9675 = n1565 & n5806 ;
  assign n9676 = n4841 & n9675 ;
  assign n9677 = ( n7104 & n7430 ) | ( n7104 & ~n9104 ) | ( n7430 & ~n9104 ) ;
  assign n9678 = ( n1641 & n2597 ) | ( n1641 & ~n9677 ) | ( n2597 & ~n9677 ) ;
  assign n9679 = ( n3481 & n9676 ) | ( n3481 & ~n9678 ) | ( n9676 & ~n9678 ) ;
  assign n9685 = ( n1599 & n5237 ) | ( n1599 & ~n9619 ) | ( n5237 & ~n9619 ) ;
  assign n9683 = n5874 ^ n3506 ^ n1562 ;
  assign n9680 = ( n3819 & n4224 ) | ( n3819 & ~n6117 ) | ( n4224 & ~n6117 ) ;
  assign n9681 = n9680 ^ n1113 ^ 1'b0 ;
  assign n9682 = n6485 & n9681 ;
  assign n9684 = n9683 ^ n9682 ^ n8850 ;
  assign n9686 = n9685 ^ n9684 ^ n7384 ;
  assign n9697 = ( n2097 & n4134 ) | ( n2097 & n5367 ) | ( n4134 & n5367 ) ;
  assign n9687 = n5207 ^ n3653 ^ 1'b0 ;
  assign n9688 = n7613 & ~n9687 ;
  assign n9689 = n6539 ^ n4082 ^ n3552 ;
  assign n9693 = n1810 ^ n963 ^ 1'b0 ;
  assign n9690 = n1707 & ~n3484 ;
  assign n9691 = n9690 ^ x25 ^ 1'b0 ;
  assign n9692 = n9691 ^ n3162 ^ n1505 ;
  assign n9694 = n9693 ^ n9692 ^ n3898 ;
  assign n9695 = ~n9689 & n9694 ;
  assign n9696 = ( n9252 & n9688 ) | ( n9252 & ~n9695 ) | ( n9688 & ~n9695 ) ;
  assign n9698 = n9697 ^ n9696 ^ n503 ;
  assign n9699 = n6966 ^ n5994 ^ n1343 ;
  assign n9700 = n9699 ^ n3810 ^ 1'b0 ;
  assign n9701 = n9576 & n9700 ;
  assign n9702 = n9173 ^ n5854 ^ n3236 ;
  assign n9703 = n3750 & n7467 ;
  assign n9704 = n673 & n6330 ;
  assign n9705 = ~n9703 & n9704 ;
  assign n9706 = n6371 ^ n5929 ^ n4084 ;
  assign n9707 = n2145 & ~n5531 ;
  assign n9708 = ~n9706 & n9707 ;
  assign n9709 = ( n1272 & n5307 ) | ( n1272 & n5840 ) | ( n5307 & n5840 ) ;
  assign n9712 = n4077 ^ n3749 ^ 1'b0 ;
  assign n9713 = ( ~n6223 & n6910 ) | ( ~n6223 & n9712 ) | ( n6910 & n9712 ) ;
  assign n9714 = n9713 ^ n3939 ^ n1418 ;
  assign n9710 = ( n694 & n2379 ) | ( n694 & ~n8438 ) | ( n2379 & ~n8438 ) ;
  assign n9711 = n9710 ^ n5759 ^ n3087 ;
  assign n9715 = n9714 ^ n9711 ^ 1'b0 ;
  assign n9716 = n4391 & ~n4481 ;
  assign n9717 = n9716 ^ n1295 ^ 1'b0 ;
  assign n9718 = n9717 ^ n4959 ^ 1'b0 ;
  assign n9719 = ( ~n7883 & n9057 ) | ( ~n7883 & n9718 ) | ( n9057 & n9718 ) ;
  assign n9720 = ( ~n914 & n1499 ) | ( ~n914 & n2031 ) | ( n1499 & n2031 ) ;
  assign n9721 = ~n5007 & n9177 ;
  assign n9722 = n9720 & n9721 ;
  assign n9723 = n3792 ^ n1402 ^ n1066 ;
  assign n9724 = n1233 & ~n2050 ;
  assign n9725 = n9724 ^ n6519 ^ 1'b0 ;
  assign n9726 = n997 & ~n2319 ;
  assign n9727 = ~n4759 & n9726 ;
  assign n9728 = n9727 ^ n4812 ^ x108 ;
  assign n9729 = ( n3118 & n9725 ) | ( n3118 & ~n9728 ) | ( n9725 & ~n9728 ) ;
  assign n9730 = ( n9722 & n9723 ) | ( n9722 & n9729 ) | ( n9723 & n9729 ) ;
  assign n9731 = n8216 ^ n655 ^ x34 ;
  assign n9732 = n5668 ^ n1872 ^ 1'b0 ;
  assign n9733 = n9732 ^ n9231 ^ n5971 ;
  assign n9734 = ( n394 & ~n5251 ) | ( n394 & n6621 ) | ( ~n5251 & n6621 ) ;
  assign n9735 = n9734 ^ n1796 ^ n1009 ;
  assign n9736 = x92 & n1534 ;
  assign n9737 = ~n9735 & n9736 ;
  assign n9738 = ( n5398 & ~n5640 ) | ( n5398 & n7385 ) | ( ~n5640 & n7385 ) ;
  assign n9744 = n7059 ^ n993 ^ 1'b0 ;
  assign n9740 = n1809 & n2731 ;
  assign n9741 = n9740 ^ n2520 ^ 1'b0 ;
  assign n9739 = ~n2099 & n2747 ;
  assign n9742 = n9741 ^ n9739 ^ 1'b0 ;
  assign n9743 = x179 & n9742 ;
  assign n9745 = n9744 ^ n9743 ^ n5102 ;
  assign n9746 = ( n9737 & ~n9738 ) | ( n9737 & n9745 ) | ( ~n9738 & n9745 ) ;
  assign n9747 = x95 & ~n9564 ;
  assign n9748 = n9747 ^ n3300 ^ 1'b0 ;
  assign n9749 = ~n1581 & n9748 ;
  assign n9750 = ( n628 & n1635 ) | ( n628 & n5230 ) | ( n1635 & n5230 ) ;
  assign n9751 = n2388 | n8907 ;
  assign n9752 = n9751 ^ n3930 ^ 1'b0 ;
  assign n9753 = n3576 ^ n2162 ^ n1710 ;
  assign n9754 = ( n6306 & n9699 ) | ( n6306 & n9753 ) | ( n9699 & n9753 ) ;
  assign n9755 = ( n9750 & n9752 ) | ( n9750 & ~n9754 ) | ( n9752 & ~n9754 ) ;
  assign n9756 = n8501 ^ n4478 ^ n2789 ;
  assign n9757 = n9756 ^ n861 ^ 1'b0 ;
  assign n9758 = n3203 & ~n9757 ;
  assign n9759 = n9758 ^ n7090 ^ 1'b0 ;
  assign n9760 = n2590 ^ n2035 ^ n1706 ;
  assign n9761 = n9760 ^ n5470 ^ x241 ;
  assign n9762 = x157 & n9761 ;
  assign n9765 = x87 & ~n912 ;
  assign n9766 = n9765 ^ n5150 ^ 1'b0 ;
  assign n9767 = n6237 ^ n3188 ^ n785 ;
  assign n9768 = n9767 ^ n974 ^ 1'b0 ;
  assign n9769 = n9766 & n9768 ;
  assign n9763 = n5000 ^ n1651 ^ n1636 ;
  assign n9764 = n9763 ^ n7021 ^ 1'b0 ;
  assign n9770 = n9769 ^ n9764 ^ n1550 ;
  assign n9781 = ~x5 & n1059 ;
  assign n9778 = n1486 | n6194 ;
  assign n9779 = n272 | n9778 ;
  assign n9780 = ( n838 & n4057 ) | ( n838 & n9779 ) | ( n4057 & n9779 ) ;
  assign n9782 = n9781 ^ n9780 ^ n1583 ;
  assign n9775 = n1620 | n6775 ;
  assign n9776 = n385 & ~n9775 ;
  assign n9771 = ( n1463 & n1623 ) | ( n1463 & ~n3852 ) | ( n1623 & ~n3852 ) ;
  assign n9772 = n9771 ^ n6549 ^ n5724 ;
  assign n9773 = ( n3618 & n5128 ) | ( n3618 & n9772 ) | ( n5128 & n9772 ) ;
  assign n9774 = n4637 & n9773 ;
  assign n9777 = n9776 ^ n9774 ^ 1'b0 ;
  assign n9783 = n9782 ^ n9777 ^ n9331 ;
  assign n9784 = ~n1082 & n9783 ;
  assign n9785 = ~n1282 & n9784 ;
  assign n9786 = n4010 | n6410 ;
  assign n9787 = ( n4341 & n5110 ) | ( n4341 & n9786 ) | ( n5110 & n9786 ) ;
  assign n9788 = n9787 ^ n6164 ^ n4730 ;
  assign n9791 = n5722 ^ n2102 ^ n1971 ;
  assign n9789 = n2919 & n9206 ;
  assign n9790 = n9789 ^ n6533 ^ n4739 ;
  assign n9792 = n9791 ^ n9790 ^ n578 ;
  assign n9793 = ( n5080 & ~n9788 ) | ( n5080 & n9792 ) | ( ~n9788 & n9792 ) ;
  assign n9794 = n9793 ^ n6024 ^ x151 ;
  assign n9795 = n7829 ^ n3029 ^ n654 ;
  assign n9796 = n7168 | n9629 ;
  assign n9797 = n9796 ^ n5335 ^ n3015 ;
  assign n9798 = n4745 ^ n2255 ^ 1'b0 ;
  assign n9799 = ( n6452 & n8121 ) | ( n6452 & n9798 ) | ( n8121 & n9798 ) ;
  assign n9800 = ( n6364 & n9797 ) | ( n6364 & ~n9799 ) | ( n9797 & ~n9799 ) ;
  assign n9805 = n3104 ^ n3079 ^ n1118 ;
  assign n9801 = ~x36 & n1381 ;
  assign n9802 = ~n6235 & n6248 ;
  assign n9803 = n9801 & n9802 ;
  assign n9804 = n9803 ^ n3702 ^ n1811 ;
  assign n9806 = n9805 ^ n9804 ^ 1'b0 ;
  assign n9809 = n3395 ^ n3390 ^ n2635 ;
  assign n9810 = ( n3797 & n5987 ) | ( n3797 & ~n9809 ) | ( n5987 & ~n9809 ) ;
  assign n9811 = ( n1240 & n2012 ) | ( n1240 & ~n9810 ) | ( n2012 & ~n9810 ) ;
  assign n9807 = n6946 & ~n7104 ;
  assign n9808 = n9807 ^ n7494 ^ n1553 ;
  assign n9812 = n9811 ^ n9808 ^ x189 ;
  assign n9813 = n3777 ^ n1910 ^ 1'b0 ;
  assign n9814 = n9813 ^ n948 ^ 1'b0 ;
  assign n9815 = n3119 & n9814 ;
  assign n9816 = n9166 ^ n4389 ^ n1616 ;
  assign n9817 = n7598 ^ n4362 ^ n2593 ;
  assign n9818 = n5246 & n9817 ;
  assign n9819 = ( x236 & n2561 ) | ( x236 & n3083 ) | ( n2561 & n3083 ) ;
  assign n9820 = ( n1017 & n3361 ) | ( n1017 & ~n9819 ) | ( n3361 & ~n9819 ) ;
  assign n9821 = n9820 ^ n2656 ^ n1964 ;
  assign n9822 = ( n4335 & ~n9372 ) | ( n4335 & n9821 ) | ( ~n9372 & n9821 ) ;
  assign n9823 = n9822 ^ n8968 ^ 1'b0 ;
  assign n9824 = ( ~n1701 & n9818 ) | ( ~n1701 & n9823 ) | ( n9818 & n9823 ) ;
  assign n9828 = n7765 ^ n704 ^ n641 ;
  assign n9825 = ( ~x254 & n1395 ) | ( ~x254 & n5634 ) | ( n1395 & n5634 ) ;
  assign n9826 = n9825 ^ n3605 ^ n952 ;
  assign n9827 = n9826 ^ n7489 ^ n1937 ;
  assign n9829 = n9828 ^ n9827 ^ n8396 ;
  assign n9830 = ( ~n9816 & n9824 ) | ( ~n9816 & n9829 ) | ( n9824 & n9829 ) ;
  assign n9831 = n7568 ^ n3291 ^ 1'b0 ;
  assign n9832 = n9831 ^ n1986 ^ n277 ;
  assign n9833 = ~n1792 & n2330 ;
  assign n9834 = n9833 ^ n4020 ^ n3938 ;
  assign n9835 = ( ~n647 & n7718 ) | ( ~n647 & n9834 ) | ( n7718 & n9834 ) ;
  assign n9836 = n9835 ^ n9161 ^ n7040 ;
  assign n9837 = n6936 ^ n359 ^ n296 ;
  assign n9838 = ( n5054 & n5698 ) | ( n5054 & n9837 ) | ( n5698 & n9837 ) ;
  assign n9844 = n3433 ^ n1987 ^ 1'b0 ;
  assign n9841 = n4061 ^ n2850 ^ n2563 ;
  assign n9842 = ( n652 & n1015 ) | ( n652 & ~n4665 ) | ( n1015 & ~n4665 ) ;
  assign n9843 = ( ~n5711 & n9841 ) | ( ~n5711 & n9842 ) | ( n9841 & n9842 ) ;
  assign n9845 = n9844 ^ n9843 ^ n3604 ;
  assign n9839 = n2248 | n6809 ;
  assign n9840 = n8013 | n9839 ;
  assign n9846 = n9845 ^ n9840 ^ 1'b0 ;
  assign n9847 = ( n768 & n5882 ) | ( n768 & n8150 ) | ( n5882 & n8150 ) ;
  assign n9848 = n2970 ^ n508 ^ 1'b0 ;
  assign n9849 = ( n3287 & ~n3377 ) | ( n3287 & n9848 ) | ( ~n3377 & n9848 ) ;
  assign n9850 = n9849 ^ n7168 ^ n4061 ;
  assign n9853 = ( x135 & n1289 ) | ( x135 & ~n2312 ) | ( n1289 & ~n2312 ) ;
  assign n9851 = ( ~n3922 & n4115 ) | ( ~n3922 & n5017 ) | ( n4115 & n5017 ) ;
  assign n9852 = ( n6424 & ~n7940 ) | ( n6424 & n9851 ) | ( ~n7940 & n9851 ) ;
  assign n9854 = n9853 ^ n9852 ^ 1'b0 ;
  assign n9855 = n9850 | n9854 ;
  assign n9856 = n9855 ^ n7094 ^ n1956 ;
  assign n9857 = n6754 ^ n3825 ^ n1410 ;
  assign n9858 = ( n3126 & ~n6413 ) | ( n3126 & n9857 ) | ( ~n6413 & n9857 ) ;
  assign n9859 = n3591 | n9858 ;
  assign n9860 = n1394 & n7706 ;
  assign n9861 = ~n7039 & n9860 ;
  assign n9862 = n9859 & ~n9861 ;
  assign n9863 = n9469 & n9862 ;
  assign n9864 = n5094 & n5128 ;
  assign n9865 = ~n2929 & n9864 ;
  assign n9866 = n6154 & ~n9865 ;
  assign n9867 = n9866 ^ n6336 ^ x63 ;
  assign n9877 = ~n306 & n1635 ;
  assign n9878 = n9877 ^ n9111 ^ 1'b0 ;
  assign n9879 = ~n1077 & n9878 ;
  assign n9880 = ( ~x201 & n3428 ) | ( ~x201 & n9879 ) | ( n3428 & n9879 ) ;
  assign n9873 = ( x199 & n1062 ) | ( x199 & n7399 ) | ( n1062 & n7399 ) ;
  assign n9871 = n5950 ^ n3523 ^ n432 ;
  assign n9872 = n9871 ^ n4701 ^ n1822 ;
  assign n9874 = n9873 ^ n9872 ^ n576 ;
  assign n9875 = n9874 ^ n9209 ^ 1'b0 ;
  assign n9869 = n6955 ^ n3678 ^ 1'b0 ;
  assign n9870 = ~n8117 & n9869 ;
  assign n9876 = n9875 ^ n9870 ^ n1649 ;
  assign n9868 = n6232 ^ n2250 ^ 1'b0 ;
  assign n9881 = n9880 ^ n9876 ^ n9868 ;
  assign n9884 = n4307 ^ n3109 ^ x53 ;
  assign n9885 = n9884 ^ n6740 ^ n3933 ;
  assign n9886 = n9885 ^ n1619 ^ x8 ;
  assign n9882 = n2922 ^ n1916 ^ n1242 ;
  assign n9883 = n9882 ^ n1698 ^ 1'b0 ;
  assign n9887 = n9886 ^ n9883 ^ n5251 ;
  assign n9888 = n9887 ^ n9769 ^ 1'b0 ;
  assign n9889 = n2100 | n9888 ;
  assign n9890 = ( x221 & n1769 ) | ( x221 & ~n3570 ) | ( n1769 & ~n3570 ) ;
  assign n9891 = ~n6425 & n9890 ;
  assign n9892 = n9891 ^ n1695 ^ 1'b0 ;
  assign n9898 = n2056 & ~n3148 ;
  assign n9899 = n6399 ^ n1414 ^ x160 ;
  assign n9900 = n9899 ^ n5891 ^ n4487 ;
  assign n9904 = n7334 ^ n5477 ^ n2971 ;
  assign n9903 = n3149 ^ n926 ^ x229 ;
  assign n9901 = ( n1968 & n3606 ) | ( n1968 & ~n3651 ) | ( n3606 & ~n3651 ) ;
  assign n9902 = ( ~n1391 & n4317 ) | ( ~n1391 & n9901 ) | ( n4317 & n9901 ) ;
  assign n9905 = n9904 ^ n9903 ^ n9902 ;
  assign n9906 = ( n9898 & n9900 ) | ( n9898 & ~n9905 ) | ( n9900 & ~n9905 ) ;
  assign n9896 = ( n867 & ~n3074 ) | ( n867 & n3478 ) | ( ~n3074 & n3478 ) ;
  assign n9895 = ~n1097 & n1135 ;
  assign n9897 = n9896 ^ n9895 ^ 1'b0 ;
  assign n9907 = n9906 ^ n9897 ^ n9195 ;
  assign n9893 = n5090 ^ n2465 ^ x25 ;
  assign n9894 = n8186 & n9893 ;
  assign n9908 = n9907 ^ n9894 ^ 1'b0 ;
  assign n9909 = ( ~n6149 & n9892 ) | ( ~n6149 & n9908 ) | ( n9892 & n9908 ) ;
  assign n9914 = ( n2247 & ~n3613 ) | ( n2247 & n6292 ) | ( ~n3613 & n6292 ) ;
  assign n9911 = n1030 ^ x100 ^ 1'b0 ;
  assign n9912 = ( n1236 & n6576 ) | ( n1236 & n9911 ) | ( n6576 & n9911 ) ;
  assign n9913 = ( n2296 & n7034 ) | ( n2296 & n9912 ) | ( n7034 & n9912 ) ;
  assign n9915 = n9914 ^ n9913 ^ n2700 ;
  assign n9910 = n9341 ^ n7836 ^ 1'b0 ;
  assign n9916 = n9915 ^ n9910 ^ 1'b0 ;
  assign n9917 = n9571 ^ n6393 ^ n3722 ;
  assign n9918 = n9917 ^ n8992 ^ n1577 ;
  assign n9919 = ( n685 & ~n2046 ) | ( n685 & n3106 ) | ( ~n2046 & n3106 ) ;
  assign n9920 = ( n3789 & n4307 ) | ( n3789 & n9646 ) | ( n4307 & n9646 ) ;
  assign n9921 = n7450 | n9920 ;
  assign n9924 = n8007 ^ n3693 ^ n3282 ;
  assign n9922 = n8147 ^ n6752 ^ n6387 ;
  assign n9923 = n5274 & ~n9922 ;
  assign n9925 = n9924 ^ n9923 ^ n8617 ;
  assign n9926 = n6326 | n8833 ;
  assign n9927 = ~n1791 & n9926 ;
  assign n9928 = n6810 ^ n6371 ^ n6110 ;
  assign n9929 = ( n4516 & ~n5178 ) | ( n4516 & n9026 ) | ( ~n5178 & n9026 ) ;
  assign n9933 = n3147 ^ n798 ^ n279 ;
  assign n9930 = n5108 ^ n3725 ^ n2741 ;
  assign n9931 = n7189 & ~n9273 ;
  assign n9932 = ( n7026 & n9930 ) | ( n7026 & n9931 ) | ( n9930 & n9931 ) ;
  assign n9934 = n9933 ^ n9932 ^ 1'b0 ;
  assign n9935 = ( n1839 & ~n4841 ) | ( n1839 & n7997 ) | ( ~n4841 & n7997 ) ;
  assign n9936 = ( n996 & ~n6752 ) | ( n996 & n9935 ) | ( ~n6752 & n9935 ) ;
  assign n9937 = n7482 ^ n5317 ^ n781 ;
  assign n9938 = ( x236 & n4454 ) | ( x236 & n9937 ) | ( n4454 & n9937 ) ;
  assign n9939 = n4109 & ~n9938 ;
  assign n9940 = ~n3035 & n9939 ;
  assign n9941 = n3041 ^ n1021 ^ x235 ;
  assign n9942 = ( n6010 & n8770 ) | ( n6010 & ~n9941 ) | ( n8770 & ~n9941 ) ;
  assign n9943 = ( n2382 & n9940 ) | ( n2382 & ~n9942 ) | ( n9940 & ~n9942 ) ;
  assign n9944 = ( x113 & n681 ) | ( x113 & n2042 ) | ( n681 & n2042 ) ;
  assign n9945 = ( n1986 & ~n5171 ) | ( n1986 & n9944 ) | ( ~n5171 & n9944 ) ;
  assign n9946 = n9945 ^ n5724 ^ 1'b0 ;
  assign n9947 = n3437 & ~n9946 ;
  assign n9949 = ( n1016 & n1923 ) | ( n1016 & n4687 ) | ( n1923 & n4687 ) ;
  assign n9948 = n3533 & n9318 ;
  assign n9950 = n9949 ^ n9948 ^ 1'b0 ;
  assign n9958 = n6182 ^ n1812 ^ n1256 ;
  assign n9959 = n4443 ^ n3477 ^ 1'b0 ;
  assign n9960 = n9958 & ~n9959 ;
  assign n9957 = ~n6541 & n6979 ;
  assign n9961 = n9960 ^ n9957 ^ 1'b0 ;
  assign n9969 = n6690 ^ n724 ^ n582 ;
  assign n9970 = n9969 ^ n3458 ^ n1885 ;
  assign n9964 = n3548 | n6137 ;
  assign n9965 = n9964 ^ n5700 ^ 1'b0 ;
  assign n9966 = n9965 ^ n3083 ^ n2894 ;
  assign n9962 = ( ~n595 & n1450 ) | ( ~n595 & n1800 ) | ( n1450 & n1800 ) ;
  assign n9963 = ~n6044 & n9962 ;
  assign n9967 = n9966 ^ n9963 ^ 1'b0 ;
  assign n9968 = ~n1064 & n9967 ;
  assign n9971 = n9970 ^ n9968 ^ 1'b0 ;
  assign n9972 = n9961 | n9971 ;
  assign n9951 = ( n996 & ~n1034 ) | ( n996 & n3168 ) | ( ~n1034 & n3168 ) ;
  assign n9952 = ( ~n2577 & n7331 ) | ( ~n2577 & n9951 ) | ( n7331 & n9951 ) ;
  assign n9954 = ( ~n2609 & n5162 ) | ( ~n2609 & n9418 ) | ( n5162 & n9418 ) ;
  assign n9953 = ( x31 & n5048 ) | ( x31 & ~n7306 ) | ( n5048 & ~n7306 ) ;
  assign n9955 = n9954 ^ n9953 ^ n2092 ;
  assign n9956 = n9952 & ~n9955 ;
  assign n9973 = n9972 ^ n9956 ^ 1'b0 ;
  assign n9974 = n4159 & n4988 ;
  assign n9975 = n4029 ^ n811 ^ 1'b0 ;
  assign n9976 = n9974 | n9975 ;
  assign n9977 = ( n4289 & n7222 ) | ( n4289 & ~n9976 ) | ( n7222 & ~n9976 ) ;
  assign n9978 = n3542 ^ x37 ^ 1'b0 ;
  assign n9979 = x59 & n9978 ;
  assign n9980 = n9979 ^ n464 ^ 1'b0 ;
  assign n9981 = ( x161 & n951 ) | ( x161 & ~n7887 ) | ( n951 & ~n7887 ) ;
  assign n9982 = n6843 ^ n2448 ^ n2339 ;
  assign n9983 = ~n480 & n1586 ;
  assign n9984 = n9983 ^ n5519 ^ 1'b0 ;
  assign n9985 = n9984 ^ n1784 ^ 1'b0 ;
  assign n9986 = ~n9982 & n9985 ;
  assign n9987 = ~n3439 & n8260 ;
  assign n9988 = ~n9986 & n9987 ;
  assign n9989 = ( n9980 & n9981 ) | ( n9980 & ~n9988 ) | ( n9981 & ~n9988 ) ;
  assign n9991 = n3798 ^ n2179 ^ n952 ;
  assign n9990 = n4862 ^ n2690 ^ n1179 ;
  assign n9992 = n9991 ^ n9990 ^ n5077 ;
  assign n9993 = n9550 ^ n6543 ^ n5757 ;
  assign n9994 = n9993 ^ n9157 ^ n4188 ;
  assign n9995 = ~n3612 & n8871 ;
  assign n9996 = n9995 ^ n4635 ^ n1710 ;
  assign n9997 = ( ~n7757 & n8247 ) | ( ~n7757 & n9996 ) | ( n8247 & n9996 ) ;
  assign n9998 = n1062 | n9997 ;
  assign n10001 = n2129 ^ n800 ^ 1'b0 ;
  assign n10000 = n7921 ^ n7819 ^ n2530 ;
  assign n10002 = n10001 ^ n10000 ^ n3726 ;
  assign n9999 = ( n973 & n4970 ) | ( n973 & ~n9685 ) | ( n4970 & ~n9685 ) ;
  assign n10003 = n10002 ^ n9999 ^ n2235 ;
  assign n10004 = ( ~n647 & n2606 ) | ( ~n647 & n7992 ) | ( n2606 & n7992 ) ;
  assign n10005 = ( ~n904 & n3200 ) | ( ~n904 & n10004 ) | ( n3200 & n10004 ) ;
  assign n10014 = ( n2738 & n3999 ) | ( n2738 & n8784 ) | ( n3999 & n8784 ) ;
  assign n10015 = ( ~n2744 & n3682 ) | ( ~n2744 & n5706 ) | ( n3682 & n5706 ) ;
  assign n10016 = n10014 | n10015 ;
  assign n10017 = n5107 & ~n10016 ;
  assign n10018 = ( n1872 & n6829 ) | ( n1872 & n10017 ) | ( n6829 & n10017 ) ;
  assign n10006 = n6121 ^ n4204 ^ n2946 ;
  assign n10008 = n1048 & n4903 ;
  assign n10009 = n10008 ^ n8034 ^ 1'b0 ;
  assign n10010 = n3370 & ~n10009 ;
  assign n10007 = ( n3294 & ~n4157 ) | ( n3294 & n7156 ) | ( ~n4157 & n7156 ) ;
  assign n10011 = n10010 ^ n10007 ^ n1405 ;
  assign n10012 = ( n2615 & ~n3629 ) | ( n2615 & n10011 ) | ( ~n3629 & n10011 ) ;
  assign n10013 = n10006 & ~n10012 ;
  assign n10019 = n10018 ^ n10013 ^ 1'b0 ;
  assign n10020 = ~n5696 & n10019 ;
  assign n10021 = n10005 & n10020 ;
  assign n10022 = n7168 ^ n3298 ^ n3167 ;
  assign n10023 = n4874 ^ n4375 ^ n964 ;
  assign n10024 = n8920 & ~n10023 ;
  assign n10025 = ( n3356 & n10022 ) | ( n3356 & n10024 ) | ( n10022 & n10024 ) ;
  assign n10026 = ( n1169 & n6907 ) | ( n1169 & ~n7913 ) | ( n6907 & ~n7913 ) ;
  assign n10028 = ( x97 & ~n1459 ) | ( x97 & n2330 ) | ( ~n1459 & n2330 ) ;
  assign n10029 = n10028 ^ n4874 ^ n669 ;
  assign n10027 = ~n7471 & n8914 ;
  assign n10030 = n10029 ^ n10027 ^ 1'b0 ;
  assign n10032 = n3557 & ~n8428 ;
  assign n10033 = ~n4227 & n10032 ;
  assign n10034 = n868 | n10033 ;
  assign n10035 = n4840 | n10034 ;
  assign n10031 = n7363 ^ n795 ^ x174 ;
  assign n10036 = n10035 ^ n10031 ^ n3200 ;
  assign n10037 = ~n1610 & n5812 ;
  assign n10038 = n6822 ^ n3901 ^ n864 ;
  assign n10039 = ( ~n10036 & n10037 ) | ( ~n10036 & n10038 ) | ( n10037 & n10038 ) ;
  assign n10040 = n821 & n5985 ;
  assign n10041 = n10040 ^ n9653 ^ n7423 ;
  assign n10055 = n7245 ^ n2521 ^ n1501 ;
  assign n10043 = n6562 ^ n1198 ^ 1'b0 ;
  assign n10044 = ( n2988 & n9524 ) | ( n2988 & n10043 ) | ( n9524 & n10043 ) ;
  assign n10051 = n4980 ^ n2962 ^ 1'b0 ;
  assign n10052 = n4391 & n10051 ;
  assign n10046 = ( x4 & n1827 ) | ( x4 & n8760 ) | ( n1827 & n8760 ) ;
  assign n10047 = n10046 ^ n4775 ^ 1'b0 ;
  assign n10048 = n6213 ^ n6207 ^ n1435 ;
  assign n10049 = ( n3300 & n10047 ) | ( n3300 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10050 = n10049 ^ n5894 ^ 1'b0 ;
  assign n10045 = n2831 | n3396 ;
  assign n10053 = n10052 ^ n10050 ^ n10045 ;
  assign n10054 = ( n5641 & ~n10044 ) | ( n5641 & n10053 ) | ( ~n10044 & n10053 ) ;
  assign n10042 = ( n4520 & n7174 ) | ( n4520 & ~n8629 ) | ( n7174 & ~n8629 ) ;
  assign n10056 = n10055 ^ n10054 ^ n10042 ;
  assign n10057 = n4180 ^ n446 ^ 1'b0 ;
  assign n10058 = n7990 ^ n3830 ^ n1293 ;
  assign n10059 = n2285 | n6045 ;
  assign n10060 = n10058 & n10059 ;
  assign n10061 = ~n10057 & n10060 ;
  assign n10062 = n903 & ~n6408 ;
  assign n10063 = ~n8776 & n8935 ;
  assign n10064 = n7534 & n10063 ;
  assign n10065 = n10062 | n10064 ;
  assign n10066 = x67 & n3983 ;
  assign n10067 = ~n2756 & n10066 ;
  assign n10068 = ( ~n976 & n1555 ) | ( ~n976 & n10067 ) | ( n1555 & n10067 ) ;
  assign n10069 = n10068 ^ n1423 ^ x24 ;
  assign n10070 = ( ~n1443 & n1870 ) | ( ~n1443 & n7803 ) | ( n1870 & n7803 ) ;
  assign n10071 = n4177 & ~n10070 ;
  assign n10072 = n10071 ^ n6270 ^ 1'b0 ;
  assign n10074 = n7944 ^ n3606 ^ n466 ;
  assign n10075 = n2344 ^ n1275 ^ 1'b0 ;
  assign n10076 = n10075 ^ n8896 ^ 1'b0 ;
  assign n10077 = n10074 | n10076 ;
  assign n10073 = n1173 ^ n1120 ^ n859 ;
  assign n10078 = n10077 ^ n10073 ^ 1'b0 ;
  assign n10079 = n1632 & ~n10078 ;
  assign n10080 = n10079 ^ n10005 ^ 1'b0 ;
  assign n10081 = n10072 | n10080 ;
  assign n10082 = ( n1509 & ~n3050 ) | ( n1509 & n4002 ) | ( ~n3050 & n4002 ) ;
  assign n10083 = n3213 ^ n427 ^ 1'b0 ;
  assign n10084 = ~n473 & n10083 ;
  assign n10085 = ( x200 & n4957 ) | ( x200 & n10084 ) | ( n4957 & n10084 ) ;
  assign n10086 = n8880 & ~n10085 ;
  assign n10087 = n10082 | n10086 ;
  assign n10088 = n8658 | n10087 ;
  assign n10089 = n7330 ^ n2905 ^ n2191 ;
  assign n10090 = n377 | n10089 ;
  assign n10091 = n10090 ^ n4349 ^ 1'b0 ;
  assign n10092 = ( n641 & ~n778 ) | ( n641 & n5390 ) | ( ~n778 & n5390 ) ;
  assign n10093 = ( n8694 & ~n10091 ) | ( n8694 & n10092 ) | ( ~n10091 & n10092 ) ;
  assign n10097 = n582 & ~n9294 ;
  assign n10098 = n6621 & n10097 ;
  assign n10094 = n8971 ^ n3470 ^ n1608 ;
  assign n10095 = ( n719 & n3093 ) | ( n719 & n10094 ) | ( n3093 & n10094 ) ;
  assign n10096 = ( n4219 & ~n6681 ) | ( n4219 & n10095 ) | ( ~n6681 & n10095 ) ;
  assign n10099 = n10098 ^ n10096 ^ n9302 ;
  assign n10100 = n6936 ^ n2162 ^ 1'b0 ;
  assign n10101 = n8013 ^ n5074 ^ n4097 ;
  assign n10102 = ( n4105 & n10074 ) | ( n4105 & n10101 ) | ( n10074 & n10101 ) ;
  assign n10103 = n10100 | n10102 ;
  assign n10106 = n7671 ^ n5871 ^ n4899 ;
  assign n10104 = ( ~x197 & n2338 ) | ( ~x197 & n7359 ) | ( n2338 & n7359 ) ;
  assign n10105 = ( ~n4840 & n6041 ) | ( ~n4840 & n10104 ) | ( n6041 & n10104 ) ;
  assign n10107 = n10106 ^ n10105 ^ n8599 ;
  assign n10108 = n10107 ^ n1281 ^ 1'b0 ;
  assign n10109 = n10103 & n10108 ;
  assign n10110 = ( n8983 & n10099 ) | ( n8983 & n10109 ) | ( n10099 & n10109 ) ;
  assign n10116 = n3279 ^ x167 ^ 1'b0 ;
  assign n10117 = n1436 & ~n10116 ;
  assign n10115 = ~n2597 & n9501 ;
  assign n10111 = n2553 ^ x210 ^ 1'b0 ;
  assign n10112 = ~n3085 & n10111 ;
  assign n10113 = ( n2868 & ~n4520 ) | ( n2868 & n10112 ) | ( ~n4520 & n10112 ) ;
  assign n10114 = ( ~n7240 & n7464 ) | ( ~n7240 & n10113 ) | ( n7464 & n10113 ) ;
  assign n10118 = n10117 ^ n10115 ^ n10114 ;
  assign n10124 = n8440 ^ n2735 ^ 1'b0 ;
  assign n10125 = ( ~n587 & n5353 ) | ( ~n587 & n10124 ) | ( n5353 & n10124 ) ;
  assign n10119 = n2759 ^ n2294 ^ n934 ;
  assign n10120 = n3204 | n10119 ;
  assign n10121 = n561 & ~n10120 ;
  assign n10122 = ( ~n832 & n6394 ) | ( ~n832 & n9587 ) | ( n6394 & n9587 ) ;
  assign n10123 = ( n1909 & n10121 ) | ( n1909 & ~n10122 ) | ( n10121 & ~n10122 ) ;
  assign n10126 = n10125 ^ n10123 ^ n3444 ;
  assign n10127 = n6649 | n10126 ;
  assign n10137 = n7660 ^ n5227 ^ n2739 ;
  assign n10133 = n2950 ^ n568 ^ 1'b0 ;
  assign n10134 = n8713 & ~n10133 ;
  assign n10135 = n3428 ^ n2319 ^ n1571 ;
  assign n10136 = ( n6293 & ~n10134 ) | ( n6293 & n10135 ) | ( ~n10134 & n10135 ) ;
  assign n10128 = n4523 ^ n3627 ^ 1'b0 ;
  assign n10130 = ( n2216 & ~n2303 ) | ( n2216 & n5194 ) | ( ~n2303 & n5194 ) ;
  assign n10129 = ( ~n4358 & n6158 ) | ( ~n4358 & n7348 ) | ( n6158 & n7348 ) ;
  assign n10131 = n10130 ^ n10129 ^ n5787 ;
  assign n10132 = ( n6945 & n10128 ) | ( n6945 & ~n10131 ) | ( n10128 & ~n10131 ) ;
  assign n10138 = n10137 ^ n10136 ^ n10132 ;
  assign n10139 = n1588 ^ n639 ^ 1'b0 ;
  assign n10140 = n10139 ^ n6600 ^ n1071 ;
  assign n10141 = n4270 ^ n890 ^ 1'b0 ;
  assign n10142 = ~n10140 & n10141 ;
  assign n10143 = ( n3271 & n6413 ) | ( n3271 & n10142 ) | ( n6413 & n10142 ) ;
  assign n10144 = n10143 ^ n8562 ^ n7549 ;
  assign n10145 = ~n508 & n6707 ;
  assign n10146 = n9666 ^ n1897 ^ 1'b0 ;
  assign n10147 = n10145 & ~n10146 ;
  assign n10148 = ~n8053 & n10147 ;
  assign n10149 = n10148 ^ n614 ^ 1'b0 ;
  assign n10150 = x39 & x168 ;
  assign n10151 = n10150 ^ n4836 ^ 1'b0 ;
  assign n10152 = n10151 ^ n4064 ^ 1'b0 ;
  assign n10153 = ~n2681 & n10152 ;
  assign n10154 = n10153 ^ n5833 ^ n2560 ;
  assign n10155 = n7693 ^ n3545 ^ n2770 ;
  assign n10156 = n8650 & n10155 ;
  assign n10157 = ~n10154 & n10156 ;
  assign n10158 = n7156 ^ n5991 ^ n3317 ;
  assign n10159 = n8910 ^ n2733 ^ 1'b0 ;
  assign n10160 = n10158 & ~n10159 ;
  assign n10161 = ( ~n313 & n8833 ) | ( ~n313 & n9149 ) | ( n8833 & n9149 ) ;
  assign n10162 = x18 & n5547 ;
  assign n10163 = n10161 & n10162 ;
  assign n10164 = n9017 ^ n2481 ^ n1211 ;
  assign n10165 = n6839 ^ n6395 ^ n5556 ;
  assign n10166 = n7058 ^ n6398 ^ 1'b0 ;
  assign n10167 = n6034 ^ n680 ^ n576 ;
  assign n10168 = n10167 ^ n8104 ^ n4685 ;
  assign n10170 = ( n588 & ~n3554 ) | ( n588 & n5459 ) | ( ~n3554 & n5459 ) ;
  assign n10169 = n3253 ^ n2127 ^ 1'b0 ;
  assign n10171 = n10170 ^ n10169 ^ n3167 ;
  assign n10172 = n10171 ^ n9771 ^ n2528 ;
  assign n10173 = n1013 | n5583 ;
  assign n10174 = n7195 ^ n407 ^ 1'b0 ;
  assign n10175 = ( n944 & ~n10173 ) | ( n944 & n10174 ) | ( ~n10173 & n10174 ) ;
  assign n10176 = n10175 ^ n7513 ^ n6177 ;
  assign n10177 = ( n8615 & n10172 ) | ( n8615 & ~n10176 ) | ( n10172 & ~n10176 ) ;
  assign n10178 = n10168 & ~n10177 ;
  assign n10179 = n7286 | n9798 ;
  assign n10180 = n10179 ^ n1467 ^ x114 ;
  assign n10181 = n318 | n1705 ;
  assign n10182 = n10181 ^ n1394 ^ 1'b0 ;
  assign n10183 = n8288 ^ n3522 ^ x223 ;
  assign n10184 = n10183 ^ n2931 ^ 1'b0 ;
  assign n10185 = ( ~x170 & n10182 ) | ( ~x170 & n10184 ) | ( n10182 & n10184 ) ;
  assign n10186 = n4293 ^ n3277 ^ n2902 ;
  assign n10187 = ( ~n683 & n2261 ) | ( ~n683 & n9844 ) | ( n2261 & n9844 ) ;
  assign n10188 = ( n4679 & n10186 ) | ( n4679 & n10187 ) | ( n10186 & n10187 ) ;
  assign n10194 = ( n3776 & n4977 ) | ( n3776 & ~n6109 ) | ( n4977 & ~n6109 ) ;
  assign n10189 = ( ~n1779 & n3492 ) | ( ~n1779 & n4122 ) | ( n3492 & n4122 ) ;
  assign n10190 = n9144 | n10189 ;
  assign n10191 = n10190 ^ n5082 ^ 1'b0 ;
  assign n10192 = n6584 | n10191 ;
  assign n10193 = n9779 | n10192 ;
  assign n10195 = n10194 ^ n10193 ^ n7204 ;
  assign n10196 = ( n434 & n785 ) | ( n434 & n6083 ) | ( n785 & n6083 ) ;
  assign n10197 = n5207 ^ n2622 ^ 1'b0 ;
  assign n10198 = n10197 ^ n5433 ^ n1731 ;
  assign n10199 = n10196 & ~n10198 ;
  assign n10200 = n10199 ^ n6140 ^ 1'b0 ;
  assign n10201 = ~n1009 & n3155 ;
  assign n10202 = n6303 & n10201 ;
  assign n10203 = n10202 ^ n5525 ^ n4410 ;
  assign n10204 = n1207 & n10203 ;
  assign n10205 = ~n10200 & n10204 ;
  assign n10206 = n3729 & ~n10205 ;
  assign n10207 = n6588 & n10206 ;
  assign n10208 = n8728 ^ n8545 ^ n8080 ;
  assign n10215 = n4253 ^ n2169 ^ n564 ;
  assign n10213 = n1108 | n6454 ;
  assign n10214 = n10213 ^ n1922 ^ 1'b0 ;
  assign n10216 = n10215 ^ n10214 ^ n1282 ;
  assign n10209 = ( n2665 & n4960 ) | ( n2665 & n6352 ) | ( n4960 & n6352 ) ;
  assign n10210 = n10209 ^ n3621 ^ n1782 ;
  assign n10211 = n7798 ^ n6067 ^ n4525 ;
  assign n10212 = n10210 & ~n10211 ;
  assign n10217 = n10216 ^ n10212 ^ n9660 ;
  assign n10222 = ( x144 & ~n1723 ) | ( x144 & n3037 ) | ( ~n1723 & n3037 ) ;
  assign n10218 = n3672 ^ n2935 ^ 1'b0 ;
  assign n10219 = n5339 & n10218 ;
  assign n10220 = ~n9873 & n10219 ;
  assign n10221 = n10220 ^ n2623 ^ 1'b0 ;
  assign n10223 = n10222 ^ n10221 ^ n2499 ;
  assign n10224 = n8505 ^ n2553 ^ 1'b0 ;
  assign n10225 = n8767 ^ n1937 ^ n957 ;
  assign n10226 = ( n4703 & n7073 ) | ( n4703 & n10225 ) | ( n7073 & n10225 ) ;
  assign n10227 = ~n1325 & n7801 ;
  assign n10228 = n10227 ^ n2617 ^ 1'b0 ;
  assign n10229 = n10228 ^ n7299 ^ n3898 ;
  assign n10230 = ( n10224 & n10226 ) | ( n10224 & n10229 ) | ( n10226 & n10229 ) ;
  assign n10232 = n4481 ^ n1924 ^ n1495 ;
  assign n10231 = ~n2710 & n4893 ;
  assign n10233 = n10232 ^ n10231 ^ 1'b0 ;
  assign n10234 = ( n2663 & ~n3690 ) | ( n2663 & n10233 ) | ( ~n3690 & n10233 ) ;
  assign n10235 = n1561 & n10234 ;
  assign n10236 = n1445 & n10235 ;
  assign n10237 = ( n311 & n2662 ) | ( n311 & n10236 ) | ( n2662 & n10236 ) ;
  assign n10238 = n10237 ^ n10055 ^ n2375 ;
  assign n10250 = ( ~n1105 & n1977 ) | ( ~n1105 & n3143 ) | ( n1977 & n3143 ) ;
  assign n10251 = n4469 & n10250 ;
  assign n10245 = n2602 ^ n2038 ^ x182 ;
  assign n10246 = n10245 ^ n4841 ^ 1'b0 ;
  assign n10247 = n5406 | n10246 ;
  assign n10248 = n3063 & n6426 ;
  assign n10249 = n10247 & n10248 ;
  assign n10252 = n10251 ^ n10249 ^ n3105 ;
  assign n10253 = n10252 ^ n3396 ^ 1'b0 ;
  assign n10242 = n9753 ^ n2070 ^ n530 ;
  assign n10239 = n1564 & ~n2554 ;
  assign n10240 = n938 & n10239 ;
  assign n10241 = n10240 ^ n7370 ^ n4122 ;
  assign n10243 = n10242 ^ n10241 ^ n4032 ;
  assign n10244 = n10243 ^ n6503 ^ n3608 ;
  assign n10254 = n10253 ^ n10244 ^ n9179 ;
  assign n10255 = ~n2104 & n4343 ;
  assign n10256 = n5037 & n10255 ;
  assign n10257 = n5582 ^ n5108 ^ 1'b0 ;
  assign n10267 = ( x40 & n639 ) | ( x40 & n2835 ) | ( n639 & n2835 ) ;
  assign n10268 = n10267 ^ n7806 ^ n7655 ;
  assign n10263 = n1224 | n5223 ;
  assign n10264 = n10263 ^ n8014 ^ 1'b0 ;
  assign n10265 = n10264 ^ n8928 ^ 1'b0 ;
  assign n10266 = n9082 | n10265 ;
  assign n10258 = n8787 ^ n3685 ^ n3588 ;
  assign n10259 = n1371 & n4761 ;
  assign n10260 = ( n979 & ~n10258 ) | ( n979 & n10259 ) | ( ~n10258 & n10259 ) ;
  assign n10261 = n4537 & n10260 ;
  assign n10262 = n10261 ^ n979 ^ 1'b0 ;
  assign n10269 = n10268 ^ n10266 ^ n10262 ;
  assign n10270 = ( n10256 & n10257 ) | ( n10256 & ~n10269 ) | ( n10257 & ~n10269 ) ;
  assign n10271 = ( x206 & ~n981 ) | ( x206 & n6898 ) | ( ~n981 & n6898 ) ;
  assign n10272 = ~n1073 & n5079 ;
  assign n10273 = ( n3120 & n4937 ) | ( n3120 & n5459 ) | ( n4937 & n5459 ) ;
  assign n10274 = n10273 ^ n5333 ^ n3997 ;
  assign n10275 = ( n6630 & n10272 ) | ( n6630 & ~n10274 ) | ( n10272 & ~n10274 ) ;
  assign n10277 = n3629 ^ n1729 ^ x4 ;
  assign n10276 = ( ~n858 & n6090 ) | ( ~n858 & n7286 ) | ( n6090 & n7286 ) ;
  assign n10278 = n10277 ^ n10276 ^ 1'b0 ;
  assign n10279 = n2003 ^ n817 ^ 1'b0 ;
  assign n10280 = ~n9424 & n10279 ;
  assign n10281 = n760 | n7476 ;
  assign n10282 = n10280 | n10281 ;
  assign n10283 = n4136 & n7970 ;
  assign n10284 = ~x221 & n10283 ;
  assign n10285 = ( n8890 & n10282 ) | ( n8890 & n10284 ) | ( n10282 & n10284 ) ;
  assign n10290 = ( n3188 & n6224 ) | ( n3188 & n7793 ) | ( n6224 & n7793 ) ;
  assign n10288 = n4441 & n4540 ;
  assign n10289 = ~n4926 & n10288 ;
  assign n10286 = n1923 & n2441 ;
  assign n10287 = ( n7467 & ~n9831 ) | ( n7467 & n10286 ) | ( ~n9831 & n10286 ) ;
  assign n10291 = n10290 ^ n10289 ^ n10287 ;
  assign n10292 = n6191 ^ n3847 ^ n3098 ;
  assign n10293 = n10292 ^ n3431 ^ 1'b0 ;
  assign n10294 = n9488 ^ x216 ^ 1'b0 ;
  assign n10295 = ~n7815 & n10294 ;
  assign n10298 = ~n2098 & n3480 ;
  assign n10299 = n907 & n10298 ;
  assign n10300 = n10299 ^ n7698 ^ 1'b0 ;
  assign n10296 = ( n3223 & n7450 ) | ( n3223 & ~n7817 ) | ( n7450 & ~n7817 ) ;
  assign n10297 = ( n6582 & ~n8606 ) | ( n6582 & n10296 ) | ( ~n8606 & n10296 ) ;
  assign n10301 = n10300 ^ n10297 ^ x95 ;
  assign n10302 = ( n7734 & ~n9797 ) | ( n7734 & n10301 ) | ( ~n9797 & n10301 ) ;
  assign n10303 = n5540 ^ n4747 ^ 1'b0 ;
  assign n10304 = ( n10295 & n10302 ) | ( n10295 & ~n10303 ) | ( n10302 & ~n10303 ) ;
  assign n10306 = ~n1594 & n7438 ;
  assign n10307 = ~n8381 & n10306 ;
  assign n10305 = n3495 & n9703 ;
  assign n10308 = n10307 ^ n10305 ^ 1'b0 ;
  assign n10309 = n8035 ^ n7598 ^ n6685 ;
  assign n10310 = n7213 ^ n6208 ^ x216 ;
  assign n10311 = n10310 ^ n6361 ^ 1'b0 ;
  assign n10312 = n10309 & ~n10311 ;
  assign n10313 = ( n4178 & n4301 ) | ( n4178 & ~n6805 ) | ( n4301 & ~n6805 ) ;
  assign n10314 = ~n3349 & n7992 ;
  assign n10315 = ~n8189 & n10314 ;
  assign n10316 = n2523 & n2876 ;
  assign n10317 = ( n3978 & n4216 ) | ( n3978 & ~n8082 ) | ( n4216 & ~n8082 ) ;
  assign n10318 = ( ~n3671 & n10316 ) | ( ~n3671 & n10317 ) | ( n10316 & n10317 ) ;
  assign n10319 = ( n853 & n1410 ) | ( n853 & ~n7893 ) | ( n1410 & ~n7893 ) ;
  assign n10320 = n10319 ^ n4175 ^ 1'b0 ;
  assign n10321 = ( n2633 & n9227 ) | ( n2633 & n10320 ) | ( n9227 & n10320 ) ;
  assign n10322 = n1568 | n4373 ;
  assign n10323 = ( ~n2173 & n10321 ) | ( ~n2173 & n10322 ) | ( n10321 & n10322 ) ;
  assign n10324 = n10323 ^ n7347 ^ n6654 ;
  assign n10326 = n3078 ^ n1556 ^ n310 ;
  assign n10327 = ( x81 & n5058 ) | ( x81 & n10326 ) | ( n5058 & n10326 ) ;
  assign n10328 = ( ~n2824 & n4836 ) | ( ~n2824 & n9403 ) | ( n4836 & n9403 ) ;
  assign n10329 = ( n1393 & ~n10327 ) | ( n1393 & n10328 ) | ( ~n10327 & n10328 ) ;
  assign n10330 = ( n5115 & n7491 ) | ( n5115 & n10329 ) | ( n7491 & n10329 ) ;
  assign n10325 = n2834 ^ n1485 ^ n1282 ;
  assign n10331 = n10330 ^ n10325 ^ n3632 ;
  assign n10332 = n10014 ^ n8922 ^ n6002 ;
  assign n10333 = n10332 ^ n9236 ^ n4010 ;
  assign n10336 = n1851 ^ n1504 ^ n427 ;
  assign n10337 = n10336 ^ n3347 ^ n1389 ;
  assign n10338 = n3300 ^ x94 ^ 1'b0 ;
  assign n10339 = n2323 & ~n10338 ;
  assign n10340 = ~n10337 & n10339 ;
  assign n10341 = n10340 ^ n8126 ^ 1'b0 ;
  assign n10334 = ~n362 & n3588 ;
  assign n10335 = ( n893 & n3825 ) | ( n893 & ~n10334 ) | ( n3825 & ~n10334 ) ;
  assign n10342 = n10341 ^ n10335 ^ n9512 ;
  assign n10343 = n4785 & n7330 ;
  assign n10344 = n8178 & n10343 ;
  assign n10345 = ( n1423 & ~n3785 ) | ( n1423 & n10344 ) | ( ~n3785 & n10344 ) ;
  assign n10346 = ( n2590 & n7893 ) | ( n2590 & ~n10345 ) | ( n7893 & ~n10345 ) ;
  assign n10347 = ( n1936 & n3654 ) | ( n1936 & ~n5954 ) | ( n3654 & ~n5954 ) ;
  assign n10348 = n10347 ^ n3854 ^ 1'b0 ;
  assign n10349 = n1624 & n7467 ;
  assign n10350 = n10349 ^ n5900 ^ 1'b0 ;
  assign n10351 = ( n1396 & n1908 ) | ( n1396 & ~n10350 ) | ( n1908 & ~n10350 ) ;
  assign n10352 = n8486 ^ n3824 ^ 1'b0 ;
  assign n10353 = n3188 & ~n4807 ;
  assign n10354 = n10353 ^ n6179 ^ 1'b0 ;
  assign n10355 = ~n646 & n5306 ;
  assign n10356 = n10354 & n10355 ;
  assign n10357 = n10356 ^ n7144 ^ n6142 ;
  assign n10358 = n3143 ^ n2540 ^ n267 ;
  assign n10359 = ( n1111 & n3007 ) | ( n1111 & ~n3306 ) | ( n3007 & ~n3306 ) ;
  assign n10367 = ( ~n2082 & n4066 ) | ( ~n2082 & n10219 ) | ( n4066 & n10219 ) ;
  assign n10365 = ( n992 & ~n5043 ) | ( n992 & n8920 ) | ( ~n5043 & n8920 ) ;
  assign n10366 = n10365 ^ n9955 ^ n5554 ;
  assign n10360 = n3159 ^ n1887 ^ 1'b0 ;
  assign n10361 = ~n2319 & n10360 ;
  assign n10362 = n10361 ^ n7804 ^ n4283 ;
  assign n10363 = n567 & n10362 ;
  assign n10364 = n10363 ^ n4371 ^ n1029 ;
  assign n10368 = n10367 ^ n10366 ^ n10364 ;
  assign n10369 = ( n5988 & n8182 ) | ( n5988 & n10368 ) | ( n8182 & n10368 ) ;
  assign n10370 = ( n10358 & n10359 ) | ( n10358 & n10369 ) | ( n10359 & n10369 ) ;
  assign n10371 = n7685 ^ n1029 ^ 1'b0 ;
  assign n10372 = ~n903 & n10371 ;
  assign n10373 = n1637 & n1774 ;
  assign n10374 = n10373 ^ n4200 ^ 1'b0 ;
  assign n10375 = ( ~n3715 & n7282 ) | ( ~n3715 & n10374 ) | ( n7282 & n10374 ) ;
  assign n10376 = n10375 ^ n8648 ^ n2371 ;
  assign n10377 = n10372 & n10376 ;
  assign n10378 = n10377 ^ n8318 ^ 1'b0 ;
  assign n10379 = n10378 ^ n8039 ^ n4701 ;
  assign n10380 = n7849 ^ n5461 ^ x214 ;
  assign n10381 = n10380 ^ n9821 ^ x33 ;
  assign n10382 = ~n4544 & n10381 ;
  assign n10394 = ( n1941 & n2974 ) | ( n1941 & ~n8316 ) | ( n2974 & ~n8316 ) ;
  assign n10395 = ( n2976 & n7572 ) | ( n2976 & n10394 ) | ( n7572 & n10394 ) ;
  assign n10396 = n2391 ^ n1184 ^ n710 ;
  assign n10397 = ( n6292 & ~n10395 ) | ( n6292 & n10396 ) | ( ~n10395 & n10396 ) ;
  assign n10383 = ( x252 & n2317 ) | ( x252 & ~n4212 ) | ( n2317 & ~n4212 ) ;
  assign n10384 = x55 & n10383 ;
  assign n10385 = n3105 & n10384 ;
  assign n10386 = n10385 ^ n3976 ^ n297 ;
  assign n10387 = n8031 ^ n577 ^ 1'b0 ;
  assign n10388 = n10386 & n10387 ;
  assign n10389 = n8220 ^ n8095 ^ 1'b0 ;
  assign n10390 = ( ~n4683 & n5194 ) | ( ~n4683 & n5414 ) | ( n5194 & n5414 ) ;
  assign n10391 = n10390 ^ n6223 ^ 1'b0 ;
  assign n10392 = ( ~n4392 & n4697 ) | ( ~n4392 & n10391 ) | ( n4697 & n10391 ) ;
  assign n10393 = ( n10388 & n10389 ) | ( n10388 & ~n10392 ) | ( n10389 & ~n10392 ) ;
  assign n10398 = n10397 ^ n10393 ^ n2109 ;
  assign n10399 = ( n522 & ~n1101 ) | ( n522 & n10398 ) | ( ~n1101 & n10398 ) ;
  assign n10400 = ( n5000 & n7992 ) | ( n5000 & n8557 ) | ( n7992 & n8557 ) ;
  assign n10401 = n8226 ^ x11 ^ 1'b0 ;
  assign n10402 = n10401 ^ n6414 ^ n4494 ;
  assign n10403 = n10402 ^ n1344 ^ 1'b0 ;
  assign n10404 = n5605 & ~n10403 ;
  assign n10405 = n10404 ^ n5985 ^ n2971 ;
  assign n10407 = n1967 ^ n1611 ^ 1'b0 ;
  assign n10406 = ( n740 & n6074 ) | ( n740 & n8118 ) | ( n6074 & n8118 ) ;
  assign n10408 = n10407 ^ n10406 ^ n3005 ;
  assign n10409 = n2950 & ~n10408 ;
  assign n10410 = n10409 ^ n1919 ^ 1'b0 ;
  assign n10411 = n2127 ^ n1598 ^ 1'b0 ;
  assign n10412 = n284 & n10411 ;
  assign n10413 = n10412 ^ n1922 ^ n1538 ;
  assign n10414 = n10413 ^ x193 ^ 1'b0 ;
  assign n10415 = n10414 ^ n3892 ^ n2865 ;
  assign n10419 = n9925 ^ n5014 ^ n2770 ;
  assign n10416 = n1696 ^ n1150 ^ 1'b0 ;
  assign n10417 = ( ~n767 & n2168 ) | ( ~n767 & n7197 ) | ( n2168 & n7197 ) ;
  assign n10418 = n10416 & ~n10417 ;
  assign n10420 = n10419 ^ n10418 ^ 1'b0 ;
  assign n10421 = n7290 ^ n1069 ^ n969 ;
  assign n10422 = n10421 ^ n4538 ^ n3976 ;
  assign n10423 = ( n963 & n2697 ) | ( n963 & n6060 ) | ( n2697 & n6060 ) ;
  assign n10424 = n4479 ^ n3624 ^ n3114 ;
  assign n10425 = ( n3374 & n5521 ) | ( n3374 & ~n5679 ) | ( n5521 & ~n5679 ) ;
  assign n10426 = ( x20 & n841 ) | ( x20 & ~n10425 ) | ( n841 & ~n10425 ) ;
  assign n10427 = n4061 & ~n8881 ;
  assign n10428 = ~n2187 & n10427 ;
  assign n10429 = n10428 ^ n6048 ^ n940 ;
  assign n10430 = ( ~n10424 & n10426 ) | ( ~n10424 & n10429 ) | ( n10426 & n10429 ) ;
  assign n10431 = n1768 ^ n749 ^ 1'b0 ;
  assign n10432 = n10431 ^ n8691 ^ n5094 ;
  assign n10433 = n7022 ^ n5870 ^ x165 ;
  assign n10436 = n1007 & ~n9660 ;
  assign n10437 = ~n3096 & n10436 ;
  assign n10435 = ( x145 & n585 ) | ( x145 & n2974 ) | ( n585 & n2974 ) ;
  assign n10438 = n10437 ^ n10435 ^ n7207 ;
  assign n10434 = n475 | n7950 ;
  assign n10439 = n10438 ^ n10434 ^ 1'b0 ;
  assign n10440 = ( ~n4044 & n4382 ) | ( ~n4044 & n10439 ) | ( n4382 & n10439 ) ;
  assign n10441 = ( n9770 & n10433 ) | ( n9770 & n10440 ) | ( n10433 & n10440 ) ;
  assign n10442 = ( ~n3275 & n5247 ) | ( ~n3275 & n5822 ) | ( n5247 & n5822 ) ;
  assign n10443 = n2805 | n10442 ;
  assign n10444 = n5303 ^ n1055 ^ n313 ;
  assign n10445 = n645 & ~n10444 ;
  assign n10446 = n10445 ^ n2221 ^ n1951 ;
  assign n10447 = ( n2911 & ~n3190 ) | ( n2911 & n6524 ) | ( ~n3190 & n6524 ) ;
  assign n10448 = n10447 ^ n2574 ^ 1'b0 ;
  assign n10449 = n2845 | n10448 ;
  assign n10450 = ( n8732 & n10446 ) | ( n8732 & n10449 ) | ( n10446 & n10449 ) ;
  assign n10457 = ( n1785 & n1900 ) | ( n1785 & ~n3075 ) | ( n1900 & ~n3075 ) ;
  assign n10458 = n10457 ^ n2162 ^ 1'b0 ;
  assign n10452 = ( n1811 & n3370 ) | ( n1811 & ~n7749 ) | ( n3370 & ~n7749 ) ;
  assign n10453 = ( n722 & ~n5017 ) | ( n722 & n10452 ) | ( ~n5017 & n10452 ) ;
  assign n10454 = ( x77 & n5613 ) | ( x77 & ~n10453 ) | ( n5613 & ~n10453 ) ;
  assign n10455 = n10454 ^ n3289 ^ n2646 ;
  assign n10456 = n346 & n10455 ;
  assign n10459 = n10458 ^ n10456 ^ 1'b0 ;
  assign n10451 = n9951 ^ n6342 ^ n4638 ;
  assign n10460 = n10459 ^ n10451 ^ 1'b0 ;
  assign n10461 = n4596 & ~n10460 ;
  assign n10462 = ( ~n661 & n1983 ) | ( ~n661 & n10461 ) | ( n1983 & n10461 ) ;
  assign n10464 = ~n3878 & n4603 ;
  assign n10465 = ~x54 & n10464 ;
  assign n10466 = n3258 & ~n10465 ;
  assign n10467 = ~n6803 & n10466 ;
  assign n10463 = ( n1791 & n2117 ) | ( n1791 & ~n8980 ) | ( n2117 & ~n8980 ) ;
  assign n10468 = n10467 ^ n10463 ^ n1780 ;
  assign n10469 = n8432 ^ n7459 ^ n1907 ;
  assign n10470 = ~n3980 & n8346 ;
  assign n10471 = n10469 & n10470 ;
  assign n10472 = n5309 | n8880 ;
  assign n10473 = n9227 ^ n6266 ^ 1'b0 ;
  assign n10474 = ( n2094 & n3926 ) | ( n2094 & ~n5508 ) | ( n3926 & ~n5508 ) ;
  assign n10482 = ~n3628 & n6124 ;
  assign n10483 = n10482 ^ n5800 ^ 1'b0 ;
  assign n10484 = ( n781 & n2856 ) | ( n781 & n10483 ) | ( n2856 & n10483 ) ;
  assign n10485 = ( n4583 & n10094 ) | ( n4583 & n10484 ) | ( n10094 & n10484 ) ;
  assign n10475 = ( n1972 & n2684 ) | ( n1972 & ~n7755 ) | ( n2684 & ~n7755 ) ;
  assign n10476 = ( n883 & n4841 ) | ( n883 & ~n10475 ) | ( n4841 & ~n10475 ) ;
  assign n10477 = ( ~n755 & n3923 ) | ( ~n755 & n10476 ) | ( n3923 & n10476 ) ;
  assign n10478 = n9017 ^ n739 ^ 1'b0 ;
  assign n10479 = ( n2433 & n10477 ) | ( n2433 & ~n10478 ) | ( n10477 & ~n10478 ) ;
  assign n10480 = ( ~n2627 & n3301 ) | ( ~n2627 & n7638 ) | ( n3301 & n7638 ) ;
  assign n10481 = n10479 | n10480 ;
  assign n10486 = n10485 ^ n10481 ^ n4410 ;
  assign n10487 = ( n1114 & n5162 ) | ( n1114 & ~n6718 ) | ( n5162 & ~n6718 ) ;
  assign n10488 = n4420 & ~n10487 ;
  assign n10489 = n10488 ^ n7913 ^ 1'b0 ;
  assign n10490 = ( n3117 & n3133 ) | ( n3117 & n9896 ) | ( n3133 & n9896 ) ;
  assign n10491 = n10490 ^ n8731 ^ n3321 ;
  assign n10492 = n10491 ^ n10104 ^ n8828 ;
  assign n10499 = n1708 & ~n5526 ;
  assign n10497 = ( n1707 & ~n4559 ) | ( n1707 & n5579 ) | ( ~n4559 & n5579 ) ;
  assign n10493 = n3788 & n9478 ;
  assign n10494 = n793 & n10493 ;
  assign n10495 = n926 | n6465 ;
  assign n10496 = n10494 & ~n10495 ;
  assign n10498 = n10497 ^ n10496 ^ n4654 ;
  assign n10500 = n10499 ^ n10498 ^ n6708 ;
  assign n10501 = ( n5044 & n9723 ) | ( n5044 & ~n10500 ) | ( n9723 & ~n10500 ) ;
  assign n10506 = n1946 | n6223 ;
  assign n10503 = n3797 ^ n1430 ^ 1'b0 ;
  assign n10504 = n1879 & ~n10503 ;
  assign n10502 = ( x200 & ~n7402 ) | ( x200 & n9269 ) | ( ~n7402 & n9269 ) ;
  assign n10505 = n10504 ^ n10502 ^ n1536 ;
  assign n10507 = n10506 ^ n10505 ^ n9655 ;
  assign n10508 = x63 & x77 ;
  assign n10509 = n4197 ^ n3180 ^ 1'b0 ;
  assign n10510 = ( ~n2777 & n8990 ) | ( ~n2777 & n10509 ) | ( n8990 & n10509 ) ;
  assign n10511 = n4841 ^ n3324 ^ 1'b0 ;
  assign n10512 = ( n10508 & n10510 ) | ( n10508 & n10511 ) | ( n10510 & n10511 ) ;
  assign n10518 = n6993 ^ n1500 ^ 1'b0 ;
  assign n10516 = n1131 & n1374 ;
  assign n10517 = ( n1081 & n7457 ) | ( n1081 & n10516 ) | ( n7457 & n10516 ) ;
  assign n10513 = n6970 ^ n4628 ^ n3920 ;
  assign n10514 = ( n517 & n6977 ) | ( n517 & ~n10513 ) | ( n6977 & ~n10513 ) ;
  assign n10515 = n10514 ^ n7921 ^ 1'b0 ;
  assign n10519 = n10518 ^ n10517 ^ n10515 ;
  assign n10520 = ( x221 & n8374 ) | ( x221 & n10519 ) | ( n8374 & n10519 ) ;
  assign n10521 = n7791 ^ n4277 ^ n3354 ;
  assign n10522 = n7708 ^ n5032 ^ n4524 ;
  assign n10523 = ( n1533 & ~n3626 ) | ( n1533 & n9438 ) | ( ~n3626 & n9438 ) ;
  assign n10524 = n10523 ^ n7866 ^ n1150 ;
  assign n10525 = ( n10521 & ~n10522 ) | ( n10521 & n10524 ) | ( ~n10522 & n10524 ) ;
  assign n10526 = n2738 & n10525 ;
  assign n10527 = ~n4801 & n10526 ;
  assign n10528 = n7462 ^ n7115 ^ n1226 ;
  assign n10530 = ~n926 & n4982 ;
  assign n10531 = n10530 ^ n5204 ^ 1'b0 ;
  assign n10532 = ~n5909 & n10531 ;
  assign n10529 = ~n1296 & n9385 ;
  assign n10533 = n10532 ^ n10529 ^ 1'b0 ;
  assign n10534 = ( n2944 & n5836 ) | ( n2944 & n10208 ) | ( n5836 & n10208 ) ;
  assign n10535 = ( n4860 & ~n4987 ) | ( n4860 & n8689 ) | ( ~n4987 & n8689 ) ;
  assign n10536 = ( ~x90 & n2510 ) | ( ~x90 & n10535 ) | ( n2510 & n10535 ) ;
  assign n10537 = n10536 ^ n3870 ^ n276 ;
  assign n10538 = n4770 ^ n4616 ^ n2108 ;
  assign n10539 = ( n1630 & n2469 ) | ( n1630 & ~n2905 ) | ( n2469 & ~n2905 ) ;
  assign n10540 = n10539 ^ n5238 ^ n2617 ;
  assign n10541 = ( n7774 & n10538 ) | ( n7774 & ~n10540 ) | ( n10538 & ~n10540 ) ;
  assign n10542 = n587 | n1958 ;
  assign n10543 = n8872 | n10542 ;
  assign n10544 = ( x49 & n2815 ) | ( x49 & ~n10543 ) | ( n2815 & ~n10543 ) ;
  assign n10545 = ( n10186 & ~n10541 ) | ( n10186 & n10544 ) | ( ~n10541 & n10544 ) ;
  assign n10546 = ( n1837 & n10537 ) | ( n1837 & n10545 ) | ( n10537 & n10545 ) ;
  assign n10550 = n5542 ^ n4808 ^ n277 ;
  assign n10551 = ( x122 & ~n7348 ) | ( x122 & n10550 ) | ( ~n7348 & n10550 ) ;
  assign n10547 = ~n1690 & n7911 ;
  assign n10548 = n10547 ^ n3395 ^ n2331 ;
  assign n10549 = n10548 ^ n3002 ^ 1'b0 ;
  assign n10552 = n10551 ^ n10549 ^ 1'b0 ;
  assign n10553 = n1749 & n10552 ;
  assign n10554 = n2456 ^ n2244 ^ n1205 ;
  assign n10556 = ( x154 & ~n658 ) | ( x154 & n8319 ) | ( ~n658 & n8319 ) ;
  assign n10557 = n5559 ^ n2819 ^ n1901 ;
  assign n10558 = ( n4143 & n10556 ) | ( n4143 & ~n10557 ) | ( n10556 & ~n10557 ) ;
  assign n10559 = n10558 ^ n1108 ^ 1'b0 ;
  assign n10555 = ~n3177 & n9968 ;
  assign n10560 = n10559 ^ n10555 ^ 1'b0 ;
  assign n10561 = ~n10554 & n10560 ;
  assign n10565 = n537 & ~n5296 ;
  assign n10566 = n10565 ^ x211 ^ 1'b0 ;
  assign n10567 = ( n2443 & n6093 ) | ( n2443 & ~n10566 ) | ( n6093 & ~n10566 ) ;
  assign n10562 = n640 ^ n301 ^ x72 ;
  assign n10563 = n10562 ^ n8881 ^ n2811 ;
  assign n10564 = ( n6497 & n9813 ) | ( n6497 & ~n10563 ) | ( n9813 & ~n10563 ) ;
  assign n10568 = n10567 ^ n10564 ^ n4515 ;
  assign n10569 = ( n480 & n2042 ) | ( n480 & ~n4538 ) | ( n2042 & ~n4538 ) ;
  assign n10570 = ( ~n278 & n2597 ) | ( ~n278 & n5841 ) | ( n2597 & n5841 ) ;
  assign n10571 = n3345 & ~n10570 ;
  assign n10572 = ~n5937 & n10571 ;
  assign n10573 = n10572 ^ n9914 ^ n1903 ;
  assign n10574 = n10573 ^ n10417 ^ 1'b0 ;
  assign n10575 = ~n10569 & n10574 ;
  assign n10576 = n10575 ^ n6733 ^ 1'b0 ;
  assign n10577 = n10576 ^ n10410 ^ n10267 ;
  assign n10578 = ~n4356 & n7389 ;
  assign n10579 = ( n1027 & n5251 ) | ( n1027 & n10578 ) | ( n5251 & n10578 ) ;
  assign n10580 = n10579 ^ n3159 ^ 1'b0 ;
  assign n10581 = n7089 & ~n10580 ;
  assign n10582 = n3387 ^ n1996 ^ 1'b0 ;
  assign n10583 = n10582 ^ n4835 ^ n1221 ;
  assign n10584 = ( n3828 & ~n6574 ) | ( n3828 & n10583 ) | ( ~n6574 & n10583 ) ;
  assign n10585 = n5045 ^ n540 ^ x57 ;
  assign n10586 = n10585 ^ n9930 ^ n2410 ;
  assign n10587 = ( ~n3977 & n10584 ) | ( ~n3977 & n10586 ) | ( n10584 & n10586 ) ;
  assign n10588 = n10587 ^ n4427 ^ n1098 ;
  assign n10589 = n6154 ^ n3110 ^ n2143 ;
  assign n10590 = n359 & n2320 ;
  assign n10591 = n4962 ^ n562 ^ 1'b0 ;
  assign n10592 = n2442 & ~n10591 ;
  assign n10595 = ( ~x153 & n279 ) | ( ~x153 & n3857 ) | ( n279 & n3857 ) ;
  assign n10593 = ~n3544 & n4558 ;
  assign n10594 = n10593 ^ n2632 ^ 1'b0 ;
  assign n10596 = n10595 ^ n10594 ^ n7513 ;
  assign n10597 = ( n10590 & ~n10592 ) | ( n10590 & n10596 ) | ( ~n10592 & n10596 ) ;
  assign n10598 = ~n10589 & n10597 ;
  assign n10599 = n10598 ^ n9803 ^ n5790 ;
  assign n10600 = n4515 | n9009 ;
  assign n10601 = n10600 ^ n6933 ^ 1'b0 ;
  assign n10602 = ~n1139 & n10601 ;
  assign n10603 = ( n2516 & n4678 ) | ( n2516 & n6468 ) | ( n4678 & n6468 ) ;
  assign n10604 = ( n2032 & n10113 ) | ( n2032 & ~n10603 ) | ( n10113 & ~n10603 ) ;
  assign n10608 = n6506 ^ n2755 ^ x97 ;
  assign n10607 = ( n418 & n8945 ) | ( n418 & n9769 ) | ( n8945 & n9769 ) ;
  assign n10605 = ( ~x192 & n2623 ) | ( ~x192 & n4422 ) | ( n2623 & n4422 ) ;
  assign n10606 = n10605 ^ n8274 ^ n4512 ;
  assign n10609 = n10608 ^ n10607 ^ n10606 ;
  assign n10610 = ( n10233 & n10604 ) | ( n10233 & ~n10609 ) | ( n10604 & ~n10609 ) ;
  assign n10611 = ( n8673 & n9604 ) | ( n8673 & n9890 ) | ( n9604 & n9890 ) ;
  assign n10612 = ( n2591 & n7627 ) | ( n2591 & n9798 ) | ( n7627 & n9798 ) ;
  assign n10613 = ( ~n1492 & n9696 ) | ( ~n1492 & n10612 ) | ( n9696 & n10612 ) ;
  assign n10614 = n8233 ^ n2687 ^ n316 ;
  assign n10615 = ( ~x32 & n3160 ) | ( ~x32 & n10614 ) | ( n3160 & n10614 ) ;
  assign n10616 = ( x171 & n4044 ) | ( x171 & n4687 ) | ( n4044 & n4687 ) ;
  assign n10617 = n3174 ^ n847 ^ 1'b0 ;
  assign n10618 = ( n3610 & n5979 ) | ( n3610 & n10617 ) | ( n5979 & n10617 ) ;
  assign n10619 = ( n4104 & ~n9809 ) | ( n4104 & n10618 ) | ( ~n9809 & n10618 ) ;
  assign n10620 = ( n5731 & n10457 ) | ( n5731 & n10619 ) | ( n10457 & n10619 ) ;
  assign n10621 = n4399 & n10620 ;
  assign n10622 = ~n8094 & n10621 ;
  assign n10623 = n10622 ^ n9980 ^ n9211 ;
  assign n10624 = n1060 & ~n3109 ;
  assign n10625 = ( n3776 & n6111 ) | ( n3776 & n10624 ) | ( n6111 & n10624 ) ;
  assign n10626 = n2615 ^ n1454 ^ 1'b0 ;
  assign n10628 = ~n3679 & n6994 ;
  assign n10629 = n10628 ^ n7457 ^ n3519 ;
  assign n10627 = n4868 & ~n8278 ;
  assign n10630 = n10629 ^ n10627 ^ 1'b0 ;
  assign n10632 = x227 & n5317 ;
  assign n10631 = ( x42 & ~n1166 ) | ( x42 & n3906 ) | ( ~n1166 & n3906 ) ;
  assign n10633 = n10632 ^ n10631 ^ n742 ;
  assign n10634 = ( n7588 & n9610 ) | ( n7588 & n10633 ) | ( n9610 & n10633 ) ;
  assign n10635 = ~n10630 & n10634 ;
  assign n10636 = ( ~n1675 & n2379 ) | ( ~n1675 & n6423 ) | ( n2379 & n6423 ) ;
  assign n10637 = n10636 ^ n7912 ^ 1'b0 ;
  assign n10638 = n2640 & n10637 ;
  assign n10639 = ( x43 & n1238 ) | ( x43 & n5641 ) | ( n1238 & n5641 ) ;
  assign n10640 = n10639 ^ n2818 ^ 1'b0 ;
  assign n10641 = n10638 & ~n10640 ;
  assign n10642 = n8708 ^ n4178 ^ n976 ;
  assign n10643 = ( n5790 & n8156 ) | ( n5790 & n10642 ) | ( n8156 & n10642 ) ;
  assign n10644 = ( n2810 & n5490 ) | ( n2810 & ~n10643 ) | ( n5490 & ~n10643 ) ;
  assign n10657 = n3764 ^ n2222 ^ 1'b0 ;
  assign n10655 = n1910 & n5442 ;
  assign n10656 = n3560 & n10655 ;
  assign n10658 = n10657 ^ n10656 ^ n3750 ;
  assign n10645 = n3177 ^ n2615 ^ n2554 ;
  assign n10646 = ( x209 & ~n2034 ) | ( x209 & n2680 ) | ( ~n2034 & n2680 ) ;
  assign n10647 = ( n8080 & ~n10645 ) | ( n8080 & n10646 ) | ( ~n10645 & n10646 ) ;
  assign n10648 = n7515 ^ n5013 ^ 1'b0 ;
  assign n10649 = n2590 | n10648 ;
  assign n10650 = ( n3241 & n4698 ) | ( n3241 & n8517 ) | ( n4698 & n8517 ) ;
  assign n10651 = n2325 & n3044 ;
  assign n10652 = ( n10649 & ~n10650 ) | ( n10649 & n10651 ) | ( ~n10650 & n10651 ) ;
  assign n10653 = n10647 & ~n10652 ;
  assign n10654 = n10653 ^ n4860 ^ 1'b0 ;
  assign n10659 = n10658 ^ n10654 ^ n7171 ;
  assign n10660 = n5937 ^ n432 ^ n269 ;
  assign n10661 = n7911 ^ n4369 ^ n337 ;
  assign n10662 = n10660 | n10661 ;
  assign n10663 = ~n4457 & n8374 ;
  assign n10664 = ( n1613 & ~n1871 ) | ( n1613 & n4559 ) | ( ~n1871 & n4559 ) ;
  assign n10665 = n6904 | n10664 ;
  assign n10666 = n10663 & ~n10665 ;
  assign n10667 = n7145 ^ n6024 ^ n2336 ;
  assign n10668 = ~n1308 & n2721 ;
  assign n10669 = n10668 ^ n2655 ^ n1123 ;
  assign n10670 = n10669 ^ n5101 ^ n4541 ;
  assign n10671 = ( n4213 & ~n4795 ) | ( n4213 & n10439 ) | ( ~n4795 & n10439 ) ;
  assign n10672 = ( n3158 & n7865 ) | ( n3158 & ~n10671 ) | ( n7865 & ~n10671 ) ;
  assign n10673 = ( ~x249 & n5331 ) | ( ~x249 & n9239 ) | ( n5331 & n9239 ) ;
  assign n10674 = n7342 & ~n10673 ;
  assign n10675 = n10672 & n10674 ;
  assign n10676 = ( n2644 & n3253 ) | ( n2644 & ~n6381 ) | ( n3253 & ~n6381 ) ;
  assign n10677 = ( ~n3042 & n3496 ) | ( ~n3042 & n8139 ) | ( n3496 & n8139 ) ;
  assign n10678 = n7774 & ~n9720 ;
  assign n10679 = n4612 & ~n10678 ;
  assign n10680 = ( n2077 & n5316 ) | ( n2077 & ~n10679 ) | ( n5316 & ~n10679 ) ;
  assign n10681 = ( n974 & n2790 ) | ( n974 & n5704 ) | ( n2790 & n5704 ) ;
  assign n10682 = n3990 ^ n3604 ^ n2518 ;
  assign n10683 = n10682 ^ n7976 ^ n2275 ;
  assign n10684 = ~n3938 & n10683 ;
  assign n10685 = n10684 ^ n7719 ^ 1'b0 ;
  assign n10686 = n4504 ^ n2217 ^ 1'b0 ;
  assign n10687 = n4134 | n10686 ;
  assign n10688 = n10687 ^ n3301 ^ n2227 ;
  assign n10689 = n1308 & n5780 ;
  assign n10690 = n10689 ^ n5419 ^ 1'b0 ;
  assign n10691 = n6815 & ~n10690 ;
  assign n10692 = ~n10688 & n10691 ;
  assign n10693 = ( n10163 & n10685 ) | ( n10163 & ~n10692 ) | ( n10685 & ~n10692 ) ;
  assign n10694 = ( n567 & n1352 ) | ( n567 & n2782 ) | ( n1352 & n2782 ) ;
  assign n10695 = n622 & ~n10694 ;
  assign n10696 = n10347 & n10695 ;
  assign n10697 = n10696 ^ n3822 ^ 1'b0 ;
  assign n10698 = ( n2566 & n6446 ) | ( n2566 & ~n10697 ) | ( n6446 & ~n10697 ) ;
  assign n10699 = n8319 & n10698 ;
  assign n10702 = n2992 ^ n1377 ^ 1'b0 ;
  assign n10703 = n10702 ^ n6714 ^ x246 ;
  assign n10701 = n1197 | n8348 ;
  assign n10704 = n10703 ^ n10701 ^ 1'b0 ;
  assign n10700 = n3936 & ~n6165 ;
  assign n10705 = n10704 ^ n10700 ^ 1'b0 ;
  assign n10706 = ( n5740 & n7811 ) | ( n5740 & n10705 ) | ( n7811 & n10705 ) ;
  assign n10707 = n10706 ^ n4794 ^ n549 ;
  assign n10711 = ( n1274 & n4873 ) | ( n1274 & ~n5309 ) | ( n4873 & ~n5309 ) ;
  assign n10708 = n529 | n6544 ;
  assign n10709 = ( n4085 & ~n4351 ) | ( n4085 & n10596 ) | ( ~n4351 & n10596 ) ;
  assign n10710 = ( ~x19 & n10708 ) | ( ~x19 & n10709 ) | ( n10708 & n10709 ) ;
  assign n10712 = n10711 ^ n10710 ^ n6039 ;
  assign n10713 = n8975 ^ n6874 ^ n1091 ;
  assign n10714 = n10713 ^ n1925 ^ 1'b0 ;
  assign n10715 = n10712 & n10714 ;
  assign n10717 = n2697 ^ n1315 ^ n898 ;
  assign n10718 = ( n6284 & n8635 ) | ( n6284 & n10717 ) | ( n8635 & n10717 ) ;
  assign n10716 = n5551 ^ n2861 ^ n1212 ;
  assign n10719 = n10718 ^ n10716 ^ 1'b0 ;
  assign n10720 = n10719 ^ n9070 ^ n8686 ;
  assign n10727 = ~n2780 & n5331 ;
  assign n10728 = ~n5460 & n10727 ;
  assign n10724 = n2710 | n8573 ;
  assign n10725 = n799 | n10724 ;
  assign n10723 = ( n3764 & n3778 ) | ( n3764 & ~n7363 ) | ( n3778 & ~n7363 ) ;
  assign n10726 = n10725 ^ n10723 ^ n4644 ;
  assign n10721 = n8591 & ~n10431 ;
  assign n10722 = n10721 ^ n9813 ^ n2716 ;
  assign n10729 = n10728 ^ n10726 ^ n10722 ;
  assign n10730 = x244 & ~n5162 ;
  assign n10731 = n10730 ^ n3144 ^ 1'b0 ;
  assign n10732 = n1801 & ~n10094 ;
  assign n10733 = n10732 ^ n5027 ^ 1'b0 ;
  assign n10734 = n10731 | n10733 ;
  assign n10735 = n5624 & ~n10734 ;
  assign n10739 = n7660 ^ n4695 ^ 1'b0 ;
  assign n10736 = n6064 ^ n3254 ^ n2878 ;
  assign n10737 = n3014 ^ n596 ^ 1'b0 ;
  assign n10738 = n10736 & n10737 ;
  assign n10740 = n10739 ^ n10738 ^ 1'b0 ;
  assign n10741 = n1730 & ~n10740 ;
  assign n10742 = ( n5220 & n7904 ) | ( n5220 & ~n8374 ) | ( n7904 & ~n8374 ) ;
  assign n10743 = ( n6858 & n6958 ) | ( n6858 & n10742 ) | ( n6958 & n10742 ) ;
  assign n10744 = n7808 ^ n6301 ^ n6192 ;
  assign n10745 = ( x198 & n3080 ) | ( x198 & n10744 ) | ( n3080 & n10744 ) ;
  assign n10746 = ( ~n1445 & n10743 ) | ( ~n1445 & n10745 ) | ( n10743 & n10745 ) ;
  assign n10747 = ~n423 & n9170 ;
  assign n10748 = n3472 & ~n10747 ;
  assign n10749 = n10748 ^ n796 ^ 1'b0 ;
  assign n10750 = n655 | n10749 ;
  assign n10751 = n1614 & ~n10750 ;
  assign n10752 = ( n1796 & ~n3137 ) | ( n1796 & n6425 ) | ( ~n3137 & n6425 ) ;
  assign n10753 = ( n2859 & n7929 ) | ( n2859 & ~n10752 ) | ( n7929 & ~n10752 ) ;
  assign n10754 = ~n543 & n9309 ;
  assign n10755 = n10754 ^ n3880 ^ 1'b0 ;
  assign n10756 = n648 & n10755 ;
  assign n10757 = ~n9437 & n10756 ;
  assign n10762 = ( n2025 & ~n2730 ) | ( n2025 & n2735 ) | ( ~n2730 & n2735 ) ;
  assign n10763 = n10762 ^ n8945 ^ n1240 ;
  assign n10761 = ( n1635 & n4820 ) | ( n1635 & n5076 ) | ( n4820 & n5076 ) ;
  assign n10764 = n10763 ^ n10761 ^ x18 ;
  assign n10758 = ( n469 & ~n3725 ) | ( n469 & n5133 ) | ( ~n3725 & n5133 ) ;
  assign n10759 = ( ~n5218 & n7499 ) | ( ~n5218 & n10758 ) | ( n7499 & n10758 ) ;
  assign n10760 = ~n2396 & n10759 ;
  assign n10765 = n10764 ^ n10760 ^ n390 ;
  assign n10768 = ( n746 & n1454 ) | ( n746 & ~n1897 ) | ( n1454 & ~n1897 ) ;
  assign n10766 = ~n1873 & n9493 ;
  assign n10767 = n3020 | n10766 ;
  assign n10769 = n10768 ^ n10767 ^ 1'b0 ;
  assign n10770 = n10765 & n10769 ;
  assign n10771 = n8925 & n9301 ;
  assign n10772 = n10771 ^ n9064 ^ 1'b0 ;
  assign n10774 = n7658 ^ n5181 ^ 1'b0 ;
  assign n10775 = n973 | n10774 ;
  assign n10773 = ( ~n1440 & n2200 ) | ( ~n1440 & n3469 ) | ( n2200 & n3469 ) ;
  assign n10776 = n10775 ^ n10773 ^ n8053 ;
  assign n10777 = ( x190 & n4143 ) | ( x190 & ~n8350 ) | ( n4143 & ~n8350 ) ;
  assign n10778 = ( n2067 & n7433 ) | ( n2067 & n8647 ) | ( n7433 & n8647 ) ;
  assign n10779 = ( n8980 & n10777 ) | ( n8980 & n10778 ) | ( n10777 & n10778 ) ;
  assign n10780 = ( n3274 & ~n5233 ) | ( n3274 & n5799 ) | ( ~n5233 & n5799 ) ;
  assign n10781 = ( x127 & n10779 ) | ( x127 & ~n10780 ) | ( n10779 & ~n10780 ) ;
  assign n10782 = n4916 ^ n2385 ^ 1'b0 ;
  assign n10783 = ~n3288 & n10782 ;
  assign n10784 = n1756 & n3625 ;
  assign n10785 = n10784 ^ n7990 ^ 1'b0 ;
  assign n10786 = n10785 ^ n2727 ^ n1676 ;
  assign n10787 = n10786 ^ n8699 ^ n5039 ;
  assign n10788 = ( n8468 & ~n10783 ) | ( n8468 & n10787 ) | ( ~n10783 & n10787 ) ;
  assign n10789 = n5907 ^ n1637 ^ 1'b0 ;
  assign n10790 = n10789 ^ n8004 ^ n1371 ;
  assign n10791 = n5065 ^ n1163 ^ 1'b0 ;
  assign n10792 = n7990 & n10791 ;
  assign n10793 = n1150 & ~n5924 ;
  assign n10794 = n10793 ^ n3071 ^ 1'b0 ;
  assign n10795 = ( ~n6181 & n7410 ) | ( ~n6181 & n10794 ) | ( n7410 & n10794 ) ;
  assign n10796 = ( n522 & ~n10792 ) | ( n522 & n10795 ) | ( ~n10792 & n10795 ) ;
  assign n10798 = n714 & ~n6883 ;
  assign n10799 = n10798 ^ n339 ^ 1'b0 ;
  assign n10800 = n6723 | n10799 ;
  assign n10797 = n4543 ^ n1744 ^ 1'b0 ;
  assign n10801 = n10800 ^ n10797 ^ n4104 ;
  assign n10802 = ( n511 & n1067 ) | ( n511 & ~n4186 ) | ( n1067 & ~n4186 ) ;
  assign n10803 = n10802 ^ n3819 ^ 1'b0 ;
  assign n10804 = n4743 & n10803 ;
  assign n10805 = n10804 ^ n5418 ^ 1'b0 ;
  assign n10806 = ~x206 & n5010 ;
  assign n10807 = ~n6015 & n10806 ;
  assign n10808 = n4961 & n5483 ;
  assign n10809 = n10808 ^ n1256 ^ 1'b0 ;
  assign n10810 = n10809 ^ n7073 ^ n4792 ;
  assign n10811 = n9379 ^ n6666 ^ x191 ;
  assign n10812 = n3174 | n6349 ;
  assign n10815 = ( n1293 & n4338 ) | ( n1293 & ~n8575 ) | ( n4338 & ~n8575 ) ;
  assign n10814 = ( ~n927 & n2389 ) | ( ~n927 & n8364 ) | ( n2389 & n8364 ) ;
  assign n10813 = ( x81 & n4744 ) | ( x81 & ~n8377 ) | ( n4744 & ~n8377 ) ;
  assign n10816 = n10815 ^ n10814 ^ n10813 ;
  assign n10817 = ( ~n10811 & n10812 ) | ( ~n10811 & n10816 ) | ( n10812 & n10816 ) ;
  assign n10818 = ~n4235 & n10817 ;
  assign n10819 = n4715 & n10818 ;
  assign n10820 = ( n9841 & ~n10810 ) | ( n9841 & n10819 ) | ( ~n10810 & n10819 ) ;
  assign n10821 = n10820 ^ n6073 ^ n2877 ;
  assign n10822 = n4257 ^ n3578 ^ n3298 ;
  assign n10823 = ( n3419 & ~n8485 ) | ( n3419 & n10822 ) | ( ~n8485 & n10822 ) ;
  assign n10824 = ~n702 & n2305 ;
  assign n10825 = n10823 | n10824 ;
  assign n10826 = n5453 | n10825 ;
  assign n10827 = n809 & ~n3937 ;
  assign n10828 = ~n1470 & n10827 ;
  assign n10829 = n5712 & ~n10828 ;
  assign n10830 = n10829 ^ n6532 ^ 1'b0 ;
  assign n10831 = ( ~n4385 & n9026 ) | ( ~n4385 & n10830 ) | ( n9026 & n10830 ) ;
  assign n10832 = n10831 ^ n8111 ^ n994 ;
  assign n10833 = x68 & ~n2020 ;
  assign n10838 = n1724 ^ n742 ^ n720 ;
  assign n10834 = x32 & ~n2978 ;
  assign n10835 = n10834 ^ n3718 ^ 1'b0 ;
  assign n10836 = n2062 | n10835 ;
  assign n10837 = n10836 ^ n343 ^ 1'b0 ;
  assign n10839 = n10838 ^ n10837 ^ 1'b0 ;
  assign n10840 = n3739 & n10839 ;
  assign n10841 = n990 & n5822 ;
  assign n10842 = ~n7838 & n10841 ;
  assign n10843 = ( ~n6779 & n10840 ) | ( ~n6779 & n10842 ) | ( n10840 & n10842 ) ;
  assign n10844 = ( n2679 & n10833 ) | ( n2679 & n10843 ) | ( n10833 & n10843 ) ;
  assign n10845 = n3110 | n10844 ;
  assign n10846 = ( n7893 & n9685 ) | ( n7893 & n10845 ) | ( n9685 & n10845 ) ;
  assign n10847 = n9961 ^ n1497 ^ n947 ;
  assign n10849 = n9712 ^ n8350 ^ n4690 ;
  assign n10848 = ( n2364 & ~n3421 ) | ( n2364 & n6257 ) | ( ~n3421 & n6257 ) ;
  assign n10850 = n10849 ^ n10848 ^ n9923 ;
  assign n10851 = n3564 & n10850 ;
  assign n10852 = n10851 ^ n6879 ^ 1'b0 ;
  assign n10853 = n9466 ^ n1886 ^ n751 ;
  assign n10854 = n6601 ^ n2752 ^ 1'b0 ;
  assign n10855 = n2956 & ~n6662 ;
  assign n10858 = ( n2644 & ~n4410 ) | ( n2644 & n7792 ) | ( ~n4410 & n7792 ) ;
  assign n10856 = ( n1189 & n3212 ) | ( n1189 & ~n4122 ) | ( n3212 & ~n4122 ) ;
  assign n10857 = n10856 ^ n9475 ^ n6387 ;
  assign n10859 = n10858 ^ n10857 ^ n3455 ;
  assign n10860 = n10859 ^ n4872 ^ n1690 ;
  assign n10861 = ( n10854 & ~n10855 ) | ( n10854 & n10860 ) | ( ~n10855 & n10860 ) ;
  assign n10870 = n6313 ^ n5605 ^ n1451 ;
  assign n10871 = n10870 ^ n1826 ^ n1258 ;
  assign n10862 = ~n6206 & n8163 ;
  assign n10863 = ~n7293 & n10862 ;
  assign n10866 = ( n1682 & n3784 ) | ( n1682 & n3838 ) | ( n3784 & n3838 ) ;
  assign n10867 = ( n2821 & n7492 ) | ( n2821 & n10866 ) | ( n7492 & n10866 ) ;
  assign n10865 = ( ~n895 & n1272 ) | ( ~n895 & n3479 ) | ( n1272 & n3479 ) ;
  assign n10864 = ( n412 & n5734 ) | ( n412 & n9129 ) | ( n5734 & n9129 ) ;
  assign n10868 = n10867 ^ n10865 ^ n10864 ;
  assign n10869 = n10863 | n10868 ;
  assign n10872 = n10871 ^ n10869 ^ 1'b0 ;
  assign n10876 = n4961 ^ n1577 ^ n463 ;
  assign n10875 = n2962 & n7414 ;
  assign n10877 = n10876 ^ n10875 ^ n1725 ;
  assign n10873 = ( ~x160 & n875 ) | ( ~x160 & n3614 ) | ( n875 & n3614 ) ;
  assign n10874 = n10873 ^ n10249 ^ n3942 ;
  assign n10878 = n10877 ^ n10874 ^ n6828 ;
  assign n10879 = n10878 ^ n10196 ^ n9655 ;
  assign n10880 = n2857 ^ n2275 ^ 1'b0 ;
  assign n10881 = n774 | n10880 ;
  assign n10883 = n5328 ^ n4500 ^ n2033 ;
  assign n10882 = ( n1369 & n5904 ) | ( n1369 & ~n9660 ) | ( n5904 & ~n9660 ) ;
  assign n10884 = n10883 ^ n10882 ^ n2517 ;
  assign n10885 = ( n6820 & n10237 ) | ( n6820 & n10884 ) | ( n10237 & n10884 ) ;
  assign n10886 = ( n3932 & n10881 ) | ( n3932 & n10885 ) | ( n10881 & n10885 ) ;
  assign n10887 = ( ~n3084 & n3558 ) | ( ~n3084 & n3992 ) | ( n3558 & n3992 ) ;
  assign n10888 = ( n2383 & n2865 ) | ( n2383 & ~n5952 ) | ( n2865 & ~n5952 ) ;
  assign n10889 = ( n4007 & n8325 ) | ( n4007 & n9938 ) | ( n8325 & n9938 ) ;
  assign n10890 = ( ~n10170 & n10888 ) | ( ~n10170 & n10889 ) | ( n10888 & n10889 ) ;
  assign n10891 = ( n4572 & ~n10887 ) | ( n4572 & n10890 ) | ( ~n10887 & n10890 ) ;
  assign n10892 = ( n1562 & n5804 ) | ( n1562 & ~n9631 ) | ( n5804 & ~n9631 ) ;
  assign n10893 = n6114 ^ n5845 ^ n1669 ;
  assign n10894 = n4685 & ~n7752 ;
  assign n10895 = n10894 ^ n5582 ^ n3421 ;
  assign n10896 = ( n400 & ~n10893 ) | ( n400 & n10895 ) | ( ~n10893 & n10895 ) ;
  assign n10899 = n1156 ^ n688 ^ 1'b0 ;
  assign n10897 = ( n1103 & ~n7760 ) | ( n1103 & n10536 ) | ( ~n7760 & n10536 ) ;
  assign n10898 = n2651 & n10897 ;
  assign n10900 = n10899 ^ n10898 ^ 1'b0 ;
  assign n10901 = ( n5985 & n10896 ) | ( n5985 & n10900 ) | ( n10896 & n10900 ) ;
  assign n10902 = ( ~n7259 & n10892 ) | ( ~n7259 & n10901 ) | ( n10892 & n10901 ) ;
  assign n10903 = ~n3695 & n10047 ;
  assign n10904 = ( n1447 & n2586 ) | ( n1447 & ~n10903 ) | ( n2586 & ~n10903 ) ;
  assign n10913 = n1290 ^ n1120 ^ 1'b0 ;
  assign n10914 = ~n828 & n10913 ;
  assign n10907 = n5453 ^ n459 ^ 1'b0 ;
  assign n10908 = n4985 & ~n10907 ;
  assign n10909 = n10908 ^ n9905 ^ n8356 ;
  assign n10910 = n7635 ^ n7627 ^ 1'b0 ;
  assign n10911 = n10909 & n10910 ;
  assign n10912 = ( x216 & n8211 ) | ( x216 & ~n10911 ) | ( n8211 & ~n10911 ) ;
  assign n10905 = n8442 ^ n6565 ^ n6165 ;
  assign n10906 = ( n1830 & ~n8677 ) | ( n1830 & n10905 ) | ( ~n8677 & n10905 ) ;
  assign n10915 = n10914 ^ n10912 ^ n10906 ;
  assign n10956 = n8836 ^ n540 ^ x21 ;
  assign n10954 = n7114 ^ n1509 ^ 1'b0 ;
  assign n10941 = ( n1600 & n6247 ) | ( n1600 & n8244 ) | ( n6247 & n8244 ) ;
  assign n10950 = n3662 ^ n2155 ^ n547 ;
  assign n10947 = ( n2442 & n3067 ) | ( n2442 & ~n3235 ) | ( n3067 & ~n3235 ) ;
  assign n10945 = n3231 | n7370 ;
  assign n10946 = n10945 ^ n2197 ^ 1'b0 ;
  assign n10942 = n6884 & ~n10694 ;
  assign n10943 = ~n4654 & n10942 ;
  assign n10944 = ( n4569 & ~n5465 ) | ( n4569 & n10943 ) | ( ~n5465 & n10943 ) ;
  assign n10948 = n10947 ^ n10946 ^ n10944 ;
  assign n10949 = n10948 ^ n8888 ^ n1377 ;
  assign n10951 = n10950 ^ n10949 ^ 1'b0 ;
  assign n10952 = ~n10941 & n10951 ;
  assign n10953 = n7485 & n10952 ;
  assign n10955 = n10954 ^ n10953 ^ 1'b0 ;
  assign n10957 = n10956 ^ n10955 ^ n1182 ;
  assign n10958 = n5119 & ~n10957 ;
  assign n10959 = n10958 ^ n5017 ^ 1'b0 ;
  assign n10928 = n3855 ^ n3355 ^ x109 ;
  assign n10929 = ( n4431 & n4702 ) | ( n4431 & ~n10928 ) | ( n4702 & ~n10928 ) ;
  assign n10930 = n10929 ^ n4153 ^ 1'b0 ;
  assign n10931 = ~n6347 & n10930 ;
  assign n10925 = n2721 ^ n2255 ^ x35 ;
  assign n10926 = n10925 ^ n8214 ^ n1299 ;
  assign n10927 = n10926 ^ n1652 ^ n388 ;
  assign n10932 = n10931 ^ n10927 ^ n10854 ;
  assign n10924 = ( ~n1185 & n1289 ) | ( ~n1185 & n1441 ) | ( n1289 & n1441 ) ;
  assign n10933 = n10932 ^ n10924 ^ n1427 ;
  assign n10934 = n1497 & n10539 ;
  assign n10935 = ( n9357 & ~n10933 ) | ( n9357 & n10934 ) | ( ~n10933 & n10934 ) ;
  assign n10916 = x166 & ~n732 ;
  assign n10917 = ~x99 & n10916 ;
  assign n10918 = n6909 ^ n3441 ^ n1635 ;
  assign n10919 = ( ~n374 & n4597 ) | ( ~n374 & n10918 ) | ( n4597 & n10918 ) ;
  assign n10920 = ( n6426 & ~n10917 ) | ( n6426 & n10919 ) | ( ~n10917 & n10919 ) ;
  assign n10921 = ~n7116 & n10920 ;
  assign n10922 = n10921 ^ n7006 ^ 1'b0 ;
  assign n10923 = n10922 ^ n6977 ^ 1'b0 ;
  assign n10936 = n10935 ^ n10923 ^ n1580 ;
  assign n10937 = n1326 & n7938 ;
  assign n10938 = n10937 ^ n1053 ^ 1'b0 ;
  assign n10939 = n7423 | n10938 ;
  assign n10940 = n10936 & ~n10939 ;
  assign n10960 = n10959 ^ n10940 ^ n1988 ;
  assign n10961 = n1215 & ~n7772 ;
  assign n10962 = ( n6103 & n7799 ) | ( n6103 & ~n10961 ) | ( n7799 & ~n10961 ) ;
  assign n10963 = n8262 & ~n10962 ;
  assign n10964 = n3525 & ~n5034 ;
  assign n10965 = ( ~n3112 & n6319 ) | ( ~n3112 & n10964 ) | ( n6319 & n10964 ) ;
  assign n10970 = ( n1753 & n5264 ) | ( n1753 & ~n5724 ) | ( n5264 & ~n5724 ) ;
  assign n10966 = n5259 & n7192 ;
  assign n10967 = n4080 & ~n10966 ;
  assign n10968 = ~n4775 & n10967 ;
  assign n10969 = n10968 ^ n10484 ^ n5207 ;
  assign n10971 = n10970 ^ n10969 ^ 1'b0 ;
  assign n10972 = n9799 ^ n8711 ^ 1'b0 ;
  assign n10973 = n9660 ^ n6187 ^ 1'b0 ;
  assign n10974 = n8919 ^ n4385 ^ 1'b0 ;
  assign n10975 = n10973 | n10974 ;
  assign n10976 = n10975 ^ n5834 ^ n4460 ;
  assign n10999 = ( x89 & n1067 ) | ( x89 & ~n4978 ) | ( n1067 & ~n4978 ) ;
  assign n10991 = n3139 | n6785 ;
  assign n10992 = n5290 | n10991 ;
  assign n10993 = n9104 ^ n8258 ^ n714 ;
  assign n10994 = n10992 & ~n10993 ;
  assign n10995 = n10994 ^ n8288 ^ 1'b0 ;
  assign n10987 = n5742 ^ n5667 ^ n2180 ;
  assign n10988 = n10987 ^ n9311 ^ n2592 ;
  assign n10984 = n9600 ^ n6069 ^ n2567 ;
  assign n10985 = n953 & ~n3086 ;
  assign n10986 = n10984 | n10985 ;
  assign n10989 = n10988 ^ n10986 ^ 1'b0 ;
  assign n10990 = n6166 & ~n10989 ;
  assign n10996 = n10995 ^ n10990 ^ n1190 ;
  assign n10997 = n10996 ^ n2762 ^ x6 ;
  assign n10977 = n5401 | n10457 ;
  assign n10980 = n8575 ^ n3096 ^ 1'b0 ;
  assign n10981 = n610 & ~n10980 ;
  assign n10978 = ( n546 & ~n733 ) | ( n546 & n3906 ) | ( ~n733 & n3906 ) ;
  assign n10979 = ( n1135 & ~n9207 ) | ( n1135 & n10978 ) | ( ~n9207 & n10978 ) ;
  assign n10982 = n10981 ^ n10979 ^ 1'b0 ;
  assign n10983 = n10977 & ~n10982 ;
  assign n10998 = n10997 ^ n10983 ^ 1'b0 ;
  assign n11000 = n10999 ^ n10998 ^ 1'b0 ;
  assign n11001 = ~n10976 & n11000 ;
  assign n11004 = ( n1022 & n1763 ) | ( n1022 & ~n7204 ) | ( n1763 & ~n7204 ) ;
  assign n11005 = ( n478 & n2856 ) | ( n478 & ~n11004 ) | ( n2856 & ~n11004 ) ;
  assign n11003 = n654 & n3192 ;
  assign n11006 = n11005 ^ n11003 ^ 1'b0 ;
  assign n11007 = n11006 ^ n8412 ^ n5504 ;
  assign n11008 = ( n2718 & n6034 ) | ( n2718 & ~n11007 ) | ( n6034 & ~n11007 ) ;
  assign n11002 = n3673 ^ n2041 ^ n1560 ;
  assign n11009 = n11008 ^ n11002 ^ n8643 ;
  assign n11017 = ( ~n2296 & n4138 ) | ( ~n2296 & n5718 ) | ( n4138 & n5718 ) ;
  assign n11018 = n11017 ^ n3357 ^ n1370 ;
  assign n11011 = ~n6543 & n10380 ;
  assign n11012 = n6883 & n11011 ;
  assign n11013 = n3314 & ~n11012 ;
  assign n11014 = n11013 ^ n9691 ^ 1'b0 ;
  assign n11010 = n8011 ^ n2492 ^ n403 ;
  assign n11015 = n11014 ^ n11010 ^ 1'b0 ;
  assign n11016 = n6295 & n11015 ;
  assign n11019 = n11018 ^ n11016 ^ n4341 ;
  assign n11020 = n6294 ^ n3209 ^ 1'b0 ;
  assign n11021 = n4502 ^ n3468 ^ n1912 ;
  assign n11022 = ( n6720 & n11020 ) | ( n6720 & ~n11021 ) | ( n11020 & ~n11021 ) ;
  assign n11025 = n3311 | n5469 ;
  assign n11023 = n10421 ^ n5341 ^ n1910 ;
  assign n11024 = n9140 | n11023 ;
  assign n11026 = n11025 ^ n11024 ^ 1'b0 ;
  assign n11027 = ( n2204 & n11022 ) | ( n2204 & ~n11026 ) | ( n11022 & ~n11026 ) ;
  assign n11028 = n3794 & ~n11027 ;
  assign n11029 = n9644 & n11028 ;
  assign n11030 = ( n4640 & ~n4667 ) | ( n4640 & n11029 ) | ( ~n4667 & n11029 ) ;
  assign n11031 = n11019 | n11030 ;
  assign n11032 = ( ~n2033 & n3798 ) | ( ~n2033 & n10049 ) | ( n3798 & n10049 ) ;
  assign n11033 = n5909 ^ n448 ^ 1'b0 ;
  assign n11034 = n11033 ^ n10642 ^ 1'b0 ;
  assign n11035 = ( n6805 & n10678 ) | ( n6805 & n11034 ) | ( n10678 & n11034 ) ;
  assign n11036 = ( n1128 & ~n1310 ) | ( n1128 & n6227 ) | ( ~n1310 & n6227 ) ;
  assign n11037 = ( n5724 & n11035 ) | ( n5724 & n11036 ) | ( n11035 & n11036 ) ;
  assign n11038 = n1943 & n11037 ;
  assign n11039 = n2724 ^ n442 ^ 1'b0 ;
  assign n11040 = ( n716 & n926 ) | ( n716 & ~n1381 ) | ( n926 & ~n1381 ) ;
  assign n11041 = ( n2721 & n11039 ) | ( n2721 & n11040 ) | ( n11039 & n11040 ) ;
  assign n11042 = ( n6941 & ~n8992 ) | ( n6941 & n9289 ) | ( ~n8992 & n9289 ) ;
  assign n11043 = ~n5242 & n6833 ;
  assign n11044 = ( ~n1862 & n5940 ) | ( ~n1862 & n6737 ) | ( n5940 & n6737 ) ;
  assign n11045 = n6822 ^ n1136 ^ 1'b0 ;
  assign n11046 = ~n11044 & n11045 ;
  assign n11047 = ~n2396 & n11046 ;
  assign n11048 = n3657 & n11047 ;
  assign n11049 = n11048 ^ n2740 ^ 1'b0 ;
  assign n11050 = ~n2303 & n11049 ;
  assign n11051 = n6026 ^ n4269 ^ n4224 ;
  assign n11052 = n5786 & n11051 ;
  assign n11053 = n11052 ^ n7771 ^ 1'b0 ;
  assign n11054 = ~n5212 & n11053 ;
  assign n11055 = n2916 & n11054 ;
  assign n11056 = ( n3501 & n6497 ) | ( n3501 & ~n7518 ) | ( n6497 & ~n7518 ) ;
  assign n11057 = x181 & ~n11056 ;
  assign n11058 = n5205 ^ n5036 ^ 1'b0 ;
  assign n11059 = ( n2089 & ~n8953 ) | ( n2089 & n11058 ) | ( ~n8953 & n11058 ) ;
  assign n11061 = n6559 ^ n6010 ^ n894 ;
  assign n11060 = ~n3329 & n3924 ;
  assign n11062 = n11061 ^ n11060 ^ 1'b0 ;
  assign n11063 = n3086 & ~n11062 ;
  assign n11064 = ( ~n7112 & n11059 ) | ( ~n7112 & n11063 ) | ( n11059 & n11063 ) ;
  assign n11065 = n11057 & n11064 ;
  assign n11066 = n11055 & n11065 ;
  assign n11067 = n8078 ^ n6878 ^ n1187 ;
  assign n11068 = n5600 ^ n1824 ^ n787 ;
  assign n11069 = ( n3341 & n9231 ) | ( n3341 & ~n11068 ) | ( n9231 & ~n11068 ) ;
  assign n11070 = n2418 ^ n1559 ^ 1'b0 ;
  assign n11071 = n11070 ^ n5368 ^ n1831 ;
  assign n11072 = n3847 ^ n2243 ^ 1'b0 ;
  assign n11073 = n2197 | n11072 ;
  assign n11074 = n11073 ^ n5861 ^ n437 ;
  assign n11075 = n11074 ^ n2024 ^ n1056 ;
  assign n11076 = ( n3001 & n6672 ) | ( n3001 & n11075 ) | ( n6672 & n11075 ) ;
  assign n11077 = n11071 | n11076 ;
  assign n11078 = n11077 ^ n5859 ^ 1'b0 ;
  assign n11079 = ( n5094 & ~n11069 ) | ( n5094 & n11078 ) | ( ~n11069 & n11078 ) ;
  assign n11080 = n11067 & n11079 ;
  assign n11084 = n3583 ^ n412 ^ n353 ;
  assign n11082 = n8665 ^ x153 ^ 1'b0 ;
  assign n11083 = n3363 & n11082 ;
  assign n11081 = n8102 ^ n5462 ^ n1963 ;
  assign n11085 = n11084 ^ n11083 ^ n11081 ;
  assign n11086 = n11085 ^ n7308 ^ x143 ;
  assign n11087 = n5304 ^ n3096 ^ 1'b0 ;
  assign n11088 = n377 | n11087 ;
  assign n11089 = n11088 ^ n4109 ^ 1'b0 ;
  assign n11090 = n8092 ^ n5588 ^ n5534 ;
  assign n11091 = ( n976 & ~n4317 ) | ( n976 & n6335 ) | ( ~n4317 & n6335 ) ;
  assign n11092 = n1634 & n11091 ;
  assign n11093 = ~n11090 & n11092 ;
  assign n11101 = n2601 ^ n2408 ^ n1560 ;
  assign n11097 = n3129 ^ n345 ^ 1'b0 ;
  assign n11098 = n9771 & ~n11097 ;
  assign n11094 = n2854 ^ n1813 ^ n1422 ;
  assign n11095 = ( n2323 & n6201 ) | ( n2323 & n7293 ) | ( n6201 & n7293 ) ;
  assign n11096 = ~n11094 & n11095 ;
  assign n11099 = n11098 ^ n11096 ^ 1'b0 ;
  assign n11100 = n11099 ^ n7587 ^ n2102 ;
  assign n11102 = n11101 ^ n11100 ^ 1'b0 ;
  assign n11103 = ~n1282 & n11102 ;
  assign n11104 = n11103 ^ n7710 ^ n2554 ;
  assign n11105 = n6654 ^ n3604 ^ n1223 ;
  assign n11106 = x161 & n4070 ;
  assign n11107 = n11106 ^ n3779 ^ 1'b0 ;
  assign n11108 = n3838 & n11107 ;
  assign n11109 = n11108 ^ n4610 ^ n4126 ;
  assign n11110 = ( ~n3796 & n11105 ) | ( ~n3796 & n11109 ) | ( n11105 & n11109 ) ;
  assign n11111 = ( n2616 & ~n5346 ) | ( n2616 & n5657 ) | ( ~n5346 & n5657 ) ;
  assign n11112 = n11111 ^ n7926 ^ n7371 ;
  assign n11114 = n7482 ^ n5104 ^ 1'b0 ;
  assign n11113 = n6737 ^ n3947 ^ n2312 ;
  assign n11115 = n11114 ^ n11113 ^ n2586 ;
  assign n11116 = ( ~n9706 & n11112 ) | ( ~n9706 & n11115 ) | ( n11112 & n11115 ) ;
  assign n11117 = n2291 ^ n1574 ^ 1'b0 ;
  assign n11118 = n350 & n11117 ;
  assign n11119 = ( n3742 & ~n4186 ) | ( n3742 & n9803 ) | ( ~n4186 & n9803 ) ;
  assign n11120 = ( n2005 & n3097 ) | ( n2005 & ~n9887 ) | ( n3097 & ~n9887 ) ;
  assign n11122 = n607 & n2905 ;
  assign n11123 = n2674 & n11122 ;
  assign n11124 = ( x11 & n5463 ) | ( x11 & ~n11123 ) | ( n5463 & ~n11123 ) ;
  assign n11125 = n4572 & n11124 ;
  assign n11126 = n11125 ^ n1467 ^ 1'b0 ;
  assign n11121 = n1840 | n3784 ;
  assign n11127 = n11126 ^ n11121 ^ 1'b0 ;
  assign n11128 = ( n3095 & n6124 ) | ( n3095 & ~n11005 ) | ( n6124 & ~n11005 ) ;
  assign n11129 = n11127 & ~n11128 ;
  assign n11130 = ( n8368 & ~n9608 ) | ( n8368 & n11129 ) | ( ~n9608 & n11129 ) ;
  assign n11131 = ( n3544 & ~n4872 ) | ( n3544 & n5792 ) | ( ~n4872 & n5792 ) ;
  assign n11132 = n11131 ^ x152 ^ 1'b0 ;
  assign n11133 = n7209 ^ n1476 ^ 1'b0 ;
  assign n11134 = ~n451 & n11133 ;
  assign n11135 = n11134 ^ n9014 ^ 1'b0 ;
  assign n11136 = n9426 ^ n6179 ^ n276 ;
  assign n11137 = ( n6531 & n11135 ) | ( n6531 & n11136 ) | ( n11135 & n11136 ) ;
  assign n11138 = ~n11132 & n11137 ;
  assign n11144 = ( ~n1132 & n2505 ) | ( ~n1132 & n9732 ) | ( n2505 & n9732 ) ;
  assign n11141 = ( n2382 & n5252 ) | ( n2382 & n7352 ) | ( n5252 & n7352 ) ;
  assign n11142 = x23 | n11141 ;
  assign n11139 = n2905 & n8690 ;
  assign n11140 = n9454 & n11139 ;
  assign n11143 = n11142 ^ n11140 ^ n5783 ;
  assign n11145 = n11144 ^ n11143 ^ n2591 ;
  assign n11146 = n8615 ^ n3128 ^ n735 ;
  assign n11147 = n1266 & ~n7499 ;
  assign n11148 = n5598 & ~n11147 ;
  assign n11149 = ~n11146 & n11148 ;
  assign n11154 = n4917 ^ n1911 ^ 1'b0 ;
  assign n11152 = ( ~n1777 & n3399 ) | ( ~n1777 & n3906 ) | ( n3399 & n3906 ) ;
  assign n11150 = ~n3451 & n6237 ;
  assign n11151 = n11150 ^ n3765 ^ n1499 ;
  assign n11153 = n11152 ^ n11151 ^ n3509 ;
  assign n11155 = n11154 ^ n11153 ^ n9332 ;
  assign n11156 = n8151 ^ n5160 ^ n551 ;
  assign n11157 = ( n862 & n2291 ) | ( n862 & n4412 ) | ( n2291 & n4412 ) ;
  assign n11158 = n4677 ^ n2132 ^ 1'b0 ;
  assign n11159 = n2154 & n11158 ;
  assign n11160 = ( ~n1567 & n5209 ) | ( ~n1567 & n11159 ) | ( n5209 & n11159 ) ;
  assign n11161 = n11160 ^ n7366 ^ 1'b0 ;
  assign n11162 = n11157 & ~n11161 ;
  assign n11169 = ( n2440 & ~n3060 ) | ( n2440 & n7991 ) | ( ~n3060 & n7991 ) ;
  assign n11170 = n11169 ^ n5964 ^ n2829 ;
  assign n11163 = n3985 ^ n1465 ^ x64 ;
  assign n11164 = n4110 ^ n2929 ^ n1779 ;
  assign n11165 = ( ~n1741 & n4494 ) | ( ~n1741 & n11164 ) | ( n4494 & n11164 ) ;
  assign n11166 = ( n7781 & n11163 ) | ( n7781 & ~n11165 ) | ( n11163 & ~n11165 ) ;
  assign n11167 = n11166 ^ n3367 ^ n1136 ;
  assign n11168 = n11167 ^ n2385 ^ 1'b0 ;
  assign n11171 = n11170 ^ n11168 ^ n1567 ;
  assign n11172 = n9720 ^ n3077 ^ n2202 ;
  assign n11173 = ( n1169 & ~n9670 ) | ( n1169 & n11172 ) | ( ~n9670 & n11172 ) ;
  assign n11174 = n11173 ^ n10169 ^ 1'b0 ;
  assign n11175 = ~n1419 & n6249 ;
  assign n11176 = n11175 ^ n3494 ^ 1'b0 ;
  assign n11177 = ( n10296 & n11174 ) | ( n10296 & ~n11176 ) | ( n11174 & ~n11176 ) ;
  assign n11178 = n8242 ^ n1240 ^ 1'b0 ;
  assign n11179 = ~n5154 & n11178 ;
  assign n11180 = ( ~n1226 & n2950 ) | ( ~n1226 & n3710 ) | ( n2950 & n3710 ) ;
  assign n11181 = ( n1069 & n9495 ) | ( n1069 & n11180 ) | ( n9495 & n11180 ) ;
  assign n11182 = ( ~n4779 & n6057 ) | ( ~n4779 & n11181 ) | ( n6057 & n11181 ) ;
  assign n11183 = n6197 ^ n5183 ^ 1'b0 ;
  assign n11184 = n11183 ^ n7059 ^ n1547 ;
  assign n11185 = n9067 & ~n10716 ;
  assign n11186 = ~n8615 & n11185 ;
  assign n11187 = n8364 ^ n3944 ^ n809 ;
  assign n11188 = ( n2855 & n3250 ) | ( n2855 & ~n6858 ) | ( n3250 & ~n6858 ) ;
  assign n11189 = ( n1361 & n7963 ) | ( n1361 & ~n11188 ) | ( n7963 & ~n11188 ) ;
  assign n11190 = n11187 | n11189 ;
  assign n11191 = ( n1682 & n4280 ) | ( n1682 & n6000 ) | ( n4280 & n6000 ) ;
  assign n11192 = ( ~n6072 & n8834 ) | ( ~n6072 & n11191 ) | ( n8834 & n11191 ) ;
  assign n11193 = n3680 ^ n602 ^ 1'b0 ;
  assign n11194 = ( n1459 & ~n4502 ) | ( n1459 & n11193 ) | ( ~n4502 & n11193 ) ;
  assign n11195 = n11194 ^ n8787 ^ n8742 ;
  assign n11203 = ( n1319 & ~n4868 ) | ( n1319 & n9106 ) | ( ~n4868 & n9106 ) ;
  assign n11199 = n6423 ^ n5885 ^ n5609 ;
  assign n11200 = ~n10809 & n11199 ;
  assign n11201 = n11200 ^ n8837 ^ 1'b0 ;
  assign n11202 = ( ~n794 & n2313 ) | ( ~n794 & n11201 ) | ( n2313 & n11201 ) ;
  assign n11197 = n4064 ^ n1408 ^ 1'b0 ;
  assign n11196 = n2697 | n6588 ;
  assign n11198 = n11197 ^ n11196 ^ 1'b0 ;
  assign n11204 = n11203 ^ n11202 ^ n11198 ;
  assign n11205 = n11204 ^ n7028 ^ 1'b0 ;
  assign n11206 = ~n11195 & n11205 ;
  assign n11207 = ( n2396 & n4344 ) | ( n2396 & n4872 ) | ( n4344 & n4872 ) ;
  assign n11208 = ( n1921 & ~n6850 ) | ( n1921 & n11207 ) | ( ~n6850 & n11207 ) ;
  assign n11213 = x166 & ~n4359 ;
  assign n11214 = n1547 & n11213 ;
  assign n11209 = n1010 | n1670 ;
  assign n11210 = n11209 ^ n820 ^ 1'b0 ;
  assign n11211 = n11210 ^ n2735 ^ n264 ;
  assign n11212 = n11211 ^ n8844 ^ n5751 ;
  assign n11215 = n11214 ^ n11212 ^ n7632 ;
  assign n11216 = n2858 & n11215 ;
  assign n11217 = n9535 & n11216 ;
  assign n11218 = n1859 | n11217 ;
  assign n11219 = n6629 ^ n631 ^ 1'b0 ;
  assign n11220 = ( n2023 & ~n5204 ) | ( n2023 & n11219 ) | ( ~n5204 & n11219 ) ;
  assign n11221 = ( ~n630 & n3826 ) | ( ~n630 & n11220 ) | ( n3826 & n11220 ) ;
  assign n11222 = n11221 ^ n4411 ^ 1'b0 ;
  assign n11223 = n1973 ^ x137 ^ 1'b0 ;
  assign n11227 = ~n633 & n4549 ;
  assign n11228 = n4859 & ~n11227 ;
  assign n11229 = n11228 ^ n8225 ^ 1'b0 ;
  assign n11224 = ~x80 & n10413 ;
  assign n11225 = ( n8502 & n9070 ) | ( n8502 & ~n11224 ) | ( n9070 & ~n11224 ) ;
  assign n11226 = ( x219 & n1198 ) | ( x219 & n11225 ) | ( n1198 & n11225 ) ;
  assign n11230 = n11229 ^ n11226 ^ n9555 ;
  assign n11231 = n3445 ^ n3375 ^ n448 ;
  assign n11232 = n11231 ^ n7519 ^ n2225 ;
  assign n11233 = n6540 ^ n2348 ^ 1'b0 ;
  assign n11234 = ( n4939 & ~n11232 ) | ( n4939 & n11233 ) | ( ~n11232 & n11233 ) ;
  assign n11235 = n2351 & ~n4337 ;
  assign n11236 = n11235 ^ n3340 ^ n2510 ;
  assign n11237 = n7487 ^ n6699 ^ n5164 ;
  assign n11238 = ( n2566 & n11236 ) | ( n2566 & ~n11237 ) | ( n11236 & ~n11237 ) ;
  assign n11239 = n9348 ^ n6331 ^ 1'b0 ;
  assign n11240 = n2596 & n11239 ;
  assign n11241 = n7526 ^ n4773 ^ 1'b0 ;
  assign n11242 = n8501 & ~n11241 ;
  assign n11243 = n8822 ^ n4306 ^ n3901 ;
  assign n11244 = n10988 | n11243 ;
  assign n11245 = n11242 | n11244 ;
  assign n11246 = ~n4191 & n5877 ;
  assign n11247 = n3366 ^ n3069 ^ n1282 ;
  assign n11248 = ( n2968 & n6336 ) | ( n2968 & ~n11247 ) | ( n6336 & ~n11247 ) ;
  assign n11249 = n6955 ^ n6283 ^ n4129 ;
  assign n11250 = n312 & n7818 ;
  assign n11251 = n11249 & n11250 ;
  assign n11252 = n11251 ^ n5286 ^ 1'b0 ;
  assign n11253 = n11014 ^ n6082 ^ 1'b0 ;
  assign n11254 = n11252 | n11253 ;
  assign n11255 = n8440 ^ n3245 ^ 1'b0 ;
  assign n11256 = ( x124 & ~n8713 ) | ( x124 & n10895 ) | ( ~n8713 & n10895 ) ;
  assign n11257 = n6231 ^ n1535 ^ n531 ;
  assign n11258 = n640 | n1945 ;
  assign n11259 = n9805 | n11258 ;
  assign n11260 = ( n1491 & ~n4460 ) | ( n1491 & n8909 ) | ( ~n4460 & n8909 ) ;
  assign n11261 = n4938 | n10130 ;
  assign n11262 = ( n1392 & n2042 ) | ( n1392 & n2743 ) | ( n2042 & n2743 ) ;
  assign n11263 = n11262 ^ n7302 ^ x90 ;
  assign n11264 = ( n11260 & n11261 ) | ( n11260 & ~n11263 ) | ( n11261 & ~n11263 ) ;
  assign n11265 = ( n1787 & ~n5466 ) | ( n1787 & n7637 ) | ( ~n5466 & n7637 ) ;
  assign n11266 = n11265 ^ n6788 ^ 1'b0 ;
  assign n11267 = n11264 & n11266 ;
  assign n11268 = ( ~n5521 & n6684 ) | ( ~n5521 & n7973 ) | ( n6684 & n7973 ) ;
  assign n11269 = n11268 ^ n1909 ^ n740 ;
  assign n11270 = ( n4360 & n10824 ) | ( n4360 & ~n11269 ) | ( n10824 & ~n11269 ) ;
  assign n11271 = n3439 & ~n11270 ;
  assign n11272 = x232 & ~n2254 ;
  assign n11273 = n11272 ^ n8115 ^ 1'b0 ;
  assign n11276 = ~n4608 & n7671 ;
  assign n11277 = n11276 ^ n8652 ^ 1'b0 ;
  assign n11274 = ( n2726 & ~n3124 ) | ( n2726 & n5777 ) | ( ~n3124 & n5777 ) ;
  assign n11275 = ( n8228 & n9299 ) | ( n8228 & ~n11274 ) | ( n9299 & ~n11274 ) ;
  assign n11278 = n11277 ^ n11275 ^ n8260 ;
  assign n11279 = n11273 & n11278 ;
  assign n11287 = n9514 ^ n5886 ^ n3920 ;
  assign n11280 = n4304 ^ n4042 ^ 1'b0 ;
  assign n11281 = n11280 ^ n7167 ^ n1074 ;
  assign n11282 = n10167 | n11281 ;
  assign n11283 = n11282 ^ n7728 ^ 1'b0 ;
  assign n11284 = n11283 ^ n6114 ^ n821 ;
  assign n11285 = n11284 ^ n4697 ^ n2843 ;
  assign n11286 = n3792 & n11285 ;
  assign n11288 = n11287 ^ n11286 ^ 1'b0 ;
  assign n11289 = n6184 ^ n4989 ^ n1012 ;
  assign n11290 = ~n2041 & n3558 ;
  assign n11291 = ~n286 & n11290 ;
  assign n11292 = n11291 ^ n9217 ^ n1286 ;
  assign n11293 = n11292 ^ n5539 ^ 1'b0 ;
  assign n11294 = n9961 | n11293 ;
  assign n11295 = n11289 | n11294 ;
  assign n11296 = n1279 | n9319 ;
  assign n11297 = n11295 | n11296 ;
  assign n11298 = ( n4515 & n11288 ) | ( n4515 & n11297 ) | ( n11288 & n11297 ) ;
  assign n11303 = n4368 ^ n3361 ^ n1422 ;
  assign n11304 = ( ~n3598 & n6750 ) | ( ~n3598 & n11303 ) | ( n6750 & n11303 ) ;
  assign n11301 = n5555 ^ n2572 ^ n2491 ;
  assign n11299 = ( n4124 & n5013 ) | ( n4124 & n8263 ) | ( n5013 & n8263 ) ;
  assign n11300 = n11299 ^ n346 ^ n305 ;
  assign n11302 = n11301 ^ n11300 ^ n2015 ;
  assign n11305 = n11304 ^ n11302 ^ n846 ;
  assign n11306 = ( n1190 & n1395 ) | ( n1190 & ~n2465 ) | ( n1395 & ~n2465 ) ;
  assign n11307 = n5506 & n11306 ;
  assign n11308 = n11307 ^ n10058 ^ n7746 ;
  assign n11309 = ( n2566 & ~n3298 ) | ( n2566 & n6408 ) | ( ~n3298 & n6408 ) ;
  assign n11310 = n11309 ^ n1749 ^ x20 ;
  assign n11311 = ( ~x77 & x97 ) | ( ~x77 & n9741 ) | ( x97 & n9741 ) ;
  assign n11312 = ( n7891 & n11310 ) | ( n7891 & n11311 ) | ( n11310 & n11311 ) ;
  assign n11313 = n2730 & n4808 ;
  assign n11314 = n11313 ^ n4007 ^ 1'b0 ;
  assign n11315 = n11314 ^ n4516 ^ 1'b0 ;
  assign n11316 = n5319 | n11315 ;
  assign n11317 = n11316 ^ n3906 ^ 1'b0 ;
  assign n11318 = ~n7977 & n11317 ;
  assign n11319 = ( n687 & n11312 ) | ( n687 & n11318 ) | ( n11312 & n11318 ) ;
  assign n11320 = ( ~n766 & n11308 ) | ( ~n766 & n11319 ) | ( n11308 & n11319 ) ;
  assign n11321 = n859 | n1580 ;
  assign n11322 = ( n3746 & ~n7771 ) | ( n3746 & n11321 ) | ( ~n7771 & n11321 ) ;
  assign n11323 = n3250 & n5439 ;
  assign n11324 = n11323 ^ n6202 ^ 1'b0 ;
  assign n11325 = n7629 ^ n1694 ^ 1'b0 ;
  assign n11326 = ( n8157 & ~n11324 ) | ( n8157 & n11325 ) | ( ~n11324 & n11325 ) ;
  assign n11327 = n5880 & n8770 ;
  assign n11328 = ~n330 & n11327 ;
  assign n11329 = ( ~n5057 & n8813 ) | ( ~n5057 & n11328 ) | ( n8813 & n11328 ) ;
  assign n11330 = n10271 ^ n3969 ^ n3582 ;
  assign n11333 = n6969 ^ n6636 ^ n3629 ;
  assign n11331 = ( ~n341 & n1126 ) | ( ~n341 & n9930 ) | ( n1126 & n9930 ) ;
  assign n11332 = n11331 ^ n10516 ^ x193 ;
  assign n11334 = n11333 ^ n11332 ^ n3621 ;
  assign n11335 = ( ~n8466 & n10537 ) | ( ~n8466 & n11334 ) | ( n10537 & n11334 ) ;
  assign n11336 = n10776 ^ n8054 ^ n7847 ;
  assign n11359 = ( n1682 & ~n2782 ) | ( n1682 & n4808 ) | ( ~n2782 & n4808 ) ;
  assign n11340 = n10098 ^ n9359 ^ n4571 ;
  assign n11337 = ( x153 & n3741 ) | ( x153 & ~n7598 ) | ( n3741 & ~n7598 ) ;
  assign n11338 = n9294 ^ x155 ^ 1'b0 ;
  assign n11339 = n11337 & ~n11338 ;
  assign n11341 = n11340 ^ n11339 ^ 1'b0 ;
  assign n11342 = n1005 & n6374 ;
  assign n11343 = n9476 & n11342 ;
  assign n11344 = n364 & n989 ;
  assign n11345 = n6022 & n11344 ;
  assign n11346 = n3404 | n11345 ;
  assign n11347 = n11346 ^ n1005 ^ 1'b0 ;
  assign n11348 = ( n6151 & n11343 ) | ( n6151 & ~n11347 ) | ( n11343 & ~n11347 ) ;
  assign n11349 = ( ~x209 & n272 ) | ( ~x209 & n1791 ) | ( n272 & n1791 ) ;
  assign n11351 = n5363 ^ n3349 ^ n1238 ;
  assign n11350 = ( x159 & n1019 ) | ( x159 & n6696 ) | ( n1019 & n6696 ) ;
  assign n11352 = n11351 ^ n11350 ^ n2687 ;
  assign n11353 = ( ~n8998 & n11349 ) | ( ~n8998 & n11352 ) | ( n11349 & n11352 ) ;
  assign n11354 = ~n11348 & n11353 ;
  assign n11355 = n11341 & n11354 ;
  assign n11356 = n10214 ^ n1148 ^ 1'b0 ;
  assign n11357 = n11356 ^ n8670 ^ 1'b0 ;
  assign n11358 = ~n11355 & n11357 ;
  assign n11360 = n11359 ^ n11358 ^ n5572 ;
  assign n11361 = n10600 ^ n10010 ^ n2801 ;
  assign n11362 = n4000 ^ n1613 ^ 1'b0 ;
  assign n11363 = n11362 ^ n7577 ^ 1'b0 ;
  assign n11364 = n11361 & ~n11363 ;
  assign n11365 = n3792 ^ n3138 ^ n2807 ;
  assign n11366 = n11365 ^ n1386 ^ 1'b0 ;
  assign n11367 = n8353 ^ n5241 ^ 1'b0 ;
  assign n11368 = ~n3978 & n11367 ;
  assign n11369 = ~n2422 & n11368 ;
  assign n11375 = ( ~x35 & n2483 ) | ( ~x35 & n3875 ) | ( n2483 & n3875 ) ;
  assign n11370 = ( ~n3865 & n5723 ) | ( ~n3865 & n11299 ) | ( n5723 & n11299 ) ;
  assign n11371 = n6977 ^ n1373 ^ 1'b0 ;
  assign n11372 = ( ~n5258 & n10943 ) | ( ~n5258 & n11371 ) | ( n10943 & n11371 ) ;
  assign n11373 = n11372 ^ n7503 ^ n2175 ;
  assign n11374 = ( n1571 & ~n11370 ) | ( n1571 & n11373 ) | ( ~n11370 & n11373 ) ;
  assign n11376 = n11375 ^ n11374 ^ 1'b0 ;
  assign n11377 = ~n2081 & n11376 ;
  assign n11378 = ( x65 & n7570 ) | ( x65 & ~n8647 ) | ( n7570 & ~n8647 ) ;
  assign n11379 = n7941 | n11378 ;
  assign n11380 = ( n3999 & ~n4526 ) | ( n3999 & n9872 ) | ( ~n4526 & n9872 ) ;
  assign n11381 = ( n1515 & n11379 ) | ( n1515 & ~n11380 ) | ( n11379 & ~n11380 ) ;
  assign n11382 = n11381 ^ n7778 ^ n3887 ;
  assign n11383 = n3037 ^ x108 ^ 1'b0 ;
  assign n11384 = n7286 ^ n536 ^ 1'b0 ;
  assign n11385 = n10854 & n11384 ;
  assign n11386 = ( n4675 & ~n9331 ) | ( n4675 & n11385 ) | ( ~n9331 & n11385 ) ;
  assign n11387 = ( n6156 & n11383 ) | ( n6156 & n11386 ) | ( n11383 & n11386 ) ;
  assign n11388 = ( n11377 & ~n11382 ) | ( n11377 & n11387 ) | ( ~n11382 & n11387 ) ;
  assign n11389 = ~n5543 & n5843 ;
  assign n11390 = n3313 & n11389 ;
  assign n11391 = ( n4741 & n9898 ) | ( n4741 & ~n11390 ) | ( n9898 & ~n11390 ) ;
  assign n11392 = n6854 ^ n3560 ^ n1866 ;
  assign n11393 = n11392 ^ n4702 ^ n425 ;
  assign n11394 = n5028 ^ n1006 ^ 1'b0 ;
  assign n11395 = n340 | n11394 ;
  assign n11396 = ( n3732 & n7128 ) | ( n3732 & ~n11395 ) | ( n7128 & ~n11395 ) ;
  assign n11397 = n11393 & n11396 ;
  assign n11398 = ~n11391 & n11397 ;
  assign n11399 = n11398 ^ n2195 ^ 1'b0 ;
  assign n11400 = n2042 ^ n997 ^ x120 ;
  assign n11401 = n11400 ^ n6241 ^ n958 ;
  assign n11402 = ( n3787 & ~n7784 ) | ( n3787 & n11401 ) | ( ~n7784 & n11401 ) ;
  assign n11403 = ( n1671 & n4914 ) | ( n1671 & ~n8319 ) | ( n4914 & ~n8319 ) ;
  assign n11404 = ( ~n1229 & n2653 ) | ( ~n1229 & n11403 ) | ( n2653 & n11403 ) ;
  assign n11405 = n11404 ^ n5559 ^ n3151 ;
  assign n11406 = n7249 & n11405 ;
  assign n11407 = n2931 ^ n553 ^ 1'b0 ;
  assign n11408 = ( n5654 & n6376 ) | ( n5654 & ~n9358 ) | ( n6376 & ~n9358 ) ;
  assign n11409 = ( n8117 & n11407 ) | ( n8117 & ~n11408 ) | ( n11407 & ~n11408 ) ;
  assign n11410 = n11409 ^ n4876 ^ n2498 ;
  assign n11411 = ( n3343 & n3514 ) | ( n3343 & ~n11410 ) | ( n3514 & ~n11410 ) ;
  assign n11420 = n10401 ^ n7483 ^ n6958 ;
  assign n11416 = ( n1711 & n3180 ) | ( n1711 & n6963 ) | ( n3180 & n6963 ) ;
  assign n11417 = ~n3516 & n6674 ;
  assign n11418 = ( n2384 & n4147 ) | ( n2384 & n5151 ) | ( n4147 & n5151 ) ;
  assign n11419 = ( ~n11416 & n11417 ) | ( ~n11416 & n11418 ) | ( n11417 & n11418 ) ;
  assign n11412 = ( n1423 & n3777 ) | ( n1423 & n4887 ) | ( n3777 & n4887 ) ;
  assign n11413 = n11412 ^ n8272 ^ n1673 ;
  assign n11414 = ( n952 & n2105 ) | ( n952 & ~n9431 ) | ( n2105 & ~n9431 ) ;
  assign n11415 = ( ~n10126 & n11413 ) | ( ~n10126 & n11414 ) | ( n11413 & n11414 ) ;
  assign n11421 = n11420 ^ n11419 ^ n11415 ;
  assign n11422 = ( n11406 & n11411 ) | ( n11406 & ~n11421 ) | ( n11411 & ~n11421 ) ;
  assign n11423 = ( x138 & n2216 ) | ( x138 & n4978 ) | ( n2216 & n4978 ) ;
  assign n11424 = n11423 ^ n11095 ^ n3241 ;
  assign n11425 = n11283 ^ x188 ^ 1'b0 ;
  assign n11426 = ( n5884 & n11424 ) | ( n5884 & ~n11425 ) | ( n11424 & ~n11425 ) ;
  assign n11432 = ~n2004 & n4296 ;
  assign n11433 = n11432 ^ n5324 ^ 1'b0 ;
  assign n11434 = ( n377 & n4573 ) | ( n377 & n4860 ) | ( n4573 & n4860 ) ;
  assign n11435 = n3139 ^ n2917 ^ n1635 ;
  assign n11436 = n8426 & n11435 ;
  assign n11437 = ( n4391 & n11434 ) | ( n4391 & n11436 ) | ( n11434 & n11436 ) ;
  assign n11438 = ( ~n7733 & n11433 ) | ( ~n7733 & n11437 ) | ( n11433 & n11437 ) ;
  assign n11427 = ( n2254 & n3930 ) | ( n2254 & ~n6571 ) | ( n3930 & ~n6571 ) ;
  assign n11428 = n3739 & n4960 ;
  assign n11429 = n11427 & n11428 ;
  assign n11430 = n3648 & ~n11429 ;
  assign n11431 = n11430 ^ n10736 ^ 1'b0 ;
  assign n11439 = n11438 ^ n11431 ^ 1'b0 ;
  assign n11440 = n6655 ^ n5811 ^ n3152 ;
  assign n11441 = ( ~n2860 & n6314 ) | ( ~n2860 & n11440 ) | ( n6314 & n11440 ) ;
  assign n11442 = n2269 & n11441 ;
  assign n11443 = ~n5195 & n11442 ;
  assign n11444 = n4803 & ~n11443 ;
  assign n11445 = ~n11439 & n11444 ;
  assign n11451 = n3990 & ~n8629 ;
  assign n11452 = n11451 ^ n3317 ^ 1'b0 ;
  assign n11446 = n6639 ^ n3433 ^ n1614 ;
  assign n11447 = n5799 ^ n4293 ^ 1'b0 ;
  assign n11448 = ( n2272 & n4119 ) | ( n2272 & ~n11447 ) | ( n4119 & ~n11447 ) ;
  assign n11449 = n312 & n11448 ;
  assign n11450 = ( n7459 & n11446 ) | ( n7459 & n11449 ) | ( n11446 & n11449 ) ;
  assign n11453 = n11452 ^ n11450 ^ n3202 ;
  assign n11454 = ~n1722 & n3921 ;
  assign n11455 = ( ~n2303 & n3869 ) | ( ~n2303 & n11454 ) | ( n3869 & n11454 ) ;
  assign n11456 = n4916 & n6284 ;
  assign n11457 = n11456 ^ n8193 ^ 1'b0 ;
  assign n11458 = n11407 & n11457 ;
  assign n11459 = n5537 ^ n1706 ^ 1'b0 ;
  assign n11460 = ~n11458 & n11459 ;
  assign n11461 = n11460 ^ n2545 ^ 1'b0 ;
  assign n11462 = n7412 ^ n1557 ^ 1'b0 ;
  assign n11463 = n11462 ^ n6965 ^ n6061 ;
  assign n11464 = n11463 ^ n2823 ^ 1'b0 ;
  assign n11465 = n8025 & n11464 ;
  assign n11466 = ( n5134 & ~n8056 ) | ( n5134 & n11465 ) | ( ~n8056 & n11465 ) ;
  assign n11467 = ( n11455 & n11461 ) | ( n11455 & n11466 ) | ( n11461 & n11466 ) ;
  assign n11468 = n7303 ^ n1551 ^ n1445 ;
  assign n11469 = ( x146 & ~x252 ) | ( x146 & n11468 ) | ( ~x252 & n11468 ) ;
  assign n11470 = ( x69 & n3633 ) | ( x69 & ~n10987 ) | ( n3633 & ~n10987 ) ;
  assign n11471 = n11470 ^ n8656 ^ 1'b0 ;
  assign n11472 = n2237 ^ n990 ^ 1'b0 ;
  assign n11473 = n11472 ^ n4203 ^ n3950 ;
  assign n11474 = n2018 & n8732 ;
  assign n11475 = ( n11400 & n11473 ) | ( n11400 & n11474 ) | ( n11473 & n11474 ) ;
  assign n11476 = n11475 ^ n4444 ^ 1'b0 ;
  assign n11477 = ~n11471 & n11476 ;
  assign n11480 = n1774 & n9871 ;
  assign n11481 = n11480 ^ n2455 ^ 1'b0 ;
  assign n11482 = ( n1187 & ~n1918 ) | ( n1187 & n11481 ) | ( ~n1918 & n11481 ) ;
  assign n11478 = n5784 | n5873 ;
  assign n11479 = n7165 & n11478 ;
  assign n11483 = n11482 ^ n11479 ^ 1'b0 ;
  assign n11484 = ( ~n4162 & n4600 ) | ( ~n4162 & n9602 ) | ( n4600 & n9602 ) ;
  assign n11485 = n11484 ^ n9486 ^ 1'b0 ;
  assign n11486 = n8188 ^ n7746 ^ n4213 ;
  assign n11489 = ( ~n715 & n1705 ) | ( ~n715 & n3741 ) | ( n1705 & n3741 ) ;
  assign n11490 = n11489 ^ n4172 ^ x7 ;
  assign n11487 = n5155 ^ n1731 ^ 1'b0 ;
  assign n11488 = n11487 ^ n11299 ^ n7222 ;
  assign n11491 = n11490 ^ n11488 ^ n4234 ;
  assign n11492 = ( n10381 & n11486 ) | ( n10381 & n11491 ) | ( n11486 & n11491 ) ;
  assign n11493 = n11438 ^ n10500 ^ 1'b0 ;
  assign n11494 = n9653 ^ n5462 ^ n2876 ;
  assign n11495 = ( ~n4018 & n11493 ) | ( ~n4018 & n11494 ) | ( n11493 & n11494 ) ;
  assign n11496 = n2830 & n6426 ;
  assign n11497 = n11496 ^ n572 ^ 1'b0 ;
  assign n11498 = n11497 ^ n2631 ^ 1'b0 ;
  assign n11501 = n838 ^ n390 ^ 1'b0 ;
  assign n11502 = n5363 ^ n4968 ^ n3189 ;
  assign n11503 = ~n11501 & n11502 ;
  assign n11504 = n11503 ^ n3757 ^ 1'b0 ;
  assign n11499 = n2430 ^ n1271 ^ 1'b0 ;
  assign n11500 = n11499 ^ n3354 ^ 1'b0 ;
  assign n11505 = n11504 ^ n11500 ^ n5019 ;
  assign n11506 = n3865 | n10935 ;
  assign n11507 = n3045 | n11506 ;
  assign n11508 = n7088 ^ n4275 ^ n3930 ;
  assign n11509 = n10931 & ~n11508 ;
  assign n11510 = ~n11507 & n11509 ;
  assign n11511 = ~n5272 & n8431 ;
  assign n11512 = ( n4341 & n9764 ) | ( n4341 & n11511 ) | ( n9764 & n11511 ) ;
  assign n11516 = ( n2229 & n3085 ) | ( n2229 & ~n5845 ) | ( n3085 & ~n5845 ) ;
  assign n11517 = n1460 ^ n593 ^ 1'b0 ;
  assign n11518 = n11517 ^ n2574 ^ x9 ;
  assign n11519 = ( n1301 & n11516 ) | ( n1301 & n11518 ) | ( n11516 & n11518 ) ;
  assign n11513 = n8289 ^ n5705 ^ x116 ;
  assign n11514 = n11513 ^ n4798 ^ 1'b0 ;
  assign n11515 = ~n1113 & n11514 ;
  assign n11520 = n11519 ^ n11515 ^ n544 ;
  assign n11521 = n7484 ^ n6436 ^ n5909 ;
  assign n11522 = n10660 | n11521 ;
  assign n11533 = n6165 ^ n2491 ^ x140 ;
  assign n11531 = n3443 | n5725 ;
  assign n11530 = n7132 ^ n3266 ^ n868 ;
  assign n11532 = n11531 ^ n11530 ^ n2919 ;
  assign n11534 = n11533 ^ n11532 ^ n2580 ;
  assign n11523 = ( n2352 & n7635 ) | ( n2352 & ~n9120 ) | ( n7635 & ~n9120 ) ;
  assign n11524 = ( n2295 & ~n3021 ) | ( n2295 & n6031 ) | ( ~n3021 & n6031 ) ;
  assign n11525 = ( x16 & ~n1163 ) | ( x16 & n4745 ) | ( ~n1163 & n4745 ) ;
  assign n11526 = ~n11524 & n11525 ;
  assign n11527 = ~n3456 & n11526 ;
  assign n11528 = n11527 ^ n7412 ^ n5952 ;
  assign n11529 = n11523 & ~n11528 ;
  assign n11535 = n11534 ^ n11529 ^ 1'b0 ;
  assign n11536 = n11535 ^ n5792 ^ 1'b0 ;
  assign n11537 = n8722 & n11536 ;
  assign n11538 = n10302 ^ n10158 ^ 1'b0 ;
  assign n11539 = n8226 ^ n6199 ^ n4428 ;
  assign n11540 = ( n1126 & ~n3435 ) | ( n1126 & n5260 ) | ( ~n3435 & n5260 ) ;
  assign n11541 = ( ~n4017 & n11539 ) | ( ~n4017 & n11540 ) | ( n11539 & n11540 ) ;
  assign n11542 = n11541 ^ x110 ^ 1'b0 ;
  assign n11543 = ( n3305 & ~n5952 ) | ( n3305 & n6719 ) | ( ~n5952 & n6719 ) ;
  assign n11544 = n11543 ^ n1356 ^ 1'b0 ;
  assign n11545 = n10561 | n11544 ;
  assign n11546 = n9009 ^ n3616 ^ n2292 ;
  assign n11547 = ( n1625 & ~n4651 ) | ( n1625 & n5487 ) | ( ~n4651 & n5487 ) ;
  assign n11548 = n5180 & ~n6077 ;
  assign n11549 = ( n5943 & n10696 ) | ( n5943 & ~n11548 ) | ( n10696 & ~n11548 ) ;
  assign n11550 = ( ~n6427 & n9231 ) | ( ~n6427 & n11549 ) | ( n9231 & n11549 ) ;
  assign n11552 = n1604 | n5714 ;
  assign n11553 = n1649 & ~n11552 ;
  assign n11551 = n10583 ^ n7507 ^ n5982 ;
  assign n11554 = n11553 ^ n11551 ^ n8077 ;
  assign n11555 = ( n11245 & ~n11550 ) | ( n11245 & n11554 ) | ( ~n11550 & n11554 ) ;
  assign n11556 = ( n5858 & n11547 ) | ( n5858 & n11555 ) | ( n11547 & n11555 ) ;
  assign n11557 = n10763 ^ n6099 ^ x49 ;
  assign n11558 = n11557 ^ n3749 ^ x68 ;
  assign n11559 = n2188 & ~n11006 ;
  assign n11560 = ~n10055 & n11559 ;
  assign n11561 = n4704 ^ n3431 ^ n2575 ;
  assign n11562 = n6969 ^ n408 ^ 1'b0 ;
  assign n11563 = n11561 & ~n11562 ;
  assign n11564 = ~n2663 & n6240 ;
  assign n11565 = n882 | n899 ;
  assign n11566 = ( n548 & ~n4684 ) | ( n548 & n11565 ) | ( ~n4684 & n11565 ) ;
  assign n11567 = n11566 ^ n4701 ^ n4642 ;
  assign n11568 = n11567 ^ n1840 ^ 1'b0 ;
  assign n11569 = n11564 & n11568 ;
  assign n11570 = n5800 ^ n5253 ^ n2606 ;
  assign n11571 = n7816 ^ n636 ^ 1'b0 ;
  assign n11572 = n3835 & n11571 ;
  assign n11573 = ( n4841 & n5104 ) | ( n4841 & n11572 ) | ( n5104 & n11572 ) ;
  assign n11574 = ( n430 & n6577 ) | ( n430 & ~n11573 ) | ( n6577 & ~n11573 ) ;
  assign n11575 = n11570 & ~n11574 ;
  assign n11576 = n11035 & n11575 ;
  assign n11577 = n10447 ^ n5540 ^ n643 ;
  assign n11582 = n4257 ^ n2828 ^ n1077 ;
  assign n11580 = ( n876 & n1566 ) | ( n876 & ~n4769 ) | ( n1566 & ~n4769 ) ;
  assign n11579 = ( n1437 & n4609 ) | ( n1437 & n7082 ) | ( n4609 & n7082 ) ;
  assign n11578 = n10264 ^ n9173 ^ n938 ;
  assign n11581 = n11580 ^ n11579 ^ n11578 ;
  assign n11583 = n11582 ^ n11581 ^ n3790 ;
  assign n11584 = n9074 ^ n5875 ^ 1'b0 ;
  assign n11585 = n11583 & ~n11584 ;
  assign n11586 = ( n11576 & n11577 ) | ( n11576 & n11585 ) | ( n11577 & n11585 ) ;
  assign n11587 = n11586 ^ n8011 ^ n287 ;
  assign n11591 = ( n1623 & n3107 ) | ( n1623 & ~n5967 ) | ( n3107 & ~n5967 ) ;
  assign n11592 = ( n580 & n7058 ) | ( n580 & n10578 ) | ( n7058 & n10578 ) ;
  assign n11593 = ( n10258 & n11591 ) | ( n10258 & ~n11592 ) | ( n11591 & ~n11592 ) ;
  assign n11594 = n11593 ^ n6752 ^ 1'b0 ;
  assign n11588 = n1487 | n1562 ;
  assign n11589 = n11588 ^ n10447 ^ n5143 ;
  assign n11590 = n11237 & ~n11589 ;
  assign n11595 = n11594 ^ n11590 ^ 1'b0 ;
  assign n11619 = n8828 ^ n3207 ^ 1'b0 ;
  assign n11620 = n11619 ^ n3080 ^ 1'b0 ;
  assign n11621 = n4345 & ~n11620 ;
  assign n11597 = ( ~n1478 & n3925 ) | ( ~n1478 & n6910 ) | ( n3925 & n6910 ) ;
  assign n11598 = n4612 & ~n5777 ;
  assign n11599 = n10407 | n11598 ;
  assign n11600 = n11597 | n11599 ;
  assign n11596 = n800 & n2535 ;
  assign n11601 = n11600 ^ n11596 ^ 1'b0 ;
  assign n11602 = n11601 ^ n10292 ^ 1'b0 ;
  assign n11603 = n10057 & n11140 ;
  assign n11604 = n11603 ^ n1211 ^ 1'b0 ;
  assign n11605 = n3826 | n9353 ;
  assign n11606 = n11605 ^ n4133 ^ n4051 ;
  assign n11607 = ( n3680 & n5761 ) | ( n3680 & n6926 ) | ( n5761 & n6926 ) ;
  assign n11608 = ( x53 & n7562 ) | ( x53 & ~n11607 ) | ( n7562 & ~n11607 ) ;
  assign n11609 = ( ~n1975 & n11606 ) | ( ~n1975 & n11608 ) | ( n11606 & n11608 ) ;
  assign n11612 = ( n536 & n1007 ) | ( n536 & ~n1950 ) | ( n1007 & ~n1950 ) ;
  assign n11610 = ( n1719 & n2787 ) | ( n1719 & ~n5024 ) | ( n2787 & ~n5024 ) ;
  assign n11611 = n11610 ^ n7346 ^ n5736 ;
  assign n11613 = n11612 ^ n11611 ^ n6067 ;
  assign n11614 = ( n2141 & n6891 ) | ( n2141 & ~n11613 ) | ( n6891 & ~n11613 ) ;
  assign n11615 = n11614 ^ n1266 ^ 1'b0 ;
  assign n11616 = ( n1322 & ~n11609 ) | ( n1322 & n11615 ) | ( ~n11609 & n11615 ) ;
  assign n11617 = ( n8764 & n11604 ) | ( n8764 & n11616 ) | ( n11604 & n11616 ) ;
  assign n11618 = n11602 & ~n11617 ;
  assign n11622 = n11621 ^ n11618 ^ 1'b0 ;
  assign n11623 = ( n406 & n3894 ) | ( n406 & n5564 ) | ( n3894 & n5564 ) ;
  assign n11626 = ( n3455 & ~n5858 ) | ( n3455 & n7032 ) | ( ~n5858 & n7032 ) ;
  assign n11627 = ( ~n1690 & n7025 ) | ( ~n1690 & n11626 ) | ( n7025 & n11626 ) ;
  assign n11624 = n7880 ^ n7324 ^ n1106 ;
  assign n11625 = n11624 ^ n7377 ^ n1509 ;
  assign n11628 = n11627 ^ n11625 ^ n6069 ;
  assign n11632 = ( n792 & n7331 ) | ( n792 & ~n9399 ) | ( n7331 & ~n9399 ) ;
  assign n11633 = ( n959 & n5283 ) | ( n959 & ~n10918 ) | ( n5283 & ~n10918 ) ;
  assign n11634 = ( n1266 & n10455 ) | ( n1266 & ~n11633 ) | ( n10455 & ~n11633 ) ;
  assign n11635 = n11632 & ~n11634 ;
  assign n11636 = n11635 ^ n6103 ^ 1'b0 ;
  assign n11629 = n3355 & n6366 ;
  assign n11630 = n11629 ^ n1271 ^ 1'b0 ;
  assign n11631 = ( ~n2633 & n10785 ) | ( ~n2633 & n11630 ) | ( n10785 & n11630 ) ;
  assign n11637 = n11636 ^ n11631 ^ 1'b0 ;
  assign n11638 = n4378 & ~n11637 ;
  assign n11639 = n4703 ^ n3074 ^ x60 ;
  assign n11640 = ( n2834 & ~n4625 ) | ( n2834 & n6048 ) | ( ~n4625 & n6048 ) ;
  assign n11641 = n5142 ^ n951 ^ x130 ;
  assign n11642 = n11641 ^ n5085 ^ 1'b0 ;
  assign n11643 = ~n5962 & n11642 ;
  assign n11644 = n2757 ^ n660 ^ 1'b0 ;
  assign n11645 = n1863 & ~n11644 ;
  assign n11646 = ( n1436 & n2940 ) | ( n1436 & n11645 ) | ( n2940 & n11645 ) ;
  assign n11647 = ( n4787 & ~n5144 ) | ( n4787 & n11455 ) | ( ~n5144 & n11455 ) ;
  assign n11648 = ( n7168 & n11646 ) | ( n7168 & ~n11647 ) | ( n11646 & ~n11647 ) ;
  assign n11649 = n11648 ^ n1026 ^ 1'b0 ;
  assign n11650 = n11488 ^ n7072 ^ n2905 ;
  assign n11651 = ( n1332 & n1979 ) | ( n1332 & n7009 ) | ( n1979 & n7009 ) ;
  assign n11652 = ( ~n1935 & n11650 ) | ( ~n1935 & n11651 ) | ( n11650 & n11651 ) ;
  assign n11661 = n10161 ^ n4166 ^ 1'b0 ;
  assign n11653 = n3554 | n10656 ;
  assign n11654 = n11653 ^ n3100 ^ 1'b0 ;
  assign n11655 = n1595 | n2636 ;
  assign n11656 = n11655 ^ n480 ^ 1'b0 ;
  assign n11657 = ( n6164 & n6222 ) | ( n6164 & ~n11656 ) | ( n6222 & ~n11656 ) ;
  assign n11658 = n2566 & ~n11657 ;
  assign n11659 = n11658 ^ n3067 ^ 1'b0 ;
  assign n11660 = ( n9296 & n11654 ) | ( n9296 & ~n11659 ) | ( n11654 & ~n11659 ) ;
  assign n11662 = n11661 ^ n11660 ^ n1292 ;
  assign n11663 = n2879 & ~n4454 ;
  assign n11664 = n2134 & n11663 ;
  assign n11665 = n10946 | n11664 ;
  assign n11666 = n1104 & ~n11665 ;
  assign n11667 = n2396 | n9057 ;
  assign n11668 = n11667 ^ n11408 ^ 1'b0 ;
  assign n11669 = ( n3766 & ~n7708 ) | ( n3766 & n11668 ) | ( ~n7708 & n11668 ) ;
  assign n11670 = ( n4864 & ~n7945 ) | ( n4864 & n9384 ) | ( ~n7945 & n9384 ) ;
  assign n11674 = n10888 ^ n10694 ^ n555 ;
  assign n11675 = n11674 ^ n8871 ^ n4991 ;
  assign n11672 = n4866 ^ n2030 ^ n558 ;
  assign n11671 = n9120 ^ n2062 ^ n1475 ;
  assign n11673 = n11672 ^ n11671 ^ n785 ;
  assign n11676 = n11675 ^ n11673 ^ n9884 ;
  assign n11677 = ( n4929 & n6042 ) | ( n4929 & n7210 ) | ( n6042 & n7210 ) ;
  assign n11678 = n11677 ^ n10897 ^ 1'b0 ;
  assign n11679 = ( n1432 & n1712 ) | ( n1432 & n4405 ) | ( n1712 & n4405 ) ;
  assign n11680 = n11679 ^ n10569 ^ n1836 ;
  assign n11681 = ( n10140 & n11678 ) | ( n10140 & n11680 ) | ( n11678 & n11680 ) ;
  assign n11682 = ( n5490 & n11238 ) | ( n5490 & ~n11681 ) | ( n11238 & ~n11681 ) ;
  assign n11683 = n5583 ^ n3421 ^ n1139 ;
  assign n11684 = ( n373 & n392 ) | ( n373 & n1863 ) | ( n392 & n1863 ) ;
  assign n11685 = ( n417 & ~n1532 ) | ( n417 & n4337 ) | ( ~n1532 & n4337 ) ;
  assign n11686 = ( n1424 & ~n2029 ) | ( n1424 & n3093 ) | ( ~n2029 & n3093 ) ;
  assign n11687 = ( n932 & n7741 ) | ( n932 & ~n11686 ) | ( n7741 & ~n11686 ) ;
  assign n11688 = ( ~n11684 & n11685 ) | ( ~n11684 & n11687 ) | ( n11685 & n11687 ) ;
  assign n11689 = n3194 & ~n8350 ;
  assign n11690 = ( ~n3794 & n5326 ) | ( ~n3794 & n11689 ) | ( n5326 & n11689 ) ;
  assign n11691 = n11690 ^ n11127 ^ n3413 ;
  assign n11692 = ( n2170 & n11688 ) | ( n2170 & ~n11691 ) | ( n11688 & ~n11691 ) ;
  assign n11693 = ( ~n7105 & n11683 ) | ( ~n7105 & n11692 ) | ( n11683 & n11692 ) ;
  assign n11695 = n2895 ^ n2138 ^ 1'b0 ;
  assign n11696 = n7669 ^ n1961 ^ 1'b0 ;
  assign n11697 = ( n868 & ~n11695 ) | ( n868 & n11696 ) | ( ~n11695 & n11696 ) ;
  assign n11698 = n11697 ^ n6459 ^ x153 ;
  assign n11699 = ( n4298 & n9025 ) | ( n4298 & ~n11698 ) | ( n9025 & ~n11698 ) ;
  assign n11694 = n2472 | n8337 ;
  assign n11700 = n11699 ^ n11694 ^ 1'b0 ;
  assign n11708 = n6299 ^ n3126 ^ n1802 ;
  assign n11709 = ( n8180 & n8994 ) | ( n8180 & ~n11708 ) | ( n8994 & ~n11708 ) ;
  assign n11701 = ( n1306 & n2746 ) | ( n1306 & ~n6856 ) | ( n2746 & ~n6856 ) ;
  assign n11702 = n11701 ^ n4043 ^ n1442 ;
  assign n11703 = n607 & n5045 ;
  assign n11704 = n11703 ^ n11231 ^ 1'b0 ;
  assign n11705 = n6497 | n7519 ;
  assign n11706 = n11704 & ~n11705 ;
  assign n11707 = ( n7530 & n11702 ) | ( n7530 & ~n11706 ) | ( n11702 & ~n11706 ) ;
  assign n11710 = n11709 ^ n11707 ^ n11661 ;
  assign n11711 = n4176 | n4685 ;
  assign n11712 = n11711 ^ n464 ^ 1'b0 ;
  assign n11713 = n1557 & n11712 ;
  assign n11714 = n2082 ^ n1101 ^ 1'b0 ;
  assign n11715 = n11714 ^ n2006 ^ x107 ;
  assign n11716 = n1631 & ~n11715 ;
  assign n11717 = n11716 ^ n6158 ^ n666 ;
  assign n11718 = n10380 & n11717 ;
  assign n11719 = ~n8817 & n11718 ;
  assign n11720 = ( n1405 & n4163 ) | ( n1405 & n8734 ) | ( n4163 & n8734 ) ;
  assign n11721 = n11720 ^ n10315 ^ n7679 ;
  assign n11722 = n8213 ^ n4266 ^ n645 ;
  assign n11723 = n11722 ^ n308 ^ 1'b0 ;
  assign n11724 = n5724 | n11723 ;
  assign n11725 = ( ~n3940 & n10301 ) | ( ~n3940 & n11724 ) | ( n10301 & n11724 ) ;
  assign n11726 = ( n1517 & n2052 ) | ( n1517 & n6094 ) | ( n2052 & n6094 ) ;
  assign n11727 = n6686 & n7632 ;
  assign n11728 = ~n4559 & n11727 ;
  assign n11729 = n6625 ^ n5505 ^ n4508 ;
  assign n11730 = ( n7892 & n9440 ) | ( n7892 & ~n11729 ) | ( n9440 & ~n11729 ) ;
  assign n11731 = ( n4652 & n11728 ) | ( n4652 & ~n11730 ) | ( n11728 & ~n11730 ) ;
  assign n11734 = n5258 ^ n4252 ^ 1'b0 ;
  assign n11735 = n5880 & n11734 ;
  assign n11736 = n11735 ^ n3768 ^ 1'b0 ;
  assign n11732 = ( ~n866 & n2982 ) | ( ~n866 & n4985 ) | ( n2982 & n4985 ) ;
  assign n11733 = ( n788 & n2283 ) | ( n788 & ~n11732 ) | ( n2283 & ~n11732 ) ;
  assign n11737 = n11736 ^ n11733 ^ n10194 ;
  assign n11740 = n10214 ^ n9085 ^ n8077 ;
  assign n11741 = n8646 ^ n1029 ^ 1'b0 ;
  assign n11742 = ~n3408 & n11741 ;
  assign n11743 = ( ~n8511 & n11740 ) | ( ~n8511 & n11742 ) | ( n11740 & n11742 ) ;
  assign n11744 = ( n596 & ~n1393 ) | ( n596 & n11227 ) | ( ~n1393 & n11227 ) ;
  assign n11745 = n4681 | n11744 ;
  assign n11746 = n11743 | n11745 ;
  assign n11747 = ( n3095 & n5174 ) | ( n3095 & ~n11746 ) | ( n5174 & ~n11746 ) ;
  assign n11738 = n11702 ^ n1456 ^ 1'b0 ;
  assign n11739 = n1766 & ~n11738 ;
  assign n11748 = n11747 ^ n11739 ^ n10786 ;
  assign n11749 = n11249 ^ n4217 ^ n341 ;
  assign n11750 = n11749 ^ n5833 ^ n1477 ;
  assign n11751 = n11750 ^ n2515 ^ n735 ;
  assign n11752 = n10502 ^ n2192 ^ n1473 ;
  assign n11753 = n4907 ^ n4689 ^ n334 ;
  assign n11754 = ( n3699 & ~n4357 ) | ( n3699 & n6465 ) | ( ~n4357 & n6465 ) ;
  assign n11755 = ( n867 & n1814 ) | ( n867 & ~n11754 ) | ( n1814 & ~n11754 ) ;
  assign n11759 = n7390 ^ n3497 ^ 1'b0 ;
  assign n11760 = ~n6649 & n11759 ;
  assign n11756 = ~n6740 & n9813 ;
  assign n11757 = n11756 ^ n4523 ^ 1'b0 ;
  assign n11758 = n11757 ^ n2801 ^ 1'b0 ;
  assign n11761 = n11760 ^ n11758 ^ n1207 ;
  assign n11762 = n11755 | n11761 ;
  assign n11763 = n11762 ^ n380 ^ 1'b0 ;
  assign n11764 = n11753 | n11763 ;
  assign n11765 = n11764 ^ n10740 ^ 1'b0 ;
  assign n11766 = n6965 & ~n6993 ;
  assign n11767 = n11766 ^ n3770 ^ n2982 ;
  assign n11768 = ( ~n7499 & n9739 ) | ( ~n7499 & n11767 ) | ( n9739 & n11767 ) ;
  assign n11769 = n8687 ^ n6687 ^ x100 ;
  assign n11770 = n11769 ^ n1824 ^ n1582 ;
  assign n11771 = n11770 ^ n8391 ^ n961 ;
  assign n11773 = ~x214 & n9585 ;
  assign n11772 = ( n1131 & n1135 ) | ( n1131 & n8127 ) | ( n1135 & n8127 ) ;
  assign n11774 = n11773 ^ n11772 ^ n4642 ;
  assign n11775 = n391 & n1839 ;
  assign n11776 = n10845 & n11775 ;
  assign n11777 = ( x99 & n1620 ) | ( x99 & ~n11776 ) | ( n1620 & ~n11776 ) ;
  assign n11778 = ~n3978 & n5140 ;
  assign n11779 = n11778 ^ n5966 ^ 1'b0 ;
  assign n11780 = n4014 ^ n1190 ^ n269 ;
  assign n11781 = n11780 ^ n10431 ^ n3539 ;
  assign n11782 = ( ~n1342 & n10705 ) | ( ~n1342 & n11781 ) | ( n10705 & n11781 ) ;
  assign n11783 = n4072 ^ n3807 ^ n3493 ;
  assign n11784 = ( n3459 & ~n3929 ) | ( n3459 & n7613 ) | ( ~n3929 & n7613 ) ;
  assign n11785 = ( x62 & n2459 ) | ( x62 & ~n8896 ) | ( n2459 & ~n8896 ) ;
  assign n11786 = n3646 & n11785 ;
  assign n11787 = n11786 ^ n6399 ^ n4685 ;
  assign n11788 = ~n3422 & n11787 ;
  assign n11789 = n11788 ^ n8352 ^ 1'b0 ;
  assign n11790 = ( ~n11783 & n11784 ) | ( ~n11783 & n11789 ) | ( n11784 & n11789 ) ;
  assign n11791 = ( n3063 & n3634 ) | ( n3063 & ~n8250 ) | ( n3634 & ~n8250 ) ;
  assign n11792 = n1148 & n2499 ;
  assign n11793 = ~n11791 & n11792 ;
  assign n11794 = n7979 ^ n5224 ^ 1'b0 ;
  assign n11795 = n11794 ^ n10698 ^ n1112 ;
  assign n11796 = ( ~n5667 & n7747 ) | ( ~n5667 & n7838 ) | ( n7747 & n7838 ) ;
  assign n11797 = n11796 ^ n3174 ^ n2978 ;
  assign n11798 = ~n3796 & n7251 ;
  assign n11799 = ( n4520 & ~n10372 ) | ( n4520 & n11798 ) | ( ~n10372 & n11798 ) ;
  assign n11800 = n1654 | n1828 ;
  assign n11801 = n10840 | n11800 ;
  assign n11802 = n11801 ^ n5800 ^ n3982 ;
  assign n11803 = ( ~n336 & n11799 ) | ( ~n336 & n11802 ) | ( n11799 & n11802 ) ;
  assign n11804 = ( n599 & n4095 ) | ( n599 & ~n7669 ) | ( n4095 & ~n7669 ) ;
  assign n11805 = ( n7445 & n10335 ) | ( n7445 & ~n11804 ) | ( n10335 & ~n11804 ) ;
  assign n11806 = n1733 & ~n2017 ;
  assign n11807 = ( ~n4713 & n5000 ) | ( ~n4713 & n11806 ) | ( n5000 & n11806 ) ;
  assign n11808 = ( n3948 & n10728 ) | ( n3948 & n11807 ) | ( n10728 & n11807 ) ;
  assign n11809 = ( n1912 & n2950 ) | ( n1912 & ~n7319 ) | ( n2950 & ~n7319 ) ;
  assign n11810 = n11809 ^ n7600 ^ 1'b0 ;
  assign n11811 = n11808 | n11810 ;
  assign n11812 = n10046 ^ n2305 ^ n2289 ;
  assign n11813 = ( n5937 & n8169 ) | ( n5937 & ~n11057 ) | ( n8169 & ~n11057 ) ;
  assign n11814 = ( ~n4705 & n11812 ) | ( ~n4705 & n11813 ) | ( n11812 & n11813 ) ;
  assign n11815 = ( n4684 & n6312 ) | ( n4684 & n11814 ) | ( n6312 & n11814 ) ;
  assign n11816 = n8930 ^ n7141 ^ n2536 ;
  assign n11817 = ~n5871 & n11816 ;
  assign n11825 = n1492 ^ n1353 ^ n1204 ;
  assign n11826 = n11825 ^ n3759 ^ n2762 ;
  assign n11818 = n10067 ^ n2235 ^ n682 ;
  assign n11819 = n3644 ^ n1405 ^ 1'b0 ;
  assign n11820 = n11818 & n11819 ;
  assign n11821 = n11820 ^ n7685 ^ n3884 ;
  assign n11822 = ( n5999 & ~n9556 ) | ( n5999 & n11821 ) | ( ~n9556 & n11821 ) ;
  assign n11823 = n1325 | n11822 ;
  assign n11824 = n8118 | n11823 ;
  assign n11827 = n11826 ^ n11824 ^ n1959 ;
  assign n11828 = n8470 ^ n4335 ^ n3631 ;
  assign n11829 = n4694 | n11828 ;
  assign n11830 = ( ~n1851 & n9481 ) | ( ~n1851 & n11829 ) | ( n9481 & n11829 ) ;
  assign n11831 = n11830 ^ n8000 ^ n6302 ;
  assign n11832 = ( ~n3375 & n6494 ) | ( ~n3375 & n6621 ) | ( n6494 & n6621 ) ;
  assign n11833 = ( n4207 & n8806 ) | ( n4207 & ~n11832 ) | ( n8806 & ~n11832 ) ;
  assign n11834 = n635 & ~n11833 ;
  assign n11835 = n6313 ^ n5584 ^ n2863 ;
  assign n11836 = ~n10257 & n11835 ;
  assign n11837 = ( n11822 & ~n11834 ) | ( n11822 & n11836 ) | ( ~n11834 & n11836 ) ;
  assign n11838 = ( n1695 & n2849 ) | ( n1695 & ~n11783 ) | ( n2849 & ~n11783 ) ;
  assign n11839 = ( ~n1979 & n2688 ) | ( ~n1979 & n11838 ) | ( n2688 & n11838 ) ;
  assign n11840 = ~n1344 & n6195 ;
  assign n11841 = n11840 ^ n8359 ^ n4397 ;
  assign n11842 = n11841 ^ n2024 ^ 1'b0 ;
  assign n11843 = n11839 & n11842 ;
  assign n11844 = ( n1169 & n4159 ) | ( n1169 & ~n5630 ) | ( n4159 & ~n5630 ) ;
  assign n11845 = ( n635 & n4164 ) | ( n635 & n11084 ) | ( n4164 & n11084 ) ;
  assign n11846 = n1879 ^ n1541 ^ n282 ;
  assign n11847 = ~n8405 & n11846 ;
  assign n11849 = ( n5924 & ~n6110 ) | ( n5924 & n10843 ) | ( ~n6110 & n10843 ) ;
  assign n11848 = n7354 ^ n6971 ^ 1'b0 ;
  assign n11850 = n11849 ^ n11848 ^ n1598 ;
  assign n11851 = ( ~n2147 & n11847 ) | ( ~n2147 & n11850 ) | ( n11847 & n11850 ) ;
  assign n11852 = n11851 ^ n7581 ^ 1'b0 ;
  assign n11853 = ( n6294 & n11845 ) | ( n6294 & n11852 ) | ( n11845 & n11852 ) ;
  assign n11854 = n5251 ^ n455 ^ 1'b0 ;
  assign n11855 = n8087 & ~n11854 ;
  assign n11856 = n9033 ^ n2521 ^ 1'b0 ;
  assign n11857 = n542 & ~n11856 ;
  assign n11858 = ( n290 & n2883 ) | ( n290 & n11857 ) | ( n2883 & n11857 ) ;
  assign n11859 = n11855 | n11858 ;
  assign n11860 = x130 & ~n5660 ;
  assign n11861 = n1163 & n11860 ;
  assign n11862 = n11861 ^ n3425 ^ 1'b0 ;
  assign n11867 = ( n1916 & n2467 ) | ( n1916 & ~n2923 ) | ( n2467 & ~n2923 ) ;
  assign n11863 = n4878 ^ n4142 ^ 1'b0 ;
  assign n11864 = ~n6223 & n11863 ;
  assign n11865 = n378 & ~n11864 ;
  assign n11866 = ( n3883 & ~n5028 ) | ( n3883 & n11865 ) | ( ~n5028 & n11865 ) ;
  assign n11868 = n11867 ^ n11866 ^ n6821 ;
  assign n11869 = ( n7687 & n11862 ) | ( n7687 & ~n11868 ) | ( n11862 & ~n11868 ) ;
  assign n11870 = n2744 ^ n2664 ^ n2217 ;
  assign n11871 = ( n1379 & n6938 ) | ( n1379 & n7570 ) | ( n6938 & n7570 ) ;
  assign n11872 = ( ~n839 & n3408 ) | ( ~n839 & n11871 ) | ( n3408 & n11871 ) ;
  assign n11873 = ( n4674 & ~n9097 ) | ( n4674 & n11872 ) | ( ~n9097 & n11872 ) ;
  assign n11874 = n6917 ^ n5834 ^ n4379 ;
  assign n11875 = n2334 | n4181 ;
  assign n11876 = n4403 & ~n11875 ;
  assign n11877 = n1153 & ~n6549 ;
  assign n11891 = n10619 ^ n2276 ^ 1'b0 ;
  assign n11892 = ~n1882 & n11891 ;
  assign n11890 = ( n3924 & n4348 ) | ( n3924 & ~n5324 ) | ( n4348 & ~n5324 ) ;
  assign n11878 = n3996 ^ n286 ^ 1'b0 ;
  assign n11879 = n1787 & ~n11878 ;
  assign n11880 = n1132 ^ n790 ^ n336 ;
  assign n11881 = n1845 & ~n7282 ;
  assign n11882 = ( n1225 & n11880 ) | ( n1225 & n11881 ) | ( n11880 & n11881 ) ;
  assign n11883 = ( n3229 & n6317 ) | ( n3229 & ~n11882 ) | ( n6317 & ~n11882 ) ;
  assign n11884 = ~n1009 & n2341 ;
  assign n11885 = n11884 ^ n413 ^ 1'b0 ;
  assign n11886 = ( n838 & n11883 ) | ( n838 & n11885 ) | ( n11883 & n11885 ) ;
  assign n11887 = n4854 ^ n4821 ^ n1310 ;
  assign n11888 = n11887 ^ n6951 ^ n6022 ;
  assign n11889 = ( n11879 & ~n11886 ) | ( n11879 & n11888 ) | ( ~n11886 & n11888 ) ;
  assign n11893 = n11892 ^ n11890 ^ n11889 ;
  assign n11894 = ( n11876 & n11877 ) | ( n11876 & ~n11893 ) | ( n11877 & ~n11893 ) ;
  assign n11902 = n7667 ^ n5547 ^ 1'b0 ;
  assign n11903 = ( ~n5127 & n5899 ) | ( ~n5127 & n11902 ) | ( n5899 & n11902 ) ;
  assign n11899 = ( ~n2052 & n2917 ) | ( ~n2052 & n5162 ) | ( n2917 & n5162 ) ;
  assign n11898 = n8503 ^ n1588 ^ 1'b0 ;
  assign n11900 = n11899 ^ n11898 ^ n10421 ;
  assign n11895 = ( ~n1048 & n2517 ) | ( ~n1048 & n3709 ) | ( n2517 & n3709 ) ;
  assign n11896 = n11895 ^ n10196 ^ 1'b0 ;
  assign n11897 = n9010 & n11896 ;
  assign n11901 = n11900 ^ n11897 ^ n8120 ;
  assign n11904 = n11903 ^ n11901 ^ n5418 ;
  assign n11905 = n551 & n7562 ;
  assign n11906 = n9020 ^ n4152 ^ n3204 ;
  assign n11907 = ( n5844 & ~n7040 ) | ( n5844 & n11906 ) | ( ~n7040 & n11906 ) ;
  assign n11908 = ~n3028 & n3345 ;
  assign n11909 = n11908 ^ n4597 ^ 1'b0 ;
  assign n11910 = n1012 | n11909 ;
  assign n11911 = n4375 | n11910 ;
  assign n11912 = n11911 ^ n7572 ^ n1194 ;
  assign n11913 = ( n7433 & n11907 ) | ( n7433 & n11912 ) | ( n11907 & n11912 ) ;
  assign n11916 = n3563 ^ n3364 ^ 1'b0 ;
  assign n11917 = n686 & n11916 ;
  assign n11918 = n11917 ^ n5559 ^ n307 ;
  assign n11919 = ( n465 & ~n1585 ) | ( n465 & n11918 ) | ( ~n1585 & n11918 ) ;
  assign n11914 = n10072 ^ n5531 ^ n4999 ;
  assign n11915 = n11914 ^ n7762 ^ n6991 ;
  assign n11920 = n11919 ^ n11915 ^ n5652 ;
  assign n11921 = n2209 ^ n1686 ^ n1519 ;
  assign n11922 = ( ~n413 & n5829 ) | ( ~n413 & n10119 ) | ( n5829 & n10119 ) ;
  assign n11923 = ( ~n7166 & n11921 ) | ( ~n7166 & n11922 ) | ( n11921 & n11922 ) ;
  assign n11924 = n11923 ^ n11128 ^ n1737 ;
  assign n11925 = n5194 ^ n2899 ^ n2132 ;
  assign n11926 = ( ~n2227 & n5357 ) | ( ~n2227 & n10084 ) | ( n5357 & n10084 ) ;
  assign n11927 = ~n3938 & n11926 ;
  assign n11928 = ~n272 & n11927 ;
  assign n11929 = ( n2176 & n7168 ) | ( n2176 & ~n11928 ) | ( n7168 & ~n11928 ) ;
  assign n11930 = n10337 ^ n4254 ^ n3867 ;
  assign n11931 = ( n4987 & n11929 ) | ( n4987 & ~n11930 ) | ( n11929 & ~n11930 ) ;
  assign n11932 = ( n9821 & n11925 ) | ( n9821 & n11931 ) | ( n11925 & n11931 ) ;
  assign n11933 = ( ~n1462 & n3322 ) | ( ~n1462 & n7497 ) | ( n3322 & n7497 ) ;
  assign n11934 = n8283 & ~n11933 ;
  assign n11935 = ~n295 & n11934 ;
  assign n11936 = n10723 ^ n10209 ^ n4511 ;
  assign n11937 = ( n464 & n2383 ) | ( n464 & ~n11936 ) | ( n2383 & ~n11936 ) ;
  assign n11938 = ( n2500 & n11935 ) | ( n2500 & n11937 ) | ( n11935 & n11937 ) ;
  assign n11939 = ~x150 & n11645 ;
  assign n11940 = ( n1617 & n8439 ) | ( n1617 & ~n11939 ) | ( n8439 & ~n11939 ) ;
  assign n11941 = n578 ^ x174 ^ 1'b0 ;
  assign n11942 = n11940 | n11941 ;
  assign n11943 = n11942 ^ n2835 ^ 1'b0 ;
  assign n11944 = n5812 & n11943 ;
  assign n11945 = n4997 ^ n412 ^ 1'b0 ;
  assign n11946 = n11944 & ~n11945 ;
  assign n11948 = n10309 ^ n9804 ^ n3376 ;
  assign n11949 = n7209 ^ n3884 ^ n2231 ;
  assign n11950 = ( n1626 & n7139 ) | ( n1626 & n11949 ) | ( n7139 & n11949 ) ;
  assign n11951 = n11950 ^ n3174 ^ n1686 ;
  assign n11952 = n7957 ^ n7394 ^ n1765 ;
  assign n11953 = ( n1860 & n4843 ) | ( n1860 & ~n11952 ) | ( n4843 & ~n11952 ) ;
  assign n11954 = ( n11948 & n11951 ) | ( n11948 & ~n11953 ) | ( n11951 & ~n11953 ) ;
  assign n11947 = n1133 & ~n8010 ;
  assign n11955 = n11954 ^ n11947 ^ 1'b0 ;
  assign n11956 = n11683 ^ n9875 ^ n6458 ;
  assign n11957 = n6218 ^ n2612 ^ 1'b0 ;
  assign n11958 = n766 | n11957 ;
  assign n11959 = n11958 ^ n3324 ^ 1'b0 ;
  assign n11960 = n3544 ^ n2509 ^ 1'b0 ;
  assign n11966 = n11433 ^ n10893 ^ n3924 ;
  assign n11963 = n10439 ^ n5507 ^ x209 ;
  assign n11964 = ( x198 & n1310 ) | ( x198 & n11963 ) | ( n1310 & n11963 ) ;
  assign n11965 = n11964 ^ n11311 ^ n5890 ;
  assign n11961 = x192 & n8737 ;
  assign n11962 = n11961 ^ n5887 ^ n3187 ;
  assign n11967 = n11966 ^ n11965 ^ n11962 ;
  assign n11973 = n6709 ^ n1264 ^ n761 ;
  assign n11974 = n11973 ^ n3838 ^ n600 ;
  assign n11968 = n2907 ^ n2105 ^ 1'b0 ;
  assign n11969 = n11968 ^ n3805 ^ 1'b0 ;
  assign n11970 = n6562 | n11969 ;
  assign n11971 = n2672 & ~n11970 ;
  assign n11972 = ( ~n3428 & n6411 ) | ( ~n3428 & n11971 ) | ( n6411 & n11971 ) ;
  assign n11975 = n11974 ^ n11972 ^ n7858 ;
  assign n11977 = ( n2679 & n5638 ) | ( n2679 & ~n9767 ) | ( n5638 & ~n9767 ) ;
  assign n11978 = n11977 ^ n7387 ^ n1476 ;
  assign n11979 = n11978 ^ n8178 ^ n6025 ;
  assign n11980 = ~n8112 & n11979 ;
  assign n11976 = x10 & n2988 ;
  assign n11981 = n11980 ^ n11976 ^ 1'b0 ;
  assign n11982 = n7975 ^ n7152 ^ 1'b0 ;
  assign n11983 = n8004 | n11982 ;
  assign n11984 = ( n4251 & n5372 ) | ( n4251 & n11983 ) | ( n5372 & n11983 ) ;
  assign n11985 = ( x53 & ~n4694 ) | ( x53 & n11984 ) | ( ~n4694 & n11984 ) ;
  assign n11986 = n11985 ^ n7958 ^ n2871 ;
  assign n11987 = n10516 ^ n3556 ^ n2901 ;
  assign n11988 = ( n366 & ~n1340 ) | ( n366 & n9796 ) | ( ~n1340 & n9796 ) ;
  assign n11989 = n5175 ^ n862 ^ n366 ;
  assign n11990 = n11989 ^ n4659 ^ 1'b0 ;
  assign n11991 = n11988 & n11990 ;
  assign n11992 = ( ~n3921 & n11987 ) | ( ~n3921 & n11991 ) | ( n11987 & n11991 ) ;
  assign n11993 = ( n1963 & n2537 ) | ( n1963 & n3981 ) | ( n2537 & n3981 ) ;
  assign n11994 = ( n5704 & ~n8440 ) | ( n5704 & n11993 ) | ( ~n8440 & n11993 ) ;
  assign n11995 = n7615 ^ n6299 ^ n2862 ;
  assign n11996 = ( n7025 & n7537 ) | ( n7025 & n11995 ) | ( n7537 & n11995 ) ;
  assign n11997 = n3141 & ~n11961 ;
  assign n11998 = n4043 & n11997 ;
  assign n11999 = ( n1129 & n2911 ) | ( n1129 & ~n11998 ) | ( n2911 & ~n11998 ) ;
  assign n12000 = ( n2366 & n7588 ) | ( n2366 & ~n9598 ) | ( n7588 & ~n9598 ) ;
  assign n12001 = n749 & n5625 ;
  assign n12002 = n12001 ^ n1629 ^ 1'b0 ;
  assign n12003 = n7989 ^ n5519 ^ n2696 ;
  assign n12004 = ( ~n8153 & n12002 ) | ( ~n8153 & n12003 ) | ( n12002 & n12003 ) ;
  assign n12005 = n1156 & n4662 ;
  assign n12006 = n1191 & n12005 ;
  assign n12007 = ~n12004 & n12006 ;
  assign n12008 = n8107 ^ n5228 ^ n569 ;
  assign n12009 = ( n2713 & ~n10706 ) | ( n2713 & n12008 ) | ( ~n10706 & n12008 ) ;
  assign n12010 = n11471 ^ n10348 ^ 1'b0 ;
  assign n12011 = ~n4541 & n12010 ;
  assign n12012 = ( n2014 & n7538 ) | ( n2014 & n7955 ) | ( n7538 & n7955 ) ;
  assign n12013 = ( n4624 & ~n8728 ) | ( n4624 & n9426 ) | ( ~n8728 & n9426 ) ;
  assign n12014 = ( n898 & n3328 ) | ( n898 & ~n12013 ) | ( n3328 & ~n12013 ) ;
  assign n12015 = ( n885 & n3122 ) | ( n885 & ~n12014 ) | ( n3122 & ~n12014 ) ;
  assign n12016 = ( ~n4485 & n12012 ) | ( ~n4485 & n12015 ) | ( n12012 & n12015 ) ;
  assign n12017 = n1731 ^ n1063 ^ n479 ;
  assign n12018 = n12017 ^ n4131 ^ n1698 ;
  assign n12019 = n12018 ^ n10173 ^ n9717 ;
  assign n12020 = n1608 & ~n10171 ;
  assign n12021 = n12020 ^ n5127 ^ n1270 ;
  assign n12022 = n12019 | n12021 ;
  assign n12024 = n3298 & n7504 ;
  assign n12025 = ~n3365 & n12024 ;
  assign n12023 = ( ~n4681 & n7302 ) | ( ~n4681 & n7317 ) | ( n7302 & n7317 ) ;
  assign n12026 = n12025 ^ n12023 ^ x92 ;
  assign n12027 = n12026 ^ n5523 ^ n4036 ;
  assign n12028 = n6803 & n12027 ;
  assign n12029 = n12022 & n12028 ;
  assign n12030 = ( n281 & n4040 ) | ( n281 & n4408 ) | ( n4040 & n4408 ) ;
  assign n12031 = ~n2000 & n12030 ;
  assign n12032 = n12031 ^ n8731 ^ n733 ;
  assign n12033 = ( n3216 & n6538 ) | ( n3216 & ~n9003 ) | ( n6538 & ~n9003 ) ;
  assign n12034 = n3223 ^ n2623 ^ n805 ;
  assign n12035 = ( n1254 & n6134 ) | ( n1254 & ~n12034 ) | ( n6134 & ~n12034 ) ;
  assign n12036 = n4108 & ~n5632 ;
  assign n12037 = n12036 ^ n5861 ^ 1'b0 ;
  assign n12038 = n9402 & ~n12037 ;
  assign n12039 = n1071 | n5889 ;
  assign n12040 = n12039 ^ n1454 ^ 1'b0 ;
  assign n12041 = n12038 & ~n12040 ;
  assign n12042 = n3989 ^ n3255 ^ n645 ;
  assign n12043 = n12042 ^ n11598 ^ 1'b0 ;
  assign n12044 = n3342 & n12043 ;
  assign n12045 = ( ~n3216 & n9431 ) | ( ~n3216 & n12044 ) | ( n9431 & n12044 ) ;
  assign n12046 = ( ~n5584 & n6531 ) | ( ~n5584 & n10153 ) | ( n6531 & n10153 ) ;
  assign n12047 = n12046 ^ n6153 ^ n3182 ;
  assign n12048 = ( n5661 & ~n9192 ) | ( n5661 & n12047 ) | ( ~n9192 & n12047 ) ;
  assign n12049 = n12048 ^ n462 ^ 1'b0 ;
  assign n12050 = ( n7618 & n12045 ) | ( n7618 & n12049 ) | ( n12045 & n12049 ) ;
  assign n12051 = n487 & ~n10817 ;
  assign n12052 = n11392 ^ n3311 ^ 1'b0 ;
  assign n12053 = n6179 & n12052 ;
  assign n12054 = n6990 ^ n6154 ^ n3937 ;
  assign n12055 = ( n2260 & n12053 ) | ( n2260 & ~n12054 ) | ( n12053 & ~n12054 ) ;
  assign n12056 = ( n854 & n3599 ) | ( n854 & ~n4327 ) | ( n3599 & ~n4327 ) ;
  assign n12057 = n5987 & ~n12056 ;
  assign n12058 = ~n12055 & n12057 ;
  assign n12059 = n8908 ^ n744 ^ n399 ;
  assign n12060 = n12059 ^ n6002 ^ 1'b0 ;
  assign n12061 = n10783 & ~n12060 ;
  assign n12071 = n3605 ^ n321 ^ 1'b0 ;
  assign n12072 = n6302 ^ n5377 ^ 1'b0 ;
  assign n12073 = n8233 & ~n12072 ;
  assign n12074 = ( n5804 & n12071 ) | ( n5804 & n12073 ) | ( n12071 & n12073 ) ;
  assign n12070 = ( n868 & n1986 ) | ( n868 & n11429 ) | ( n1986 & n11429 ) ;
  assign n12062 = ( n2169 & n2812 ) | ( n2169 & n4965 ) | ( n2812 & n4965 ) ;
  assign n12063 = n12062 ^ n5994 ^ n3618 ;
  assign n12064 = n7669 ^ n5927 ^ n5052 ;
  assign n12065 = n12063 | n12064 ;
  assign n12066 = n2809 | n12065 ;
  assign n12067 = ~n1678 & n11436 ;
  assign n12068 = n12067 ^ n4943 ^ 1'b0 ;
  assign n12069 = ( n11362 & n12066 ) | ( n11362 & n12068 ) | ( n12066 & n12068 ) ;
  assign n12075 = n12074 ^ n12070 ^ n12069 ;
  assign n12076 = n7149 ^ n363 ^ 1'b0 ;
  assign n12077 = n6988 | n12076 ;
  assign n12078 = n12077 ^ n9974 ^ n6000 ;
  assign n12079 = ( n3484 & ~n8318 ) | ( n3484 & n12078 ) | ( ~n8318 & n12078 ) ;
  assign n12080 = ( n5185 & ~n6993 ) | ( n5185 & n12079 ) | ( ~n6993 & n12079 ) ;
  assign n12081 = n12080 ^ x116 ^ 1'b0 ;
  assign n12087 = ( ~x45 & n4247 ) | ( ~x45 & n8713 ) | ( n4247 & n8713 ) ;
  assign n12082 = n5310 & ~n6235 ;
  assign n12083 = n1645 & n12082 ;
  assign n12084 = n4779 & n12083 ;
  assign n12085 = n12084 ^ n9125 ^ n5445 ;
  assign n12086 = n4033 & ~n12085 ;
  assign n12088 = n12087 ^ n12086 ^ 1'b0 ;
  assign n12089 = ( n4528 & n5848 ) | ( n4528 & n9353 ) | ( n5848 & n9353 ) ;
  assign n12090 = ( n270 & n643 ) | ( n270 & n3060 ) | ( n643 & n3060 ) ;
  assign n12091 = n8590 | n12090 ;
  assign n12092 = n8973 & ~n12091 ;
  assign n12093 = ( n4122 & ~n5539 ) | ( n4122 & n12092 ) | ( ~n5539 & n12092 ) ;
  assign n12094 = n12089 & ~n12093 ;
  assign n12095 = ( n2917 & n8542 ) | ( n2917 & n12094 ) | ( n8542 & n12094 ) ;
  assign n12097 = n9297 ^ n7735 ^ n6035 ;
  assign n12096 = n5957 ^ n2511 ^ 1'b0 ;
  assign n12098 = n12097 ^ n12096 ^ n8679 ;
  assign n12101 = n1923 & ~n8317 ;
  assign n12099 = ~n4842 & n5276 ;
  assign n12100 = n12099 ^ n7316 ^ n4756 ;
  assign n12102 = n12101 ^ n12100 ^ 1'b0 ;
  assign n12104 = ( n842 & ~n2324 ) | ( n842 & n10134 ) | ( ~n2324 & n10134 ) ;
  assign n12105 = n12104 ^ n6571 ^ n1655 ;
  assign n12103 = n10447 ^ n10045 ^ x146 ;
  assign n12106 = n12105 ^ n12103 ^ n8808 ;
  assign n12107 = n4687 ^ n1752 ^ x157 ;
  assign n12108 = n8934 ^ n7444 ^ n2729 ;
  assign n12109 = n4942 & n12108 ;
  assign n12110 = n9382 | n12109 ;
  assign n12111 = n8455 & ~n12110 ;
  assign n12112 = n11237 & ~n12111 ;
  assign n12113 = ( n11311 & n12107 ) | ( n11311 & ~n12112 ) | ( n12107 & ~n12112 ) ;
  assign n12114 = n6415 ^ n531 ^ 1'b0 ;
  assign n12115 = x20 & n12114 ;
  assign n12116 = n2693 | n12115 ;
  assign n12117 = ( n4428 & ~n5465 ) | ( n4428 & n7251 ) | ( ~n5465 & n7251 ) ;
  assign n12118 = n3907 ^ n2201 ^ 1'b0 ;
  assign n12119 = ( ~n3773 & n12117 ) | ( ~n3773 & n12118 ) | ( n12117 & n12118 ) ;
  assign n12120 = n10786 ^ n6134 ^ 1'b0 ;
  assign n12121 = n6531 | n12120 ;
  assign n12122 = n1522 | n12121 ;
  assign n12123 = ~n2523 & n7811 ;
  assign n12124 = n12123 ^ x9 ^ 1'b0 ;
  assign n12125 = n4581 ^ n2746 ^ n724 ;
  assign n12126 = ( n3033 & ~n7129 ) | ( n3033 & n12125 ) | ( ~n7129 & n12125 ) ;
  assign n12127 = ( ~n4917 & n12124 ) | ( ~n4917 & n12126 ) | ( n12124 & n12126 ) ;
  assign n12133 = n11457 ^ n1191 ^ n720 ;
  assign n12130 = n2431 ^ n1182 ^ 1'b0 ;
  assign n12131 = x65 & n12130 ;
  assign n12128 = ~n1030 & n8960 ;
  assign n12129 = n12128 ^ n2342 ^ 1'b0 ;
  assign n12132 = n12131 ^ n12129 ^ n5614 ;
  assign n12134 = n12133 ^ n12132 ^ n4545 ;
  assign n12141 = n7796 ^ n2795 ^ n2219 ;
  assign n12137 = n5371 ^ x86 ^ 1'b0 ;
  assign n12138 = ~n1990 & n12137 ;
  assign n12139 = ( ~n3681 & n5181 ) | ( ~n3681 & n5441 ) | ( n5181 & n5441 ) ;
  assign n12140 = n12138 & n12139 ;
  assign n12142 = n12141 ^ n12140 ^ 1'b0 ;
  assign n12135 = ( n1809 & ~n7231 ) | ( n1809 & n10865 ) | ( ~n7231 & n10865 ) ;
  assign n12136 = n12135 ^ n7260 ^ n3379 ;
  assign n12143 = n12142 ^ n12136 ^ n1477 ;
  assign n12144 = ( n3727 & n6397 ) | ( n3727 & n12143 ) | ( n6397 & n12143 ) ;
  assign n12145 = n7540 ^ n1007 ^ 1'b0 ;
  assign n12146 = n2267 & ~n12145 ;
  assign n12147 = ( n2524 & n6766 ) | ( n2524 & ~n12146 ) | ( n6766 & ~n12146 ) ;
  assign n12151 = n5893 ^ n2046 ^ n1140 ;
  assign n12152 = n12151 ^ n4035 ^ n3552 ;
  assign n12148 = ( n6092 & n8219 ) | ( n6092 & ~n8687 ) | ( n8219 & ~n8687 ) ;
  assign n12149 = n12148 ^ n5271 ^ n3448 ;
  assign n12150 = n12149 ^ n11237 ^ n536 ;
  assign n12153 = n12152 ^ n12150 ^ n1445 ;
  assign n12154 = n12153 ^ n2889 ^ 1'b0 ;
  assign n12155 = ~x200 & n12154 ;
  assign n12158 = n8933 ^ n5217 ^ n3523 ;
  assign n12156 = n11490 ^ n2667 ^ 1'b0 ;
  assign n12157 = n1295 & n12156 ;
  assign n12159 = n12158 ^ n12157 ^ n4294 ;
  assign n12160 = n12159 ^ n8158 ^ 1'b0 ;
  assign n12161 = ( n1179 & ~n5459 ) | ( n1179 & n6321 ) | ( ~n5459 & n6321 ) ;
  assign n12162 = n9893 ^ n8629 ^ n3257 ;
  assign n12163 = ( n2729 & ~n9938 ) | ( n2729 & n12162 ) | ( ~n9938 & n12162 ) ;
  assign n12164 = ( n532 & n1576 ) | ( n532 & ~n12163 ) | ( n1576 & ~n12163 ) ;
  assign n12165 = n5693 ^ n2080 ^ 1'b0 ;
  assign n12166 = n3386 | n12165 ;
  assign n12167 = n6056 & ~n12062 ;
  assign n12168 = n12166 & n12167 ;
  assign n12169 = ~n8887 & n12168 ;
  assign n12170 = ~n1364 & n1908 ;
  assign n12171 = ( n2853 & ~n9694 ) | ( n2853 & n10452 ) | ( ~n9694 & n10452 ) ;
  assign n12172 = ( n7258 & n12170 ) | ( n7258 & n12171 ) | ( n12170 & n12171 ) ;
  assign n12174 = n7940 ^ n7755 ^ n1873 ;
  assign n12173 = n7715 ^ n5464 ^ 1'b0 ;
  assign n12175 = n12174 ^ n12173 ^ n10998 ;
  assign n12176 = n264 & ~n5655 ;
  assign n12177 = ~n3608 & n12176 ;
  assign n12178 = n11918 ^ n3633 ^ 1'b0 ;
  assign n12179 = n7192 ^ n4887 ^ x24 ;
  assign n12180 = n12179 ^ n9829 ^ 1'b0 ;
  assign n12181 = ( n10570 & n12178 ) | ( n10570 & n12180 ) | ( n12178 & n12180 ) ;
  assign n12187 = n362 & ~n5370 ;
  assign n12188 = n6898 & n12187 ;
  assign n12182 = n556 & ~n3016 ;
  assign n12183 = n4887 & n12182 ;
  assign n12184 = ( n948 & ~n3180 ) | ( n948 & n12183 ) | ( ~n3180 & n12183 ) ;
  assign n12185 = n12184 ^ n5734 ^ n4702 ;
  assign n12186 = n12185 ^ n7591 ^ n2135 ;
  assign n12189 = n12188 ^ n12186 ^ n1033 ;
  assign n12190 = n11433 ^ n2073 ^ 1'b0 ;
  assign n12191 = n12190 ^ n4712 ^ n2701 ;
  assign n12192 = n12191 ^ n2676 ^ 1'b0 ;
  assign n12193 = n11654 | n12192 ;
  assign n12194 = ( ~n6614 & n12174 ) | ( ~n6614 & n12193 ) | ( n12174 & n12193 ) ;
  assign n12196 = n2600 ^ n2581 ^ n828 ;
  assign n12195 = n4089 & ~n9677 ;
  assign n12197 = n12196 ^ n12195 ^ 1'b0 ;
  assign n12205 = x231 & n1937 ;
  assign n12202 = n11780 ^ n7955 ^ n3318 ;
  assign n12203 = n12202 ^ n6448 ^ n1605 ;
  assign n12198 = n2873 ^ x144 ^ 1'b0 ;
  assign n12199 = n6938 & n12198 ;
  assign n12200 = ( n2947 & n8736 ) | ( n2947 & n12199 ) | ( n8736 & n12199 ) ;
  assign n12201 = n12200 ^ n3534 ^ 1'b0 ;
  assign n12204 = n12203 ^ n12201 ^ n5077 ;
  assign n12206 = n12205 ^ n12204 ^ n2432 ;
  assign n12207 = n11849 ^ n9231 ^ n1316 ;
  assign n12208 = ( n4686 & n10745 ) | ( n4686 & n12207 ) | ( n10745 & n12207 ) ;
  assign n12209 = n12208 ^ n5918 ^ n2213 ;
  assign n12210 = ( ~n485 & n3395 ) | ( ~n485 & n5317 ) | ( n3395 & n5317 ) ;
  assign n12214 = ( n3726 & ~n8404 ) | ( n3726 & n8438 ) | ( ~n8404 & n8438 ) ;
  assign n12211 = n3705 ^ n711 ^ 1'b0 ;
  assign n12212 = n9308 & n12211 ;
  assign n12213 = n12212 ^ n9152 ^ n4184 ;
  assign n12215 = n12214 ^ n12213 ^ n3076 ;
  assign n12216 = n547 & ~n3069 ;
  assign n12217 = ~n12215 & n12216 ;
  assign n12218 = n2856 ^ n2507 ^ n330 ;
  assign n12219 = n5218 & n12218 ;
  assign n12220 = ( n5801 & n7816 ) | ( n5801 & n12219 ) | ( n7816 & n12219 ) ;
  assign n12221 = ( n2421 & n3380 ) | ( n2421 & ~n6390 ) | ( n3380 & ~n6390 ) ;
  assign n12222 = x208 & n2094 ;
  assign n12223 = ~n5782 & n12222 ;
  assign n12224 = n12223 ^ n10266 ^ n8050 ;
  assign n12225 = ( n5463 & n12221 ) | ( n5463 & n12224 ) | ( n12221 & n12224 ) ;
  assign n12226 = ( n4026 & n9609 ) | ( n4026 & ~n12111 ) | ( n9609 & ~n12111 ) ;
  assign n12227 = n2977 | n10354 ;
  assign n12228 = n8036 ^ n5090 ^ n3681 ;
  assign n12229 = n12228 ^ n11391 ^ n631 ;
  assign n12230 = ( x112 & n345 ) | ( x112 & ~n4355 ) | ( n345 & ~n4355 ) ;
  assign n12231 = ( n884 & n11473 ) | ( n884 & ~n12230 ) | ( n11473 & ~n12230 ) ;
  assign n12241 = ( n1212 & ~n5156 ) | ( n1212 & n7171 ) | ( ~n5156 & n7171 ) ;
  assign n12237 = ~n2472 & n4244 ;
  assign n12238 = ~n2059 & n12237 ;
  assign n12239 = n12238 ^ n7159 ^ n1960 ;
  assign n12232 = n7047 ^ n1829 ^ x245 ;
  assign n12233 = n6984 ^ n4556 ^ n2906 ;
  assign n12234 = n12233 ^ n3940 ^ 1'b0 ;
  assign n12235 = n3127 & ~n12234 ;
  assign n12236 = ~n12232 & n12235 ;
  assign n12240 = n12239 ^ n12236 ^ n4315 ;
  assign n12242 = n12241 ^ n12240 ^ n7431 ;
  assign n12258 = n866 ^ n804 ^ 1'b0 ;
  assign n12259 = n1519 & ~n12258 ;
  assign n12260 = n2521 & ~n12259 ;
  assign n12261 = n12260 ^ n2518 ^ n1623 ;
  assign n12255 = n974 | n7793 ;
  assign n12256 = n12255 ^ n912 ^ 1'b0 ;
  assign n12253 = n8438 ^ n7994 ^ n6240 ;
  assign n12254 = n12253 ^ n9767 ^ n500 ;
  assign n12250 = n506 | n6636 ;
  assign n12251 = n11798 ^ n10439 ^ n10385 ;
  assign n12252 = ( ~n5119 & n12250 ) | ( ~n5119 & n12251 ) | ( n12250 & n12251 ) ;
  assign n12257 = n12256 ^ n12254 ^ n12252 ;
  assign n12262 = n12261 ^ n12257 ^ n1747 ;
  assign n12244 = n366 & ~n9429 ;
  assign n12245 = n7648 ^ n3145 ^ 1'b0 ;
  assign n12246 = n4503 ^ n1557 ^ n428 ;
  assign n12247 = ( n5035 & ~n7811 ) | ( n5035 & n12246 ) | ( ~n7811 & n12246 ) ;
  assign n12248 = ( n9366 & ~n12245 ) | ( n9366 & n12247 ) | ( ~n12245 & n12247 ) ;
  assign n12249 = ( n415 & n12244 ) | ( n415 & ~n12248 ) | ( n12244 & ~n12248 ) ;
  assign n12263 = n12262 ^ n12249 ^ n1942 ;
  assign n12243 = n1965 & ~n2496 ;
  assign n12264 = n12263 ^ n12243 ^ n1343 ;
  assign n12265 = n1782 & n4336 ;
  assign n12266 = ( n354 & ~n2739 ) | ( n354 & n4408 ) | ( ~n2739 & n4408 ) ;
  assign n12267 = n7120 ^ n6082 ^ n4156 ;
  assign n12268 = n12267 ^ n10654 ^ 1'b0 ;
  assign n12269 = n6798 & ~n12268 ;
  assign n12270 = ( n12265 & n12266 ) | ( n12265 & ~n12269 ) | ( n12266 & ~n12269 ) ;
  assign n12273 = ( n697 & n2474 ) | ( n697 & n2636 ) | ( n2474 & n2636 ) ;
  assign n12274 = n12273 ^ n8835 ^ n1971 ;
  assign n12271 = n7554 | n8229 ;
  assign n12272 = n12271 ^ n11281 ^ n4629 ;
  assign n12275 = n12274 ^ n12272 ^ n11018 ;
  assign n12276 = n7515 | n8888 ;
  assign n12277 = n12276 ^ n3200 ^ 1'b0 ;
  assign n12278 = n1538 & n2196 ;
  assign n12279 = ( n7465 & n9090 ) | ( n7465 & n12278 ) | ( n9090 & n12278 ) ;
  assign n12282 = n6248 ^ n4301 ^ 1'b0 ;
  assign n12283 = ( ~n1595 & n4424 ) | ( ~n1595 & n12282 ) | ( n4424 & n12282 ) ;
  assign n12280 = x125 & n5529 ;
  assign n12281 = ~n457 & n12280 ;
  assign n12284 = n12283 ^ n12281 ^ n10395 ;
  assign n12285 = n12284 ^ n9269 ^ n9060 ;
  assign n12286 = n1085 ^ n335 ^ x227 ;
  assign n12287 = ( n4916 & n6811 ) | ( n4916 & n12286 ) | ( n6811 & n12286 ) ;
  assign n12288 = n12287 ^ n6324 ^ n1224 ;
  assign n12289 = n12288 ^ n1106 ^ 1'b0 ;
  assign n12293 = ~n3371 & n7544 ;
  assign n12294 = n12293 ^ n5681 ^ 1'b0 ;
  assign n12291 = n4752 ^ n4091 ^ n2484 ;
  assign n12290 = n11911 ^ n3132 ^ 1'b0 ;
  assign n12292 = n12291 ^ n12290 ^ n4710 ;
  assign n12295 = n12294 ^ n12292 ^ n8604 ;
  assign n12296 = n1760 ^ n1116 ^ x90 ;
  assign n12297 = ( n1288 & n12295 ) | ( n1288 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12298 = n11349 ^ n9827 ^ n4149 ;
  assign n12299 = n3259 ^ n2436 ^ n599 ;
  assign n12300 = n12299 ^ n4701 ^ n2361 ;
  assign n12301 = n3854 & n6752 ;
  assign n12302 = n12301 ^ n5429 ^ 1'b0 ;
  assign n12303 = ( n3560 & n12300 ) | ( n3560 & n12302 ) | ( n12300 & n12302 ) ;
  assign n12304 = n12303 ^ n11396 ^ n4719 ;
  assign n12315 = ( n7810 & ~n8674 ) | ( n7810 & n9951 ) | ( ~n8674 & n9951 ) ;
  assign n12310 = ~n1384 & n2101 ;
  assign n12311 = n2800 & n12310 ;
  assign n12312 = ( n1455 & ~n3360 ) | ( n1455 & n12311 ) | ( ~n3360 & n12311 ) ;
  assign n12313 = n12312 ^ n4023 ^ n971 ;
  assign n12314 = ( ~n552 & n4835 ) | ( ~n552 & n12313 ) | ( n4835 & n12313 ) ;
  assign n12305 = n5918 | n6587 ;
  assign n12306 = n6953 | n12305 ;
  assign n12307 = ( n4017 & n9345 ) | ( n4017 & ~n11025 ) | ( n9345 & ~n11025 ) ;
  assign n12308 = n4999 | n12307 ;
  assign n12309 = ( n10035 & n12306 ) | ( n10035 & ~n12308 ) | ( n12306 & ~n12308 ) ;
  assign n12316 = n12315 ^ n12314 ^ n12309 ;
  assign n12317 = ( ~n1760 & n3334 ) | ( ~n1760 & n10232 ) | ( n3334 & n10232 ) ;
  assign n12318 = ( n1365 & n2232 ) | ( n1365 & n12317 ) | ( n2232 & n12317 ) ;
  assign n12320 = ( ~n1202 & n6364 ) | ( ~n1202 & n7064 ) | ( n6364 & n7064 ) ;
  assign n12321 = ( n2942 & ~n3629 ) | ( n2942 & n12320 ) | ( ~n3629 & n12320 ) ;
  assign n12322 = ( ~n3630 & n11106 ) | ( ~n3630 & n12321 ) | ( n11106 & n12321 ) ;
  assign n12319 = ( ~n362 & n1774 ) | ( ~n362 & n2680 ) | ( n1774 & n2680 ) ;
  assign n12323 = n12322 ^ n12319 ^ 1'b0 ;
  assign n12324 = ~n7114 & n12323 ;
  assign n12325 = n12324 ^ n12174 ^ n2372 ;
  assign n12326 = n4637 & ~n12325 ;
  assign n12327 = ~n9769 & n12326 ;
  assign n12328 = n6701 ^ n3354 ^ n2897 ;
  assign n12329 = n4608 ^ n2135 ^ 1'b0 ;
  assign n12330 = n3496 | n12329 ;
  assign n12331 = ( ~n5840 & n11173 ) | ( ~n5840 & n12069 ) | ( n11173 & n12069 ) ;
  assign n12340 = n10914 ^ n2587 ^ 1'b0 ;
  assign n12338 = ( n884 & n1666 ) | ( n884 & ~n4626 ) | ( n1666 & ~n4626 ) ;
  assign n12339 = ~n998 & n12338 ;
  assign n12341 = n12340 ^ n12339 ^ 1'b0 ;
  assign n12332 = ( n6045 & ~n6416 ) | ( n6045 & n9401 ) | ( ~n6416 & n9401 ) ;
  assign n12334 = ~n4936 & n5895 ;
  assign n12333 = n5636 ^ n4894 ^ n3191 ;
  assign n12335 = n12334 ^ n12333 ^ n8792 ;
  assign n12336 = ( n2315 & n8964 ) | ( n2315 & n12335 ) | ( n8964 & n12335 ) ;
  assign n12337 = ( n1610 & n12332 ) | ( n1610 & ~n12336 ) | ( n12332 & ~n12336 ) ;
  assign n12342 = n12341 ^ n12337 ^ n538 ;
  assign n12343 = n12146 ^ n8818 ^ n4321 ;
  assign n12348 = n8554 ^ n2602 ^ 1'b0 ;
  assign n12349 = n11722 | n12348 ;
  assign n12350 = n3412 & ~n5353 ;
  assign n12351 = ~n6312 & n12350 ;
  assign n12352 = n12349 & n12351 ;
  assign n12345 = n3727 ^ n2170 ^ n1807 ;
  assign n12344 = ( x224 & ~n2159 ) | ( x224 & n6368 ) | ( ~n2159 & n6368 ) ;
  assign n12346 = n12345 ^ n12344 ^ n6314 ;
  assign n12347 = n7067 & n12346 ;
  assign n12353 = n12352 ^ n12347 ^ 1'b0 ;
  assign n12354 = ( n7196 & n12343 ) | ( n7196 & n12353 ) | ( n12343 & n12353 ) ;
  assign n12358 = ( ~n4807 & n7876 ) | ( ~n4807 & n9485 ) | ( n7876 & n9485 ) ;
  assign n12355 = n3055 | n7843 ;
  assign n12356 = n1821 & ~n12355 ;
  assign n12357 = ( n3761 & ~n4406 ) | ( n3761 & n12356 ) | ( ~n4406 & n12356 ) ;
  assign n12359 = n12358 ^ n12357 ^ 1'b0 ;
  assign n12360 = x170 & n3670 ;
  assign n12361 = n11349 & n12360 ;
  assign n12362 = n2129 | n8640 ;
  assign n12363 = n12361 & ~n12362 ;
  assign n12364 = ~n7285 & n10035 ;
  assign n12365 = ~n662 & n12364 ;
  assign n12366 = ( n9877 & ~n12363 ) | ( n9877 & n12365 ) | ( ~n12363 & n12365 ) ;
  assign n12371 = n1968 ^ x20 ^ 1'b0 ;
  assign n12372 = n2229 & n12371 ;
  assign n12373 = n3800 ^ n464 ^ 1'b0 ;
  assign n12374 = n11880 & ~n12373 ;
  assign n12375 = ( n11524 & n12372 ) | ( n11524 & n12374 ) | ( n12372 & n12374 ) ;
  assign n12376 = n10799 ^ n2036 ^ n1611 ;
  assign n12377 = n12375 & ~n12376 ;
  assign n12367 = ( n4323 & n6950 ) | ( n4323 & n10401 ) | ( n6950 & n10401 ) ;
  assign n12368 = ( n901 & ~n4177 ) | ( n901 & n12367 ) | ( ~n4177 & n12367 ) ;
  assign n12369 = n2559 & ~n6771 ;
  assign n12370 = ~n12368 & n12369 ;
  assign n12378 = n12377 ^ n12370 ^ n11219 ;
  assign n12379 = ( n6786 & ~n8350 ) | ( n6786 & n10208 ) | ( ~n8350 & n10208 ) ;
  assign n12380 = ( n1162 & ~n2581 ) | ( n1162 & n12265 ) | ( ~n2581 & n12265 ) ;
  assign n12386 = n6620 ^ n4207 ^ n2439 ;
  assign n12383 = n472 & ~n10210 ;
  assign n12384 = n12383 ^ n1980 ^ 1'b0 ;
  assign n12385 = n12384 ^ n5026 ^ n595 ;
  assign n12381 = n6282 ^ n5058 ^ n998 ;
  assign n12382 = n12381 ^ n5562 ^ n1984 ;
  assign n12387 = n12386 ^ n12385 ^ n12382 ;
  assign n12389 = n4274 ^ n2450 ^ n2379 ;
  assign n12390 = n12389 ^ n3519 ^ 1'b0 ;
  assign n12388 = ( n1282 & n2790 ) | ( n1282 & n7484 ) | ( n2790 & n7484 ) ;
  assign n12391 = n12390 ^ n12388 ^ n9269 ;
  assign n12394 = n7260 ^ n6319 ^ n2437 ;
  assign n12395 = n12394 ^ n7114 ^ n4951 ;
  assign n12396 = n12395 ^ n6361 ^ 1'b0 ;
  assign n12397 = n12396 ^ n5649 ^ n2313 ;
  assign n12392 = n4567 ^ n4059 ^ 1'b0 ;
  assign n12393 = n4169 & n12392 ;
  assign n12398 = n12397 ^ n12393 ^ 1'b0 ;
  assign n12399 = n12391 & n12398 ;
  assign n12400 = ( n2391 & ~n12387 ) | ( n2391 & n12399 ) | ( ~n12387 & n12399 ) ;
  assign n12401 = ( n1895 & ~n9267 ) | ( n1895 & n9576 ) | ( ~n9267 & n9576 ) ;
  assign n12402 = ( ~n2231 & n6673 ) | ( ~n2231 & n12401 ) | ( n6673 & n12401 ) ;
  assign n12404 = n11812 ^ n2088 ^ x62 ;
  assign n12405 = n5066 & n12404 ;
  assign n12403 = ( n6034 & ~n6559 ) | ( n6034 & n11755 ) | ( ~n6559 & n11755 ) ;
  assign n12406 = n12405 ^ n12403 ^ n4421 ;
  assign n12407 = n2938 ^ n1372 ^ x4 ;
  assign n12408 = ( ~n1787 & n10031 ) | ( ~n1787 & n12291 ) | ( n10031 & n12291 ) ;
  assign n12409 = ~n12407 & n12408 ;
  assign n12410 = ~n10626 & n12409 ;
  assign n12411 = n8881 ^ n5247 ^ x220 ;
  assign n12412 = ( n952 & n5875 ) | ( n952 & n12411 ) | ( n5875 & n12411 ) ;
  assign n12413 = n6086 ^ n4784 ^ n675 ;
  assign n12414 = n6554 & n12413 ;
  assign n12415 = n12412 & n12414 ;
  assign n12416 = n11880 ^ n6277 ^ n5385 ;
  assign n12417 = ( n2977 & ~n4149 ) | ( n2977 & n9239 ) | ( ~n4149 & n9239 ) ;
  assign n12420 = n4020 ^ x23 ^ 1'b0 ;
  assign n12418 = n8482 ^ n6026 ^ 1'b0 ;
  assign n12419 = n7268 & ~n12418 ;
  assign n12421 = n12420 ^ n12419 ^ 1'b0 ;
  assign n12422 = ~n6807 & n12421 ;
  assign n12423 = ( n363 & n12417 ) | ( n363 & n12422 ) | ( n12417 & n12422 ) ;
  assign n12429 = ( n4648 & ~n5041 ) | ( n4648 & n5220 ) | ( ~n5041 & n5220 ) ;
  assign n12424 = n3324 ^ n1770 ^ 1'b0 ;
  assign n12425 = ( n841 & ~n4223 ) | ( n841 & n11164 ) | ( ~n4223 & n11164 ) ;
  assign n12426 = ( n3400 & n5556 ) | ( n3400 & ~n12425 ) | ( n5556 & ~n12425 ) ;
  assign n12427 = n12426 ^ n7605 ^ n4636 ;
  assign n12428 = ( ~n7897 & n12424 ) | ( ~n7897 & n12427 ) | ( n12424 & n12427 ) ;
  assign n12430 = n12429 ^ n12428 ^ 1'b0 ;
  assign n12431 = ( ~n623 & n810 ) | ( ~n623 & n11497 ) | ( n810 & n11497 ) ;
  assign n12432 = n12208 ^ n2941 ^ x1 ;
  assign n12433 = n2455 ^ n1405 ^ 1'b0 ;
  assign n12434 = n12432 | n12433 ;
  assign n12435 = n12431 & ~n12434 ;
  assign n12436 = n5331 & ~n6559 ;
  assign n12437 = n12436 ^ n766 ^ 1'b0 ;
  assign n12438 = n3329 ^ n2629 ^ 1'b0 ;
  assign n12439 = n12438 ^ n5290 ^ n1519 ;
  assign n12440 = n12437 & n12439 ;
  assign n12441 = n3942 ^ n3165 ^ n571 ;
  assign n12442 = ( n4392 & n9615 ) | ( n4392 & n12441 ) | ( n9615 & n12441 ) ;
  assign n12443 = ( ~n3792 & n4432 ) | ( ~n3792 & n6450 ) | ( n4432 & n6450 ) ;
  assign n12444 = n5020 & n12443 ;
  assign n12445 = n4704 | n12444 ;
  assign n12446 = n3084 | n12445 ;
  assign n12447 = n407 & ~n2167 ;
  assign n12448 = n12447 ^ n1854 ^ 1'b0 ;
  assign n12449 = ( n5382 & ~n9430 ) | ( n5382 & n12448 ) | ( ~n9430 & n12448 ) ;
  assign n12450 = n5815 & n12449 ;
  assign n12452 = n8603 ^ n1193 ^ 1'b0 ;
  assign n12453 = n12452 ^ n3128 ^ 1'b0 ;
  assign n12454 = n7442 & ~n12453 ;
  assign n12455 = ( n8938 & n10926 ) | ( n8938 & n12454 ) | ( n10926 & n12454 ) ;
  assign n12456 = x8 | n12455 ;
  assign n12451 = ( n3454 & n5822 ) | ( n3454 & n10950 ) | ( n5822 & n10950 ) ;
  assign n12457 = n12456 ^ n12451 ^ 1'b0 ;
  assign n12458 = n10711 ^ n8462 ^ n6023 ;
  assign n12459 = n12458 ^ n6672 ^ 1'b0 ;
  assign n12460 = ~n2607 & n3425 ;
  assign n12461 = n12460 ^ n1923 ^ 1'b0 ;
  assign n12470 = ( ~n1033 & n1536 ) | ( ~n1033 & n1943 ) | ( n1536 & n1943 ) ;
  assign n12471 = n12470 ^ n6329 ^ n803 ;
  assign n12472 = ( n6790 & ~n9927 ) | ( n6790 & n12471 ) | ( ~n9927 & n12471 ) ;
  assign n12466 = n5309 ^ n960 ^ 1'b0 ;
  assign n12467 = n12466 ^ n8462 ^ 1'b0 ;
  assign n12465 = n6988 ^ n5710 ^ n1863 ;
  assign n12462 = n5354 ^ n3846 ^ n1871 ;
  assign n12463 = n12462 ^ n6706 ^ n3311 ;
  assign n12464 = n12463 ^ n8027 ^ n7613 ;
  assign n12468 = n12467 ^ n12465 ^ n12464 ;
  assign n12469 = n9306 & ~n12468 ;
  assign n12473 = n12472 ^ n12469 ^ 1'b0 ;
  assign n12474 = n12473 ^ n1719 ^ x203 ;
  assign n12475 = ( n566 & n1767 ) | ( n566 & ~n12474 ) | ( n1767 & ~n12474 ) ;
  assign n12476 = ( ~n2486 & n4511 ) | ( ~n2486 & n7544 ) | ( n4511 & n7544 ) ;
  assign n12477 = ( ~n2939 & n9529 ) | ( ~n2939 & n12476 ) | ( n9529 & n12476 ) ;
  assign n12478 = n12477 ^ n2003 ^ x128 ;
  assign n12479 = ( n3718 & n5904 ) | ( n3718 & n12278 ) | ( n5904 & n12278 ) ;
  assign n12480 = ( n3998 & ~n10224 ) | ( n3998 & n12479 ) | ( ~n10224 & n12479 ) ;
  assign n12481 = n1685 & n6197 ;
  assign n12482 = n12481 ^ n441 ^ 1'b0 ;
  assign n12483 = n297 & n12482 ;
  assign n12484 = n12480 & n12483 ;
  assign n12493 = n2914 & ~n4958 ;
  assign n12485 = n7099 ^ n5358 ^ n4161 ;
  assign n12486 = ~n2205 & n12485 ;
  assign n12487 = n12486 ^ n3792 ^ 1'b0 ;
  assign n12488 = n12487 ^ n12184 ^ n4048 ;
  assign n12489 = ( n2768 & ~n7156 ) | ( n2768 & n10809 ) | ( ~n7156 & n10809 ) ;
  assign n12490 = n9896 ^ n1499 ^ 1'b0 ;
  assign n12491 = ( n8246 & n12489 ) | ( n8246 & n12490 ) | ( n12489 & n12490 ) ;
  assign n12492 = ( n2936 & n12488 ) | ( n2936 & n12491 ) | ( n12488 & n12491 ) ;
  assign n12494 = n12493 ^ n12492 ^ n9678 ;
  assign n12495 = n10222 ^ n6477 ^ 1'b0 ;
  assign n12496 = n3076 & n12495 ;
  assign n12497 = n12496 ^ n9604 ^ n4941 ;
  assign n12498 = n3526 | n11292 ;
  assign n12499 = n7150 & ~n12109 ;
  assign n12500 = ~n6122 & n12499 ;
  assign n12501 = n11420 ^ n6433 ^ n5336 ;
  assign n12502 = ( n5878 & ~n12500 ) | ( n5878 & n12501 ) | ( ~n12500 & n12501 ) ;
  assign n12503 = ( n3521 & n4730 ) | ( n3521 & ~n12502 ) | ( n4730 & ~n12502 ) ;
  assign n12504 = n7237 ^ n2698 ^ 1'b0 ;
  assign n12505 = ~n12503 & n12504 ;
  assign n12506 = n11231 ^ n11044 ^ x94 ;
  assign n12507 = n12506 ^ n4674 ^ n1156 ;
  assign n12508 = n12507 ^ n6749 ^ n3530 ;
  assign n12509 = n12508 ^ n3960 ^ 1'b0 ;
  assign n12510 = n10079 & n12509 ;
  assign n12511 = n11722 ^ n3258 ^ n3069 ;
  assign n12512 = ( n284 & ~n2939 ) | ( n284 & n12511 ) | ( ~n2939 & n12511 ) ;
  assign n12513 = n980 ^ x160 ^ 1'b0 ;
  assign n12514 = ~n1654 & n12513 ;
  assign n12515 = n3822 ^ n3180 ^ n1675 ;
  assign n12516 = n12515 ^ n10845 ^ n5813 ;
  assign n12517 = ( n7883 & n12514 ) | ( n7883 & n12516 ) | ( n12514 & n12516 ) ;
  assign n12518 = n5060 | n9378 ;
  assign n12520 = n11714 ^ n6875 ^ n1757 ;
  assign n12521 = n12520 ^ n9717 ^ n3681 ;
  assign n12519 = n11902 ^ n11747 ^ n4988 ;
  assign n12522 = n12521 ^ n12519 ^ n2037 ;
  assign n12523 = n11678 ^ n4175 ^ n1528 ;
  assign n12524 = n12523 ^ n9358 ^ n614 ;
  assign n12525 = n3694 ^ n2059 ^ n1582 ;
  assign n12526 = ( ~n577 & n7020 ) | ( ~n577 & n12525 ) | ( n7020 & n12525 ) ;
  assign n12527 = n12526 ^ n6530 ^ 1'b0 ;
  assign n12528 = n4560 & n6171 ;
  assign n12529 = n7213 ^ n4921 ^ x242 ;
  assign n12530 = ~n7646 & n7796 ;
  assign n12531 = ~n12529 & n12530 ;
  assign n12532 = n12531 ^ n8190 ^ n744 ;
  assign n12537 = ( ~n299 & n5035 ) | ( ~n299 & n9424 ) | ( n5035 & n9424 ) ;
  assign n12538 = n12537 ^ n5459 ^ n2383 ;
  assign n12533 = ( n2966 & n4134 ) | ( n2966 & ~n8055 ) | ( n4134 & ~n8055 ) ;
  assign n12534 = ( ~n2177 & n4654 ) | ( ~n2177 & n12533 ) | ( n4654 & n12533 ) ;
  assign n12535 = n12534 ^ n3376 ^ 1'b0 ;
  assign n12536 = n857 & ~n12535 ;
  assign n12539 = n12538 ^ n12536 ^ n503 ;
  assign n12540 = ( n1245 & ~n12532 ) | ( n1245 & n12539 ) | ( ~n12532 & n12539 ) ;
  assign n12544 = n2845 ^ n1714 ^ n505 ;
  assign n12545 = n9843 ^ n3807 ^ n742 ;
  assign n12546 = ( ~n662 & n2596 ) | ( ~n662 & n12545 ) | ( n2596 & n12545 ) ;
  assign n12547 = ( ~n4484 & n12544 ) | ( ~n4484 & n12546 ) | ( n12544 & n12546 ) ;
  assign n12541 = n6131 ^ n2635 ^ n1614 ;
  assign n12542 = n12541 ^ n943 ^ x38 ;
  assign n12543 = ( n517 & n8771 ) | ( n517 & ~n12542 ) | ( n8771 & ~n12542 ) ;
  assign n12548 = n12547 ^ n12543 ^ n7479 ;
  assign n12549 = n4101 ^ n2430 ^ 1'b0 ;
  assign n12550 = ~n2375 & n12549 ;
  assign n12551 = ~n1491 & n12550 ;
  assign n12552 = n12551 ^ n11364 ^ 1'b0 ;
  assign n12553 = n12462 & ~n12552 ;
  assign n12559 = n1864 & ~n3547 ;
  assign n12560 = n3546 & n12559 ;
  assign n12561 = n12560 ^ n7455 ^ 1'b0 ;
  assign n12554 = n4299 | n12284 ;
  assign n12555 = n12554 ^ n9198 ^ 1'b0 ;
  assign n12556 = ( ~n380 & n600 ) | ( ~n380 & n2831 ) | ( n600 & n2831 ) ;
  assign n12557 = n12556 ^ n1564 ^ 1'b0 ;
  assign n12558 = n12555 & n12557 ;
  assign n12562 = n12561 ^ n12558 ^ n1585 ;
  assign n12563 = n12562 ^ n11352 ^ n385 ;
  assign n12564 = ( n537 & ~n2145 ) | ( n537 & n2246 ) | ( ~n2145 & n2246 ) ;
  assign n12565 = ( n1862 & n5579 ) | ( n1862 & ~n12564 ) | ( n5579 & ~n12564 ) ;
  assign n12566 = ( ~n2932 & n12146 ) | ( ~n2932 & n12565 ) | ( n12146 & n12565 ) ;
  assign n12569 = ( ~n2169 & n6874 ) | ( ~n2169 & n7141 ) | ( n6874 & n7141 ) ;
  assign n12567 = n8484 & n12453 ;
  assign n12568 = n12567 ^ n11834 ^ 1'b0 ;
  assign n12570 = n12569 ^ n12568 ^ n11331 ;
  assign n12571 = n12570 ^ n3715 ^ 1'b0 ;
  assign n12572 = n3222 & ~n12571 ;
  assign n12573 = ( n7370 & n7845 ) | ( n7370 & ~n11672 ) | ( n7845 & ~n11672 ) ;
  assign n12574 = n9809 & n12573 ;
  assign n12575 = ~n12572 & n12574 ;
  assign n12576 = ~n5676 & n7596 ;
  assign n12577 = n12576 ^ n3487 ^ 1'b0 ;
  assign n12578 = ( n392 & n1030 ) | ( n392 & n1543 ) | ( n1030 & n1543 ) ;
  assign n12579 = n12577 & ~n12578 ;
  assign n12580 = ~n2183 & n12579 ;
  assign n12581 = n12580 ^ n10642 ^ n5967 ;
  assign n12582 = n10731 ^ n7632 ^ n2687 ;
  assign n12583 = n565 & ~n2751 ;
  assign n12584 = n12583 ^ n2942 ^ 1'b0 ;
  assign n12585 = ( n988 & n12582 ) | ( n988 & ~n12584 ) | ( n12582 & ~n12584 ) ;
  assign n12586 = ( n12575 & ~n12581 ) | ( n12575 & n12585 ) | ( ~n12581 & n12585 ) ;
  assign n12588 = n3469 ^ n2727 ^ 1'b0 ;
  assign n12587 = n3900 ^ n2838 ^ n1250 ;
  assign n12589 = n12588 ^ n12587 ^ n1827 ;
  assign n12600 = n3938 ^ n2710 ^ x188 ;
  assign n12598 = n5528 & n6773 ;
  assign n12596 = n8393 ^ n2581 ^ x48 ;
  assign n12594 = n1284 ^ n1161 ^ n385 ;
  assign n12593 = n3076 ^ n1319 ^ n294 ;
  assign n12591 = n5887 ^ n3813 ^ n1056 ;
  assign n12592 = ( n5095 & n6221 ) | ( n5095 & n12591 ) | ( n6221 & n12591 ) ;
  assign n12595 = n12594 ^ n12593 ^ n12592 ;
  assign n12597 = n12596 ^ n12595 ^ n5190 ;
  assign n12599 = n12598 ^ n12597 ^ n5601 ;
  assign n12590 = n9102 ^ n7211 ^ n2051 ;
  assign n12601 = n12600 ^ n12599 ^ n12590 ;
  assign n12617 = n6935 ^ n3777 ^ n858 ;
  assign n12618 = n7048 ^ n5698 ^ 1'b0 ;
  assign n12619 = ~n12617 & n12618 ;
  assign n12620 = n12619 ^ n3612 ^ n908 ;
  assign n12621 = ~n382 & n12620 ;
  assign n12622 = n12621 ^ n3833 ^ 1'b0 ;
  assign n12612 = n2931 & n7159 ;
  assign n12613 = n6787 ^ n3318 ^ 1'b0 ;
  assign n12614 = n2060 & ~n12613 ;
  assign n12615 = ( n2954 & n12612 ) | ( n2954 & n12614 ) | ( n12612 & n12614 ) ;
  assign n12616 = n12615 ^ n635 ^ n498 ;
  assign n12603 = n8359 & n9706 ;
  assign n12604 = n12603 ^ n7067 ^ 1'b0 ;
  assign n12605 = ~n8419 & n9527 ;
  assign n12606 = n1027 & ~n6210 ;
  assign n12607 = n12605 & n12606 ;
  assign n12608 = n7787 ^ n3479 ^ n2907 ;
  assign n12609 = n12608 ^ n5674 ^ n2002 ;
  assign n12610 = n12609 ^ n7102 ^ n832 ;
  assign n12611 = ( n12604 & ~n12607 ) | ( n12604 & n12610 ) | ( ~n12607 & n12610 ) ;
  assign n12623 = n12622 ^ n12616 ^ n12611 ;
  assign n12602 = n3516 | n10993 ;
  assign n12624 = n12623 ^ n12602 ^ 1'b0 ;
  assign n12625 = ( ~n12589 & n12601 ) | ( ~n12589 & n12624 ) | ( n12601 & n12624 ) ;
  assign n12629 = n6586 ^ n2978 ^ n2299 ;
  assign n12630 = ( n5756 & ~n9260 ) | ( n5756 & n12629 ) | ( ~n9260 & n12629 ) ;
  assign n12626 = x162 & ~n12546 ;
  assign n12627 = n3282 & n12626 ;
  assign n12628 = ( ~n7212 & n12267 ) | ( ~n7212 & n12627 ) | ( n12267 & n12627 ) ;
  assign n12631 = n12630 ^ n12628 ^ n10038 ;
  assign n12632 = n4114 ^ n1889 ^ n1840 ;
  assign n12633 = n11504 ^ n9612 ^ n5911 ;
  assign n12634 = ( n3608 & ~n11547 ) | ( n3608 & n11845 ) | ( ~n11547 & n11845 ) ;
  assign n12635 = n12634 ^ n4915 ^ n3414 ;
  assign n12636 = ( ~n855 & n8149 ) | ( ~n855 & n10383 ) | ( n8149 & n10383 ) ;
  assign n12637 = n12636 ^ n10174 ^ n337 ;
  assign n12638 = ( n1515 & n1666 ) | ( n1515 & n9272 ) | ( n1666 & n9272 ) ;
  assign n12639 = ( ~n846 & n1529 ) | ( ~n846 & n12191 ) | ( n1529 & n12191 ) ;
  assign n12640 = ( ~n11285 & n12638 ) | ( ~n11285 & n12639 ) | ( n12638 & n12639 ) ;
  assign n12641 = ( ~n3557 & n7830 ) | ( ~n3557 & n9760 ) | ( n7830 & n9760 ) ;
  assign n12642 = n12641 ^ n2911 ^ 1'b0 ;
  assign n12643 = ~n3049 & n12642 ;
  assign n12644 = ( n5058 & ~n12090 ) | ( n5058 & n12643 ) | ( ~n12090 & n12643 ) ;
  assign n12648 = x154 & ~n4521 ;
  assign n12647 = ( ~n827 & n3957 ) | ( ~n827 & n5023 ) | ( n3957 & n5023 ) ;
  assign n12649 = n12648 ^ n12647 ^ n656 ;
  assign n12645 = ( n4288 & ~n5290 ) | ( n4288 & n5777 ) | ( ~n5290 & n5777 ) ;
  assign n12646 = ( x23 & ~n12479 ) | ( x23 & n12645 ) | ( ~n12479 & n12645 ) ;
  assign n12650 = n12649 ^ n12646 ^ n4789 ;
  assign n12651 = ( x122 & n1048 ) | ( x122 & n4608 ) | ( n1048 & n4608 ) ;
  assign n12654 = n9050 ^ n2224 ^ n1937 ;
  assign n12652 = ( n365 & n8282 ) | ( n365 & ~n8907 ) | ( n8282 & ~n8907 ) ;
  assign n12653 = n12652 ^ n2894 ^ n2550 ;
  assign n12655 = n12654 ^ n12653 ^ 1'b0 ;
  assign n12656 = ( n5792 & n10590 ) | ( n5792 & n12655 ) | ( n10590 & n12655 ) ;
  assign n12657 = ( n1581 & ~n11829 ) | ( n1581 & n12656 ) | ( ~n11829 & n12656 ) ;
  assign n12658 = n12651 | n12657 ;
  assign n12659 = x57 & ~n10587 ;
  assign n12660 = n12659 ^ n7306 ^ 1'b0 ;
  assign n12663 = n2425 | n6541 ;
  assign n12662 = n4241 | n9222 ;
  assign n12664 = n12663 ^ n12662 ^ n9741 ;
  assign n12661 = ( ~x172 & x225 ) | ( ~x172 & n1092 ) | ( x225 & n1092 ) ;
  assign n12665 = n12664 ^ n12661 ^ n9140 ;
  assign n12666 = ( ~n2949 & n2994 ) | ( ~n2949 & n6237 ) | ( n2994 & n6237 ) ;
  assign n12667 = ( x51 & ~n3770 ) | ( x51 & n12666 ) | ( ~n3770 & n12666 ) ;
  assign n12668 = n12667 ^ n9409 ^ n4614 ;
  assign n12669 = ( n6743 & n9797 ) | ( n6743 & n10121 ) | ( n9797 & n10121 ) ;
  assign n12675 = ( n868 & n4836 ) | ( n868 & ~n5723 ) | ( n4836 & ~n5723 ) ;
  assign n12670 = n9720 ^ n2378 ^ x121 ;
  assign n12671 = ( x164 & n4849 ) | ( x164 & n12670 ) | ( n4849 & n12670 ) ;
  assign n12672 = n8813 & n12671 ;
  assign n12673 = n12672 ^ n4420 ^ 1'b0 ;
  assign n12674 = ( n1215 & n3345 ) | ( n1215 & n12673 ) | ( n3345 & n12673 ) ;
  assign n12676 = n12675 ^ n12674 ^ n7784 ;
  assign n12677 = ( ~n12668 & n12669 ) | ( ~n12668 & n12676 ) | ( n12669 & n12676 ) ;
  assign n12678 = ( n275 & n907 ) | ( n275 & n1590 ) | ( n907 & n1590 ) ;
  assign n12679 = n8504 & n10514 ;
  assign n12680 = ( ~n2985 & n3336 ) | ( ~n2985 & n5788 ) | ( n3336 & n5788 ) ;
  assign n12681 = n478 & n3910 ;
  assign n12682 = n12681 ^ n10098 ^ 1'b0 ;
  assign n12683 = ( n9920 & n12680 ) | ( n9920 & ~n12682 ) | ( n12680 & ~n12682 ) ;
  assign n12684 = ( n12678 & ~n12679 ) | ( n12678 & n12683 ) | ( ~n12679 & n12683 ) ;
  assign n12685 = n5670 ^ n3253 ^ n1278 ;
  assign n12686 = ( n969 & n8204 ) | ( n969 & n8903 ) | ( n8204 & n8903 ) ;
  assign n12687 = n6930 & ~n12686 ;
  assign n12688 = n12687 ^ n5799 ^ 1'b0 ;
  assign n12689 = ( n5539 & n12685 ) | ( n5539 & n12688 ) | ( n12685 & n12688 ) ;
  assign n12690 = ( ~n8912 & n10075 ) | ( ~n8912 & n12135 ) | ( n10075 & n12135 ) ;
  assign n12691 = n12690 ^ n1942 ^ x18 ;
  assign n12692 = n9761 ^ n7990 ^ n7669 ;
  assign n12693 = n12692 ^ n8647 ^ n3421 ;
  assign n12695 = n4454 ^ n4032 ^ n1505 ;
  assign n12694 = n2551 | n3657 ;
  assign n12696 = n12695 ^ n12694 ^ 1'b0 ;
  assign n12697 = ~n12693 & n12696 ;
  assign n12698 = ( n1204 & ~n5840 ) | ( n1204 & n7646 ) | ( ~n5840 & n7646 ) ;
  assign n12699 = ( ~n485 & n6259 ) | ( ~n485 & n10619 ) | ( n6259 & n10619 ) ;
  assign n12700 = ( ~n3579 & n7347 ) | ( ~n3579 & n7495 ) | ( n7347 & n7495 ) ;
  assign n12701 = n7333 ^ n4573 ^ n1678 ;
  assign n12702 = ~n5875 & n12634 ;
  assign n12703 = ~n12701 & n12702 ;
  assign n12704 = n12703 ^ n884 ^ 1'b0 ;
  assign n12705 = n12704 ^ n12408 ^ n2983 ;
  assign n12706 = n5739 ^ n498 ^ 1'b0 ;
  assign n12707 = n4099 & n12706 ;
  assign n12708 = n12707 ^ n7595 ^ n4060 ;
  assign n12709 = n12708 ^ n6718 ^ n3764 ;
  assign n12710 = n10272 ^ n10266 ^ n8976 ;
  assign n12711 = n11398 ^ n7568 ^ n2138 ;
  assign n12712 = n12711 ^ n12269 ^ n1840 ;
  assign n12727 = ( n1385 & n3824 ) | ( n1385 & ~n11695 ) | ( n3824 & ~n11695 ) ;
  assign n12723 = n5115 ^ n3613 ^ n1558 ;
  assign n12720 = ( n7849 & n10870 ) | ( n7849 & ~n11083 ) | ( n10870 & ~n11083 ) ;
  assign n12721 = n12720 ^ n9454 ^ n5086 ;
  assign n12719 = n1987 | n6262 ;
  assign n12722 = n12721 ^ n12719 ^ 1'b0 ;
  assign n12724 = n12723 ^ n12722 ^ n4440 ;
  assign n12716 = ( n417 & n8905 ) | ( n417 & n12218 ) | ( n8905 & n12218 ) ;
  assign n12713 = ( ~n379 & n3707 ) | ( ~n379 & n8848 ) | ( n3707 & n8848 ) ;
  assign n12714 = n12713 ^ n5845 ^ n1082 ;
  assign n12715 = ( n5756 & n8786 ) | ( n5756 & n12714 ) | ( n8786 & n12714 ) ;
  assign n12717 = n12716 ^ n12715 ^ n3949 ;
  assign n12718 = n12717 ^ n9104 ^ n335 ;
  assign n12725 = n12724 ^ n12718 ^ n6275 ;
  assign n12726 = n4464 & n12725 ;
  assign n12728 = n12727 ^ n12726 ^ 1'b0 ;
  assign n12729 = n12728 ^ n11746 ^ n8925 ;
  assign n12731 = n6720 ^ n6439 ^ n3327 ;
  assign n12730 = ( n505 & ~n7341 ) | ( n505 & n8043 ) | ( ~n7341 & n8043 ) ;
  assign n12732 = n12731 ^ n12730 ^ 1'b0 ;
  assign n12733 = n4414 & n12732 ;
  assign n12734 = n12733 ^ n11772 ^ n9993 ;
  assign n12735 = n2757 ^ n1281 ^ 1'b0 ;
  assign n12736 = n696 & n12735 ;
  assign n12737 = n9267 ^ n2677 ^ n420 ;
  assign n12738 = ( n1529 & ~n4798 ) | ( n1529 & n6530 ) | ( ~n4798 & n6530 ) ;
  assign n12739 = ( n7771 & ~n12737 ) | ( n7771 & n12738 ) | ( ~n12737 & n12738 ) ;
  assign n12740 = ( n7402 & n10473 ) | ( n7402 & n12739 ) | ( n10473 & n12739 ) ;
  assign n12741 = n8484 ^ n1183 ^ n323 ;
  assign n12742 = ( n7798 & n8133 ) | ( n7798 & n12741 ) | ( n8133 & n12741 ) ;
  assign n12743 = n12515 ^ n4406 ^ n1512 ;
  assign n12744 = n12743 ^ n2647 ^ 1'b0 ;
  assign n12745 = n12742 & ~n12744 ;
  assign n12746 = n8802 & n12745 ;
  assign n12747 = n12746 ^ n9695 ^ 1'b0 ;
  assign n12748 = ~n6045 & n10092 ;
  assign n12749 = n6530 ^ n3007 ^ n2455 ;
  assign n12750 = n2401 ^ n1834 ^ 1'b0 ;
  assign n12753 = n2853 | n3562 ;
  assign n12754 = n12753 ^ n2486 ^ 1'b0 ;
  assign n12751 = n6444 ^ n3942 ^ n1774 ;
  assign n12752 = n12751 ^ n10554 ^ n7085 ;
  assign n12755 = n12754 ^ n12752 ^ n4296 ;
  assign n12756 = ( n12749 & n12750 ) | ( n12749 & ~n12755 ) | ( n12750 & ~n12755 ) ;
  assign n12757 = n4884 ^ n4189 ^ n3478 ;
  assign n12758 = n11123 ^ n8692 ^ 1'b0 ;
  assign n12759 = n9341 ^ n642 ^ 1'b0 ;
  assign n12760 = ~n5689 & n12759 ;
  assign n12761 = ( n1724 & ~n3609 ) | ( n1724 & n12760 ) | ( ~n3609 & n12760 ) ;
  assign n12762 = ( n12757 & ~n12758 ) | ( n12757 & n12761 ) | ( ~n12758 & n12761 ) ;
  assign n12763 = n4072 & n12762 ;
  assign n12764 = n6804 ^ n5246 ^ 1'b0 ;
  assign n12765 = n9587 & ~n12764 ;
  assign n12766 = n11675 ^ n5368 ^ n4603 ;
  assign n12767 = ( n2750 & n5324 ) | ( n2750 & n6358 ) | ( n5324 & n6358 ) ;
  assign n12768 = ( n7627 & ~n12766 ) | ( n7627 & n12767 ) | ( ~n12766 & n12767 ) ;
  assign n12769 = n8318 & ~n10035 ;
  assign n12770 = n6948 ^ n4026 ^ 1'b0 ;
  assign n12771 = n1893 | n2093 ;
  assign n12772 = n12770 & ~n12771 ;
  assign n12773 = n1431 & ~n3000 ;
  assign n12774 = n12773 ^ n2515 ^ 1'b0 ;
  assign n12775 = n12774 ^ n8459 ^ n4039 ;
  assign n12776 = n8167 ^ n2655 ^ n2362 ;
  assign n12777 = n5319 | n12776 ;
  assign n12778 = n12777 ^ n5319 ^ 1'b0 ;
  assign n12779 = ( n5925 & ~n12775 ) | ( n5925 & n12778 ) | ( ~n12775 & n12778 ) ;
  assign n12780 = n7102 & n12779 ;
  assign n12781 = ( ~n12769 & n12772 ) | ( ~n12769 & n12780 ) | ( n12772 & n12780 ) ;
  assign n12784 = n473 | n3079 ;
  assign n12785 = n2212 & ~n12784 ;
  assign n12782 = n8571 ^ n5424 ^ n2717 ;
  assign n12783 = n3471 & n12782 ;
  assign n12786 = n12785 ^ n12783 ^ 1'b0 ;
  assign n12787 = n7410 ^ n3112 ^ n2292 ;
  assign n12788 = ( n711 & n846 ) | ( n711 & n2107 ) | ( n846 & n2107 ) ;
  assign n12789 = n12788 ^ n2343 ^ n936 ;
  assign n12790 = ( n3021 & n12787 ) | ( n3021 & n12789 ) | ( n12787 & n12789 ) ;
  assign n12791 = ( ~n1745 & n12786 ) | ( ~n1745 & n12790 ) | ( n12786 & n12790 ) ;
  assign n12792 = n10347 ^ n8427 ^ n968 ;
  assign n12793 = ( n2664 & n10546 ) | ( n2664 & ~n12792 ) | ( n10546 & ~n12792 ) ;
  assign n12794 = ( n7974 & ~n11615 ) | ( n7974 & n12793 ) | ( ~n11615 & n12793 ) ;
  assign n12795 = n10537 ^ n9499 ^ n702 ;
  assign n12796 = n12795 ^ n7532 ^ n3114 ;
  assign n12797 = ( n8324 & n10649 ) | ( n8324 & n11977 ) | ( n10649 & n11977 ) ;
  assign n12798 = ( x79 & n6108 ) | ( x79 & ~n6456 ) | ( n6108 & ~n6456 ) ;
  assign n12799 = n12798 ^ n12544 ^ n3051 ;
  assign n12800 = n3559 ^ n1427 ^ n567 ;
  assign n12801 = n12238 ^ n5127 ^ 1'b0 ;
  assign n12802 = n12801 ^ n3744 ^ 1'b0 ;
  assign n12803 = ( n8286 & n12800 ) | ( n8286 & n12802 ) | ( n12800 & n12802 ) ;
  assign n12804 = n9980 ^ n5373 ^ n2472 ;
  assign n12805 = n6445 ^ n6241 ^ n2170 ;
  assign n12806 = n12804 & n12805 ;
  assign n12807 = n9943 & n12806 ;
  assign n12808 = n4428 ^ n2498 ^ 1'b0 ;
  assign n12809 = n10136 & n12808 ;
  assign n12810 = n12809 ^ n11937 ^ n8283 ;
  assign n12813 = n3994 ^ n2845 ^ n1455 ;
  assign n12811 = ( ~n3551 & n6070 ) | ( ~n3551 & n7922 ) | ( n6070 & n7922 ) ;
  assign n12812 = n12811 ^ n7795 ^ n5303 ;
  assign n12814 = n12813 ^ n12812 ^ n12294 ;
  assign n12815 = ( n5536 & n5709 ) | ( n5536 & ~n6303 ) | ( n5709 & ~n6303 ) ;
  assign n12816 = n4188 | n12648 ;
  assign n12817 = n2949 | n12816 ;
  assign n12818 = n12815 & n12817 ;
  assign n12819 = ( n3893 & n5703 ) | ( n3893 & n10875 ) | ( n5703 & n10875 ) ;
  assign n12820 = n262 & ~n1897 ;
  assign n12821 = n12820 ^ n1940 ^ 1'b0 ;
  assign n12822 = n12821 ^ n6299 ^ n4233 ;
  assign n12823 = ( n2577 & ~n12819 ) | ( n2577 & n12822 ) | ( ~n12819 & n12822 ) ;
  assign n12824 = n2272 ^ n950 ^ x95 ;
  assign n12825 = ( n3793 & ~n9041 ) | ( n3793 & n12824 ) | ( ~n9041 & n12824 ) ;
  assign n12826 = ( n3114 & n6098 ) | ( n3114 & ~n11989 ) | ( n6098 & ~n11989 ) ;
  assign n12827 = n12826 ^ n1031 ^ n848 ;
  assign n12828 = ( n5466 & n5706 ) | ( n5466 & ~n12827 ) | ( n5706 & ~n12827 ) ;
  assign n12829 = ( ~n7055 & n12825 ) | ( ~n7055 & n12828 ) | ( n12825 & n12828 ) ;
  assign n12830 = n8432 ^ n7776 ^ n4702 ;
  assign n12835 = ( ~n680 & n736 ) | ( ~n680 & n3375 ) | ( n736 & n3375 ) ;
  assign n12832 = n6714 ^ n729 ^ n533 ;
  assign n12833 = n12832 ^ n3379 ^ 1'b0 ;
  assign n12834 = ( n2216 & n7433 ) | ( n2216 & ~n12833 ) | ( n7433 & ~n12833 ) ;
  assign n12831 = ( n3048 & n6666 ) | ( n3048 & n7559 ) | ( n6666 & n7559 ) ;
  assign n12836 = n12835 ^ n12834 ^ n12831 ;
  assign n12837 = n12836 ^ n10385 ^ n5813 ;
  assign n12843 = n2183 ^ n1454 ^ 1'b0 ;
  assign n12841 = n9529 ^ n8546 ^ n2395 ;
  assign n12842 = n12841 ^ n9422 ^ 1'b0 ;
  assign n12838 = n4688 ^ n3608 ^ n2036 ;
  assign n12839 = n12838 ^ n5388 ^ n3888 ;
  assign n12840 = n12839 ^ n12821 ^ n3199 ;
  assign n12844 = n12843 ^ n12842 ^ n12840 ;
  assign n12845 = ( ~n1783 & n4401 ) | ( ~n1783 & n10344 ) | ( n4401 & n10344 ) ;
  assign n12846 = ( n302 & n7792 ) | ( n302 & ~n12845 ) | ( n7792 & ~n12845 ) ;
  assign n12847 = n7658 ^ n7334 ^ n5564 ;
  assign n12848 = n9703 & ~n12847 ;
  assign n12849 = n8096 & ~n12848 ;
  assign n12850 = n12849 ^ n11464 ^ 1'b0 ;
  assign n12852 = ( n5180 & n5191 ) | ( n5180 & ~n8374 ) | ( n5191 & ~n8374 ) ;
  assign n12856 = n5618 ^ n990 ^ x208 ;
  assign n12853 = ( x27 & ~x198 ) | ( x27 & n2106 ) | ( ~x198 & n2106 ) ;
  assign n12854 = ( n519 & n654 ) | ( n519 & ~n9654 ) | ( n654 & ~n9654 ) ;
  assign n12855 = n12853 & n12854 ;
  assign n12857 = n12856 ^ n12855 ^ 1'b0 ;
  assign n12858 = ( n3693 & n11277 ) | ( n3693 & n12857 ) | ( n11277 & n12857 ) ;
  assign n12859 = ( n12273 & n12852 ) | ( n12273 & ~n12858 ) | ( n12852 & ~n12858 ) ;
  assign n12851 = n11032 ^ n3353 ^ 1'b0 ;
  assign n12860 = n12859 ^ n12851 ^ n10252 ;
  assign n12869 = ~n3932 & n4110 ;
  assign n12867 = x80 & n5067 ;
  assign n12861 = n6917 ^ n1515 ^ n571 ;
  assign n12862 = ( n2505 & ~n3828 ) | ( n2505 & n12861 ) | ( ~n3828 & n12861 ) ;
  assign n12863 = n12862 ^ n3796 ^ 1'b0 ;
  assign n12864 = ~n1509 & n12863 ;
  assign n12865 = ( ~n1742 & n5316 ) | ( ~n1742 & n12864 ) | ( n5316 & n12864 ) ;
  assign n12866 = ~n5723 & n12865 ;
  assign n12868 = n12867 ^ n12866 ^ 1'b0 ;
  assign n12870 = n12869 ^ n12868 ^ n10332 ;
  assign n12871 = n10134 ^ n7523 ^ n4189 ;
  assign n12872 = ( ~n7100 & n7492 ) | ( ~n7100 & n8042 ) | ( n7492 & n8042 ) ;
  assign n12873 = ( n3524 & n10439 ) | ( n3524 & n12872 ) | ( n10439 & n12872 ) ;
  assign n12874 = n12873 ^ n5088 ^ 1'b0 ;
  assign n12875 = ~n12871 & n12874 ;
  assign n12880 = n3708 ^ n1208 ^ 1'b0 ;
  assign n12881 = n12880 ^ n7274 ^ 1'b0 ;
  assign n12877 = ( n849 & ~n4904 ) | ( n849 & n7217 ) | ( ~n4904 & n7217 ) ;
  assign n12878 = n5579 & ~n12877 ;
  assign n12879 = ~n10455 & n12878 ;
  assign n12876 = n9445 ^ n8430 ^ n666 ;
  assign n12882 = n12881 ^ n12879 ^ n12876 ;
  assign n12883 = n12882 ^ n3231 ^ 1'b0 ;
  assign n12889 = x144 & ~n1090 ;
  assign n12890 = ~x206 & n12889 ;
  assign n12891 = n1701 & ~n5476 ;
  assign n12892 = ( n10140 & n12890 ) | ( n10140 & n12891 ) | ( n12890 & n12891 ) ;
  assign n12887 = n12578 ^ n4743 ^ n2610 ;
  assign n12888 = ~n2179 & n12887 ;
  assign n12893 = n12892 ^ n12888 ^ 1'b0 ;
  assign n12884 = ( ~n1795 & n1881 ) | ( ~n1795 & n2773 ) | ( n1881 & n2773 ) ;
  assign n12885 = ~n2928 & n12884 ;
  assign n12886 = n6229 | n12885 ;
  assign n12894 = n12893 ^ n12886 ^ 1'b0 ;
  assign n12895 = n12476 ^ n10554 ^ 1'b0 ;
  assign n12897 = n6299 ^ n4074 ^ n566 ;
  assign n12896 = n12317 ^ n6078 ^ n4896 ;
  assign n12898 = n12897 ^ n12896 ^ 1'b0 ;
  assign n12903 = n1224 | n5275 ;
  assign n12904 = n7177 & ~n12903 ;
  assign n12899 = ( n8618 & n12648 ) | ( n8618 & ~n12853 ) | ( n12648 & ~n12853 ) ;
  assign n12900 = n1582 & n2912 ;
  assign n12901 = n12900 ^ n4122 ^ 1'b0 ;
  assign n12902 = n12899 | n12901 ;
  assign n12905 = n12904 ^ n12902 ^ n371 ;
  assign n12906 = ( ~n7949 & n12898 ) | ( ~n7949 & n12905 ) | ( n12898 & n12905 ) ;
  assign n12908 = ( n8737 & ~n9085 ) | ( n8737 & n12221 ) | ( ~n9085 & n12221 ) ;
  assign n12907 = n10949 ^ n2050 ^ n426 ;
  assign n12909 = n12908 ^ n12907 ^ 1'b0 ;
  assign n12910 = n7797 ^ n4712 ^ 1'b0 ;
  assign n12911 = ( n1600 & ~n2255 ) | ( n1600 & n12910 ) | ( ~n2255 & n12910 ) ;
  assign n12912 = n5542 ^ n2467 ^ 1'b0 ;
  assign n12913 = ~n12911 & n12912 ;
  assign n12914 = n12913 ^ n6045 ^ 1'b0 ;
  assign n12915 = n12909 | n12914 ;
  assign n12916 = n12915 ^ n8786 ^ 1'b0 ;
  assign n12917 = n11038 ^ n3047 ^ n2440 ;
  assign n12918 = n10947 ^ n9712 ^ n4453 ;
  assign n12919 = n12918 ^ n11781 ^ n3298 ;
  assign n12920 = n12919 ^ n12203 ^ n9737 ;
  assign n12921 = n8088 ^ n995 ^ 1'b0 ;
  assign n12922 = n12921 ^ n11079 ^ n8534 ;
  assign n12923 = ( n2505 & n10311 ) | ( n2505 & n12922 ) | ( n10311 & n12922 ) ;
  assign n12924 = n8831 ^ n5506 ^ n2640 ;
  assign n12933 = n521 | n7662 ;
  assign n12934 = n12933 ^ x223 ^ 1'b0 ;
  assign n12925 = n4115 ^ n2543 ^ 1'b0 ;
  assign n12926 = n1138 & n12925 ;
  assign n12927 = ( ~x64 & n2430 ) | ( ~x64 & n3576 ) | ( n2430 & n3576 ) ;
  assign n12928 = n12927 ^ x62 ^ 1'b0 ;
  assign n12929 = n12926 & ~n12928 ;
  assign n12930 = ( n4883 & n5933 ) | ( n4883 & n12929 ) | ( n5933 & n12929 ) ;
  assign n12931 = ( n3793 & ~n5451 ) | ( n3793 & n12930 ) | ( ~n5451 & n12930 ) ;
  assign n12932 = n12931 ^ n10426 ^ n7521 ;
  assign n12935 = n12934 ^ n12932 ^ n8985 ;
  assign n12936 = ( n1399 & n5910 ) | ( n1399 & n7451 ) | ( n5910 & n7451 ) ;
  assign n12937 = n12936 ^ n3274 ^ 1'b0 ;
  assign n12938 = n9231 & n12937 ;
  assign n12939 = n4344 & ~n12938 ;
  assign n12942 = x215 & n4198 ;
  assign n12943 = n12942 ^ n9192 ^ n3796 ;
  assign n12944 = n12943 ^ n8096 ^ n2482 ;
  assign n12945 = ( n9284 & n9450 ) | ( n9284 & ~n12944 ) | ( n9450 & ~n12944 ) ;
  assign n12940 = n10143 ^ n8836 ^ n3844 ;
  assign n12941 = n12940 ^ n7182 ^ n5954 ;
  assign n12946 = n12945 ^ n12941 ^ n687 ;
  assign n12947 = n6975 ^ n2071 ^ 1'b0 ;
  assign n12948 = n9555 ^ n6468 ^ n2327 ;
  assign n12949 = n11917 ^ n3525 ^ n2876 ;
  assign n12950 = n12949 ^ n8505 ^ n5454 ;
  assign n12951 = n12950 ^ n11715 ^ n9126 ;
  assign n12952 = ( n12947 & ~n12948 ) | ( n12947 & n12951 ) | ( ~n12948 & n12951 ) ;
  assign n12953 = ( n1423 & n5088 ) | ( n1423 & n9306 ) | ( n5088 & n9306 ) ;
  assign n12954 = n12390 ^ n1320 ^ 1'b0 ;
  assign n12955 = n11016 & n12954 ;
  assign n12956 = n12955 ^ n11769 ^ 1'b0 ;
  assign n12957 = ( n7359 & n10584 ) | ( n7359 & ~n12956 ) | ( n10584 & ~n12956 ) ;
  assign n12958 = ( n2371 & ~n5716 ) | ( n2371 & n12957 ) | ( ~n5716 & n12957 ) ;
  assign n12959 = ( n5422 & n10100 ) | ( n5422 & ~n12390 ) | ( n10100 & ~n12390 ) ;
  assign n12960 = n11289 ^ n9706 ^ n3247 ;
  assign n12961 = n12959 & ~n12960 ;
  assign n12962 = n9319 & n12961 ;
  assign n12963 = ( x160 & ~n2054 ) | ( x160 & n4216 ) | ( ~n2054 & n4216 ) ;
  assign n12964 = n12963 ^ n6680 ^ n1399 ;
  assign n12965 = ( x3 & n2773 ) | ( x3 & n3862 ) | ( n2773 & n3862 ) ;
  assign n12966 = n12965 ^ n6467 ^ n3759 ;
  assign n12967 = n4209 | n12966 ;
  assign n12968 = n12964 & ~n12967 ;
  assign n12969 = ( n3867 & ~n4913 ) | ( n3867 & n10285 ) | ( ~n4913 & n10285 ) ;
  assign n12970 = n5347 ^ n3551 ^ 1'b0 ;
  assign n12971 = n4578 ^ n4214 ^ 1'b0 ;
  assign n12972 = n10273 | n12971 ;
  assign n12973 = ( ~n822 & n884 ) | ( ~n822 & n12972 ) | ( n884 & n12972 ) ;
  assign n12978 = n4323 & ~n12580 ;
  assign n12979 = n12978 ^ n6649 ^ 1'b0 ;
  assign n12974 = ( x150 & n5323 ) | ( x150 & ~n8434 ) | ( n5323 & ~n8434 ) ;
  assign n12975 = ( n3927 & ~n4861 ) | ( n3927 & n12974 ) | ( ~n4861 & n12974 ) ;
  assign n12976 = n12975 ^ n6086 ^ 1'b0 ;
  assign n12977 = ~n6229 & n12976 ;
  assign n12980 = n12979 ^ n12977 ^ 1'b0 ;
  assign n12981 = ( n3405 & n12973 ) | ( n3405 & ~n12980 ) | ( n12973 & ~n12980 ) ;
  assign n12982 = ( n4749 & n12970 ) | ( n4749 & ~n12981 ) | ( n12970 & ~n12981 ) ;
  assign n12983 = n11129 ^ n7606 ^ 1'b0 ;
  assign n12984 = ( ~x106 & n2154 ) | ( ~x106 & n2517 ) | ( n2154 & n2517 ) ;
  assign n12985 = n9325 ^ n3221 ^ 1'b0 ;
  assign n12986 = n12984 & n12985 ;
  assign n12987 = ( ~n2310 & n2677 ) | ( ~n2310 & n12986 ) | ( n2677 & n12986 ) ;
  assign n12988 = ( n2156 & ~n2484 ) | ( n2156 & n5006 ) | ( ~n2484 & n5006 ) ;
  assign n12989 = ( ~n1662 & n2212 ) | ( ~n1662 & n12988 ) | ( n2212 & n12988 ) ;
  assign n12990 = ( n1944 & n2071 ) | ( n1944 & n12989 ) | ( n2071 & n12989 ) ;
  assign n12991 = n7843 ^ n5769 ^ 1'b0 ;
  assign n12992 = n12990 & n12991 ;
  assign n12993 = n12992 ^ n5343 ^ n3820 ;
  assign n13005 = n6644 ^ n1018 ^ n334 ;
  assign n13006 = n13005 ^ n7887 ^ n2263 ;
  assign n13007 = n13006 ^ n6567 ^ n3825 ;
  assign n13003 = n3079 ^ n898 ^ 1'b0 ;
  assign n13000 = n6312 ^ n3627 ^ 1'b0 ;
  assign n12994 = n6915 ^ n5294 ^ n4981 ;
  assign n12995 = ( n284 & ~n885 ) | ( n284 & n2507 ) | ( ~n885 & n2507 ) ;
  assign n12996 = ( n3355 & n3779 ) | ( n3355 & n8346 ) | ( n3779 & n8346 ) ;
  assign n12997 = ( n3015 & n3715 ) | ( n3015 & n12996 ) | ( n3715 & n12996 ) ;
  assign n12998 = ( n1942 & n12995 ) | ( n1942 & ~n12997 ) | ( n12995 & ~n12997 ) ;
  assign n12999 = n12994 & ~n12998 ;
  assign n13001 = n13000 ^ n12999 ^ 1'b0 ;
  assign n13002 = ( n3209 & n12891 ) | ( n3209 & n13001 ) | ( n12891 & n13001 ) ;
  assign n13004 = n13003 ^ n13002 ^ n4211 ;
  assign n13008 = n13007 ^ n13004 ^ n1646 ;
  assign n13009 = n13008 ^ n12625 ^ 1'b0 ;
  assign n13010 = n862 & ~n5967 ;
  assign n13011 = n13010 ^ n6383 ^ 1'b0 ;
  assign n13012 = n10736 ^ n9555 ^ 1'b0 ;
  assign n13013 = n9834 & ~n13012 ;
  assign n13014 = n10978 & n12306 ;
  assign n13015 = n13014 ^ n11850 ^ n686 ;
  assign n13016 = ( n12721 & n13013 ) | ( n12721 & n13015 ) | ( n13013 & n13015 ) ;
  assign n13017 = n4873 ^ n3843 ^ n1495 ;
  assign n13018 = ( ~n1099 & n6656 ) | ( ~n1099 & n13017 ) | ( n6656 & n13017 ) ;
  assign n13019 = n13018 ^ n7457 ^ n5352 ;
  assign n13020 = n13019 ^ n11828 ^ x246 ;
  assign n13021 = n11572 ^ n9689 ^ n7455 ;
  assign n13022 = n13021 ^ n6549 ^ n1164 ;
  assign n13023 = ( n319 & ~n3897 ) | ( n319 & n13022 ) | ( ~n3897 & n13022 ) ;
  assign n13024 = ~n7395 & n11050 ;
  assign n13025 = n3498 & n3691 ;
  assign n13026 = ~n12712 & n13025 ;
  assign n13027 = ~n11740 & n13026 ;
  assign n13028 = n5012 & n7695 ;
  assign n13042 = ( n1177 & n1249 ) | ( n1177 & n3904 ) | ( n1249 & n3904 ) ;
  assign n13043 = n13042 ^ n11152 ^ n8358 ;
  assign n13035 = ( n5233 & ~n8968 ) | ( n5233 & n9819 ) | ( ~n8968 & n9819 ) ;
  assign n13036 = n4666 & n4861 ;
  assign n13037 = n13035 & n13036 ;
  assign n13038 = n311 & ~n4243 ;
  assign n13039 = ~n5745 & n13038 ;
  assign n13040 = ( ~n3027 & n13037 ) | ( ~n3027 & n13039 ) | ( n13037 & n13039 ) ;
  assign n13032 = n9530 ^ n6573 ^ n3776 ;
  assign n13033 = n10490 ^ n2006 ^ n944 ;
  assign n13034 = ( n8269 & n13032 ) | ( n8269 & n13033 ) | ( n13032 & n13033 ) ;
  assign n13041 = n13040 ^ n13034 ^ n10626 ;
  assign n13029 = n11440 ^ n4559 ^ n2643 ;
  assign n13030 = ( ~n1941 & n6625 ) | ( ~n1941 & n13029 ) | ( n6625 & n13029 ) ;
  assign n13031 = n13030 ^ n6632 ^ n1226 ;
  assign n13044 = n13043 ^ n13041 ^ n13031 ;
  assign n13045 = ( n1325 & n2105 ) | ( n1325 & n2613 ) | ( n2105 & n2613 ) ;
  assign n13046 = n13045 ^ n936 ^ 1'b0 ;
  assign n13047 = n4257 & n13046 ;
  assign n13048 = n315 & n12372 ;
  assign n13049 = n13048 ^ n3824 ^ 1'b0 ;
  assign n13050 = n13049 ^ n10388 ^ n4423 ;
  assign n13051 = ( n8019 & n11040 ) | ( n8019 & ~n13050 ) | ( n11040 & ~n13050 ) ;
  assign n13052 = ( ~n375 & n7816 ) | ( ~n375 & n9382 ) | ( n7816 & n9382 ) ;
  assign n13053 = ( ~n5614 & n7832 ) | ( ~n5614 & n13052 ) | ( n7832 & n13052 ) ;
  assign n13054 = ~n2083 & n2967 ;
  assign n13055 = ( ~n612 & n823 ) | ( ~n612 & n13054 ) | ( n823 & n13054 ) ;
  assign n13056 = n13053 & ~n13055 ;
  assign n13057 = n13051 & n13056 ;
  assign n13058 = n5421 & n12206 ;
  assign n13074 = n10132 ^ n2923 ^ 1'b0 ;
  assign n13069 = n5701 | n5997 ;
  assign n13070 = ( ~n1020 & n5930 ) | ( ~n1020 & n13069 ) | ( n5930 & n13069 ) ;
  assign n13071 = ~n936 & n13070 ;
  assign n13066 = n3497 ^ x132 ^ 1'b0 ;
  assign n13067 = n2310 & ~n8793 ;
  assign n13068 = n13066 & n13067 ;
  assign n13062 = n5148 ^ n4877 ^ n4020 ;
  assign n13063 = ( n850 & n2588 ) | ( n850 & ~n5326 ) | ( n2588 & ~n5326 ) ;
  assign n13064 = n13063 ^ n9642 ^ 1'b0 ;
  assign n13065 = n13062 | n13064 ;
  assign n13072 = n13071 ^ n13068 ^ n13065 ;
  assign n13073 = n13072 ^ n3490 ^ n2391 ;
  assign n13059 = ( n959 & n3725 ) | ( n959 & n7403 ) | ( n3725 & n7403 ) ;
  assign n13060 = n13059 ^ n11147 ^ n4172 ;
  assign n13061 = n13060 ^ n10919 ^ n9418 ;
  assign n13075 = n13074 ^ n13073 ^ n13061 ;
  assign n13076 = n7079 ^ n2156 ^ 1'b0 ;
  assign n13077 = x18 & ~n13076 ;
  assign n13078 = ~n11848 & n12819 ;
  assign n13079 = ~n9151 & n13078 ;
  assign n13080 = n4674 & ~n13079 ;
  assign n13081 = ~n11801 & n13080 ;
  assign n13082 = ( n10168 & n13077 ) | ( n10168 & n13081 ) | ( n13077 & n13081 ) ;
  assign n13083 = n9418 ^ x196 ^ 1'b0 ;
  assign n13084 = n13083 ^ n10877 ^ 1'b0 ;
  assign n13085 = n7204 ^ n6341 ^ n4233 ;
  assign n13086 = ( n567 & ~n5368 ) | ( n567 & n10158 ) | ( ~n5368 & n10158 ) ;
  assign n13087 = ( ~n7706 & n13085 ) | ( ~n7706 & n13086 ) | ( n13085 & n13086 ) ;
  assign n13088 = n12286 ^ n4638 ^ n4604 ;
  assign n13089 = n11504 & ~n13088 ;
  assign n13090 = n13089 ^ n12350 ^ 1'b0 ;
  assign n13091 = n11437 | n13090 ;
  assign n13092 = n13087 | n13091 ;
  assign n13093 = n13092 ^ n7229 ^ 1'b0 ;
  assign n13094 = n9777 ^ n2649 ^ n659 ;
  assign n13095 = ( ~n4365 & n9635 ) | ( ~n4365 & n11078 ) | ( n9635 & n11078 ) ;
  assign n13102 = ( n1129 & n5628 ) | ( n1129 & n6577 ) | ( n5628 & n6577 ) ;
  assign n13098 = n1165 | n2762 ;
  assign n13099 = n13098 ^ n2525 ^ n525 ;
  assign n13100 = n13099 ^ n4401 ^ x235 ;
  assign n13096 = ( n1258 & n3150 ) | ( n1258 & n6366 ) | ( n3150 & n6366 ) ;
  assign n13097 = n4946 & ~n13096 ;
  assign n13101 = n13100 ^ n13097 ^ 1'b0 ;
  assign n13103 = n13102 ^ n13101 ^ n5438 ;
  assign n13104 = n13021 ^ n508 ^ 1'b0 ;
  assign n13105 = n9270 & ~n13104 ;
  assign n13106 = n10894 ^ n396 ^ 1'b0 ;
  assign n13107 = n13105 & n13106 ;
  assign n13108 = n1761 ^ n1758 ^ n693 ;
  assign n13109 = n13108 ^ n4637 ^ 1'b0 ;
  assign n13110 = n13109 ^ n10589 ^ n7675 ;
  assign n13111 = n10345 & n13110 ;
  assign n13112 = ( n828 & n6504 ) | ( n828 & n12350 ) | ( n6504 & n12350 ) ;
  assign n13114 = n4347 ^ n3968 ^ x242 ;
  assign n13115 = n13114 ^ n4275 ^ n3871 ;
  assign n13113 = n11935 ^ n10463 ^ x131 ;
  assign n13116 = n13115 ^ n13113 ^ 1'b0 ;
  assign n13117 = n6426 & ~n13116 ;
  assign n13118 = n13117 ^ n2711 ^ 1'b0 ;
  assign n13119 = n6299 ^ n5450 ^ n332 ;
  assign n13120 = ( x13 & ~n2060 ) | ( x13 & n4108 ) | ( ~n2060 & n4108 ) ;
  assign n13121 = n13120 ^ n7047 ^ 1'b0 ;
  assign n13122 = ~n13119 & n13121 ;
  assign n13123 = n13122 ^ n9257 ^ n2909 ;
  assign n13124 = ( n13112 & ~n13118 ) | ( n13112 & n13123 ) | ( ~n13118 & n13123 ) ;
  assign n13125 = n8551 ^ n1985 ^ 1'b0 ;
  assign n13126 = ~n2107 & n13125 ;
  assign n13127 = ( x16 & n1739 ) | ( x16 & n2858 ) | ( n1739 & n2858 ) ;
  assign n13128 = n13127 ^ n4205 ^ n3058 ;
  assign n13129 = n8710 ^ n3883 ^ 1'b0 ;
  assign n13130 = ~n13128 & n13129 ;
  assign n13131 = n13130 ^ n3557 ^ 1'b0 ;
  assign n13132 = n13126 & n13131 ;
  assign n13133 = n13132 ^ n11288 ^ n3476 ;
  assign n13136 = ( n365 & ~n417 ) | ( n365 & n1724 ) | ( ~n417 & n1724 ) ;
  assign n13134 = n1324 & n7542 ;
  assign n13135 = n10202 & n13134 ;
  assign n13137 = n13136 ^ n13135 ^ n10965 ;
  assign n13138 = n10272 ^ n5648 ^ n1622 ;
  assign n13139 = ( ~n7894 & n8116 ) | ( ~n7894 & n13138 ) | ( n8116 & n13138 ) ;
  assign n13140 = ( n407 & n3587 ) | ( n407 & n13139 ) | ( n3587 & n13139 ) ;
  assign n13141 = n13140 ^ n4028 ^ 1'b0 ;
  assign n13142 = n5780 & ~n13141 ;
  assign n13143 = ~n5769 & n13142 ;
  assign n13144 = n13143 ^ n2088 ^ 1'b0 ;
  assign n13145 = ( ~n3989 & n9930 ) | ( ~n3989 & n13144 ) | ( n9930 & n13144 ) ;
  assign n13146 = n10702 ^ n8791 ^ n1279 ;
  assign n13147 = n11828 ^ n7548 ^ n5613 ;
  assign n13148 = ( ~n7206 & n8447 ) | ( ~n7206 & n13147 ) | ( n8447 & n13147 ) ;
  assign n13149 = ( ~n6777 & n13146 ) | ( ~n6777 & n13148 ) | ( n13146 & n13148 ) ;
  assign n13152 = n11685 ^ n5980 ^ n1932 ;
  assign n13150 = ( x66 & n295 ) | ( x66 & n2242 ) | ( n295 & n2242 ) ;
  assign n13151 = ( n5170 & n8191 ) | ( n5170 & ~n13150 ) | ( n8191 & ~n13150 ) ;
  assign n13153 = n13152 ^ n13151 ^ n4412 ;
  assign n13154 = ( x27 & ~n5546 ) | ( x27 & n13153 ) | ( ~n5546 & n13153 ) ;
  assign n13155 = n5485 & n13154 ;
  assign n13156 = n6047 & n13155 ;
  assign n13157 = n12107 ^ n9609 ^ 1'b0 ;
  assign n13158 = ( n3013 & n7872 ) | ( n3013 & n11887 ) | ( n7872 & n11887 ) ;
  assign n13159 = n8034 ^ n1956 ^ 1'b0 ;
  assign n13160 = n13159 ^ n8315 ^ n8167 ;
  assign n13161 = n13160 ^ n4568 ^ n3689 ;
  assign n13162 = ( ~x94 & n6853 ) | ( ~x94 & n13161 ) | ( n6853 & n13161 ) ;
  assign n13167 = n7468 ^ n2922 ^ n1438 ;
  assign n13168 = ~n633 & n13167 ;
  assign n13169 = ~n8651 & n13168 ;
  assign n13166 = n5065 | n5870 ;
  assign n13163 = n2536 & n3841 ;
  assign n13164 = ~n2981 & n13163 ;
  assign n13165 = n13164 ^ n8901 ^ 1'b0 ;
  assign n13170 = n13169 ^ n13166 ^ n13165 ;
  assign n13171 = ( n1030 & ~n5090 ) | ( n1030 & n13170 ) | ( ~n5090 & n13170 ) ;
  assign n13173 = n10326 ^ n937 ^ x200 ;
  assign n13174 = n13173 ^ x101 ^ 1'b0 ;
  assign n13175 = n12117 | n13174 ;
  assign n13176 = n13175 ^ n2889 ^ n864 ;
  assign n13177 = n6323 ^ n4518 ^ 1'b0 ;
  assign n13178 = ~n11370 & n13177 ;
  assign n13179 = n12149 & n13178 ;
  assign n13180 = ~n13176 & n13179 ;
  assign n13172 = x158 & n1289 ;
  assign n13181 = n13180 ^ n13172 ^ 1'b0 ;
  assign n13182 = n4981 | n6936 ;
  assign n13185 = n11926 & ~n13108 ;
  assign n13186 = ~n418 & n13185 ;
  assign n13183 = n4801 & ~n7098 ;
  assign n13184 = n13183 ^ n632 ^ 1'b0 ;
  assign n13187 = n13186 ^ n13184 ^ n8581 ;
  assign n13188 = ( ~n9270 & n9635 ) | ( ~n9270 & n10117 ) | ( n9635 & n10117 ) ;
  assign n13189 = ( n2733 & n3563 ) | ( n2733 & n5380 ) | ( n3563 & n5380 ) ;
  assign n13190 = ( n4198 & n8219 ) | ( n4198 & n13189 ) | ( n8219 & n13189 ) ;
  assign n13191 = n13190 ^ n3174 ^ 1'b0 ;
  assign n13192 = n13191 ^ n4683 ^ 1'b0 ;
  assign n13193 = ~n13188 & n13192 ;
  assign n13194 = n13187 & n13193 ;
  assign n13196 = n11812 ^ n3236 ^ n2222 ;
  assign n13195 = n7341 & ~n10987 ;
  assign n13197 = n13196 ^ n13195 ^ 1'b0 ;
  assign n13198 = n8728 ^ x68 ^ 1'b0 ;
  assign n13199 = ~x156 & n13198 ;
  assign n13200 = ( n1414 & n1441 ) | ( n1414 & n3578 ) | ( n1441 & n3578 ) ;
  assign n13201 = ( n1863 & ~n2269 ) | ( n1863 & n3288 ) | ( ~n2269 & n3288 ) ;
  assign n13202 = n13201 ^ n9545 ^ n5417 ;
  assign n13203 = ( n3071 & n13200 ) | ( n3071 & n13202 ) | ( n13200 & n13202 ) ;
  assign n13204 = n13203 ^ n4545 ^ 1'b0 ;
  assign n13205 = n10033 | n13204 ;
  assign n13206 = n1355 & n2550 ;
  assign n13207 = n13206 ^ n11502 ^ 1'b0 ;
  assign n13208 = n2110 & ~n13207 ;
  assign n13209 = ( ~n3258 & n6687 ) | ( ~n3258 & n9229 ) | ( n6687 & n9229 ) ;
  assign n13210 = ( n2205 & n11901 ) | ( n2205 & n13209 ) | ( n11901 & n13209 ) ;
  assign n13211 = ( ~n6878 & n7735 ) | ( ~n6878 & n11533 ) | ( n7735 & n11533 ) ;
  assign n13212 = x83 & ~n5997 ;
  assign n13213 = n13212 ^ n1412 ^ 1'b0 ;
  assign n13214 = n13213 ^ n6975 ^ n6929 ;
  assign n13215 = ~n4543 & n4647 ;
  assign n13216 = ~n13214 & n13215 ;
  assign n13217 = ( n7750 & n13211 ) | ( n7750 & ~n13216 ) | ( n13211 & ~n13216 ) ;
  assign n13218 = n12635 ^ n5797 ^ 1'b0 ;
  assign n13219 = n3648 & n13218 ;
  assign n13221 = ( n1481 & ~n5873 ) | ( n1481 & n9662 ) | ( ~n5873 & n9662 ) ;
  assign n13220 = ~n5285 & n7999 ;
  assign n13222 = n13221 ^ n13220 ^ n11553 ;
  assign n13223 = ( n1323 & ~n4693 ) | ( n1323 & n13222 ) | ( ~n4693 & n13222 ) ;
  assign n13224 = n3767 | n11740 ;
  assign n13225 = n9224 ^ n4341 ^ 1'b0 ;
  assign n13226 = n13225 ^ n10966 ^ n7821 ;
  assign n13233 = ( n1959 & n5538 ) | ( n1959 & n7596 ) | ( n5538 & n7596 ) ;
  assign n13234 = n13233 ^ n6191 ^ n2484 ;
  assign n13235 = n9834 ^ n8305 ^ n6898 ;
  assign n13236 = ( n845 & n11427 ) | ( n845 & ~n13235 ) | ( n11427 & ~n13235 ) ;
  assign n13237 = ( n6543 & ~n13234 ) | ( n6543 & n13236 ) | ( ~n13234 & n13236 ) ;
  assign n13229 = x67 & n8191 ;
  assign n13230 = n13229 ^ n6772 ^ 1'b0 ;
  assign n13227 = n2556 & ~n6497 ;
  assign n13228 = n13227 ^ n6917 ^ 1'b0 ;
  assign n13231 = n13230 ^ n13228 ^ n6326 ;
  assign n13232 = ~n7431 & n13231 ;
  assign n13238 = n13237 ^ n13232 ^ 1'b0 ;
  assign n13239 = n13238 ^ n12233 ^ 1'b0 ;
  assign n13240 = n1912 | n13239 ;
  assign n13241 = ( ~n1599 & n4419 ) | ( ~n1599 & n12556 ) | ( n4419 & n12556 ) ;
  assign n13242 = ( ~n466 & n5288 ) | ( ~n466 & n13241 ) | ( n5288 & n13241 ) ;
  assign n13244 = n3997 ^ n3563 ^ 1'b0 ;
  assign n13243 = n9420 & ~n11848 ;
  assign n13245 = n13244 ^ n13243 ^ 1'b0 ;
  assign n13246 = ( n5889 & n7781 ) | ( n5889 & n12930 ) | ( n7781 & n12930 ) ;
  assign n13252 = ~n5636 & n8608 ;
  assign n13249 = ( n3441 & n3992 ) | ( n3441 & n4712 ) | ( n3992 & n4712 ) ;
  assign n13250 = n13249 ^ n5089 ^ n525 ;
  assign n13247 = n644 | n2024 ;
  assign n13248 = n13247 ^ n5502 ^ 1'b0 ;
  assign n13251 = n13250 ^ n13248 ^ n2142 ;
  assign n13253 = n13252 ^ n13251 ^ n3417 ;
  assign n13254 = ( n3674 & n5243 ) | ( n3674 & n13253 ) | ( n5243 & n13253 ) ;
  assign n13255 = ( ~n4489 & n13246 ) | ( ~n4489 & n13254 ) | ( n13246 & n13254 ) ;
  assign n13256 = n5012 | n6227 ;
  assign n13257 = x124 | n13256 ;
  assign n13258 = n12148 ^ n3293 ^ 1'b0 ;
  assign n13259 = n11285 ^ n7456 ^ n2167 ;
  assign n13260 = n2625 & ~n13259 ;
  assign n13261 = ~n13258 & n13260 ;
  assign n13262 = n13261 ^ n9677 ^ 1'b0 ;
  assign n13263 = ( n3537 & n6891 ) | ( n3537 & ~n6943 ) | ( n6891 & ~n6943 ) ;
  assign n13264 = ( n5331 & ~n12023 ) | ( n5331 & n13263 ) | ( ~n12023 & n13263 ) ;
  assign n13265 = ( n1745 & n3541 ) | ( n1745 & ~n4694 ) | ( n3541 & ~n4694 ) ;
  assign n13268 = ~n6905 & n8755 ;
  assign n13269 = ~n9429 & n13268 ;
  assign n13266 = n5133 ^ n2620 ^ n501 ;
  assign n13267 = n13266 ^ n6275 ^ n2474 ;
  assign n13270 = n13269 ^ n13267 ^ 1'b0 ;
  assign n13271 = n13265 & ~n13270 ;
  assign n13272 = n3185 & ~n4003 ;
  assign n13273 = n13272 ^ n4430 ^ 1'b0 ;
  assign n13274 = ~x33 & n11687 ;
  assign n13275 = n12983 | n13274 ;
  assign n13276 = n7003 & ~n13275 ;
  assign n13282 = n1491 ^ n1172 ^ x231 ;
  assign n13277 = n8773 ^ n3951 ^ 1'b0 ;
  assign n13278 = ~n5966 & n13277 ;
  assign n13279 = ( n735 & n5790 ) | ( n735 & ~n11881 ) | ( n5790 & ~n11881 ) ;
  assign n13280 = n2331 | n13279 ;
  assign n13281 = ( n2783 & n13278 ) | ( n2783 & ~n13280 ) | ( n13278 & ~n13280 ) ;
  assign n13283 = n13282 ^ n13281 ^ n538 ;
  assign n13284 = n5247 & ~n6060 ;
  assign n13285 = n13284 ^ n7106 ^ n854 ;
  assign n13286 = n3714 ^ n2996 ^ n2737 ;
  assign n13287 = n13286 ^ n9924 ^ n4997 ;
  assign n13297 = ( n1236 & n4325 ) | ( n1236 & n8240 ) | ( n4325 & n8240 ) ;
  assign n13294 = ~n5374 & n8651 ;
  assign n13295 = n13294 ^ n5910 ^ 1'b0 ;
  assign n13296 = n13295 ^ n10881 ^ n2383 ;
  assign n13292 = ( ~n2018 & n3996 ) | ( ~n2018 & n8655 ) | ( n3996 & n8655 ) ;
  assign n13293 = n13292 ^ n1274 ^ x105 ;
  assign n13298 = n13297 ^ n13296 ^ n13293 ;
  assign n13289 = ( n1776 & ~n4841 ) | ( n1776 & n6378 ) | ( ~n4841 & n6378 ) ;
  assign n13290 = n13289 ^ n6392 ^ n4698 ;
  assign n13288 = n13225 ^ n12815 ^ x31 ;
  assign n13291 = n13290 ^ n13288 ^ n11706 ;
  assign n13299 = n13298 ^ n13291 ^ n12898 ;
  assign n13300 = n10992 & n12592 ;
  assign n13301 = n13300 ^ n12516 ^ 1'b0 ;
  assign n13302 = n13301 ^ n6632 ^ 1'b0 ;
  assign n13303 = ( ~n4948 & n6110 ) | ( ~n4948 & n13302 ) | ( n6110 & n13302 ) ;
  assign n13304 = ( ~x211 & n1505 ) | ( ~x211 & n7938 ) | ( n1505 & n7938 ) ;
  assign n13314 = ( n1778 & ~n2034 ) | ( n1778 & n7436 ) | ( ~n2034 & n7436 ) ;
  assign n13310 = ~n6288 & n7047 ;
  assign n13311 = ~n4452 & n13310 ;
  assign n13307 = n4301 | n4317 ;
  assign n13308 = n13307 ^ n6578 ^ 1'b0 ;
  assign n13309 = n4256 & n13308 ;
  assign n13312 = n13311 ^ n13309 ^ 1'b0 ;
  assign n13313 = ( n4230 & n7689 ) | ( n4230 & ~n13312 ) | ( n7689 & ~n13312 ) ;
  assign n13305 = x230 & n5546 ;
  assign n13306 = n13305 ^ n5557 ^ n1605 ;
  assign n13315 = n13314 ^ n13313 ^ n13306 ;
  assign n13322 = n6086 ^ n4242 ^ 1'b0 ;
  assign n13316 = ( n3386 & n3616 ) | ( n3386 & n10358 ) | ( n3616 & n10358 ) ;
  assign n13317 = ( n804 & n3557 ) | ( n804 & n6601 ) | ( n3557 & n6601 ) ;
  assign n13318 = n13317 ^ n7175 ^ n4550 ;
  assign n13319 = ( n2559 & n13316 ) | ( n2559 & ~n13318 ) | ( n13316 & ~n13318 ) ;
  assign n13320 = n13319 ^ n10589 ^ n1319 ;
  assign n13321 = n3669 & n13320 ;
  assign n13323 = n13322 ^ n13321 ^ 1'b0 ;
  assign n13325 = ( n3094 & ~n5238 ) | ( n3094 & n12124 ) | ( ~n5238 & n12124 ) ;
  assign n13324 = ( n3563 & ~n4481 ) | ( n3563 & n5627 ) | ( ~n4481 & n5627 ) ;
  assign n13326 = n13325 ^ n13324 ^ 1'b0 ;
  assign n13337 = ( n296 & n746 ) | ( n296 & n7755 ) | ( n746 & n7755 ) ;
  assign n13330 = ( n4391 & n4685 ) | ( n4391 & ~n7953 ) | ( n4685 & ~n7953 ) ;
  assign n13333 = n13136 ^ n4695 ^ n4353 ;
  assign n13334 = ( n11606 & n11876 ) | ( n11606 & ~n13333 ) | ( n11876 & ~n13333 ) ;
  assign n13331 = n8804 ^ n3463 ^ 1'b0 ;
  assign n13332 = n4031 | n13331 ;
  assign n13335 = n13334 ^ n13332 ^ 1'b0 ;
  assign n13336 = ( n3792 & ~n13330 ) | ( n3792 & n13335 ) | ( ~n13330 & n13335 ) ;
  assign n13327 = n7300 ^ n1278 ^ n536 ;
  assign n13328 = n4166 | n13327 ;
  assign n13329 = ~n1491 & n13328 ;
  assign n13338 = n13337 ^ n13336 ^ n13329 ;
  assign n13339 = ~n4606 & n12525 ;
  assign n13340 = ( n5053 & n6200 ) | ( n5053 & ~n12890 ) | ( n6200 & ~n12890 ) ;
  assign n13341 = ( n7581 & ~n13339 ) | ( n7581 & n13340 ) | ( ~n13339 & n13340 ) ;
  assign n13342 = ( n2162 & n3336 ) | ( n2162 & ~n13341 ) | ( n3336 & ~n13341 ) ;
  assign n13343 = n1032 | n2343 ;
  assign n13344 = n13343 ^ n3479 ^ n1499 ;
  assign n13345 = ( n2691 & n5962 ) | ( n2691 & ~n13344 ) | ( n5962 & ~n13344 ) ;
  assign n13346 = n4386 ^ n4129 ^ n1811 ;
  assign n13352 = n2433 | n3581 ;
  assign n13348 = n4887 ^ n3546 ^ x34 ;
  assign n13347 = n11566 ^ n1130 ^ 1'b0 ;
  assign n13349 = n13348 ^ n13347 ^ n4791 ;
  assign n13350 = n12275 & n13349 ;
  assign n13351 = n13350 ^ n8775 ^ 1'b0 ;
  assign n13353 = n13352 ^ n13351 ^ n5655 ;
  assign n13354 = ~n1733 & n13297 ;
  assign n13355 = n13354 ^ n10401 ^ n5467 ;
  assign n13356 = n10987 ^ n3203 ^ n465 ;
  assign n13357 = n10646 ^ n10380 ^ 1'b0 ;
  assign n13358 = n11949 & n13357 ;
  assign n13359 = ( n2388 & n13356 ) | ( n2388 & n13358 ) | ( n13356 & n13358 ) ;
  assign n13360 = n11169 ^ n8695 ^ n4774 ;
  assign n13361 = ( ~n2124 & n3214 ) | ( ~n2124 & n13360 ) | ( n3214 & n13360 ) ;
  assign n13362 = ~n1492 & n7804 ;
  assign n13363 = n13362 ^ n6394 ^ 1'b0 ;
  assign n13364 = n12166 ^ n11164 ^ n9038 ;
  assign n13365 = ( n3977 & n13363 ) | ( n3977 & ~n13364 ) | ( n13363 & ~n13364 ) ;
  assign n13366 = n9186 ^ n6358 ^ 1'b0 ;
  assign n13367 = ~n12120 & n13366 ;
  assign n13368 = n2162 | n13367 ;
  assign n13369 = n3661 ^ n1695 ^ 1'b0 ;
  assign n13370 = n5252 ^ n4432 ^ n1926 ;
  assign n13371 = n7376 ^ n5255 ^ 1'b0 ;
  assign n13372 = ~n1798 & n13371 ;
  assign n13373 = ( n10803 & n12424 ) | ( n10803 & ~n13372 ) | ( n12424 & ~n13372 ) ;
  assign n13374 = n8097 ^ n7787 ^ n5532 ;
  assign n13375 = ( n8411 & n10198 ) | ( n8411 & ~n11696 ) | ( n10198 & ~n11696 ) ;
  assign n13376 = ( ~n3883 & n13374 ) | ( ~n3883 & n13375 ) | ( n13374 & n13375 ) ;
  assign n13377 = n13376 ^ n12916 ^ n6965 ;
  assign n13378 = n5224 ^ x191 ^ 1'b0 ;
  assign n13379 = ( n680 & n4521 ) | ( n680 & n6602 ) | ( n4521 & n6602 ) ;
  assign n13380 = ( n8175 & n11801 ) | ( n8175 & n13379 ) | ( n11801 & n13379 ) ;
  assign n13381 = ( n5276 & ~n6520 ) | ( n5276 & n13380 ) | ( ~n6520 & n13380 ) ;
  assign n13382 = ( n1919 & n12407 ) | ( n1919 & n13381 ) | ( n12407 & n13381 ) ;
  assign n13383 = n13378 | n13382 ;
  assign n13384 = n11289 | n13383 ;
  assign n13385 = n4835 ^ n4565 ^ 1'b0 ;
  assign n13386 = n3450 & ~n4429 ;
  assign n13387 = ~n5442 & n13386 ;
  assign n13388 = ( n11973 & ~n13385 ) | ( n11973 & n13387 ) | ( ~n13385 & n13387 ) ;
  assign n13389 = n8624 ^ n5074 ^ 1'b0 ;
  assign n13390 = n13388 | n13389 ;
  assign n13391 = n13390 ^ n9239 ^ x220 ;
  assign n13392 = n792 & ~n1369 ;
  assign n13393 = n13392 ^ n5193 ^ 1'b0 ;
  assign n13394 = n9462 | n13393 ;
  assign n13395 = n13394 ^ n706 ^ 1'b0 ;
  assign n13396 = n3093 & ~n13395 ;
  assign n13397 = n13396 ^ n12649 ^ n4739 ;
  assign n13400 = n8364 ^ n4313 ^ n1429 ;
  assign n13398 = ( n1774 & n8430 ) | ( n1774 & ~n9646 ) | ( n8430 & ~n9646 ) ;
  assign n13399 = n13398 ^ n3742 ^ n2717 ;
  assign n13401 = n13400 ^ n13399 ^ n10602 ;
  assign n13402 = n10212 ^ x223 ^ 1'b0 ;
  assign n13410 = n2262 & n5268 ;
  assign n13411 = n13410 ^ n2394 ^ 1'b0 ;
  assign n13412 = ( n2877 & ~n7975 ) | ( n2877 & n13411 ) | ( ~n7975 & n13411 ) ;
  assign n13413 = ( n1678 & ~n5343 ) | ( n1678 & n13412 ) | ( ~n5343 & n13412 ) ;
  assign n13407 = n6754 ^ n2687 ^ n701 ;
  assign n13403 = n10516 ^ n6456 ^ n2468 ;
  assign n13404 = ~n2609 & n13403 ;
  assign n13405 = n6624 ^ n3796 ^ n3294 ;
  assign n13406 = ( ~n2835 & n13404 ) | ( ~n2835 & n13405 ) | ( n13404 & n13405 ) ;
  assign n13408 = n13407 ^ n13406 ^ n1525 ;
  assign n13409 = n13408 ^ n6203 ^ n3782 ;
  assign n13414 = n13413 ^ n13409 ^ n4092 ;
  assign n13415 = n6178 ^ n2087 ^ n553 ;
  assign n13416 = n13415 ^ n1152 ^ 1'b0 ;
  assign n13417 = n1814 & n13416 ;
  assign n13418 = n11381 & n13417 ;
  assign n13419 = n13418 ^ n10646 ^ 1'b0 ;
  assign n13420 = n3060 ^ n2774 ^ n2432 ;
  assign n13421 = n10333 & ~n13420 ;
  assign n13422 = ~n9871 & n13421 ;
  assign n13433 = ( n4066 & ~n9152 ) | ( n4066 & n11056 ) | ( ~n9152 & n11056 ) ;
  assign n13432 = n7709 ^ n5812 ^ 1'b0 ;
  assign n13423 = ~n6531 & n8839 ;
  assign n13427 = ( ~n2312 & n2656 ) | ( ~n2312 & n3761 ) | ( n2656 & n3761 ) ;
  assign n13428 = n8714 ^ n8340 ^ n4824 ;
  assign n13429 = ( ~n10657 & n13427 ) | ( ~n10657 & n13428 ) | ( n13427 & n13428 ) ;
  assign n13424 = n7048 ^ n6625 ^ n3979 ;
  assign n13425 = n13424 ^ n5894 ^ n1817 ;
  assign n13426 = ~n6830 & n13425 ;
  assign n13430 = n13429 ^ n13426 ^ 1'b0 ;
  assign n13431 = ( n8202 & n13423 ) | ( n8202 & n13430 ) | ( n13423 & n13430 ) ;
  assign n13434 = n13433 ^ n13432 ^ n13431 ;
  assign n13435 = n9059 ^ n8840 ^ 1'b0 ;
  assign n13436 = ~n8628 & n13435 ;
  assign n13437 = n2426 & n3784 ;
  assign n13439 = n5770 ^ n4663 ^ n1497 ;
  assign n13438 = ( ~n4077 & n5450 ) | ( ~n4077 & n10590 ) | ( n5450 & n10590 ) ;
  assign n13440 = n13439 ^ n13438 ^ n6206 ;
  assign n13441 = ( n1666 & ~n11371 ) | ( n1666 & n13440 ) | ( ~n11371 & n13440 ) ;
  assign n13442 = ( n4951 & n13437 ) | ( n4951 & n13441 ) | ( n13437 & n13441 ) ;
  assign n13443 = n9510 ^ n6746 ^ 1'b0 ;
  assign n13444 = ( ~n2937 & n4211 ) | ( ~n2937 & n11892 ) | ( n4211 & n11892 ) ;
  assign n13445 = ~n8534 & n13444 ;
  assign n13446 = n9294 ^ n3429 ^ 1'b0 ;
  assign n13447 = n5909 | n13446 ;
  assign n13448 = ~n2210 & n5803 ;
  assign n13449 = n7539 ^ n4350 ^ n992 ;
  assign n13456 = ~n2983 & n3782 ;
  assign n13457 = n13456 ^ n1266 ^ 1'b0 ;
  assign n13451 = n4437 & n6691 ;
  assign n13452 = ~n4810 & n13451 ;
  assign n13453 = n5252 | n7786 ;
  assign n13454 = n2962 & ~n13453 ;
  assign n13455 = n13452 | n13454 ;
  assign n13450 = n4156 ^ n1504 ^ 1'b0 ;
  assign n13458 = n13457 ^ n13455 ^ n13450 ;
  assign n13459 = n13458 ^ n6767 ^ n4327 ;
  assign n13460 = ( n5155 & n10442 ) | ( n5155 & n13459 ) | ( n10442 & n13459 ) ;
  assign n13461 = ( ~n11462 & n13449 ) | ( ~n11462 & n13460 ) | ( n13449 & n13460 ) ;
  assign n13462 = n12146 & n12617 ;
  assign n13463 = ( n2213 & ~n6321 ) | ( n2213 & n8082 ) | ( ~n6321 & n8082 ) ;
  assign n13464 = ( n5573 & n13462 ) | ( n5573 & ~n13463 ) | ( n13462 & ~n13463 ) ;
  assign n13465 = n13464 ^ n7022 ^ 1'b0 ;
  assign n13466 = ( n6031 & ~n6290 ) | ( n6031 & n12425 ) | ( ~n6290 & n12425 ) ;
  assign n13467 = n13466 ^ n5036 ^ n4030 ;
  assign n13472 = ( n543 & n3453 ) | ( n543 & ~n3742 ) | ( n3453 & ~n3742 ) ;
  assign n13470 = n5717 | n7274 ;
  assign n13471 = ( n2129 & ~n5653 ) | ( n2129 & n13470 ) | ( ~n5653 & n13470 ) ;
  assign n13468 = n1986 ^ n1914 ^ n1862 ;
  assign n13469 = n13468 ^ n1301 ^ n547 ;
  assign n13473 = n13472 ^ n13471 ^ n13469 ;
  assign n13474 = ( ~n13465 & n13467 ) | ( ~n13465 & n13473 ) | ( n13467 & n13473 ) ;
  assign n13475 = n1056 & n4168 ;
  assign n13476 = ~n3525 & n13475 ;
  assign n13477 = n13476 ^ n11223 ^ n8972 ;
  assign n13478 = n1181 & ~n10137 ;
  assign n13479 = n6029 & n13478 ;
  assign n13480 = n13479 ^ n3341 ^ n2885 ;
  assign n13481 = n7078 ^ n3428 ^ n2609 ;
  assign n13482 = n10278 & n13481 ;
  assign n13483 = ( ~n13122 & n13480 ) | ( ~n13122 & n13482 ) | ( n13480 & n13482 ) ;
  assign n13484 = n11657 ^ n5997 ^ n3671 ;
  assign n13485 = n13484 ^ n5897 ^ 1'b0 ;
  assign n13486 = n7470 ^ n5439 ^ 1'b0 ;
  assign n13487 = n9209 | n13486 ;
  assign n13488 = n13380 | n13487 ;
  assign n13491 = n5658 ^ n2811 ^ n1896 ;
  assign n13489 = n7854 & n9257 ;
  assign n13490 = ( n7413 & ~n11396 ) | ( n7413 & n13489 ) | ( ~n11396 & n13489 ) ;
  assign n13492 = n13491 ^ n13490 ^ n9491 ;
  assign n13493 = n730 ^ x228 ^ x132 ;
  assign n13494 = n13493 ^ n2351 ^ n614 ;
  assign n13495 = ~n2580 & n6232 ;
  assign n13496 = n13495 ^ x190 ^ 1'b0 ;
  assign n13497 = n2824 & ~n13496 ;
  assign n13498 = n5071 & n13497 ;
  assign n13499 = ~n1641 & n3124 ;
  assign n13500 = ( n5156 & ~n13498 ) | ( n5156 & n13499 ) | ( ~n13498 & n13499 ) ;
  assign n13501 = ( ~n2253 & n7834 ) | ( ~n2253 & n13500 ) | ( n7834 & n13500 ) ;
  assign n13502 = ( x246 & n13494 ) | ( x246 & ~n13501 ) | ( n13494 & ~n13501 ) ;
  assign n13503 = ( n1699 & ~n11822 ) | ( n1699 & n13354 ) | ( ~n11822 & n13354 ) ;
  assign n13507 = ( n1889 & n3785 ) | ( n1889 & ~n6226 ) | ( n3785 & ~n6226 ) ;
  assign n13504 = ~n2583 & n5306 ;
  assign n13505 = ~n558 & n13504 ;
  assign n13506 = n13505 ^ n3965 ^ x185 ;
  assign n13508 = n13507 ^ n13506 ^ n3395 ;
  assign n13509 = n13508 ^ n9698 ^ n4525 ;
  assign n13511 = n3565 & n5968 ;
  assign n13512 = n13511 ^ n576 ^ 1'b0 ;
  assign n13513 = ( n465 & ~n7298 ) | ( n465 & n13512 ) | ( ~n7298 & n13512 ) ;
  assign n13510 = ( x234 & n1657 ) | ( x234 & ~n9299 ) | ( n1657 & ~n9299 ) ;
  assign n13514 = n13513 ^ n13510 ^ n2182 ;
  assign n13515 = n9160 ^ n7944 ^ n2734 ;
  assign n13516 = n5201 ^ n5088 ^ 1'b0 ;
  assign n13517 = n13516 ^ n5905 ^ n3504 ;
  assign n13518 = ( n2412 & n13515 ) | ( n2412 & ~n13517 ) | ( n13515 & ~n13517 ) ;
  assign n13519 = n5173 | n13266 ;
  assign n13520 = ( n12791 & ~n13518 ) | ( n12791 & n13519 ) | ( ~n13518 & n13519 ) ;
  assign n13521 = ( n348 & n706 ) | ( n348 & ~n13520 ) | ( n706 & ~n13520 ) ;
  assign n13522 = n8433 ^ n6957 ^ n2659 ;
  assign n13523 = n8890 & n13522 ;
  assign n13524 = n7088 ^ n2051 ^ n482 ;
  assign n13525 = n13524 ^ n5865 ^ n5184 ;
  assign n13526 = n4846 ^ n4521 ^ n394 ;
  assign n13527 = n13526 ^ n7008 ^ 1'b0 ;
  assign n13528 = n6687 & n13527 ;
  assign n13529 = ( n4945 & n13525 ) | ( n4945 & n13528 ) | ( n13525 & n13528 ) ;
  assign n13530 = ( n2473 & n6980 ) | ( n2473 & ~n13529 ) | ( n6980 & ~n13529 ) ;
  assign n13531 = n12730 ^ n8239 ^ 1'b0 ;
  assign n13532 = n13531 ^ n2052 ^ n1572 ;
  assign n13533 = n9267 ^ n6128 ^ 1'b0 ;
  assign n13534 = n13532 | n13533 ;
  assign n13535 = n1078 | n5929 ;
  assign n13536 = n13535 ^ n346 ^ 1'b0 ;
  assign n13537 = ( n284 & n6171 ) | ( n284 & ~n13536 ) | ( n6171 & ~n13536 ) ;
  assign n13542 = n2520 ^ n1723 ^ 1'b0 ;
  assign n13543 = ~n11214 & n13542 ;
  assign n13544 = ( n3472 & n6958 ) | ( n3472 & ~n8080 ) | ( n6958 & ~n8080 ) ;
  assign n13545 = n11991 ^ n4020 ^ n3430 ;
  assign n13546 = ( n13543 & n13544 ) | ( n13543 & ~n13545 ) | ( n13544 & ~n13545 ) ;
  assign n13538 = ~n1666 & n10889 ;
  assign n13539 = n13538 ^ n3523 ^ n3293 ;
  assign n13540 = n2440 & n10579 ;
  assign n13541 = n13539 & n13540 ;
  assign n13547 = n13546 ^ n13541 ^ n12064 ;
  assign n13548 = ( ~n777 & n8655 ) | ( ~n777 & n9617 ) | ( n8655 & n9617 ) ;
  assign n13549 = ( n4837 & n8869 ) | ( n4837 & n13548 ) | ( n8869 & n13548 ) ;
  assign n13550 = ( n3380 & n8604 ) | ( n3380 & n11573 ) | ( n8604 & n11573 ) ;
  assign n13551 = n2797 ^ n1491 ^ x38 ;
  assign n13562 = n8482 ^ n2478 ^ 1'b0 ;
  assign n13563 = n2840 & n13562 ;
  assign n13558 = n12593 ^ n7870 ^ n3889 ;
  assign n13559 = n3830 ^ n2333 ^ n2299 ;
  assign n13560 = ~n3679 & n13559 ;
  assign n13561 = n13558 & n13560 ;
  assign n13556 = n3750 & n7505 ;
  assign n13555 = n530 & n2276 ;
  assign n13557 = n13556 ^ n13555 ^ n7082 ;
  assign n13564 = n13563 ^ n13561 ^ n13557 ;
  assign n13552 = ( ~n5724 & n6438 ) | ( ~n5724 & n6472 ) | ( n6438 & n6472 ) ;
  assign n13553 = n13552 ^ n5963 ^ 1'b0 ;
  assign n13554 = ~n9053 & n13553 ;
  assign n13565 = n13564 ^ n13554 ^ n10790 ;
  assign n13569 = ( x7 & n5615 ) | ( x7 & n6500 ) | ( n5615 & n6500 ) ;
  assign n13570 = ~n2331 & n8061 ;
  assign n13571 = n13569 & n13570 ;
  assign n13566 = n7692 ^ n6483 ^ n2920 ;
  assign n13567 = n13566 ^ n1565 ^ n377 ;
  assign n13568 = n13567 ^ n12482 ^ 1'b0 ;
  assign n13572 = n13571 ^ n13568 ^ n6833 ;
  assign n13576 = n4758 ^ n4055 ^ 1'b0 ;
  assign n13577 = n669 & n13576 ;
  assign n13578 = ( x160 & ~n8339 ) | ( x160 & n13577 ) | ( ~n8339 & n13577 ) ;
  assign n13573 = n2394 & n12838 ;
  assign n13574 = ( n3146 & ~n3520 ) | ( n3146 & n13573 ) | ( ~n3520 & n13573 ) ;
  assign n13575 = n13574 ^ n793 ^ 1'b0 ;
  assign n13579 = n13578 ^ n13575 ^ n2504 ;
  assign n13585 = n4322 & ~n13439 ;
  assign n13586 = ~n431 & n13585 ;
  assign n13587 = ( ~n6763 & n8247 ) | ( ~n6763 & n13586 ) | ( n8247 & n13586 ) ;
  assign n13583 = n9318 ^ n2894 ^ 1'b0 ;
  assign n13581 = n7284 ^ n5453 ^ n3698 ;
  assign n13580 = n4794 & n12767 ;
  assign n13582 = n13581 ^ n13580 ^ n1953 ;
  assign n13584 = n13583 ^ n13582 ^ n2706 ;
  assign n13588 = n13587 ^ n13584 ^ n1028 ;
  assign n13596 = ~n10153 & n11549 ;
  assign n13594 = ( n1624 & n4550 ) | ( n1624 & ~n4878 ) | ( n4550 & ~n4878 ) ;
  assign n13595 = ( n487 & ~n10068 ) | ( n487 & n13594 ) | ( ~n10068 & n13594 ) ;
  assign n13589 = n8083 ^ n7384 ^ n548 ;
  assign n13590 = n2092 | n9612 ;
  assign n13591 = n459 & ~n13590 ;
  assign n13592 = ( n8315 & ~n13589 ) | ( n8315 & n13591 ) | ( ~n13589 & n13591 ) ;
  assign n13593 = n13592 ^ n7716 ^ n1877 ;
  assign n13597 = n13596 ^ n13595 ^ n13593 ;
  assign n13598 = n2138 & ~n6378 ;
  assign n13599 = n13598 ^ n9424 ^ 1'b0 ;
  assign n13600 = n13599 ^ n3371 ^ x49 ;
  assign n13601 = n13600 ^ n3882 ^ n3708 ;
  assign n13602 = ( n2090 & n11268 ) | ( n2090 & ~n13601 ) | ( n11268 & ~n13601 ) ;
  assign n13603 = n4863 ^ n1034 ^ 1'b0 ;
  assign n13604 = n13603 ^ n10856 ^ n4358 ;
  assign n13606 = n13173 ^ n4128 ^ 1'b0 ;
  assign n13607 = n3021 & n13606 ;
  assign n13605 = ( ~n461 & n1333 ) | ( ~n461 & n8956 ) | ( n1333 & n8956 ) ;
  assign n13608 = n13607 ^ n13605 ^ n10882 ;
  assign n13624 = n5961 ^ n5908 ^ n4068 ;
  assign n13625 = n13624 ^ n4452 ^ n2520 ;
  assign n13610 = n4757 ^ n4537 ^ n2260 ;
  assign n13611 = n13610 ^ n6248 ^ n703 ;
  assign n13612 = ~n1724 & n2787 ;
  assign n13613 = ( n1147 & n10031 ) | ( n1147 & ~n13612 ) | ( n10031 & ~n13612 ) ;
  assign n13614 = n661 & n13613 ;
  assign n13615 = ( n4234 & ~n13611 ) | ( n4234 & n13614 ) | ( ~n13611 & n13614 ) ;
  assign n13609 = n11176 ^ n7331 ^ n3725 ;
  assign n13616 = n13615 ^ n13609 ^ n11332 ;
  assign n13619 = ~n1769 & n8087 ;
  assign n13620 = n4135 & n13619 ;
  assign n13617 = n12671 ^ n5904 ^ 1'b0 ;
  assign n13618 = n1306 & ~n13617 ;
  assign n13621 = n13620 ^ n13618 ^ n662 ;
  assign n13622 = ~n5893 & n13621 ;
  assign n13623 = n13616 & n13622 ;
  assign n13626 = n13625 ^ n13623 ^ n7907 ;
  assign n13627 = ( x194 & ~n3623 ) | ( x194 & n4729 ) | ( ~n3623 & n4729 ) ;
  assign n13628 = n13627 ^ n9457 ^ n2891 ;
  assign n13629 = n2536 ^ n1845 ^ n346 ;
  assign n13630 = n13629 ^ n10887 ^ n9094 ;
  assign n13631 = ( ~n4629 & n10179 ) | ( ~n4629 & n13630 ) | ( n10179 & n13630 ) ;
  assign n13634 = ( n1763 & ~n1983 ) | ( n1763 & n5639 ) | ( ~n1983 & n5639 ) ;
  assign n13635 = ( n2620 & n2892 ) | ( n2620 & n13634 ) | ( n2892 & n13634 ) ;
  assign n13636 = n13635 ^ n5162 ^ n940 ;
  assign n13637 = ( n1945 & n2185 ) | ( n1945 & ~n13636 ) | ( n2185 & ~n13636 ) ;
  assign n13632 = ( x226 & ~n952 ) | ( x226 & n1712 ) | ( ~n952 & n1712 ) ;
  assign n13633 = n1363 & n13632 ;
  assign n13638 = n13637 ^ n13633 ^ 1'b0 ;
  assign n13639 = ( n7772 & n8656 ) | ( n7772 & ~n13638 ) | ( n8656 & ~n13638 ) ;
  assign n13640 = ( n7100 & n12545 ) | ( n7100 & ~n13639 ) | ( n12545 & ~n13639 ) ;
  assign n13641 = n13640 ^ n8398 ^ n2441 ;
  assign n13642 = ~n814 & n12340 ;
  assign n13643 = n13642 ^ n1682 ^ n1652 ;
  assign n13644 = n3013 ^ n2693 ^ n1284 ;
  assign n13645 = ( n1840 & n5878 ) | ( n1840 & ~n13644 ) | ( n5878 & ~n13644 ) ;
  assign n13646 = n13645 ^ n9642 ^ n1869 ;
  assign n13647 = ( ~n5578 & n8133 ) | ( ~n5578 & n9475 ) | ( n8133 & n9475 ) ;
  assign n13648 = ~n6721 & n13525 ;
  assign n13649 = n13647 & n13648 ;
  assign n13650 = ~n746 & n13649 ;
  assign n13651 = n13021 ^ n10061 ^ n5702 ;
  assign n13652 = n1611 & n3998 ;
  assign n13653 = ~n8060 & n13652 ;
  assign n13654 = n13653 ^ n6682 ^ n5115 ;
  assign n13655 = ~n4551 & n13654 ;
  assign n13656 = n8102 ^ n4545 ^ 1'b0 ;
  assign n13663 = ( n2119 & n2681 ) | ( n2119 & n7439 ) | ( n2681 & n7439 ) ;
  assign n13664 = ( n3142 & n9606 ) | ( n3142 & n13663 ) | ( n9606 & n13663 ) ;
  assign n13657 = n1365 ^ n1103 ^ n974 ;
  assign n13658 = ( n1053 & n2977 ) | ( n1053 & ~n13657 ) | ( n2977 & ~n13657 ) ;
  assign n13659 = ~n521 & n4803 ;
  assign n13660 = n6256 & n13659 ;
  assign n13661 = n13660 ^ n2738 ^ 1'b0 ;
  assign n13662 = n13658 & ~n13661 ;
  assign n13665 = n13664 ^ n13662 ^ 1'b0 ;
  assign n13666 = n13656 & n13665 ;
  assign n13672 = n6062 ^ n3733 ^ 1'b0 ;
  assign n13673 = n4613 ^ n3579 ^ 1'b0 ;
  assign n13674 = n13673 ^ n5991 ^ 1'b0 ;
  assign n13675 = ~n13672 & n13674 ;
  assign n13676 = ( n587 & n13486 ) | ( n587 & n13675 ) | ( n13486 & n13675 ) ;
  assign n13667 = n3421 ^ n2164 ^ n1286 ;
  assign n13668 = n13667 ^ x183 ^ 1'b0 ;
  assign n13669 = ( x61 & ~x66 ) | ( x61 & n316 ) | ( ~x66 & n316 ) ;
  assign n13670 = ( n1961 & ~n7418 ) | ( n1961 & n13669 ) | ( ~n7418 & n13669 ) ;
  assign n13671 = ( n12151 & ~n13668 ) | ( n12151 & n13670 ) | ( ~n13668 & n13670 ) ;
  assign n13677 = n13676 ^ n13671 ^ n2043 ;
  assign n13678 = n9988 ^ n6565 ^ n5080 ;
  assign n13681 = n2889 & n3376 ;
  assign n13682 = n13681 ^ n4754 ^ 1'b0 ;
  assign n13683 = n1515 & n13682 ;
  assign n13679 = n7341 ^ n5701 ^ n3443 ;
  assign n13680 = n13679 ^ n9713 ^ n2404 ;
  assign n13684 = n13683 ^ n13680 ^ 1'b0 ;
  assign n13691 = n5016 & ~n5309 ;
  assign n13692 = n13691 ^ n1296 ^ 1'b0 ;
  assign n13693 = n13692 ^ n4808 ^ n662 ;
  assign n13690 = ( n1062 & n2033 ) | ( n1062 & n2704 ) | ( n2033 & n2704 ) ;
  assign n13694 = n13693 ^ n13690 ^ n7776 ;
  assign n13688 = n11111 ^ n9353 ^ n7489 ;
  assign n13689 = n13688 ^ n6226 ^ n1804 ;
  assign n13686 = n8964 ^ n3872 ^ n3309 ;
  assign n13685 = ( n6188 & n9299 ) | ( n6188 & n13295 ) | ( n9299 & n13295 ) ;
  assign n13687 = n13686 ^ n13685 ^ n3487 ;
  assign n13695 = n13694 ^ n13689 ^ n13687 ;
  assign n13700 = n535 & ~n8394 ;
  assign n13701 = n11187 & n13700 ;
  assign n13702 = n13701 ^ n12079 ^ n8637 ;
  assign n13696 = ( n3406 & n6293 ) | ( n3406 & ~n10604 ) | ( n6293 & ~n10604 ) ;
  assign n13697 = n13696 ^ n4694 ^ 1'b0 ;
  assign n13698 = n11070 & n13697 ;
  assign n13699 = n13698 ^ n1965 ^ 1'b0 ;
  assign n13703 = n13702 ^ n13699 ^ 1'b0 ;
  assign n13704 = n13703 ^ n9441 ^ n3373 ;
  assign n13705 = ~n6146 & n10618 ;
  assign n13706 = n10499 & n13705 ;
  assign n13707 = n6447 & ~n13706 ;
  assign n13708 = n7858 & n13707 ;
  assign n13709 = n13708 ^ n7777 ^ n2804 ;
  assign n13710 = n13709 ^ n13249 ^ n3074 ;
  assign n13711 = n10685 ^ n6726 ^ n4299 ;
  assign n13712 = ~n1087 & n1756 ;
  assign n13713 = n13712 ^ n6425 ^ n4661 ;
  assign n13714 = ( n412 & n3380 ) | ( n412 & n13713 ) | ( n3380 & n13713 ) ;
  assign n13715 = n13714 ^ n4509 ^ 1'b0 ;
  assign n13716 = ( n4221 & ~n6902 ) | ( n4221 & n13715 ) | ( ~n6902 & n13715 ) ;
  assign n13717 = n13063 ^ n4699 ^ n4685 ;
  assign n13718 = ( n7803 & ~n8899 ) | ( n7803 & n13717 ) | ( ~n8899 & n13717 ) ;
  assign n13719 = n5247 ^ n3318 ^ n612 ;
  assign n13720 = n628 & ~n13719 ;
  assign n13721 = ~n11301 & n13720 ;
  assign n13722 = n13721 ^ n1677 ^ 1'b0 ;
  assign n13723 = n13718 & n13722 ;
  assign n13727 = n13657 ^ n2612 ^ n773 ;
  assign n13726 = n479 | n3507 ;
  assign n13728 = n13727 ^ n13726 ^ 1'b0 ;
  assign n13725 = n2261 & n3737 ;
  assign n13724 = n2387 & ~n12185 ;
  assign n13729 = n13728 ^ n13725 ^ n13724 ;
  assign n13730 = n9223 ^ n8521 ^ n395 ;
  assign n13731 = n13730 ^ n11383 ^ n863 ;
  assign n13732 = n7511 ^ n6287 ^ n5615 ;
  assign n13734 = ~n6993 & n8984 ;
  assign n13735 = n13734 ^ n5946 ^ 1'b0 ;
  assign n13733 = ( ~n3480 & n7273 ) | ( ~n3480 & n12008 ) | ( n7273 & n12008 ) ;
  assign n13736 = n13735 ^ n13733 ^ 1'b0 ;
  assign n13737 = n13732 | n13736 ;
  assign n13738 = n11864 ^ n1444 ^ 1'b0 ;
  assign n13739 = n7394 ^ n3094 ^ 1'b0 ;
  assign n13740 = n11262 | n13739 ;
  assign n13741 = ( n5654 & n9974 ) | ( n5654 & n13740 ) | ( n9974 & n13740 ) ;
  assign n13742 = n13741 ^ n7929 ^ n7674 ;
  assign n13743 = n615 ^ x153 ^ 1'b0 ;
  assign n13744 = ~n5034 & n13743 ;
  assign n13745 = ( n1390 & n1756 ) | ( n1390 & ~n7796 ) | ( n1756 & ~n7796 ) ;
  assign n13746 = ( n2297 & n3722 ) | ( n2297 & ~n13745 ) | ( n3722 & ~n13745 ) ;
  assign n13747 = ( n4961 & ~n8609 ) | ( n4961 & n9681 ) | ( ~n8609 & n9681 ) ;
  assign n13748 = n13747 ^ n2805 ^ n1710 ;
  assign n13749 = ( ~n13744 & n13746 ) | ( ~n13744 & n13748 ) | ( n13746 & n13748 ) ;
  assign n13757 = n12533 ^ n5722 ^ n1873 ;
  assign n13755 = ( ~n407 & n956 ) | ( ~n407 & n6537 ) | ( n956 & n6537 ) ;
  assign n13756 = n13755 ^ n4252 ^ n2818 ;
  assign n13758 = n13757 ^ n13756 ^ n4560 ;
  assign n13759 = ( ~n5260 & n13556 ) | ( ~n5260 & n13758 ) | ( n13556 & n13758 ) ;
  assign n13751 = n2809 & ~n2862 ;
  assign n13752 = n8483 & n13751 ;
  assign n13750 = n9694 ^ n5926 ^ n908 ;
  assign n13753 = n13752 ^ n13750 ^ n5166 ;
  assign n13754 = n13753 ^ n4464 ^ n371 ;
  assign n13760 = n13759 ^ n13754 ^ 1'b0 ;
  assign n13761 = n13749 & ~n13760 ;
  assign n13762 = n9974 ^ n6364 ^ n1606 ;
  assign n13767 = n3056 ^ n959 ^ x244 ;
  assign n13763 = n9958 ^ n9692 ^ n4980 ;
  assign n13764 = n7474 & n13763 ;
  assign n13765 = ~n7427 & n13764 ;
  assign n13766 = ( n1281 & n4219 ) | ( n1281 & n13765 ) | ( n4219 & n13765 ) ;
  assign n13768 = n13767 ^ n13766 ^ n8747 ;
  assign n13769 = ~n6544 & n10659 ;
  assign n13770 = ( n3530 & n3727 ) | ( n3530 & n12238 ) | ( n3727 & n12238 ) ;
  assign n13771 = n13770 ^ n8084 ^ n7605 ;
  assign n13772 = ( n4236 & n4765 ) | ( n4236 & n11885 ) | ( n4765 & n11885 ) ;
  assign n13773 = ( n7327 & n10303 ) | ( n7327 & n13772 ) | ( n10303 & n13772 ) ;
  assign n13774 = ( n1925 & n5749 ) | ( n1925 & n7371 ) | ( n5749 & n7371 ) ;
  assign n13780 = ( n871 & n3908 ) | ( n871 & ~n6297 ) | ( n3908 & ~n6297 ) ;
  assign n13781 = n13780 ^ n10245 ^ n7309 ;
  assign n13776 = n2979 ^ n1285 ^ n561 ;
  assign n13777 = ( n3811 & n4230 ) | ( n3811 & ~n13776 ) | ( n4230 & ~n13776 ) ;
  assign n13778 = ( n1186 & ~n11178 ) | ( n1186 & n13777 ) | ( ~n11178 & n13777 ) ;
  assign n13775 = ( n5539 & ~n7453 ) | ( n5539 & n12695 ) | ( ~n7453 & n12695 ) ;
  assign n13779 = n13778 ^ n13775 ^ n13603 ;
  assign n13782 = n13781 ^ n13779 ^ n6550 ;
  assign n13784 = n8542 | n12256 ;
  assign n13785 = n9980 & ~n13784 ;
  assign n13786 = n8115 ^ n4030 ^ 1'b0 ;
  assign n13787 = n13785 | n13786 ;
  assign n13783 = n9569 ^ n7684 ^ n463 ;
  assign n13788 = n13787 ^ n13783 ^ x227 ;
  assign n13789 = x69 & n12591 ;
  assign n13790 = ~x235 & n13789 ;
  assign n13791 = n13790 ^ n8444 ^ n5258 ;
  assign n13793 = n5325 ^ n3404 ^ x247 ;
  assign n13794 = ( ~n4885 & n6450 ) | ( ~n4885 & n13793 ) | ( n6450 & n13793 ) ;
  assign n13795 = ( n6123 & n11589 ) | ( n6123 & n13794 ) | ( n11589 & n13794 ) ;
  assign n13796 = n13795 ^ n8049 ^ n6180 ;
  assign n13792 = n7672 ^ n2891 ^ 1'b0 ;
  assign n13797 = n13796 ^ n13792 ^ n11977 ;
  assign n13801 = n6576 ^ n3712 ^ 1'b0 ;
  assign n13802 = n324 & n13801 ;
  assign n13800 = n10873 ^ n7796 ^ n4468 ;
  assign n13803 = n13802 ^ n13800 ^ n1256 ;
  assign n13804 = n13803 ^ n7181 ^ n888 ;
  assign n13805 = n12073 & ~n13804 ;
  assign n13806 = n13805 ^ n1236 ^ 1'b0 ;
  assign n13798 = ( n4330 & n8253 ) | ( n4330 & ~n12487 ) | ( n8253 & ~n12487 ) ;
  assign n13799 = ( n9305 & n10742 ) | ( n9305 & n13798 ) | ( n10742 & n13798 ) ;
  assign n13807 = n13806 ^ n13799 ^ n10056 ;
  assign n13808 = ( n4158 & n6503 ) | ( n4158 & ~n6509 ) | ( n6503 & ~n6509 ) ;
  assign n13809 = n9375 ^ n4282 ^ n2830 ;
  assign n13810 = n13809 ^ n12059 ^ n6763 ;
  assign n13811 = n776 & ~n1116 ;
  assign n13812 = n4066 & n13811 ;
  assign n13813 = n13812 ^ n6228 ^ n3061 ;
  assign n13814 = n1745 ^ n1471 ^ 1'b0 ;
  assign n13815 = n3026 & n13814 ;
  assign n13816 = ( n7957 & n8613 ) | ( n7957 & n13815 ) | ( n8613 & n13815 ) ;
  assign n13817 = n8538 ^ n7946 ^ n3050 ;
  assign n13818 = n3824 ^ n3190 ^ 1'b0 ;
  assign n13819 = n13818 ^ n8389 ^ n1557 ;
  assign n13822 = n3824 ^ n2783 ^ 1'b0 ;
  assign n13823 = ( n1902 & ~n4537 ) | ( n1902 & n9641 ) | ( ~n4537 & n9641 ) ;
  assign n13824 = n4749 | n13823 ;
  assign n13825 = n7322 ^ n6922 ^ n3549 ;
  assign n13826 = ( n6977 & n12142 ) | ( n6977 & n13825 ) | ( n12142 & n13825 ) ;
  assign n13827 = n13826 ^ n9917 ^ 1'b0 ;
  assign n13828 = ~n13824 & n13827 ;
  assign n13829 = ( n4122 & n13822 ) | ( n4122 & ~n13828 ) | ( n13822 & ~n13828 ) ;
  assign n13820 = n5730 ^ n3053 ^ n721 ;
  assign n13821 = n10546 | n13820 ;
  assign n13830 = n13829 ^ n13821 ^ 1'b0 ;
  assign n13831 = n10209 ^ n7145 ^ n2851 ;
  assign n13832 = n13831 ^ n12827 ^ 1'b0 ;
  assign n13833 = n1266 | n13832 ;
  assign n13834 = n13833 ^ n7564 ^ 1'b0 ;
  assign n13835 = ( ~n6287 & n7797 ) | ( ~n6287 & n12203 ) | ( n7797 & n12203 ) ;
  assign n13836 = n13835 ^ n4504 ^ 1'b0 ;
  assign n13837 = n5834 & n13836 ;
  assign n13838 = ( n755 & n1040 ) | ( n755 & ~n1362 ) | ( n1040 & ~n1362 ) ;
  assign n13839 = ( n2379 & ~n12578 ) | ( n2379 & n13838 ) | ( ~n12578 & n13838 ) ;
  assign n13840 = n4307 ^ n805 ^ 1'b0 ;
  assign n13841 = n13415 & ~n13840 ;
  assign n13842 = n13841 ^ n7084 ^ 1'b0 ;
  assign n13843 = n4431 & ~n12417 ;
  assign n13844 = ( n1066 & ~n4618 ) | ( n1066 & n13843 ) | ( ~n4618 & n13843 ) ;
  assign n13845 = ( n4204 & n13842 ) | ( n4204 & ~n13844 ) | ( n13842 & ~n13844 ) ;
  assign n13846 = ( n1814 & n13839 ) | ( n1814 & ~n13845 ) | ( n13839 & ~n13845 ) ;
  assign n13847 = ( ~n1522 & n7867 ) | ( ~n1522 & n8080 ) | ( n7867 & n8080 ) ;
  assign n13848 = n8746 & ~n13847 ;
  assign n13849 = ( n496 & n4599 ) | ( n496 & ~n13848 ) | ( n4599 & ~n13848 ) ;
  assign n13850 = ( n4655 & n6846 ) | ( n4655 & ~n9521 ) | ( n6846 & ~n9521 ) ;
  assign n13851 = n10435 ^ n6417 ^ n3846 ;
  assign n13852 = n5021 & n13851 ;
  assign n13853 = n13852 ^ n10057 ^ 1'b0 ;
  assign n13854 = n5204 & ~n13853 ;
  assign n13855 = n7921 ^ n7891 ^ n1278 ;
  assign n13859 = n1110 & n2343 ;
  assign n13860 = n13859 ^ n4004 ^ 1'b0 ;
  assign n13857 = n6438 ^ n1229 ^ n793 ;
  assign n13856 = ( n3007 & n3300 ) | ( n3007 & ~n11095 ) | ( n3300 & ~n11095 ) ;
  assign n13858 = n13857 ^ n13856 ^ n1024 ;
  assign n13861 = n13860 ^ n13858 ^ n5200 ;
  assign n13862 = ( n8687 & n9589 ) | ( n8687 & n13861 ) | ( n9589 & n13861 ) ;
  assign n13863 = n13380 ^ n3813 ^ n334 ;
  assign n13864 = n13863 ^ n5234 ^ 1'b0 ;
  assign n13865 = n5213 | n13864 ;
  assign n13866 = ( n4404 & n10616 ) | ( n4404 & n13865 ) | ( n10616 & n13865 ) ;
  assign n13867 = n2830 ^ n751 ^ n572 ;
  assign n13868 = n10202 ^ n9220 ^ 1'b0 ;
  assign n13869 = ~n13867 & n13868 ;
  assign n13870 = ~n11403 & n13869 ;
  assign n13871 = n1055 & n13870 ;
  assign n13872 = ~n6047 & n11134 ;
  assign n13873 = ~n10996 & n13872 ;
  assign n13874 = ( n6991 & ~n11079 ) | ( n6991 & n13873 ) | ( ~n11079 & n13873 ) ;
  assign n13875 = ( n1694 & n2316 ) | ( n1694 & ~n6212 ) | ( n2316 & ~n6212 ) ;
  assign n13876 = n8006 & n13875 ;
  assign n13880 = n2159 | n5967 ;
  assign n13881 = n13880 ^ n4075 ^ n2015 ;
  assign n13878 = ( ~n2300 & n3134 ) | ( ~n2300 & n10161 ) | ( n3134 & n10161 ) ;
  assign n13877 = n10089 ^ n4285 ^ n2383 ;
  assign n13879 = n13878 ^ n13877 ^ n7832 ;
  assign n13882 = n13881 ^ n13879 ^ n6275 ;
  assign n13883 = n3681 ^ n818 ^ 1'b0 ;
  assign n13884 = n9162 | n13883 ;
  assign n13885 = ( n10392 & n12751 ) | ( n10392 & ~n13884 ) | ( n12751 & ~n13884 ) ;
  assign n13886 = ( ~n9272 & n13882 ) | ( ~n9272 & n13885 ) | ( n13882 & n13885 ) ;
  assign n13889 = n9202 ^ n3732 ^ n1703 ;
  assign n13890 = ( n3991 & ~n5922 ) | ( n3991 & n13889 ) | ( ~n5922 & n13889 ) ;
  assign n13887 = ( n2439 & n4530 ) | ( n2439 & ~n8145 ) | ( n4530 & ~n8145 ) ;
  assign n13888 = n13887 ^ n12721 ^ 1'b0 ;
  assign n13891 = n13890 ^ n13888 ^ n7443 ;
  assign n13892 = n10617 ^ n10017 ^ 1'b0 ;
  assign n13893 = n6639 ^ n5693 ^ n2406 ;
  assign n13894 = n3913 ^ n3148 ^ 1'b0 ;
  assign n13895 = ~n3504 & n12005 ;
  assign n13896 = n13895 ^ n9676 ^ 1'b0 ;
  assign n13897 = ( n4150 & n5401 ) | ( n4150 & ~n13896 ) | ( n5401 & ~n13896 ) ;
  assign n13898 = n13897 ^ n12141 ^ n9042 ;
  assign n13899 = n399 | n1299 ;
  assign n13900 = n4764 | n13899 ;
  assign n13901 = ( ~n13894 & n13898 ) | ( ~n13894 & n13900 ) | ( n13898 & n13900 ) ;
  assign n13906 = ( n533 & n1030 ) | ( n533 & ~n2316 ) | ( n1030 & ~n2316 ) ;
  assign n13905 = n2897 & n7371 ;
  assign n13902 = n1509 | n2209 ;
  assign n13903 = n13902 ^ n2799 ^ n2585 ;
  assign n13904 = n13903 ^ n10378 ^ n6783 ;
  assign n13907 = n13906 ^ n13905 ^ n13904 ;
  assign n13908 = n3525 ^ n2258 ^ n1614 ;
  assign n13909 = n13908 ^ n7217 ^ n2731 ;
  assign n13910 = ( n2420 & n4109 ) | ( n2420 & ~n13909 ) | ( n4109 & ~n13909 ) ;
  assign n13914 = n3001 ^ n2232 ^ n593 ;
  assign n13911 = n747 & ~n10347 ;
  assign n13912 = n3134 & n13911 ;
  assign n13913 = ( n1344 & ~n6681 ) | ( n1344 & n13912 ) | ( ~n6681 & n13912 ) ;
  assign n13915 = n13914 ^ n13913 ^ 1'b0 ;
  assign n13916 = ( n8650 & n10736 ) | ( n8650 & n12910 ) | ( n10736 & n12910 ) ;
  assign n13917 = ~n8113 & n9758 ;
  assign n13918 = ~n6938 & n13917 ;
  assign n13919 = n13918 ^ n6249 ^ n644 ;
  assign n13920 = ( n12213 & n12868 ) | ( n12213 & n13919 ) | ( n12868 & n13919 ) ;
  assign n13921 = n1137 & n1231 ;
  assign n13928 = ( n1989 & n6177 ) | ( n1989 & ~n12695 ) | ( n6177 & ~n12695 ) ;
  assign n13929 = ( x120 & n7660 ) | ( x120 & ~n13928 ) | ( n7660 & ~n13928 ) ;
  assign n13930 = ( ~n10264 & n10806 ) | ( ~n10264 & n13929 ) | ( n10806 & n13929 ) ;
  assign n13923 = n5923 & n10504 ;
  assign n13922 = x176 & n6042 ;
  assign n13924 = n13923 ^ n13922 ^ 1'b0 ;
  assign n13925 = ( ~n1785 & n2883 ) | ( ~n1785 & n5301 ) | ( n2883 & n5301 ) ;
  assign n13926 = n13925 ^ n7603 ^ n580 ;
  assign n13927 = n13924 & ~n13926 ;
  assign n13931 = n13930 ^ n13927 ^ 1'b0 ;
  assign n13932 = n13921 & n13931 ;
  assign n13933 = n13932 ^ n1337 ^ 1'b0 ;
  assign n13934 = n13933 ^ n4773 ^ 1'b0 ;
  assign n13935 = n13558 ^ n10505 ^ n8384 ;
  assign n13936 = n3838 & ~n13167 ;
  assign n13937 = ( n1165 & n13935 ) | ( n1165 & n13936 ) | ( n13935 & n13936 ) ;
  assign n13941 = n11511 ^ n6108 ^ 1'b0 ;
  assign n13942 = n13941 ^ n6146 ^ n1093 ;
  assign n13943 = ~n4141 & n13942 ;
  assign n13938 = n2909 ^ n1765 ^ n582 ;
  assign n13939 = ( ~n1302 & n10442 ) | ( ~n1302 & n13938 ) | ( n10442 & n13938 ) ;
  assign n13940 = n13939 ^ n7990 ^ n744 ;
  assign n13944 = n13943 ^ n13940 ^ n4060 ;
  assign n13945 = ( ~n1102 & n1724 ) | ( ~n1102 & n8805 ) | ( n1724 & n8805 ) ;
  assign n13946 = ( n1389 & n7857 ) | ( n1389 & n10421 ) | ( n7857 & n10421 ) ;
  assign n13947 = ( n1945 & n3182 ) | ( n1945 & n8736 ) | ( n3182 & n8736 ) ;
  assign n13948 = ( n2721 & n6526 ) | ( n2721 & ~n13947 ) | ( n6526 & ~n13947 ) ;
  assign n13949 = ~n2238 & n13948 ;
  assign n13950 = n13946 & n13949 ;
  assign n13951 = n4685 ^ n2083 ^ 1'b0 ;
  assign n13952 = n10196 ^ n8839 ^ n2231 ;
  assign n13953 = n13952 ^ n8463 ^ n7578 ;
  assign n13954 = ( n1324 & n10887 ) | ( n1324 & n13953 ) | ( n10887 & n13953 ) ;
  assign n13955 = ( n7379 & n13951 ) | ( n7379 & n13954 ) | ( n13951 & n13954 ) ;
  assign n13956 = ( ~n3463 & n13950 ) | ( ~n3463 & n13955 ) | ( n13950 & n13955 ) ;
  assign n13958 = n6554 ^ n2124 ^ 1'b0 ;
  assign n13957 = n980 & n10704 ;
  assign n13959 = n13958 ^ n13957 ^ n11413 ;
  assign n13960 = n4251 ^ n1269 ^ n660 ;
  assign n13961 = ( n340 & ~n6986 ) | ( n340 & n13960 ) | ( ~n6986 & n13960 ) ;
  assign n13962 = n1975 & ~n13961 ;
  assign n13963 = n13962 ^ n6521 ^ 1'b0 ;
  assign n13964 = ( n2323 & ~n5718 ) | ( n2323 & n13963 ) | ( ~n5718 & n13963 ) ;
  assign n13965 = ( n1477 & n2356 ) | ( n1477 & n2656 ) | ( n2356 & n2656 ) ;
  assign n13966 = n13965 ^ n9962 ^ n2103 ;
  assign n13967 = n13966 ^ n6062 ^ n1094 ;
  assign n13968 = n12827 ^ n12695 ^ n9348 ;
  assign n13969 = ( n1213 & n8454 ) | ( n1213 & n13968 ) | ( n8454 & n13968 ) ;
  assign n13970 = ( n10313 & ~n13967 ) | ( n10313 & n13969 ) | ( ~n13967 & n13969 ) ;
  assign n13971 = n12374 ^ n5217 ^ n369 ;
  assign n13972 = n13971 ^ n8679 ^ n5048 ;
  assign n13973 = ( ~n1398 & n3788 ) | ( ~n1398 & n10673 ) | ( n3788 & n10673 ) ;
  assign n13974 = ( x26 & n11299 ) | ( x26 & ~n13973 ) | ( n11299 & ~n13973 ) ;
  assign n13975 = ( n2664 & n5396 ) | ( n2664 & n12695 ) | ( n5396 & n12695 ) ;
  assign n13976 = ( n2804 & n6654 ) | ( n2804 & n13975 ) | ( n6654 & n13975 ) ;
  assign n13977 = n13976 ^ n2946 ^ n2482 ;
  assign n13978 = ( n2036 & n13974 ) | ( n2036 & n13977 ) | ( n13974 & n13977 ) ;
  assign n13979 = ( n3609 & n9350 ) | ( n3609 & ~n13191 ) | ( n9350 & ~n13191 ) ;
  assign n13980 = ( ~n904 & n13114 ) | ( ~n904 & n13230 ) | ( n13114 & n13230 ) ;
  assign n13981 = ( n3116 & ~n5657 ) | ( n3116 & n13980 ) | ( ~n5657 & n13980 ) ;
  assign n13983 = n5131 ^ n4577 ^ x42 ;
  assign n13984 = n1372 & n13983 ;
  assign n13985 = ( ~n5296 & n13148 ) | ( ~n5296 & n13984 ) | ( n13148 & n13984 ) ;
  assign n13982 = n12031 ^ n10366 ^ n3629 ;
  assign n13986 = n13985 ^ n13982 ^ 1'b0 ;
  assign n13991 = n2458 & ~n9589 ;
  assign n13992 = n13991 ^ n12573 ^ n4002 ;
  assign n13987 = n11387 ^ n10183 ^ n6500 ;
  assign n13988 = ( n7373 & ~n10328 ) | ( n7373 & n10696 ) | ( ~n10328 & n10696 ) ;
  assign n13989 = n13988 ^ n5794 ^ n5108 ;
  assign n13990 = n13987 & n13989 ;
  assign n13993 = n13992 ^ n13990 ^ 1'b0 ;
  assign n13994 = n3969 ^ n3938 ^ n3701 ;
  assign n13995 = n5472 ^ n1144 ^ 1'b0 ;
  assign n13996 = ( n7462 & ~n8580 ) | ( n7462 & n13995 ) | ( ~n8580 & n13995 ) ;
  assign n13997 = n13996 ^ n7507 ^ n1827 ;
  assign n13998 = ( n13029 & n13994 ) | ( n13029 & n13997 ) | ( n13994 & n13997 ) ;
  assign n13999 = ( n1085 & n8913 ) | ( n1085 & ~n13998 ) | ( n8913 & ~n13998 ) ;
  assign n14000 = ( x182 & n4946 ) | ( x182 & n5629 ) | ( n4946 & n5629 ) ;
  assign n14001 = ( n1916 & ~n12853 ) | ( n1916 & n14000 ) | ( ~n12853 & n14000 ) ;
  assign n14002 = n9030 ^ n4181 ^ n1180 ;
  assign n14003 = n7815 ^ n7013 ^ n3672 ;
  assign n14004 = n14003 ^ n8750 ^ n8700 ;
  assign n14005 = ( n10451 & n14002 ) | ( n10451 & n14004 ) | ( n14002 & n14004 ) ;
  assign n14007 = ( n427 & n1599 ) | ( n427 & n2967 ) | ( n1599 & n2967 ) ;
  assign n14008 = ( ~n2453 & n10881 ) | ( ~n2453 & n14007 ) | ( n10881 & n14007 ) ;
  assign n14006 = ( ~n5964 & n6136 ) | ( ~n5964 & n9188 ) | ( n6136 & n9188 ) ;
  assign n14009 = n14008 ^ n14006 ^ n331 ;
  assign n14010 = ( ~n2870 & n4376 ) | ( ~n2870 & n5194 ) | ( n4376 & n5194 ) ;
  assign n14011 = n2814 ^ n2219 ^ 1'b0 ;
  assign n14012 = n1492 | n14011 ;
  assign n14013 = ( ~n5076 & n10504 ) | ( ~n5076 & n14012 ) | ( n10504 & n14012 ) ;
  assign n14014 = n14013 ^ n7003 ^ n6084 ;
  assign n14015 = n9602 ^ n9521 ^ n6432 ;
  assign n14016 = n6723 ^ n2499 ^ 1'b0 ;
  assign n14017 = ( ~n1896 & n3799 ) | ( ~n1896 & n7845 ) | ( n3799 & n7845 ) ;
  assign n14018 = n14017 ^ n11678 ^ n4858 ;
  assign n14019 = ( n9732 & n14016 ) | ( n9732 & ~n14018 ) | ( n14016 & ~n14018 ) ;
  assign n14020 = n6845 & ~n9616 ;
  assign n14021 = ~n12833 & n14020 ;
  assign n14022 = ~n1510 & n8888 ;
  assign n14023 = ( n9539 & n14021 ) | ( n9539 & ~n14022 ) | ( n14021 & ~n14022 ) ;
  assign n14024 = ( n831 & n13897 ) | ( n831 & n14023 ) | ( n13897 & n14023 ) ;
  assign n14027 = ~n2871 & n9381 ;
  assign n14025 = n5147 ^ n2560 ^ 1'b0 ;
  assign n14026 = ( n8285 & n11609 ) | ( n8285 & n14025 ) | ( n11609 & n14025 ) ;
  assign n14028 = n14027 ^ n14026 ^ n13286 ;
  assign n14029 = n13340 ^ n7676 ^ n6835 ;
  assign n14030 = n10828 ^ n2237 ^ 1'b0 ;
  assign n14031 = ~n14029 & n14030 ;
  assign n14032 = n2395 ^ n2358 ^ n1462 ;
  assign n14033 = ( ~n5056 & n5542 ) | ( ~n5056 & n14032 ) | ( n5542 & n14032 ) ;
  assign n14034 = ( n2985 & ~n6180 ) | ( n2985 & n14033 ) | ( ~n6180 & n14033 ) ;
  assign n14035 = n8365 | n14034 ;
  assign n14036 = n10961 & ~n14035 ;
  assign n14037 = n14036 ^ n10117 ^ n3004 ;
  assign n14038 = ( n1624 & n3122 ) | ( n1624 & n8652 ) | ( n3122 & n8652 ) ;
  assign n14039 = ( n890 & ~n2065 ) | ( n890 & n14038 ) | ( ~n2065 & n14038 ) ;
  assign n14040 = ~n739 & n14039 ;
  assign n14041 = n7082 & n14040 ;
  assign n14042 = ( n1959 & n6828 ) | ( n1959 & n14041 ) | ( n6828 & n14041 ) ;
  assign n14043 = n14042 ^ n10626 ^ n337 ;
  assign n14044 = n7141 ^ n4626 ^ n2435 ;
  assign n14045 = n5172 & ~n14044 ;
  assign n14046 = n14045 ^ n7589 ^ 1'b0 ;
  assign n14047 = ~n5161 & n9360 ;
  assign n14048 = n14047 ^ n12835 ^ 1'b0 ;
  assign n14049 = n14048 ^ n6835 ^ 1'b0 ;
  assign n14050 = n1303 & n14049 ;
  assign n14051 = ( n4142 & n13014 ) | ( n4142 & n14050 ) | ( n13014 & n14050 ) ;
  assign n14052 = ~n2312 & n6473 ;
  assign n14053 = ( ~n14046 & n14051 ) | ( ~n14046 & n14052 ) | ( n14051 & n14052 ) ;
  assign n14056 = n3377 ^ n1418 ^ 1'b0 ;
  assign n14057 = ~n11486 & n14056 ;
  assign n14058 = ( n2814 & n6675 ) | ( n2814 & n14057 ) | ( n6675 & n14057 ) ;
  assign n14054 = n1049 & n4113 ;
  assign n14055 = n14054 ^ n4004 ^ 1'b0 ;
  assign n14059 = n14058 ^ n14055 ^ n6349 ;
  assign n14060 = ~n10570 & n12614 ;
  assign n14061 = n14060 ^ n6589 ^ 1'b0 ;
  assign n14062 = ( n8138 & n13406 ) | ( n8138 & ~n14061 ) | ( n13406 & ~n14061 ) ;
  assign n14063 = n14062 ^ n12136 ^ 1'b0 ;
  assign n14064 = n8161 ^ n6813 ^ 1'b0 ;
  assign n14065 = n14064 ^ n3738 ^ 1'b0 ;
  assign n14066 = ( n2629 & ~n7729 ) | ( n2629 & n9631 ) | ( ~n7729 & n9631 ) ;
  assign n14067 = n14066 ^ n5794 ^ 1'b0 ;
  assign n14068 = n14065 & n14067 ;
  assign n14069 = n3835 & ~n13128 ;
  assign n14070 = n12839 ^ n6961 ^ n1530 ;
  assign n14071 = n14069 & ~n14070 ;
  assign n14072 = n14071 ^ n9809 ^ 1'b0 ;
  assign n14073 = n2628 & n3918 ;
  assign n14074 = ( n4103 & n9230 ) | ( n4103 & n14073 ) | ( n9230 & n14073 ) ;
  assign n14077 = ~n7194 & n7217 ;
  assign n14078 = n14077 ^ n4700 ^ 1'b0 ;
  assign n14075 = n5762 ^ n1571 ^ n612 ;
  assign n14076 = n14075 ^ n6659 ^ 1'b0 ;
  assign n14079 = n14078 ^ n14076 ^ n12334 ;
  assign n14082 = ( ~n3857 & n6024 ) | ( ~n3857 & n6592 ) | ( n6024 & n6592 ) ;
  assign n14083 = ( ~n1075 & n5772 ) | ( ~n1075 & n14082 ) | ( n5772 & n14082 ) ;
  assign n14084 = n14083 ^ n8957 ^ n620 ;
  assign n14080 = n2339 | n4105 ;
  assign n14081 = n13216 & ~n14080 ;
  assign n14085 = n14084 ^ n14081 ^ 1'b0 ;
  assign n14086 = n2912 & ~n14085 ;
  assign n14087 = n9666 ^ n392 ^ n313 ;
  assign n14088 = n14087 ^ n12769 ^ n3211 ;
  assign n14089 = n14088 ^ n3004 ^ x114 ;
  assign n14090 = n8813 ^ n783 ^ 1'b0 ;
  assign n14091 = ~n5200 & n11889 ;
  assign n14092 = n6958 ^ n2191 ^ n1825 ;
  assign n14093 = n14092 ^ n12346 ^ n6094 ;
  assign n14094 = n6062 & n6365 ;
  assign n14095 = n14094 ^ n12109 ^ n2112 ;
  assign n14100 = n3012 & ~n7780 ;
  assign n14101 = n14100 ^ n2501 ^ 1'b0 ;
  assign n14096 = n3579 & n3847 ;
  assign n14097 = ~n8698 & n14096 ;
  assign n14098 = n14097 ^ n2948 ^ 1'b0 ;
  assign n14099 = n14098 ^ n8397 ^ n2400 ;
  assign n14102 = n14101 ^ n14099 ^ x204 ;
  assign n14103 = n7293 ^ n3484 ^ 1'b0 ;
  assign n14104 = n8048 | n14103 ;
  assign n14105 = n3898 | n13213 ;
  assign n14106 = n14104 & ~n14105 ;
  assign n14107 = n11696 ^ n4388 ^ n2363 ;
  assign n14108 = n3750 & ~n14107 ;
  assign n14109 = n9540 & n14108 ;
  assign n14110 = ~n4576 & n11126 ;
  assign n14111 = n14109 & n14110 ;
  assign n14112 = n14111 ^ n11921 ^ n1118 ;
  assign n14113 = ( ~n2977 & n8617 ) | ( ~n2977 & n12792 ) | ( n8617 & n12792 ) ;
  assign n14114 = n10358 ^ n5183 ^ n1280 ;
  assign n14115 = n2068 ^ n296 ^ 1'b0 ;
  assign n14116 = n14114 & ~n14115 ;
  assign n14117 = n2731 & n14116 ;
  assign n14118 = ( ~n3222 & n10514 ) | ( ~n3222 & n14117 ) | ( n10514 & n14117 ) ;
  assign n14119 = n838 & ~n14118 ;
  assign n14120 = n14119 ^ n12314 ^ 1'b0 ;
  assign n14121 = n5907 ^ n5064 ^ n451 ;
  assign n14122 = ( n2271 & n7771 ) | ( n2271 & n14121 ) | ( n7771 & n14121 ) ;
  assign n14123 = ( ~n9454 & n12115 ) | ( ~n9454 & n14122 ) | ( n12115 & n14122 ) ;
  assign n14124 = ( n4863 & ~n6601 ) | ( n4863 & n8607 ) | ( ~n6601 & n8607 ) ;
  assign n14125 = n14124 ^ n9714 ^ n7752 ;
  assign n14126 = ( n8359 & n14123 ) | ( n8359 & n14125 ) | ( n14123 & n14125 ) ;
  assign n14127 = n3536 & n11303 ;
  assign n14128 = n3305 | n5309 ;
  assign n14129 = n12219 & ~n14128 ;
  assign n14130 = n14129 ^ n8123 ^ 1'b0 ;
  assign n14131 = n14130 ^ n6546 ^ n5744 ;
  assign n14132 = ~n3358 & n9760 ;
  assign n14133 = ~n7801 & n14132 ;
  assign n14134 = n14133 ^ n13280 ^ n5537 ;
  assign n14135 = n8046 ^ n4337 ^ n554 ;
  assign n14136 = ( ~n700 & n5688 ) | ( ~n700 & n12419 ) | ( n5688 & n12419 ) ;
  assign n14137 = ( x135 & n1797 ) | ( x135 & n10435 ) | ( n1797 & n10435 ) ;
  assign n14138 = ( n3828 & ~n9714 ) | ( n3828 & n13030 ) | ( ~n9714 & n13030 ) ;
  assign n14139 = ( n14136 & ~n14137 ) | ( n14136 & n14138 ) | ( ~n14137 & n14138 ) ;
  assign n14142 = ~n3879 & n9206 ;
  assign n14143 = n14142 ^ n3560 ^ 1'b0 ;
  assign n14140 = ( n9491 & ~n10429 ) | ( n9491 & n13835 ) | ( ~n10429 & n13835 ) ;
  assign n14141 = ( n402 & n10328 ) | ( n402 & ~n14140 ) | ( n10328 & ~n14140 ) ;
  assign n14144 = n14143 ^ n14141 ^ x97 ;
  assign n14147 = n8922 ^ n2804 ^ n1635 ;
  assign n14145 = ( n5279 & ~n6266 ) | ( n5279 & n8682 ) | ( ~n6266 & n8682 ) ;
  assign n14146 = n5811 & ~n14145 ;
  assign n14148 = n14147 ^ n14146 ^ 1'b0 ;
  assign n14149 = n14148 ^ n12896 ^ n5572 ;
  assign n14152 = n2631 ^ n1691 ^ 1'b0 ;
  assign n14153 = n14152 ^ n9898 ^ n8008 ;
  assign n14154 = n1525 ^ n1316 ^ 1'b0 ;
  assign n14155 = n6641 | n14154 ;
  assign n14156 = ( n8581 & n14153 ) | ( n8581 & ~n14155 ) | ( n14153 & ~n14155 ) ;
  assign n14150 = n7269 & n7644 ;
  assign n14151 = ( n8270 & n13472 ) | ( n8270 & ~n14150 ) | ( n13472 & ~n14150 ) ;
  assign n14157 = n14156 ^ n14151 ^ n8059 ;
  assign n14158 = ( ~n2358 & n3093 ) | ( ~n2358 & n12596 ) | ( n3093 & n12596 ) ;
  assign n14159 = ( ~n1001 & n4394 ) | ( ~n1001 & n6221 ) | ( n4394 & n6221 ) ;
  assign n14160 = n14159 ^ n5998 ^ 1'b0 ;
  assign n14163 = n1659 | n9510 ;
  assign n14164 = n2952 & ~n14163 ;
  assign n14165 = n7371 ^ n2102 ^ n1965 ;
  assign n14166 = ( n5238 & ~n14164 ) | ( n5238 & n14165 ) | ( ~n14164 & n14165 ) ;
  assign n14161 = n3128 ^ n2704 ^ n356 ;
  assign n14162 = n14161 ^ n2454 ^ n1954 ;
  assign n14167 = n14166 ^ n14162 ^ n3311 ;
  assign n14168 = ~n11989 & n14167 ;
  assign n14169 = n14160 & n14168 ;
  assign n14170 = n13627 ^ n11141 ^ n6074 ;
  assign n14171 = n14170 ^ n9221 ^ n8286 ;
  assign n14172 = n11350 ^ n10284 ^ n3375 ;
  assign n14173 = ( n6665 & n10629 ) | ( n6665 & ~n14172 ) | ( n10629 & ~n14172 ) ;
  assign n14174 = n901 | n3939 ;
  assign n14175 = ( x191 & ~n4640 ) | ( x191 & n14174 ) | ( ~n4640 & n14174 ) ;
  assign n14176 = ( n3284 & n5893 ) | ( n3284 & ~n14175 ) | ( n5893 & ~n14175 ) ;
  assign n14177 = ~n13223 & n14176 ;
  assign n14178 = n6530 & n14177 ;
  assign n14186 = n4747 ^ n3957 ^ n2729 ;
  assign n14183 = ( n997 & n3639 ) | ( n997 & n4026 ) | ( n3639 & n4026 ) ;
  assign n14184 = ( n1662 & ~n6788 ) | ( n1662 & n13500 ) | ( ~n6788 & n13500 ) ;
  assign n14185 = ( n1049 & n14183 ) | ( n1049 & n14184 ) | ( n14183 & n14184 ) ;
  assign n14181 = ( n434 & n8260 ) | ( n434 & ~n9085 ) | ( n8260 & ~n9085 ) ;
  assign n14182 = n4735 & n14181 ;
  assign n14187 = n14186 ^ n14185 ^ n14182 ;
  assign n14179 = ( ~n760 & n4293 ) | ( ~n760 & n7667 ) | ( n4293 & n7667 ) ;
  assign n14180 = n14179 ^ n9743 ^ n5216 ;
  assign n14188 = n14187 ^ n14180 ^ n10760 ;
  assign n14189 = ( n3679 & n11525 ) | ( n3679 & ~n13433 ) | ( n11525 & ~n13433 ) ;
  assign n14190 = ( ~n2303 & n4941 ) | ( ~n2303 & n8309 ) | ( n4941 & n8309 ) ;
  assign n14191 = ( n701 & n5335 ) | ( n701 & n14190 ) | ( n5335 & n14190 ) ;
  assign n14192 = ( ~n3629 & n5355 ) | ( ~n3629 & n8199 ) | ( n5355 & n8199 ) ;
  assign n14193 = n9378 ^ n5333 ^ n1918 ;
  assign n14194 = n8404 & ~n14193 ;
  assign n14195 = n3548 ^ n1364 ^ 1'b0 ;
  assign n14196 = ( n806 & n8507 ) | ( n806 & ~n10533 ) | ( n8507 & ~n10533 ) ;
  assign n14197 = ( n1837 & n7540 ) | ( n1837 & n14196 ) | ( n7540 & n14196 ) ;
  assign n14198 = ( ~n2049 & n3672 ) | ( ~n2049 & n9713 ) | ( n3672 & n9713 ) ;
  assign n14199 = n4760 ^ n448 ^ 1'b0 ;
  assign n14200 = ( ~n10522 & n14198 ) | ( ~n10522 & n14199 ) | ( n14198 & n14199 ) ;
  assign n14201 = ( n10650 & n14197 ) | ( n10650 & ~n14200 ) | ( n14197 & ~n14200 ) ;
  assign n14210 = n9267 ^ n8599 ^ n4090 ;
  assign n14205 = n3563 & n9029 ;
  assign n14206 = n14205 ^ n9734 ^ 1'b0 ;
  assign n14207 = ~n1724 & n14206 ;
  assign n14208 = n14207 ^ x192 ^ 1'b0 ;
  assign n14202 = n7169 | n7646 ;
  assign n14203 = n2593 | n14202 ;
  assign n14204 = n4090 & n14203 ;
  assign n14209 = n14208 ^ n14204 ^ 1'b0 ;
  assign n14211 = n14210 ^ n14209 ^ 1'b0 ;
  assign n14212 = ( n5189 & n9375 ) | ( n5189 & ~n10668 ) | ( n9375 & ~n10668 ) ;
  assign n14213 = ( n2918 & ~n4365 ) | ( n2918 & n14212 ) | ( ~n4365 & n14212 ) ;
  assign n14214 = ( n6886 & ~n8543 ) | ( n6886 & n11879 ) | ( ~n8543 & n11879 ) ;
  assign n14215 = n14214 ^ n9963 ^ n4524 ;
  assign n14216 = ( ~n5270 & n14213 ) | ( ~n5270 & n14215 ) | ( n14213 & n14215 ) ;
  assign n14217 = n8355 ^ n2715 ^ n1756 ;
  assign n14218 = ( x181 & ~n11472 ) | ( x181 & n14217 ) | ( ~n11472 & n14217 ) ;
  assign n14219 = n2665 & ~n3875 ;
  assign n14220 = n14219 ^ n1199 ^ 1'b0 ;
  assign n14221 = n4581 ^ n824 ^ 1'b0 ;
  assign n14222 = ( ~n7615 & n7765 ) | ( ~n7615 & n14221 ) | ( n7765 & n14221 ) ;
  assign n14223 = ( ~n11364 & n14220 ) | ( ~n11364 & n14222 ) | ( n14220 & n14222 ) ;
  assign n14224 = n14218 & ~n14223 ;
  assign n14226 = n13139 ^ n5772 ^ n4841 ;
  assign n14227 = ( ~n3261 & n9940 ) | ( ~n3261 & n14226 ) | ( n9940 & n14226 ) ;
  assign n14228 = ( n1202 & n1889 ) | ( n1202 & n14227 ) | ( n1889 & n14227 ) ;
  assign n14225 = x198 & n10036 ;
  assign n14229 = n14228 ^ n14225 ^ 1'b0 ;
  assign n14230 = n7289 ^ n1528 ^ x224 ;
  assign n14231 = ( n5429 & ~n8145 ) | ( n5429 & n14230 ) | ( ~n8145 & n14230 ) ;
  assign n14232 = n4409 & ~n12620 ;
  assign n14233 = n14232 ^ n10209 ^ n3011 ;
  assign n14234 = n14231 & n14233 ;
  assign n14235 = ( n442 & ~n1779 ) | ( n442 & n6562 ) | ( ~n1779 & n6562 ) ;
  assign n14236 = n7519 | n14235 ;
  assign n14240 = n5909 ^ n4571 ^ n1667 ;
  assign n14237 = n2081 & n2851 ;
  assign n14238 = ( ~n1229 & n2339 ) | ( ~n1229 & n14237 ) | ( n2339 & n14237 ) ;
  assign n14239 = ( n7130 & n8168 ) | ( n7130 & ~n14238 ) | ( n8168 & ~n14238 ) ;
  assign n14241 = n14240 ^ n14239 ^ n2462 ;
  assign n14242 = n12728 | n12812 ;
  assign n14243 = n14242 ^ n7100 ^ 1'b0 ;
  assign n14244 = ( n2212 & n8426 ) | ( n2212 & ~n13152 ) | ( n8426 & ~n13152 ) ;
  assign n14245 = n3119 & ~n11173 ;
  assign n14246 = n14245 ^ n7341 ^ 1'b0 ;
  assign n14247 = ( n336 & n6970 ) | ( n336 & n14246 ) | ( n6970 & n14246 ) ;
  assign n14248 = n11411 & n14247 ;
  assign n14249 = n14248 ^ n12147 ^ 1'b0 ;
  assign n14257 = ( ~n2903 & n3992 ) | ( ~n2903 & n4392 ) | ( n3992 & n4392 ) ;
  assign n14258 = ( n6143 & ~n10130 ) | ( n6143 & n14257 ) | ( ~n10130 & n14257 ) ;
  assign n14255 = ( n423 & n4033 ) | ( n423 & n6290 ) | ( n4033 & n6290 ) ;
  assign n14251 = n890 & ~n1679 ;
  assign n14252 = n2734 & n14251 ;
  assign n14253 = ( n368 & n4469 ) | ( n368 & n14252 ) | ( n4469 & n14252 ) ;
  assign n14254 = n14253 ^ n3385 ^ 1'b0 ;
  assign n14256 = n14255 ^ n14254 ^ n10735 ;
  assign n14250 = n12488 ^ n9379 ^ n2056 ;
  assign n14259 = n14258 ^ n14256 ^ n14250 ;
  assign n14262 = ( x163 & n2957 ) | ( x163 & ~n3693 ) | ( n2957 & ~n3693 ) ;
  assign n14260 = n11020 ^ n4712 ^ 1'b0 ;
  assign n14261 = n7922 & n14260 ;
  assign n14263 = n14262 ^ n14261 ^ n14057 ;
  assign n14264 = n14263 ^ n7572 ^ n4213 ;
  assign n14265 = x104 & ~n10438 ;
  assign n14266 = n14265 ^ x15 ^ 1'b0 ;
  assign n14267 = n14266 ^ n11212 ^ n5349 ;
  assign n14273 = ( ~n517 & n1049 ) | ( ~n517 & n3921 ) | ( n1049 & n3921 ) ;
  assign n14268 = n11945 ^ n3390 ^ n2183 ;
  assign n14269 = n11073 ^ n7633 ^ n1454 ;
  assign n14270 = n3770 & n14269 ;
  assign n14271 = n3398 & n14270 ;
  assign n14272 = ( n6613 & n14268 ) | ( n6613 & ~n14271 ) | ( n14268 & ~n14271 ) ;
  assign n14274 = n14273 ^ n14272 ^ n12612 ;
  assign n14275 = ( n1997 & ~n11739 ) | ( n1997 & n14274 ) | ( ~n11739 & n14274 ) ;
  assign n14276 = n3493 & n14222 ;
  assign n14278 = n4597 ^ n1796 ^ n1531 ;
  assign n14279 = ( ~n413 & n8466 ) | ( ~n413 & n14278 ) | ( n8466 & n14278 ) ;
  assign n14277 = n1127 | n7536 ;
  assign n14280 = n14279 ^ n14277 ^ 1'b0 ;
  assign n14281 = n14280 ^ n4641 ^ x220 ;
  assign n14282 = n14281 ^ n3269 ^ n2571 ;
  assign n14283 = n14282 ^ n6782 ^ 1'b0 ;
  assign n14284 = n4172 | n14283 ;
  assign n14285 = n9207 ^ n8013 ^ n4230 ;
  assign n14286 = ( n5570 & ~n6240 ) | ( n5570 & n14285 ) | ( ~n6240 & n14285 ) ;
  assign n14287 = n14286 ^ n12218 ^ n10445 ;
  assign n14288 = n4619 ^ n3990 ^ 1'b0 ;
  assign n14289 = n14288 ^ n1909 ^ 1'b0 ;
  assign n14290 = ~n12812 & n14289 ;
  assign n14291 = n14290 ^ n2272 ^ 1'b0 ;
  assign n14292 = ~n14287 & n14291 ;
  assign n14293 = ~n2422 & n14292 ;
  assign n14294 = n14293 ^ n11512 ^ n7687 ;
  assign n14295 = n3409 ^ n2051 ^ n1972 ;
  assign n14296 = n7874 ^ n4849 ^ n2111 ;
  assign n14297 = n14295 & ~n14296 ;
  assign n14298 = ~n947 & n14297 ;
  assign n14299 = n14298 ^ n3229 ^ 1'b0 ;
  assign n14300 = n3550 & n7023 ;
  assign n14301 = ( n2093 & ~n5856 ) | ( n2093 & n14124 ) | ( ~n5856 & n14124 ) ;
  assign n14302 = ( n8527 & ~n14300 ) | ( n8527 & n14301 ) | ( ~n14300 & n14301 ) ;
  assign n14303 = n397 & n2581 ;
  assign n14304 = n3208 & n14303 ;
  assign n14305 = ( ~n8481 & n8820 ) | ( ~n8481 & n14304 ) | ( n8820 & n14304 ) ;
  assign n14306 = n14305 ^ n13820 ^ 1'b0 ;
  assign n14308 = x173 & n2338 ;
  assign n14309 = n14308 ^ n10119 ^ n2180 ;
  assign n14307 = n12588 ^ n10437 ^ n2757 ;
  assign n14310 = n14309 ^ n14307 ^ n2467 ;
  assign n14311 = ~n3640 & n5439 ;
  assign n14312 = n14311 ^ n4613 ^ 1'b0 ;
  assign n14317 = n4554 & ~n5689 ;
  assign n14313 = n10828 ^ n5679 ^ x181 ;
  assign n14314 = n7363 ^ n5595 ^ n5170 ;
  assign n14315 = ( n7599 & n7695 ) | ( n7599 & n14314 ) | ( n7695 & n14314 ) ;
  assign n14316 = ( n9783 & n14313 ) | ( n9783 & n14315 ) | ( n14313 & n14315 ) ;
  assign n14318 = n14317 ^ n14316 ^ n14148 ;
  assign n14319 = ( n14310 & n14312 ) | ( n14310 & n14318 ) | ( n14312 & n14318 ) ;
  assign n14320 = x158 | n14319 ;
  assign n14322 = ( n2064 & n3143 ) | ( n2064 & ~n5688 ) | ( n3143 & ~n5688 ) ;
  assign n14323 = n14322 ^ n9283 ^ 1'b0 ;
  assign n14321 = n4576 | n13610 ;
  assign n14324 = n14323 ^ n14321 ^ 1'b0 ;
  assign n14326 = n3267 | n3689 ;
  assign n14325 = n10202 ^ n4962 ^ n2172 ;
  assign n14327 = n14326 ^ n14325 ^ 1'b0 ;
  assign n14328 = n14324 & n14327 ;
  assign n14329 = x160 & x189 ;
  assign n14330 = ( n3072 & n14328 ) | ( n3072 & n14329 ) | ( n14328 & n14329 ) ;
  assign n14331 = n9555 & n10179 ;
  assign n14332 = ( n1223 & ~n6687 ) | ( n1223 & n14331 ) | ( ~n6687 & n14331 ) ;
  assign n14333 = n8794 ^ n5294 ^ 1'b0 ;
  assign n14334 = n8573 & n14333 ;
  assign n14335 = n14334 ^ n4089 ^ 1'b0 ;
  assign n14336 = n2725 & n14335 ;
  assign n14338 = n8575 & ~n14217 ;
  assign n14339 = ( ~n1851 & n3812 ) | ( ~n1851 & n14338 ) | ( n3812 & n14338 ) ;
  assign n14340 = n4403 & ~n13128 ;
  assign n14341 = n8294 ^ n7348 ^ n1893 ;
  assign n14342 = ( ~n14339 & n14340 ) | ( ~n14339 & n14341 ) | ( n14340 & n14341 ) ;
  assign n14337 = n4031 ^ n2610 ^ n1447 ;
  assign n14343 = n14342 ^ n14337 ^ n13638 ;
  assign n14344 = n14343 ^ n1062 ^ 1'b0 ;
  assign n14345 = n7943 ^ n7055 ^ n4219 ;
  assign n14346 = n14345 ^ n8485 ^ 1'b0 ;
  assign n14350 = n8011 ^ n6769 ^ 1'b0 ;
  assign n14351 = n13574 | n14350 ;
  assign n14352 = n6084 & ~n14351 ;
  assign n14347 = ( ~n3484 & n7828 ) | ( ~n3484 & n13464 ) | ( n7828 & n13464 ) ;
  assign n14348 = ( n4239 & n9366 ) | ( n4239 & n14347 ) | ( n9366 & n14347 ) ;
  assign n14349 = n14348 ^ n12115 ^ n8669 ;
  assign n14353 = n14352 ^ n14349 ^ n10471 ;
  assign n14354 = ( ~n4853 & n13486 ) | ( ~n4853 & n14353 ) | ( n13486 & n14353 ) ;
  assign n14355 = n2504 & n4042 ;
  assign n14356 = n14355 ^ n8906 ^ 1'b0 ;
  assign n14357 = n12826 & n14356 ;
  assign n14358 = n14357 ^ n1602 ^ n1391 ;
  assign n14359 = n7047 ^ n3861 ^ 1'b0 ;
  assign n14360 = n14359 ^ n5977 ^ n4556 ;
  assign n14361 = n9075 ^ n6426 ^ n2595 ;
  assign n14362 = ( ~n8553 & n14360 ) | ( ~n8553 & n14361 ) | ( n14360 & n14361 ) ;
  assign n14363 = ( n6273 & n6789 ) | ( n6273 & ~n7337 ) | ( n6789 & ~n7337 ) ;
  assign n14364 = n3870 ^ x191 ^ 1'b0 ;
  assign n14365 = n14364 ^ n10989 ^ 1'b0 ;
  assign n14366 = n4399 & ~n14365 ;
  assign n14367 = ( n1063 & ~n11009 ) | ( n1063 & n14366 ) | ( ~n11009 & n14366 ) ;
  assign n14371 = n4641 ^ n1460 ^ n593 ;
  assign n14372 = ( n6890 & n7289 ) | ( n6890 & ~n14371 ) | ( n7289 & ~n14371 ) ;
  assign n14373 = n14372 ^ n7741 ^ 1'b0 ;
  assign n14374 = n14373 ^ n14198 ^ n12760 ;
  assign n14375 = n8175 ^ n5469 ^ 1'b0 ;
  assign n14376 = ~n14374 & n14375 ;
  assign n14368 = n9637 ^ n5282 ^ n2647 ;
  assign n14369 = n6933 ^ n2290 ^ 1'b0 ;
  assign n14370 = n14368 & n14369 ;
  assign n14377 = n14376 ^ n14370 ^ n10956 ;
  assign n14378 = n13860 ^ n5538 ^ 1'b0 ;
  assign n14379 = ( ~n1769 & n3825 ) | ( ~n1769 & n14378 ) | ( n3825 & n14378 ) ;
  assign n14380 = ( n1225 & n5771 ) | ( n1225 & ~n14379 ) | ( n5771 & ~n14379 ) ;
  assign n14381 = n13516 ^ n11152 ^ n6621 ;
  assign n14382 = n14381 ^ n12138 ^ n8209 ;
  assign n14383 = ( x153 & ~n948 ) | ( x153 & n6349 ) | ( ~n948 & n6349 ) ;
  assign n14384 = n747 & ~n12776 ;
  assign n14385 = ~n3118 & n14384 ;
  assign n14386 = n1123 & ~n14385 ;
  assign n14387 = n14386 ^ n5599 ^ 1'b0 ;
  assign n14388 = n14387 ^ n548 ^ x3 ;
  assign n14389 = n14383 & ~n14388 ;
  assign n14390 = ~n1101 & n14389 ;
  assign n14391 = ( n1701 & n14382 ) | ( n1701 & n14390 ) | ( n14382 & n14390 ) ;
  assign n14392 = ( ~n2234 & n12657 ) | ( ~n2234 & n13412 ) | ( n12657 & n13412 ) ;
  assign n14393 = n4624 | n7413 ;
  assign n14394 = n2580 ^ n1915 ^ 1'b0 ;
  assign n14395 = n11457 & n14394 ;
  assign n14396 = ( ~n8942 & n9204 ) | ( ~n8942 & n11957 ) | ( n9204 & n11957 ) ;
  assign n14397 = n580 & ~n14396 ;
  assign n14398 = ~n14395 & n14397 ;
  assign n14399 = n14393 & ~n14398 ;
  assign n14400 = n14399 ^ n9366 ^ 1'b0 ;
  assign n14401 = ( n6537 & n10633 ) | ( n6537 & ~n11367 ) | ( n10633 & ~n11367 ) ;
  assign n14402 = ( n7345 & n12318 ) | ( n7345 & n14401 ) | ( n12318 & n14401 ) ;
  assign n14403 = n1328 ^ n259 ^ 1'b0 ;
  assign n14404 = n1804 & ~n14403 ;
  assign n14405 = n14404 ^ n12308 ^ n3756 ;
  assign n14406 = n13886 ^ n11949 ^ 1'b0 ;
  assign n14407 = n10844 ^ n3960 ^ n2024 ;
  assign n14408 = n4182 | n14407 ;
  assign n14409 = n9462 | n14408 ;
  assign n14410 = n4471 | n9820 ;
  assign n14411 = n14410 ^ n12396 ^ n6855 ;
  assign n14412 = ( n554 & n12037 ) | ( n554 & n12092 ) | ( n12037 & n12092 ) ;
  assign n14413 = n6536 ^ n6432 ^ n1790 ;
  assign n14414 = n14413 ^ n6444 ^ 1'b0 ;
  assign n14415 = n14414 ^ n3376 ^ 1'b0 ;
  assign n14416 = n14412 | n14415 ;
  assign n14417 = ( n2378 & ~n4313 ) | ( n2378 & n5771 ) | ( ~n4313 & n5771 ) ;
  assign n14418 = ( n1809 & n6549 ) | ( n1809 & n12080 ) | ( n6549 & n12080 ) ;
  assign n14419 = ( n2336 & n2445 ) | ( n2336 & ~n2475 ) | ( n2445 & ~n2475 ) ;
  assign n14420 = n14419 ^ n10438 ^ n607 ;
  assign n14421 = ( n1509 & ~n2474 ) | ( n1509 & n4757 ) | ( ~n2474 & n4757 ) ;
  assign n14422 = n14421 ^ n3550 ^ n2738 ;
  assign n14423 = ( n6937 & ~n10041 ) | ( n6937 & n14422 ) | ( ~n10041 & n14422 ) ;
  assign n14424 = ( n11531 & ~n14420 ) | ( n11531 & n14423 ) | ( ~n14420 & n14423 ) ;
  assign n14425 = ( n14417 & n14418 ) | ( n14417 & n14424 ) | ( n14418 & n14424 ) ;
  assign n14426 = ( n3765 & n4238 ) | ( n3765 & ~n12287 ) | ( n4238 & ~n12287 ) ;
  assign n14427 = ~n13333 & n14426 ;
  assign n14428 = n14427 ^ n10599 ^ 1'b0 ;
  assign n14429 = n10931 & n13574 ;
  assign n14430 = n8384 ^ n3136 ^ 1'b0 ;
  assign n14431 = n14430 ^ n9284 ^ n3955 ;
  assign n14432 = n6715 & n14431 ;
  assign n14433 = n7536 ^ n7283 ^ n5775 ;
  assign n14434 = ( n4742 & n7342 ) | ( n4742 & n14433 ) | ( n7342 & n14433 ) ;
  assign n14435 = n12639 ^ n1318 ^ n316 ;
  assign n14436 = n14435 ^ n2298 ^ 1'b0 ;
  assign n14437 = ( ~n7357 & n7830 ) | ( ~n7357 & n12452 ) | ( n7830 & n12452 ) ;
  assign n14438 = n11763 ^ n11459 ^ n5653 ;
  assign n14439 = n2848 ^ n800 ^ 1'b0 ;
  assign n14440 = ~n8406 & n14439 ;
  assign n14441 = ~n9302 & n14440 ;
  assign n14444 = ~n3462 & n10918 ;
  assign n14442 = n2974 ^ n634 ^ 1'b0 ;
  assign n14443 = n11181 | n14442 ;
  assign n14445 = n14444 ^ n14443 ^ 1'b0 ;
  assign n14446 = n3826 & ~n14445 ;
  assign n14447 = n2374 ^ n571 ^ 1'b0 ;
  assign n14448 = n3319 & ~n14447 ;
  assign n14449 = ( ~n1392 & n3595 ) | ( ~n1392 & n8020 ) | ( n3595 & n8020 ) ;
  assign n14450 = n7901 ^ n5249 ^ n2191 ;
  assign n14451 = ( n985 & n8384 ) | ( n985 & ~n14450 ) | ( n8384 & ~n14450 ) ;
  assign n14452 = n14451 ^ n7582 ^ n1263 ;
  assign n14453 = n14449 & n14452 ;
  assign n14454 = ~n14448 & n14453 ;
  assign n14455 = n7433 ^ x72 ^ 1'b0 ;
  assign n14456 = n2755 & n14455 ;
  assign n14462 = n5669 ^ n2352 ^ n1706 ;
  assign n14463 = ( n3925 & n6056 ) | ( n3925 & ~n14462 ) | ( n6056 & ~n14462 ) ;
  assign n14464 = ( ~n2201 & n9467 ) | ( ~n2201 & n14463 ) | ( n9467 & n14463 ) ;
  assign n14465 = ( ~n604 & n7182 ) | ( ~n604 & n8760 ) | ( n7182 & n8760 ) ;
  assign n14466 = ( n3357 & n5777 ) | ( n3357 & ~n14465 ) | ( n5777 & ~n14465 ) ;
  assign n14467 = n14466 ^ n6486 ^ 1'b0 ;
  assign n14468 = n6378 ^ n2848 ^ n660 ;
  assign n14469 = n14468 ^ n1865 ^ 1'b0 ;
  assign n14470 = n9072 & n14469 ;
  assign n14471 = n14470 ^ n5711 ^ 1'b0 ;
  assign n14472 = n14467 & n14471 ;
  assign n14473 = ( n1723 & n14464 ) | ( n1723 & ~n14472 ) | ( n14464 & ~n14472 ) ;
  assign n14457 = ~n6832 & n10375 ;
  assign n14458 = ( n5581 & n11098 ) | ( n5581 & n14457 ) | ( n11098 & n14457 ) ;
  assign n14459 = ( n3980 & ~n5061 ) | ( n3980 & n11458 ) | ( ~n5061 & n11458 ) ;
  assign n14460 = n14459 ^ n7299 ^ 1'b0 ;
  assign n14461 = n14458 & n14460 ;
  assign n14474 = n14473 ^ n14461 ^ n14385 ;
  assign n14475 = ( n10476 & n12632 ) | ( n10476 & ~n14401 ) | ( n12632 & ~n14401 ) ;
  assign n14476 = ( ~n2760 & n5766 ) | ( ~n2760 & n13147 ) | ( n5766 & n13147 ) ;
  assign n14480 = n14268 ^ n1959 ^ n476 ;
  assign n14481 = ( ~n424 & n2577 ) | ( ~n424 & n14480 ) | ( n2577 & n14480 ) ;
  assign n14477 = n1903 ^ n1627 ^ 1'b0 ;
  assign n14478 = n7606 & ~n14477 ;
  assign n14479 = n2106 & n14478 ;
  assign n14482 = n14481 ^ n14479 ^ 1'b0 ;
  assign n14483 = n1463 & ~n8462 ;
  assign n14484 = n14483 ^ n7700 ^ 1'b0 ;
  assign n14485 = ( x71 & n1956 ) | ( x71 & n14484 ) | ( n1956 & n14484 ) ;
  assign n14486 = ( n4158 & n4509 ) | ( n4158 & ~n7909 ) | ( n4509 & ~n7909 ) ;
  assign n14487 = n13594 ^ n4241 ^ 1'b0 ;
  assign n14488 = n8586 & n9671 ;
  assign n14489 = ( ~n10321 & n14487 ) | ( ~n10321 & n14488 ) | ( n14487 & n14488 ) ;
  assign n14490 = ( n675 & ~n9799 ) | ( n675 & n12620 ) | ( ~n9799 & n12620 ) ;
  assign n14491 = n546 & ~n4820 ;
  assign n14492 = n4179 | n11020 ;
  assign n14493 = n14491 & ~n14492 ;
  assign n14494 = n6628 ^ n3598 ^ 1'b0 ;
  assign n14495 = n14494 ^ n6102 ^ n3477 ;
  assign n14496 = n4190 ^ n3700 ^ n2250 ;
  assign n14497 = n976 & ~n14496 ;
  assign n14498 = ( n8806 & ~n14495 ) | ( n8806 & n14497 ) | ( ~n14495 & n14497 ) ;
  assign n14499 = n14493 | n14498 ;
  assign n14500 = n12821 & ~n14499 ;
  assign n14502 = n2672 & ~n8732 ;
  assign n14503 = ~n4525 & n14502 ;
  assign n14501 = n2042 ^ n1015 ^ 1'b0 ;
  assign n14504 = n14503 ^ n14501 ^ n683 ;
  assign n14505 = ( n14490 & ~n14500 ) | ( n14490 & n14504 ) | ( ~n14500 & n14504 ) ;
  assign n14518 = n6509 ^ n3699 ^ n2161 ;
  assign n14519 = n14518 ^ n13653 ^ n12861 ;
  assign n14520 = n14519 ^ n7391 ^ n2901 ;
  assign n14513 = ( x200 & n3845 ) | ( x200 & ~n9062 ) | ( n3845 & ~n9062 ) ;
  assign n14514 = ~n3451 & n14513 ;
  assign n14515 = n14514 ^ n12422 ^ 1'b0 ;
  assign n14516 = n4804 & ~n14515 ;
  assign n14517 = n14516 ^ n2307 ^ 1'b0 ;
  assign n14506 = ( ~n2542 & n3494 ) | ( ~n2542 & n3776 ) | ( n3494 & n3776 ) ;
  assign n14510 = ( ~n2720 & n3304 ) | ( ~n2720 & n5087 ) | ( n3304 & n5087 ) ;
  assign n14508 = n1590 & n3103 ;
  assign n14509 = n3554 & n14508 ;
  assign n14507 = n10563 ^ n10165 ^ 1'b0 ;
  assign n14511 = n14510 ^ n14509 ^ n14507 ;
  assign n14512 = ( ~n7012 & n14506 ) | ( ~n7012 & n14511 ) | ( n14506 & n14511 ) ;
  assign n14521 = n14520 ^ n14517 ^ n14512 ;
  assign n14522 = ~n1009 & n1355 ;
  assign n14523 = n14522 ^ n3414 ^ 1'b0 ;
  assign n14524 = ( n1204 & ~n4808 ) | ( n1204 & n14523 ) | ( ~n4808 & n14523 ) ;
  assign n14525 = n14524 ^ n6361 ^ n2589 ;
  assign n14526 = n14525 ^ n4726 ^ n3004 ;
  assign n14527 = n3371 & ~n10384 ;
  assign n14528 = ( n842 & n7512 ) | ( n842 & n14527 ) | ( n7512 & n14527 ) ;
  assign n14533 = ( n2196 & n4597 ) | ( n2196 & ~n6285 ) | ( n4597 & ~n6285 ) ;
  assign n14534 = ( n1420 & ~n4286 ) | ( n1420 & n12259 ) | ( ~n4286 & n12259 ) ;
  assign n14535 = ( n5064 & n13858 ) | ( n5064 & ~n14534 ) | ( n13858 & ~n14534 ) ;
  assign n14536 = ( n6180 & ~n14533 ) | ( n6180 & n14535 ) | ( ~n14533 & n14535 ) ;
  assign n14537 = n9067 ^ n6369 ^ 1'b0 ;
  assign n14538 = n3376 | n14537 ;
  assign n14539 = ( n5053 & ~n12693 ) | ( n5053 & n14538 ) | ( ~n12693 & n14538 ) ;
  assign n14540 = ( n1517 & ~n14536 ) | ( n1517 & n14539 ) | ( ~n14536 & n14539 ) ;
  assign n14530 = ( n521 & n2892 ) | ( n521 & ~n12238 ) | ( n2892 & ~n12238 ) ;
  assign n14531 = ( ~x16 & n12071 ) | ( ~x16 & n14530 ) | ( n12071 & n14530 ) ;
  assign n14529 = n6228 ^ n4834 ^ n1431 ;
  assign n14532 = n14531 ^ n14529 ^ 1'b0 ;
  assign n14541 = n14540 ^ n14532 ^ n2165 ;
  assign n14546 = n5799 ^ n2580 ^ n1438 ;
  assign n14544 = n11588 ^ n3813 ^ 1'b0 ;
  assign n14545 = ~n12424 & n14544 ;
  assign n14542 = x69 & n359 ;
  assign n14543 = ~n11739 & n14542 ;
  assign n14547 = n14546 ^ n14545 ^ n14543 ;
  assign n14548 = n7197 & n7349 ;
  assign n14549 = n14548 ^ n8357 ^ 1'b0 ;
  assign n14550 = ( n718 & n4517 ) | ( n718 & ~n6509 ) | ( n4517 & ~n6509 ) ;
  assign n14551 = n14550 ^ n6575 ^ n2206 ;
  assign n14552 = n14549 & n14551 ;
  assign n14553 = n14552 ^ n4780 ^ 1'b0 ;
  assign n14554 = n9972 ^ n6463 ^ n826 ;
  assign n14555 = n10072 ^ n4942 ^ n4931 ;
  assign n14556 = n7567 | n14555 ;
  assign n14557 = n14554 | n14556 ;
  assign n14558 = ( n1798 & ~n8915 ) | ( n1798 & n14557 ) | ( ~n8915 & n14557 ) ;
  assign n14559 = n14558 ^ n12910 ^ n12103 ;
  assign n14560 = n2337 | n12944 ;
  assign n14561 = n14560 ^ n9304 ^ n6454 ;
  assign n14562 = n14561 ^ n1018 ^ 1'b0 ;
  assign n14563 = n7509 | n14562 ;
  assign n14564 = n10119 ^ n6477 ^ n5976 ;
  assign n14565 = ( n6082 & ~n6301 ) | ( n6082 & n14564 ) | ( ~n6301 & n14564 ) ;
  assign n14566 = n10191 ^ n798 ^ 1'b0 ;
  assign n14569 = ( ~x158 & n3735 ) | ( ~x158 & n4700 ) | ( n3735 & n4700 ) ;
  assign n14570 = ( n5043 & n7864 ) | ( n5043 & ~n7938 ) | ( n7864 & ~n7938 ) ;
  assign n14571 = n14570 ^ n3189 ^ n1252 ;
  assign n14572 = ( ~n5792 & n14569 ) | ( ~n5792 & n14571 ) | ( n14569 & n14571 ) ;
  assign n14567 = n11101 ^ n2556 ^ n1006 ;
  assign n14568 = n14567 ^ n552 ^ 1'b0 ;
  assign n14573 = n14572 ^ n14568 ^ n6688 ;
  assign n14574 = n14573 ^ n10271 ^ 1'b0 ;
  assign n14575 = n14566 | n14574 ;
  assign n14582 = n6991 & n13903 ;
  assign n14583 = n14582 ^ n1571 ^ 1'b0 ;
  assign n14576 = n10383 ^ n4217 ^ x35 ;
  assign n14577 = n14576 ^ n2402 ^ n783 ;
  assign n14578 = n6228 ^ n2485 ^ n401 ;
  assign n14579 = n14578 ^ n5055 ^ 1'b0 ;
  assign n14580 = n10608 & n14579 ;
  assign n14581 = ~n14577 & n14580 ;
  assign n14584 = n14583 ^ n14581 ^ n4589 ;
  assign n14585 = n9594 ^ n6581 ^ n2183 ;
  assign n14586 = n10649 ^ n9911 ^ n8320 ;
  assign n14587 = ( ~n3883 & n7368 ) | ( ~n3883 & n10124 ) | ( n7368 & n10124 ) ;
  assign n14588 = ( n10095 & n14586 ) | ( n10095 & n14587 ) | ( n14586 & n14587 ) ;
  assign n14589 = n14588 ^ n13415 ^ n1387 ;
  assign n14590 = n14589 ^ n11081 ^ 1'b0 ;
  assign n14595 = n11728 ^ n4685 ^ n2828 ;
  assign n14596 = ( n10386 & n13388 ) | ( n10386 & ~n14595 ) | ( n13388 & ~n14595 ) ;
  assign n14597 = ( n3297 & ~n8072 ) | ( n3297 & n14596 ) | ( ~n8072 & n14596 ) ;
  assign n14591 = n14278 ^ n3274 ^ 1'b0 ;
  assign n14592 = n7024 ^ x104 ^ 1'b0 ;
  assign n14593 = n14591 & ~n14592 ;
  assign n14594 = ( n3008 & n10336 ) | ( n3008 & ~n14593 ) | ( n10336 & ~n14593 ) ;
  assign n14598 = n14597 ^ n14594 ^ 1'b0 ;
  assign n14599 = ( x116 & n1248 ) | ( x116 & ~n1499 ) | ( n1248 & ~n1499 ) ;
  assign n14600 = n1753 | n14599 ;
  assign n14601 = n5041 & ~n14600 ;
  assign n14602 = ~n12865 & n14601 ;
  assign n14603 = ~n6213 & n10556 ;
  assign n14604 = n14603 ^ n7771 ^ 1'b0 ;
  assign n14605 = n292 & ~n5312 ;
  assign n14606 = n14605 ^ n5391 ^ n3769 ;
  assign n14607 = ( n11716 & ~n14604 ) | ( n11716 & n14606 ) | ( ~n14604 & n14606 ) ;
  assign n14608 = n569 & ~n5950 ;
  assign n14609 = n10702 ^ n491 ^ 1'b0 ;
  assign n14610 = ~n4600 & n14609 ;
  assign n14611 = n4072 & n14610 ;
  assign n14612 = ~n8153 & n14611 ;
  assign n14613 = ( n3230 & ~n6980 ) | ( n3230 & n14612 ) | ( ~n6980 & n14612 ) ;
  assign n14614 = ( n1774 & n2410 ) | ( n1774 & ~n4447 ) | ( n2410 & ~n4447 ) ;
  assign n14615 = n7073 & n14614 ;
  assign n14616 = n14615 ^ n9013 ^ 1'b0 ;
  assign n14617 = ( n14608 & n14613 ) | ( n14608 & ~n14616 ) | ( n14613 & ~n14616 ) ;
  assign n14618 = n4063 & ~n14309 ;
  assign n14619 = n14618 ^ n14551 ^ n13480 ;
  assign n14625 = n5246 | n6497 ;
  assign n14626 = n3378 | n14625 ;
  assign n14620 = n4849 ^ n2551 ^ n2544 ;
  assign n14621 = ~n5283 & n6910 ;
  assign n14622 = n14621 ^ n4956 ^ n2213 ;
  assign n14623 = n14620 | n14622 ;
  assign n14624 = n14623 ^ n1807 ^ 1'b0 ;
  assign n14627 = n14626 ^ n14624 ^ n1770 ;
  assign n14634 = n280 | n1882 ;
  assign n14630 = n5329 ^ n4862 ^ n4513 ;
  assign n14631 = n14630 ^ n9767 ^ n7745 ;
  assign n14632 = n14631 ^ n10262 ^ n8807 ;
  assign n14633 = ~n13555 & n14632 ;
  assign n14635 = n14634 ^ n14633 ^ 1'b0 ;
  assign n14628 = ( n2229 & ~n3176 ) | ( n2229 & n11443 ) | ( ~n3176 & n11443 ) ;
  assign n14629 = n14628 ^ n12594 ^ n9755 ;
  assign n14636 = n14635 ^ n14629 ^ n1814 ;
  assign n14637 = n1641 | n10656 ;
  assign n14638 = ( n1286 & n7043 ) | ( n1286 & n14637 ) | ( n7043 & n14637 ) ;
  assign n14639 = n2630 & ~n14638 ;
  assign n14640 = n14639 ^ n2170 ^ 1'b0 ;
  assign n14641 = n8934 & n10215 ;
  assign n14642 = n14641 ^ n1055 ^ 1'b0 ;
  assign n14645 = ( n1095 & n6321 ) | ( n1095 & n8674 ) | ( n6321 & n8674 ) ;
  assign n14643 = n13672 ^ n9292 ^ 1'b0 ;
  assign n14644 = n2291 & ~n14643 ;
  assign n14646 = n14645 ^ n14644 ^ 1'b0 ;
  assign n14647 = n7074 & ~n14646 ;
  assign n14648 = n14647 ^ n14253 ^ 1'b0 ;
  assign n14649 = n14642 & ~n14648 ;
  assign n14650 = n4841 ^ n1371 ^ x128 ;
  assign n14651 = n14650 ^ n8871 ^ n5173 ;
  assign n14652 = n14651 ^ n5235 ^ n926 ;
  assign n14653 = ( ~n2637 & n4974 ) | ( ~n2637 & n13013 ) | ( n4974 & n13013 ) ;
  assign n14654 = n911 & ~n1001 ;
  assign n14655 = ~n3335 & n14654 ;
  assign n14656 = ( n5559 & ~n6365 ) | ( n5559 & n14655 ) | ( ~n6365 & n14655 ) ;
  assign n14657 = n12599 & n14656 ;
  assign n14658 = n8019 & n8607 ;
  assign n14659 = ~n1302 & n14658 ;
  assign n14660 = ( n778 & n13186 ) | ( n778 & ~n14388 ) | ( n13186 & ~n14388 ) ;
  assign n14661 = ( n2101 & n10584 ) | ( n2101 & ~n14660 ) | ( n10584 & ~n14660 ) ;
  assign n14663 = n3093 | n7431 ;
  assign n14664 = n5463 & ~n14663 ;
  assign n14662 = n9637 ^ n7635 ^ n2973 ;
  assign n14665 = n14664 ^ n14662 ^ n11002 ;
  assign n14666 = n14661 & ~n14665 ;
  assign n14667 = ( n5367 & n9649 ) | ( n5367 & ~n14666 ) | ( n9649 & ~n14666 ) ;
  assign n14668 = n14667 ^ n11418 ^ n3379 ;
  assign n14669 = ( n6549 & n14659 ) | ( n6549 & ~n14668 ) | ( n14659 & ~n14668 ) ;
  assign n14670 = n6629 ^ n4439 ^ 1'b0 ;
  assign n14671 = n4937 | n14670 ;
  assign n14672 = n14671 ^ n5088 ^ n1017 ;
  assign n14673 = n11931 ^ n5860 ^ n3822 ;
  assign n14674 = ( n8707 & ~n14672 ) | ( n8707 & n14673 ) | ( ~n14672 & n14673 ) ;
  assign n14676 = n2841 | n9735 ;
  assign n14675 = ( ~n2972 & n13532 ) | ( ~n2972 & n14586 ) | ( n13532 & n14586 ) ;
  assign n14677 = n14676 ^ n14675 ^ n5975 ;
  assign n14678 = ( ~n3960 & n11977 ) | ( ~n3960 & n14677 ) | ( n11977 & n14677 ) ;
  assign n14683 = n9104 ^ n8577 ^ n4241 ;
  assign n14680 = ( ~n295 & n4014 ) | ( ~n295 & n8172 ) | ( n4014 & n8172 ) ;
  assign n14679 = n12367 ^ n4529 ^ n1427 ;
  assign n14681 = n14680 ^ n14679 ^ n280 ;
  assign n14682 = n14681 ^ n5466 ^ 1'b0 ;
  assign n14684 = n14683 ^ n14682 ^ n5274 ;
  assign n14685 = n6036 ^ n1434 ^ n1391 ;
  assign n14686 = n10532 ^ n6052 ^ 1'b0 ;
  assign n14687 = n14546 ^ n13558 ^ n13042 ;
  assign n14688 = n14687 ^ n7599 ^ 1'b0 ;
  assign n14689 = ~n14686 & n14688 ;
  assign n14690 = ( n4347 & n14685 ) | ( n4347 & ~n14689 ) | ( n14685 & ~n14689 ) ;
  assign n14691 = n14421 ^ n11182 ^ n10845 ;
  assign n14694 = n7354 ^ n683 ^ 1'b0 ;
  assign n14692 = n3365 ^ n2555 ^ 1'b0 ;
  assign n14693 = n4765 | n14692 ;
  assign n14695 = n14694 ^ n14693 ^ n1405 ;
  assign n14696 = ( n5828 & n10556 ) | ( n5828 & n14695 ) | ( n10556 & n14695 ) ;
  assign n14697 = ( ~n3629 & n3660 ) | ( ~n3629 & n8618 ) | ( n3660 & n8618 ) ;
  assign n14698 = ( n3864 & n9551 ) | ( n3864 & n14697 ) | ( n9551 & n14697 ) ;
  assign n14699 = ( n3927 & n9472 ) | ( n3927 & ~n14698 ) | ( n9472 & ~n14698 ) ;
  assign n14700 = n4915 | n6878 ;
  assign n14701 = n14700 ^ n3872 ^ 1'b0 ;
  assign n14702 = n7322 & n14701 ;
  assign n14703 = n8738 & n10358 ;
  assign n14704 = n14702 & n14703 ;
  assign n14707 = n14462 ^ n1938 ^ n378 ;
  assign n14705 = n10961 ^ n4384 ^ n1182 ;
  assign n14706 = ( n8493 & ~n10949 ) | ( n8493 & n14705 ) | ( ~n10949 & n14705 ) ;
  assign n14708 = n14707 ^ n14706 ^ n1363 ;
  assign n14709 = n5446 ^ n3195 ^ 1'b0 ;
  assign n14710 = n14709 ^ n9425 ^ n7539 ;
  assign n14711 = ( ~n2956 & n10785 ) | ( ~n2956 & n14710 ) | ( n10785 & n14710 ) ;
  assign n14712 = n6145 ^ n4298 ^ n2247 ;
  assign n14713 = n8442 & ~n14712 ;
  assign n14714 = n3843 & n14713 ;
  assign n14715 = n5349 ^ n4788 ^ n3054 ;
  assign n14716 = ( n6376 & n11427 ) | ( n6376 & n13938 ) | ( n11427 & n13938 ) ;
  assign n14717 = n14715 & ~n14716 ;
  assign n14718 = n14714 & n14717 ;
  assign n14719 = ( n4384 & n4841 ) | ( n4384 & n6811 ) | ( n4841 & n6811 ) ;
  assign n14720 = ~n11688 & n11840 ;
  assign n14721 = n12250 ^ n11378 ^ n3614 ;
  assign n14722 = n6628 & n9553 ;
  assign n14723 = ( ~n4962 & n14721 ) | ( ~n4962 & n14722 ) | ( n14721 & n14722 ) ;
  assign n14724 = ( n14719 & n14720 ) | ( n14719 & n14723 ) | ( n14720 & n14723 ) ;
  assign n14725 = n10173 ^ n8426 ^ n5187 ;
  assign n14726 = ~n1405 & n1666 ;
  assign n14727 = ~n5172 & n14726 ;
  assign n14728 = ( ~n8340 & n8358 ) | ( ~n8340 & n12930 ) | ( n8358 & n12930 ) ;
  assign n14729 = ( n1968 & n6279 ) | ( n1968 & ~n14728 ) | ( n6279 & ~n14728 ) ;
  assign n14730 = ( ~n3118 & n11679 ) | ( ~n3118 & n14729 ) | ( n11679 & n14729 ) ;
  assign n14731 = ~n14727 & n14730 ;
  assign n14732 = n14731 ^ n8829 ^ 1'b0 ;
  assign n14734 = n7337 ^ n6027 ^ 1'b0 ;
  assign n14735 = ( n10140 & ~n12847 ) | ( n10140 & n14734 ) | ( ~n12847 & n14734 ) ;
  assign n14733 = n9557 | n12484 ;
  assign n14736 = n14735 ^ n14733 ^ 1'b0 ;
  assign n14737 = ( n6968 & n8734 ) | ( n6968 & n11233 ) | ( n8734 & n11233 ) ;
  assign n14738 = ( ~n464 & n4135 ) | ( ~n464 & n13339 ) | ( n4135 & n13339 ) ;
  assign n14739 = n14738 ^ n6235 ^ 1'b0 ;
  assign n14740 = n14739 ^ n2307 ^ 1'b0 ;
  assign n14741 = n1597 | n14740 ;
  assign n14742 = n8771 ^ n4966 ^ 1'b0 ;
  assign n14743 = ~n372 & n14742 ;
  assign n14744 = n14743 ^ n11527 ^ n8663 ;
  assign n14745 = n14744 ^ n8197 ^ n2066 ;
  assign n14746 = n14307 ^ n13506 ^ n846 ;
  assign n14747 = ( n3820 & n11036 ) | ( n3820 & ~n14746 ) | ( n11036 & ~n14746 ) ;
  assign n14748 = ( ~n4049 & n10022 ) | ( ~n4049 & n12367 ) | ( n10022 & n12367 ) ;
  assign n14750 = ( x192 & ~n924 ) | ( x192 & n3249 ) | ( ~n924 & n3249 ) ;
  assign n14751 = n14750 ^ n7082 ^ 1'b0 ;
  assign n14749 = ( ~n2640 & n5116 ) | ( ~n2640 & n7244 ) | ( n5116 & n7244 ) ;
  assign n14752 = n14751 ^ n14749 ^ n13286 ;
  assign n14753 = ( n12419 & ~n14748 ) | ( n12419 & n14752 ) | ( ~n14748 & n14752 ) ;
  assign n14754 = ( n11124 & ~n12832 ) | ( n11124 & n13378 ) | ( ~n12832 & n13378 ) ;
  assign n14755 = ( ~n4247 & n14052 ) | ( ~n4247 & n14754 ) | ( n14052 & n14754 ) ;
  assign n14758 = n12320 ^ n7112 ^ 1'b0 ;
  assign n14759 = ~n2182 & n14758 ;
  assign n14757 = n7929 ^ n6716 ^ n5524 ;
  assign n14756 = n6270 ^ n303 ^ 1'b0 ;
  assign n14760 = n14759 ^ n14757 ^ n14756 ;
  assign n14773 = ( n5838 & n8432 ) | ( n5838 & ~n8819 ) | ( n8432 & ~n8819 ) ;
  assign n14761 = ( n5145 & ~n5179 ) | ( n5145 & n6634 ) | ( ~n5179 & n6634 ) ;
  assign n14762 = ( n7231 & n8501 ) | ( n7231 & n14761 ) | ( n8501 & n14761 ) ;
  assign n14763 = n14762 ^ n8559 ^ n7419 ;
  assign n14764 = x70 & ~n7140 ;
  assign n14765 = n6470 & n14764 ;
  assign n14766 = n14765 ^ n6963 ^ 1'b0 ;
  assign n14767 = n8071 & ~n14766 ;
  assign n14768 = ( n2176 & ~n14763 ) | ( n2176 & n14767 ) | ( ~n14763 & n14767 ) ;
  assign n14769 = n1069 & ~n6536 ;
  assign n14770 = n3187 & n14769 ;
  assign n14771 = n14770 ^ n2569 ^ 1'b0 ;
  assign n14772 = n14768 | n14771 ;
  assign n14774 = n14773 ^ n14772 ^ n411 ;
  assign n14779 = ( n2517 & n5283 ) | ( n2517 & ~n12260 ) | ( n5283 & ~n12260 ) ;
  assign n14780 = ( n4142 & n7145 ) | ( n4142 & n14779 ) | ( n7145 & n14779 ) ;
  assign n14781 = n14780 ^ n7430 ^ n1554 ;
  assign n14776 = n11657 ^ n8131 ^ 1'b0 ;
  assign n14777 = n14776 ^ n13378 ^ n10082 ;
  assign n14778 = n11985 & n14777 ;
  assign n14782 = n14781 ^ n14778 ^ 1'b0 ;
  assign n14775 = x93 & n12884 ;
  assign n14783 = n14782 ^ n14775 ^ n2243 ;
  assign n14784 = n4033 ^ n3852 ^ 1'b0 ;
  assign n14785 = n3739 & ~n14784 ;
  assign n14786 = ( n3463 & n7655 ) | ( n3463 & n14785 ) | ( n7655 & n14785 ) ;
  assign n14794 = ( n1125 & n3406 ) | ( n1125 & ~n13878 ) | ( n3406 & ~n13878 ) ;
  assign n14795 = ( n2298 & n2522 ) | ( n2298 & ~n14794 ) | ( n2522 & ~n14794 ) ;
  assign n14787 = n14012 ^ n11348 ^ n396 ;
  assign n14788 = ( n5657 & ~n10040 ) | ( n5657 & n14787 ) | ( ~n10040 & n14787 ) ;
  assign n14789 = ( ~n364 & n8404 ) | ( ~n364 & n13756 ) | ( n8404 & n13756 ) ;
  assign n14790 = n14789 ^ n5640 ^ n5531 ;
  assign n14791 = ( n12148 & n14687 ) | ( n12148 & n14790 ) | ( n14687 & n14790 ) ;
  assign n14792 = n14788 & ~n14791 ;
  assign n14793 = n14792 ^ n12541 ^ 1'b0 ;
  assign n14796 = n14795 ^ n14793 ^ n12811 ;
  assign n14801 = n10487 ^ n5415 ^ n2711 ;
  assign n14797 = n6519 & ~n7287 ;
  assign n14798 = n14797 ^ n2585 ^ 1'b0 ;
  assign n14799 = n10919 ^ n10603 ^ n2142 ;
  assign n14800 = ( ~n6814 & n14798 ) | ( ~n6814 & n14799 ) | ( n14798 & n14799 ) ;
  assign n14802 = n14801 ^ n14800 ^ n3472 ;
  assign n14803 = n4861 ^ n2267 ^ 1'b0 ;
  assign n14804 = n14803 ^ n3767 ^ n3409 ;
  assign n14805 = n3044 & n6468 ;
  assign n14806 = ~n11791 & n14805 ;
  assign n14807 = n14806 ^ n6464 ^ n2921 ;
  assign n14808 = ( n1612 & n14057 ) | ( n1612 & ~n14807 ) | ( n14057 & ~n14807 ) ;
  assign n14809 = n9843 ^ n5991 ^ 1'b0 ;
  assign n14819 = ( n826 & ~n1627 ) | ( n826 & n12141 ) | ( ~n1627 & n12141 ) ;
  assign n14812 = n353 & ~n5333 ;
  assign n14813 = n14812 ^ n9339 ^ 1'b0 ;
  assign n14810 = ( n3785 & n5041 ) | ( n3785 & n5228 ) | ( n5041 & n5228 ) ;
  assign n14811 = n11455 & ~n14810 ;
  assign n14814 = n14813 ^ n14811 ^ n7385 ;
  assign n14815 = n8333 ^ n5159 ^ 1'b0 ;
  assign n14816 = n3848 & n14815 ;
  assign n14817 = n14816 ^ n9017 ^ n4471 ;
  assign n14818 = ( ~n3317 & n14814 ) | ( ~n3317 & n14817 ) | ( n14814 & n14817 ) ;
  assign n14820 = n14819 ^ n14818 ^ n4361 ;
  assign n14821 = n14820 ^ n8744 ^ n8582 ;
  assign n14822 = ( n752 & n3444 ) | ( n752 & n14190 ) | ( n3444 & n14190 ) ;
  assign n14823 = n14822 ^ n1147 ^ 1'b0 ;
  assign n14824 = n4706 & ~n14823 ;
  assign n14825 = ( n342 & ~n14791 ) | ( n342 & n14824 ) | ( ~n14791 & n14824 ) ;
  assign n14826 = n1525 | n5663 ;
  assign n14827 = ( ~n5911 & n9715 ) | ( ~n5911 & n13406 ) | ( n9715 & n13406 ) ;
  assign n14828 = n2217 | n6740 ;
  assign n14829 = n14828 ^ n12811 ^ n4092 ;
  assign n14830 = ~n1811 & n5619 ;
  assign n14831 = n8482 & ~n14830 ;
  assign n14832 = ~n7948 & n14831 ;
  assign n14833 = n7654 & ~n8975 ;
  assign n14834 = n14833 ^ n10900 ^ n1806 ;
  assign n14835 = n14832 & ~n14834 ;
  assign n14839 = n8279 ^ n4189 ^ n1487 ;
  assign n14840 = ~n2260 & n14839 ;
  assign n14836 = n8130 ^ n4362 ^ n882 ;
  assign n14837 = n14836 ^ n1975 ^ 1'b0 ;
  assign n14838 = ~n4170 & n14837 ;
  assign n14841 = n14840 ^ n14838 ^ 1'b0 ;
  assign n14842 = n13558 | n14841 ;
  assign n14853 = ( n5458 & ~n6909 ) | ( n5458 & n7606 ) | ( ~n6909 & n7606 ) ;
  assign n14843 = ( n464 & ~n2162 ) | ( n464 & n3686 ) | ( ~n2162 & n3686 ) ;
  assign n14844 = ~n1854 & n14843 ;
  assign n14845 = n10232 & n14844 ;
  assign n14846 = ( n3352 & n4404 ) | ( n3352 & ~n12776 ) | ( n4404 & ~n12776 ) ;
  assign n14847 = n14846 ^ n9125 ^ n2563 ;
  assign n14848 = n12125 & n13115 ;
  assign n14849 = ( n4004 & n6201 ) | ( n4004 & ~n6737 ) | ( n6201 & ~n6737 ) ;
  assign n14850 = n14849 ^ n11516 ^ n3657 ;
  assign n14851 = ( ~n14847 & n14848 ) | ( ~n14847 & n14850 ) | ( n14848 & n14850 ) ;
  assign n14852 = ( n13284 & n14845 ) | ( n13284 & ~n14851 ) | ( n14845 & ~n14851 ) ;
  assign n14854 = n14853 ^ n14852 ^ n659 ;
  assign n14855 = n14854 ^ n2222 ^ n1701 ;
  assign n14861 = n2040 ^ x20 ^ 1'b0 ;
  assign n14862 = ( n2006 & ~n5897 ) | ( n2006 & n14861 ) | ( ~n5897 & n14861 ) ;
  assign n14856 = n1410 | n2599 ;
  assign n14857 = n14856 ^ n673 ^ 1'b0 ;
  assign n14858 = n12322 ^ n7193 ^ n761 ;
  assign n14859 = n5269 & n14858 ;
  assign n14860 = ~n14857 & n14859 ;
  assign n14863 = n14862 ^ n14860 ^ n6584 ;
  assign n14864 = n7850 ^ n2794 ^ n294 ;
  assign n14865 = ( n895 & n5539 ) | ( n895 & ~n6086 ) | ( n5539 & ~n6086 ) ;
  assign n14866 = n14865 ^ n13003 ^ n607 ;
  assign n14867 = ( ~n6393 & n7485 ) | ( ~n6393 & n9476 ) | ( n7485 & n9476 ) ;
  assign n14868 = n3525 & n14867 ;
  assign n14869 = n14868 ^ n12617 ^ 1'b0 ;
  assign n14870 = n13160 ^ n12765 ^ 1'b0 ;
  assign n14871 = n8407 | n14870 ;
  assign n14872 = ( n2769 & ~n4057 ) | ( n2769 & n10161 ) | ( ~n4057 & n10161 ) ;
  assign n14873 = n9354 & ~n14872 ;
  assign n14874 = n14873 ^ n13878 ^ n5575 ;
  assign n14875 = n11147 ^ n5596 ^ n4534 ;
  assign n14876 = n13400 ^ n5909 ^ n315 ;
  assign n14877 = ( ~n14306 & n14875 ) | ( ~n14306 & n14876 ) | ( n14875 & n14876 ) ;
  assign n14881 = x125 & ~n2459 ;
  assign n14878 = n2097 & ~n2884 ;
  assign n14879 = ~n6197 & n14878 ;
  assign n14880 = ( n590 & n6841 ) | ( n590 & n14879 ) | ( n6841 & n14879 ) ;
  assign n14882 = n14881 ^ n14880 ^ n6822 ;
  assign n14883 = ( n4778 & n9497 ) | ( n4778 & n14882 ) | ( n9497 & n14882 ) ;
  assign n14884 = n8938 | n11453 ;
  assign n14888 = ( n3835 & n5924 ) | ( n3835 & ~n9140 ) | ( n5924 & ~n9140 ) ;
  assign n14885 = ( n6285 & n9077 ) | ( n6285 & n9786 ) | ( n9077 & n9786 ) ;
  assign n14886 = ( ~n1943 & n3207 ) | ( ~n1943 & n5771 ) | ( n3207 & n5771 ) ;
  assign n14887 = n14885 & ~n14886 ;
  assign n14889 = n14888 ^ n14887 ^ 1'b0 ;
  assign n14890 = ( n660 & n3534 ) | ( n660 & n6653 ) | ( n3534 & n6653 ) ;
  assign n14893 = n9583 ^ x181 ^ x115 ;
  assign n14894 = n14893 ^ n1595 ^ n535 ;
  assign n14891 = ~n1558 & n5187 ;
  assign n14892 = n13912 & n14891 ;
  assign n14895 = n14894 ^ n14892 ^ n2465 ;
  assign n14896 = ( n8121 & ~n11078 ) | ( n8121 & n13079 ) | ( ~n11078 & n13079 ) ;
  assign n14897 = ~n8004 & n12273 ;
  assign n14898 = ( n14895 & ~n14896 ) | ( n14895 & n14897 ) | ( ~n14896 & n14897 ) ;
  assign n14899 = n13196 ^ n1581 ^ 1'b0 ;
  assign n14900 = ( ~n6019 & n12045 ) | ( ~n6019 & n14899 ) | ( n12045 & n14899 ) ;
  assign n14901 = ( ~x68 & n4381 ) | ( ~x68 & n4539 ) | ( n4381 & n4539 ) ;
  assign n14902 = n2435 & ~n9563 ;
  assign n14903 = n14902 ^ n8256 ^ n2151 ;
  assign n14904 = ~n11925 & n14903 ;
  assign n14905 = ~n14901 & n14904 ;
  assign n14906 = n13750 ^ n7276 ^ n4612 ;
  assign n14913 = n3000 ^ n2636 ^ n1253 ;
  assign n14914 = ( n1163 & n2208 ) | ( n1163 & n14913 ) | ( n2208 & n14913 ) ;
  assign n14915 = n8156 | n14914 ;
  assign n14907 = n14468 ^ n5218 ^ 1'b0 ;
  assign n14908 = n14907 ^ n8878 ^ n3437 ;
  assign n14909 = ( n1690 & n4015 ) | ( n1690 & n11232 ) | ( n4015 & n11232 ) ;
  assign n14910 = n14909 ^ n10389 ^ n675 ;
  assign n14911 = n14468 & n14910 ;
  assign n14912 = n14908 & n14911 ;
  assign n14916 = n14915 ^ n14912 ^ 1'b0 ;
  assign n14917 = n6564 ^ n5780 ^ 1'b0 ;
  assign n14918 = n4635 & ~n14917 ;
  assign n14919 = n14918 ^ n14656 ^ n3476 ;
  assign n14920 = n10240 ^ x231 ^ 1'b0 ;
  assign n14921 = n3033 | n14920 ;
  assign n14922 = ( n477 & n1976 ) | ( n477 & n2178 ) | ( n1976 & n2178 ) ;
  assign n14923 = n14922 ^ n7738 ^ 1'b0 ;
  assign n14924 = n4577 & ~n14923 ;
  assign n14925 = ~n14921 & n14924 ;
  assign n14926 = ~n14309 & n14925 ;
  assign n14927 = n3399 & ~n14926 ;
  assign n14928 = n14927 ^ n1961 ^ 1'b0 ;
  assign n14929 = n14928 ^ n12320 ^ n5237 ;
  assign n14930 = n771 | n9485 ;
  assign n14931 = n5316 & ~n14930 ;
  assign n14932 = ( n3576 & n7559 ) | ( n3576 & n8369 ) | ( n7559 & n8369 ) ;
  assign n14933 = n12624 ^ n11900 ^ n6715 ;
  assign n14934 = n6567 & n6842 ;
  assign n14935 = n4725 & n14934 ;
  assign n14936 = ( n281 & n6402 ) | ( n281 & n14935 ) | ( n6402 & n14935 ) ;
  assign n14937 = n14936 ^ n2563 ^ n2210 ;
  assign n14938 = n12521 ^ n11830 ^ n5472 ;
  assign n14939 = n14938 ^ n1112 ^ 1'b0 ;
  assign n14940 = n12281 ^ n5909 ^ n4628 ;
  assign n14941 = n3864 & ~n9276 ;
  assign n14942 = ( n6658 & ~n11928 ) | ( n6658 & n14941 ) | ( ~n11928 & n14941 ) ;
  assign n14943 = n14942 ^ n14661 ^ 1'b0 ;
  assign n14944 = n5574 & n14943 ;
  assign n14956 = ( n1012 & n6784 ) | ( n1012 & ~n12666 ) | ( n6784 & ~n12666 ) ;
  assign n14955 = ( n1489 & n1767 ) | ( n1489 & n5429 ) | ( n1767 & n5429 ) ;
  assign n14957 = n14956 ^ n14955 ^ n505 ;
  assign n14958 = ( n3765 & n9024 ) | ( n3765 & n14957 ) | ( n9024 & n14957 ) ;
  assign n14945 = n4491 ^ n3955 ^ n3618 ;
  assign n14946 = n14945 ^ n5150 ^ 1'b0 ;
  assign n14947 = n7944 & n14946 ;
  assign n14948 = ( ~n672 & n1599 ) | ( ~n672 & n14417 ) | ( n1599 & n14417 ) ;
  assign n14949 = n385 & ~n1907 ;
  assign n14950 = ( ~n2984 & n10447 ) | ( ~n2984 & n14949 ) | ( n10447 & n14949 ) ;
  assign n14951 = ( ~n2313 & n14948 ) | ( ~n2313 & n14950 ) | ( n14948 & n14950 ) ;
  assign n14952 = n5315 & ~n14951 ;
  assign n14953 = n14952 ^ n14843 ^ 1'b0 ;
  assign n14954 = ( ~n7657 & n14947 ) | ( ~n7657 & n14953 ) | ( n14947 & n14953 ) ;
  assign n14959 = n14958 ^ n14954 ^ n11749 ;
  assign n14960 = ( ~n2819 & n5372 ) | ( ~n2819 & n8922 ) | ( n5372 & n8922 ) ;
  assign n14961 = ( n4753 & ~n8789 ) | ( n4753 & n11806 ) | ( ~n8789 & n11806 ) ;
  assign n14962 = n11609 & ~n14961 ;
  assign n14963 = ( n3373 & n14960 ) | ( n3373 & n14962 ) | ( n14960 & n14962 ) ;
  assign n14964 = n2464 | n10062 ;
  assign n14965 = n5491 & ~n14964 ;
  assign n14967 = ( ~n707 & n3504 ) | ( ~n707 & n12466 ) | ( n3504 & n12466 ) ;
  assign n14966 = n12887 ^ n766 ^ 1'b0 ;
  assign n14968 = n14967 ^ n14966 ^ 1'b0 ;
  assign n14969 = ( n10938 & n14965 ) | ( n10938 & ~n14968 ) | ( n14965 & ~n14968 ) ;
  assign n14970 = n14969 ^ n9914 ^ n7514 ;
  assign n14971 = ( ~n452 & n2705 ) | ( ~n452 & n14970 ) | ( n2705 & n14970 ) ;
  assign n14972 = n12256 ^ n9038 ^ n4099 ;
  assign n14973 = ~n468 & n5221 ;
  assign n14974 = n14973 ^ n4809 ^ 1'b0 ;
  assign n14975 = n14974 ^ n4822 ^ 1'b0 ;
  assign n14976 = ~n10874 & n14975 ;
  assign n14977 = ( ~n889 & n1116 ) | ( ~n889 & n14976 ) | ( n1116 & n14976 ) ;
  assign n14978 = ( ~n9835 & n14972 ) | ( ~n9835 & n14977 ) | ( n14972 & n14977 ) ;
  assign n14979 = ~n5257 & n14978 ;
  assign n14980 = n4687 ^ n1694 ^ n764 ;
  assign n14981 = ( n9503 & n12660 ) | ( n9503 & ~n14980 ) | ( n12660 & ~n14980 ) ;
  assign n14982 = ( n3568 & n13431 ) | ( n3568 & n14981 ) | ( n13431 & n14981 ) ;
  assign n14983 = n5125 ^ n3385 ^ 1'b0 ;
  assign n14984 = n8168 & ~n14983 ;
  assign n14985 = n7417 ^ n2506 ^ n1736 ;
  assign n14986 = n14984 & ~n14985 ;
  assign n14987 = n14986 ^ n4272 ^ 1'b0 ;
  assign n14988 = ( n4839 & n10193 ) | ( n4839 & ~n10334 ) | ( n10193 & ~n10334 ) ;
  assign n14989 = ( x37 & n2058 ) | ( x37 & n14988 ) | ( n2058 & n14988 ) ;
  assign n14990 = ( n6397 & n8945 ) | ( n6397 & ~n14989 ) | ( n8945 & ~n14989 ) ;
  assign n14991 = n12714 ^ n12094 ^ n6182 ;
  assign n14992 = ( ~n7819 & n7959 ) | ( ~n7819 & n9630 ) | ( n7959 & n9630 ) ;
  assign n14993 = n14992 ^ n6627 ^ n3281 ;
  assign n14994 = n13563 ^ n8344 ^ n5498 ;
  assign n14995 = n14994 ^ n13815 ^ 1'b0 ;
  assign n14996 = ~n2511 & n13972 ;
  assign n14997 = n14996 ^ n7518 ^ 1'b0 ;
  assign n14998 = n7204 ^ n1514 ^ n1028 ;
  assign n14999 = ( n990 & ~n7930 ) | ( n990 & n14998 ) | ( ~n7930 & n14998 ) ;
  assign n15000 = ( n3127 & n8379 ) | ( n3127 & ~n14999 ) | ( n8379 & ~n14999 ) ;
  assign n15003 = n14148 ^ n2641 ^ 1'b0 ;
  assign n15004 = n6931 & ~n10144 ;
  assign n15005 = n15003 & n15004 ;
  assign n15001 = n2555 & n5562 ;
  assign n15002 = n15001 ^ n10455 ^ n9685 ;
  assign n15006 = n15005 ^ n15002 ^ n12132 ;
  assign n15007 = ( n6881 & ~n7741 ) | ( n6881 & n12151 ) | ( ~n7741 & n12151 ) ;
  assign n15008 = n15007 ^ n11314 ^ n10313 ;
  assign n15009 = n15008 ^ n12241 ^ n8622 ;
  assign n15010 = n2431 ^ n1220 ^ n619 ;
  assign n15011 = n15010 ^ n4195 ^ n1692 ;
  assign n15012 = ( x42 & n12869 ) | ( x42 & n15011 ) | ( n12869 & n15011 ) ;
  assign n15013 = n8849 ^ n2066 ^ n1896 ;
  assign n15014 = n15013 ^ n9146 ^ n6477 ;
  assign n15019 = n10496 ^ n8048 ^ 1'b0 ;
  assign n15020 = n15019 ^ n6848 ^ n2604 ;
  assign n15015 = ~n11728 & n12340 ;
  assign n15016 = n14083 ^ n5966 ^ n1698 ;
  assign n15017 = ( n6141 & n15015 ) | ( n6141 & ~n15016 ) | ( n15015 & ~n15016 ) ;
  assign n15018 = n9088 | n15017 ;
  assign n15021 = n15020 ^ n15018 ^ 1'b0 ;
  assign n15022 = n7717 ^ n3958 ^ 1'b0 ;
  assign n15023 = n14980 | n15022 ;
  assign n15024 = n6929 ^ n2892 ^ n1978 ;
  assign n15025 = n14164 & ~n15024 ;
  assign n15026 = ( n13580 & ~n15023 ) | ( n13580 & n15025 ) | ( ~n15023 & n15025 ) ;
  assign n15027 = n5708 ^ n5477 ^ n2815 ;
  assign n15028 = n1398 & ~n2775 ;
  assign n15029 = ( n4571 & n6380 ) | ( n4571 & ~n13209 ) | ( n6380 & ~n13209 ) ;
  assign n15030 = ( n10176 & n15028 ) | ( n10176 & n15029 ) | ( n15028 & n15029 ) ;
  assign n15031 = n15030 ^ n12199 ^ n5050 ;
  assign n15032 = n1486 | n15031 ;
  assign n15033 = n15032 ^ n8209 ^ 1'b0 ;
  assign n15040 = ( n1515 & n2393 ) | ( n1515 & ~n10605 ) | ( n2393 & ~n10605 ) ;
  assign n15041 = n7605 & n15040 ;
  assign n15042 = n7897 & n15041 ;
  assign n15043 = n15042 ^ n7905 ^ n5745 ;
  assign n15034 = n11993 ^ n8042 ^ n3991 ;
  assign n15035 = n1067 & n3720 ;
  assign n15036 = ~n9758 & n15035 ;
  assign n15037 = n15034 | n15036 ;
  assign n15038 = n811 & ~n15037 ;
  assign n15039 = ( n10634 & n14022 ) | ( n10634 & n15038 ) | ( n14022 & n15038 ) ;
  assign n15044 = n15043 ^ n15039 ^ n623 ;
  assign n15045 = n7204 | n9209 ;
  assign n15046 = n15045 ^ n10698 ^ 1'b0 ;
  assign n15047 = ( ~n5961 & n6941 ) | ( ~n5961 & n10504 ) | ( n6941 & n10504 ) ;
  assign n15048 = ( n1962 & ~n6182 ) | ( n1962 & n15047 ) | ( ~n6182 & n15047 ) ;
  assign n15049 = n12580 ^ n5322 ^ n1509 ;
  assign n15050 = n12073 ^ n10679 ^ n4032 ;
  assign n15051 = ( x170 & n2223 ) | ( x170 & n9670 ) | ( n2223 & n9670 ) ;
  assign n15052 = n15051 ^ n12564 ^ n11400 ;
  assign n15053 = n15052 ^ n14227 ^ n13498 ;
  assign n15054 = ( n514 & ~n7137 ) | ( n514 & n13543 ) | ( ~n7137 & n13543 ) ;
  assign n15055 = n2877 & ~n15054 ;
  assign n15056 = ( n10785 & n12254 ) | ( n10785 & n15055 ) | ( n12254 & n15055 ) ;
  assign n15059 = n3341 | n8784 ;
  assign n15060 = n1216 & ~n15059 ;
  assign n15057 = n5154 ^ n5150 ^ n1442 ;
  assign n15058 = n10135 & n15057 ;
  assign n15061 = n15060 ^ n15058 ^ 1'b0 ;
  assign n15062 = n15061 ^ n5690 ^ 1'b0 ;
  assign n15063 = ~n15056 & n15062 ;
  assign n15064 = n14750 ^ n11478 ^ n2304 ;
  assign n15065 = n7717 ^ n4725 ^ n2393 ;
  assign n15066 = ( n6165 & ~n11537 ) | ( n6165 & n15065 ) | ( ~n11537 & n15065 ) ;
  assign n15067 = n15066 ^ n8709 ^ n4107 ;
  assign n15068 = ( n1510 & n6495 ) | ( n1510 & n12311 ) | ( n6495 & n12311 ) ;
  assign n15069 = ( n4408 & n7722 ) | ( n4408 & ~n15068 ) | ( n7722 & ~n15068 ) ;
  assign n15070 = n346 & ~n2680 ;
  assign n15071 = n15070 ^ n14721 ^ n10433 ;
  assign n15072 = ( ~n5491 & n5672 ) | ( ~n5491 & n8849 ) | ( n5672 & n8849 ) ;
  assign n15073 = ( ~n6671 & n12813 ) | ( ~n6671 & n15072 ) | ( n12813 & n15072 ) ;
  assign n15074 = n14569 ^ n9958 ^ x7 ;
  assign n15075 = n11765 ^ n2025 ^ 1'b0 ;
  assign n15076 = ~n9882 & n15075 ;
  assign n15077 = ~n15074 & n15076 ;
  assign n15078 = n3996 ^ n3911 ^ n575 ;
  assign n15079 = n8204 | n15078 ;
  assign n15080 = ( n6917 & n7048 ) | ( n6917 & ~n15079 ) | ( n7048 & ~n15079 ) ;
  assign n15081 = ~n1044 & n10381 ;
  assign n15082 = ~n1007 & n15081 ;
  assign n15083 = ( n6652 & n6856 ) | ( n6652 & n15082 ) | ( n6856 & n15082 ) ;
  assign n15084 = n9221 ^ n7710 ^ n7534 ;
  assign n15087 = ( ~n2490 & n5354 ) | ( ~n2490 & n9825 ) | ( n5354 & n9825 ) ;
  assign n15085 = n7532 ^ n6416 ^ n6314 ;
  assign n15086 = n15085 ^ n10872 ^ n7253 ;
  assign n15088 = n15087 ^ n15086 ^ 1'b0 ;
  assign n15089 = n12507 ^ n9787 ^ n9465 ;
  assign n15090 = n14057 ^ n5723 ^ n729 ;
  assign n15091 = ( ~n879 & n4327 ) | ( ~n879 & n10132 ) | ( n4327 & n10132 ) ;
  assign n15092 = ( ~n3207 & n9020 ) | ( ~n3207 & n11021 ) | ( n9020 & n11021 ) ;
  assign n15093 = n10925 ^ n5218 ^ n5046 ;
  assign n15094 = ~n6919 & n15093 ;
  assign n15095 = n15092 & n15094 ;
  assign n15096 = n11373 ^ n7976 ^ n1978 ;
  assign n15097 = n15096 ^ n1930 ^ 1'b0 ;
  assign n15098 = ( n2815 & ~n11343 ) | ( n2815 & n11429 ) | ( ~n11343 & n11429 ) ;
  assign n15099 = n15098 ^ n9062 ^ n774 ;
  assign n15100 = n10659 & ~n15099 ;
  assign n15101 = n10866 ^ n5537 ^ n1016 ;
  assign n15102 = n15101 ^ n2234 ^ n773 ;
  assign n15103 = ( n15097 & n15100 ) | ( n15097 & ~n15102 ) | ( n15100 & ~n15102 ) ;
  assign n15104 = n10361 ^ n10186 ^ n7669 ;
  assign n15105 = ( n9681 & ~n13244 ) | ( n9681 & n15104 ) | ( ~n13244 & n15104 ) ;
  assign n15106 = n4966 ^ n4854 ^ n4043 ;
  assign n15107 = n15106 ^ n6914 ^ n1382 ;
  assign n15108 = ( n1044 & n5338 ) | ( n1044 & n15107 ) | ( n5338 & n15107 ) ;
  assign n15113 = n10580 ^ n3557 ^ n1766 ;
  assign n15116 = ( n1701 & ~n5853 ) | ( n1701 & n9042 ) | ( ~n5853 & n9042 ) ;
  assign n15114 = ~n5288 & n5800 ;
  assign n15115 = ( ~n5525 & n7125 ) | ( ~n5525 & n15114 ) | ( n7125 & n15114 ) ;
  assign n15117 = n15116 ^ n15115 ^ n2192 ;
  assign n15118 = ( n4127 & n15113 ) | ( n4127 & ~n15117 ) | ( n15113 & ~n15117 ) ;
  assign n15109 = n12947 ^ n10617 ^ n1248 ;
  assign n15110 = n5632 ^ n5460 ^ n4018 ;
  assign n15111 = ( n7086 & n15109 ) | ( n7086 & ~n15110 ) | ( n15109 & ~n15110 ) ;
  assign n15112 = n15111 ^ n6288 ^ 1'b0 ;
  assign n15119 = n15118 ^ n15112 ^ 1'b0 ;
  assign n15120 = n11664 ^ n4249 ^ 1'b0 ;
  assign n15121 = ~n2179 & n15120 ;
  assign n15122 = ( n3290 & ~n7237 ) | ( n3290 & n14967 ) | ( ~n7237 & n14967 ) ;
  assign n15123 = n2115 & ~n4481 ;
  assign n15124 = n15123 ^ n6553 ^ 1'b0 ;
  assign n15125 = ( n6340 & n9401 ) | ( n6340 & n15124 ) | ( n9401 & n15124 ) ;
  assign n15126 = n10175 ^ n766 ^ 1'b0 ;
  assign n15127 = ~n15125 & n15126 ;
  assign n15128 = ~n5196 & n15127 ;
  assign n15129 = n15122 & n15128 ;
  assign n15130 = ( n10570 & n15121 ) | ( n10570 & n15129 ) | ( n15121 & n15129 ) ;
  assign n15131 = n2901 | n5969 ;
  assign n15132 = n6093 | n7478 ;
  assign n15133 = n4189 & ~n15132 ;
  assign n15134 = n3026 & ~n15133 ;
  assign n15136 = n8580 ^ n1976 ^ x157 ;
  assign n15135 = n665 | n4253 ;
  assign n15137 = n15136 ^ n15135 ^ n7675 ;
  assign n15138 = ( ~n10113 & n15134 ) | ( ~n10113 & n15137 ) | ( n15134 & n15137 ) ;
  assign n15139 = n12942 ^ n7915 ^ n4731 ;
  assign n15140 = n15139 ^ n10385 ^ n4770 ;
  assign n15141 = ( ~n5602 & n11671 ) | ( ~n5602 & n15140 ) | ( n11671 & n15140 ) ;
  assign n15142 = n15141 ^ n5670 ^ 1'b0 ;
  assign n15143 = ~n15138 & n15142 ;
  assign n15147 = ~n11348 & n14378 ;
  assign n15144 = ( n1499 & ~n2436 ) | ( n1499 & n6988 ) | ( ~n2436 & n6988 ) ;
  assign n15145 = n15144 ^ n4388 ^ 1'b0 ;
  assign n15146 = n13639 | n15145 ;
  assign n15148 = n15147 ^ n15146 ^ 1'b0 ;
  assign n15149 = n5814 ^ n1041 ^ n779 ;
  assign n15157 = n4684 & n9624 ;
  assign n15158 = n15157 ^ n859 ^ 1'b0 ;
  assign n15159 = n15158 ^ n7216 ^ 1'b0 ;
  assign n15150 = n4307 | n7167 ;
  assign n15151 = n15150 ^ n10385 ^ 1'b0 ;
  assign n15152 = n15151 ^ n2301 ^ n755 ;
  assign n15153 = ( n5087 & ~n10646 ) | ( n5087 & n10795 ) | ( ~n10646 & n10795 ) ;
  assign n15154 = n2448 | n15153 ;
  assign n15155 = n15154 ^ n15016 ^ 1'b0 ;
  assign n15156 = ( n5978 & ~n15152 ) | ( n5978 & n15155 ) | ( ~n15152 & n15155 ) ;
  assign n15160 = n15159 ^ n15156 ^ n714 ;
  assign n15161 = ( ~n7777 & n12539 ) | ( ~n7777 & n15160 ) | ( n12539 & n15160 ) ;
  assign n15162 = ~n15149 & n15161 ;
  assign n15164 = n12963 ^ n6854 ^ n5006 ;
  assign n15163 = n11564 ^ n5663 ^ n4668 ;
  assign n15165 = n15164 ^ n15163 ^ n12715 ;
  assign n15167 = ( ~n2320 & n3628 ) | ( ~n2320 & n5510 ) | ( n3628 & n5510 ) ;
  assign n15166 = n2841 | n10385 ;
  assign n15168 = n15167 ^ n15166 ^ 1'b0 ;
  assign n15169 = ( ~n963 & n5840 ) | ( ~n963 & n15168 ) | ( n5840 & n15168 ) ;
  assign n15170 = n1675 | n7502 ;
  assign n15171 = ( n10463 & n15169 ) | ( n10463 & n15170 ) | ( n15169 & n15170 ) ;
  assign n15173 = ( n485 & n5396 ) | ( n485 & ~n11551 ) | ( n5396 & ~n11551 ) ;
  assign n15172 = n4632 ^ n1027 ^ 1'b0 ;
  assign n15174 = n15173 ^ n15172 ^ n12243 ;
  assign n15175 = ( n6359 & ~n12507 ) | ( n6359 & n13392 ) | ( ~n12507 & n13392 ) ;
  assign n15176 = n9267 ^ n7732 ^ n7180 ;
  assign n15177 = ( ~n11801 & n15175 ) | ( ~n11801 & n15176 ) | ( n15175 & n15176 ) ;
  assign n15184 = ( n2350 & ~n5612 ) | ( n2350 & n13160 ) | ( ~n5612 & n13160 ) ;
  assign n15178 = ( n5001 & ~n7190 ) | ( n5001 & n10854 ) | ( ~n7190 & n10854 ) ;
  assign n15179 = ( ~n3660 & n8563 ) | ( ~n3660 & n12869 ) | ( n8563 & n12869 ) ;
  assign n15180 = n15179 ^ n2697 ^ n1831 ;
  assign n15181 = n15180 ^ n2518 ^ 1'b0 ;
  assign n15182 = n15181 ^ n2255 ^ n590 ;
  assign n15183 = n15178 & ~n15182 ;
  assign n15185 = n15184 ^ n15183 ^ 1'b0 ;
  assign n15186 = n1550 | n11678 ;
  assign n15187 = n15186 ^ n8269 ^ 1'b0 ;
  assign n15188 = n15185 | n15187 ;
  assign n15189 = n11091 | n15188 ;
  assign n15190 = ( n711 & ~n2364 ) | ( n711 & n7185 ) | ( ~n2364 & n7185 ) ;
  assign n15191 = n2165 | n15190 ;
  assign n15192 = ( n9572 & n11007 ) | ( n9572 & n15191 ) | ( n11007 & n15191 ) ;
  assign n15193 = n14865 & ~n15192 ;
  assign n15194 = ( ~n11652 & n12200 ) | ( ~n11652 & n14798 ) | ( n12200 & n14798 ) ;
  assign n15198 = n10914 ^ n3554 ^ n2619 ;
  assign n15195 = ( n1996 & n2227 ) | ( n1996 & n5040 ) | ( n2227 & n5040 ) ;
  assign n15196 = n15195 ^ n767 ^ 1'b0 ;
  assign n15197 = n864 & n15196 ;
  assign n15199 = n15198 ^ n15197 ^ n3456 ;
  assign n15200 = n15199 ^ n13083 ^ n9041 ;
  assign n15201 = n15200 ^ n11288 ^ 1'b0 ;
  assign n15202 = n11385 ^ n9512 ^ n5409 ;
  assign n15203 = n15202 ^ n11740 ^ n10630 ;
  assign n15204 = ( ~n1507 & n5236 ) | ( ~n1507 & n15203 ) | ( n5236 & n15203 ) ;
  assign n15205 = n15204 ^ n15013 ^ n8423 ;
  assign n15206 = ( n2482 & n4309 ) | ( n2482 & ~n5425 ) | ( n4309 & ~n5425 ) ;
  assign n15207 = ( x197 & ~n522 ) | ( x197 & n15206 ) | ( ~n522 & n15206 ) ;
  assign n15208 = n15207 ^ n11945 ^ n2042 ;
  assign n15209 = n15208 ^ n6262 ^ n3826 ;
  assign n15210 = ~n868 & n15209 ;
  assign n15211 = n15210 ^ n6856 ^ 1'b0 ;
  assign n15213 = n3961 ^ x113 ^ 1'b0 ;
  assign n15214 = n15213 ^ n5622 ^ n4567 ;
  assign n15212 = ( n2619 & ~n5807 ) | ( n2619 & n7781 ) | ( ~n5807 & n7781 ) ;
  assign n15215 = n15214 ^ n15212 ^ x185 ;
  assign n15216 = n15215 ^ n4705 ^ n4048 ;
  assign n15217 = n9917 ^ n3367 ^ n1662 ;
  assign n15218 = n15217 ^ n2426 ^ n2117 ;
  assign n15219 = ( n729 & n4764 ) | ( n729 & ~n15218 ) | ( n4764 & ~n15218 ) ;
  assign n15220 = ( ~n2709 & n3798 ) | ( ~n2709 & n11684 ) | ( n3798 & n11684 ) ;
  assign n15221 = n787 & n15220 ;
  assign n15222 = ~n13018 & n15221 ;
  assign n15223 = ~n15219 & n15222 ;
  assign n15228 = ( n2271 & n6844 ) | ( n2271 & ~n10453 ) | ( n6844 & ~n10453 ) ;
  assign n15226 = ( n2076 & n3478 ) | ( n2076 & n3828 ) | ( n3478 & n3828 ) ;
  assign n15224 = n6138 ^ n655 ^ 1'b0 ;
  assign n15225 = n2619 & n15224 ;
  assign n15227 = n15226 ^ n15225 ^ n4252 ;
  assign n15229 = n15228 ^ n15227 ^ n10948 ;
  assign n15230 = ( n1141 & n1503 ) | ( n1141 & n9053 ) | ( n1503 & n9053 ) ;
  assign n15231 = ( n1826 & ~n8055 ) | ( n1826 & n15230 ) | ( ~n8055 & n15230 ) ;
  assign n15232 = n4354 & n15231 ;
  assign n15233 = n15232 ^ n6670 ^ 1'b0 ;
  assign n15234 = n15229 | n15233 ;
  assign n15235 = n12508 ^ n7561 ^ n2038 ;
  assign n15236 = n6434 ^ n6172 ^ n4523 ;
  assign n15237 = n15236 ^ n3713 ^ 1'b0 ;
  assign n15238 = n15235 | n15237 ;
  assign n15239 = n6531 ^ n2126 ^ n1308 ;
  assign n15240 = ~n1522 & n15239 ;
  assign n15245 = x166 & ~n6759 ;
  assign n15246 = ~n5564 & n15245 ;
  assign n15247 = n6673 & n7719 ;
  assign n15248 = n15246 & n15247 ;
  assign n15242 = ( n9760 & ~n13612 ) | ( n9760 & n14217 ) | ( ~n13612 & n14217 ) ;
  assign n15243 = n15242 ^ n4345 ^ n1308 ;
  assign n15241 = ( n3437 & ~n8982 ) | ( n3437 & n12890 ) | ( ~n8982 & n12890 ) ;
  assign n15244 = n15243 ^ n15241 ^ n8212 ;
  assign n15249 = n15248 ^ n15244 ^ n9799 ;
  assign n15250 = n727 | n9170 ;
  assign n15251 = ( n3400 & ~n12008 ) | ( n3400 & n15250 ) | ( ~n12008 & n15250 ) ;
  assign n15254 = ( n968 & ~n3661 ) | ( n968 & n4345 ) | ( ~n3661 & n4345 ) ;
  assign n15252 = n5072 ^ n2237 ^ 1'b0 ;
  assign n15253 = n1780 & ~n15252 ;
  assign n15255 = n15254 ^ n15253 ^ n2952 ;
  assign n15256 = n8527 ^ n6395 ^ n1963 ;
  assign n15262 = n2008 & ~n6560 ;
  assign n15263 = n15262 ^ n6514 ^ n769 ;
  assign n15257 = ( ~n2278 & n2507 ) | ( ~n2278 & n13947 ) | ( n2507 & n13947 ) ;
  assign n15258 = n15257 ^ n4349 ^ n2979 ;
  assign n15259 = n15258 ^ n3583 ^ n1371 ;
  assign n15260 = n6522 ^ n2812 ^ n757 ;
  assign n15261 = ( n3629 & ~n15259 ) | ( n3629 & n15260 ) | ( ~n15259 & n15260 ) ;
  assign n15264 = n15263 ^ n15261 ^ n6520 ;
  assign n15265 = n15264 ^ n9579 ^ n7874 ;
  assign n15266 = ( ~n910 & n15256 ) | ( ~n910 & n15265 ) | ( n15256 & n15265 ) ;
  assign n15267 = n15266 ^ n15145 ^ n13975 ;
  assign n15268 = ( n3949 & n5756 ) | ( n3949 & ~n12096 ) | ( n5756 & ~n12096 ) ;
  assign n15271 = ( n1367 & ~n4559 ) | ( n1367 & n5688 ) | ( ~n4559 & n5688 ) ;
  assign n15272 = ( n3013 & ~n4092 ) | ( n3013 & n15271 ) | ( ~n4092 & n15271 ) ;
  assign n15269 = n4074 ^ n1501 ^ 1'b0 ;
  assign n15270 = n15269 ^ n14915 ^ n10484 ;
  assign n15273 = n15272 ^ n15270 ^ n4668 ;
  assign n15274 = ( n1790 & ~n9395 ) | ( n1790 & n12139 ) | ( ~n9395 & n12139 ) ;
  assign n15275 = n15274 ^ n8503 ^ n3290 ;
  assign n15276 = n15275 ^ n2763 ^ 1'b0 ;
  assign n15277 = n15273 | n15276 ;
  assign n15279 = ( n3374 & ~n4090 ) | ( n3374 & n7161 ) | ( ~n4090 & n7161 ) ;
  assign n15278 = ( n2709 & n9034 ) | ( n2709 & n11753 ) | ( n9034 & n11753 ) ;
  assign n15280 = n15279 ^ n15278 ^ n11050 ;
  assign n15281 = ( n3216 & n3352 ) | ( n3216 & ~n4175 ) | ( n3352 & ~n4175 ) ;
  assign n15282 = ( n1474 & n2098 ) | ( n1474 & ~n15281 ) | ( n2098 & ~n15281 ) ;
  assign n15283 = n9367 | n15282 ;
  assign n15284 = n15283 ^ n14036 ^ 1'b0 ;
  assign n15285 = ( n1739 & ~n15280 ) | ( n1739 & n15284 ) | ( ~n15280 & n15284 ) ;
  assign n15286 = ( n1721 & n6179 ) | ( n1721 & n10982 ) | ( n6179 & n10982 ) ;
  assign n15287 = n5237 & n15286 ;
  assign n15288 = n15287 ^ n1146 ^ n357 ;
  assign n15289 = ( n3947 & n4460 ) | ( n3947 & n15288 ) | ( n4460 & n15288 ) ;
  assign n15290 = n2789 ^ n1962 ^ n1724 ;
  assign n15291 = n15290 ^ n12087 ^ n2237 ;
  assign n15292 = n7810 | n9217 ;
  assign n15293 = n5959 & ~n15292 ;
  assign n15294 = n15293 ^ n9277 ^ n4823 ;
  assign n15295 = n15294 ^ n12014 ^ n4025 ;
  assign n15296 = n10419 ^ n4583 ^ n403 ;
  assign n15297 = n15296 ^ n12587 ^ 1'b0 ;
  assign n15298 = n6942 & ~n8513 ;
  assign n15299 = n8090 & n15298 ;
  assign n15300 = n15299 ^ n6912 ^ 1'b0 ;
  assign n15301 = n6824 ^ n4368 ^ n2865 ;
  assign n15302 = n15301 ^ n15164 ^ n4143 ;
  assign n15303 = ( n2250 & ~n3349 ) | ( n2250 & n6933 ) | ( ~n3349 & n6933 ) ;
  assign n15304 = ( ~n8092 & n11310 ) | ( ~n8092 & n15303 ) | ( n11310 & n15303 ) ;
  assign n15305 = n15304 ^ n5275 ^ 1'b0 ;
  assign n15306 = n15302 & ~n15305 ;
  assign n15307 = ~n12698 & n15306 ;
  assign n15308 = n15307 ^ n7333 ^ 1'b0 ;
  assign n15309 = n4677 ^ x7 ^ 1'b0 ;
  assign n15310 = n15309 ^ n5028 ^ n950 ;
  assign n15311 = n12693 ^ n10569 ^ n8002 ;
  assign n15312 = n15311 ^ n5510 ^ 1'b0 ;
  assign n15313 = n11140 ^ n10879 ^ 1'b0 ;
  assign n15314 = n14218 ^ n6317 ^ 1'b0 ;
  assign n15315 = ( n12275 & n15313 ) | ( n12275 & n15314 ) | ( n15313 & n15314 ) ;
  assign n15316 = n6632 ^ n4644 ^ n666 ;
  assign n15317 = n11513 | n15316 ;
  assign n15320 = n5734 ^ n3360 ^ n3337 ;
  assign n15318 = ( n2073 & n3603 ) | ( n2073 & ~n7040 ) | ( n3603 & ~n7040 ) ;
  assign n15319 = n4298 | n15318 ;
  assign n15321 = n15320 ^ n15319 ^ 1'b0 ;
  assign n15322 = ( ~n365 & n6425 ) | ( ~n365 & n15269 ) | ( n6425 & n15269 ) ;
  assign n15323 = n3368 & n14794 ;
  assign n15324 = n15322 & n15323 ;
  assign n15325 = ( n4591 & ~n4935 ) | ( n4591 & n11872 ) | ( ~n4935 & n11872 ) ;
  assign n15326 = n11826 & ~n15325 ;
  assign n15327 = n15324 & n15326 ;
  assign n15328 = n1422 & ~n10521 ;
  assign n15329 = n4155 ^ n1337 ^ n400 ;
  assign n15330 = n361 | n8652 ;
  assign n15331 = n14152 ^ n1183 ^ x159 ;
  assign n15332 = ( n7085 & n13325 ) | ( n7085 & n15331 ) | ( n13325 & n15331 ) ;
  assign n15334 = ( n1356 & ~n6383 ) | ( n1356 & n7443 ) | ( ~n6383 & n7443 ) ;
  assign n15335 = n6904 ^ n1629 ^ 1'b0 ;
  assign n15336 = n15334 & n15335 ;
  assign n15333 = ~n4869 & n5794 ;
  assign n15337 = n15336 ^ n15333 ^ 1'b0 ;
  assign n15339 = n13176 ^ n5988 ^ x123 ;
  assign n15338 = ( n4497 & ~n5754 ) | ( n4497 & n10228 ) | ( ~n5754 & n10228 ) ;
  assign n15340 = n15339 ^ n15338 ^ n6294 ;
  assign n15341 = n5436 & n12229 ;
  assign n15342 = n12199 & n15341 ;
  assign n15343 = n12299 & ~n12375 ;
  assign n15344 = ( n1264 & n5472 ) | ( n1264 & n9781 ) | ( n5472 & n9781 ) ;
  assign n15345 = n15344 ^ n12533 ^ 1'b0 ;
  assign n15346 = n290 | n15345 ;
  assign n15347 = n6706 ^ n4415 ^ n3405 ;
  assign n15348 = ( n1029 & n7523 ) | ( n1029 & n15347 ) | ( n7523 & n15347 ) ;
  assign n15349 = n15348 ^ n4933 ^ 1'b0 ;
  assign n15350 = n15349 ^ n5571 ^ n4877 ;
  assign n15351 = ( ~n4636 & n15346 ) | ( ~n4636 & n15350 ) | ( n15346 & n15350 ) ;
  assign n15352 = ( n14090 & n15343 ) | ( n14090 & n15351 ) | ( n15343 & n15351 ) ;
  assign n15358 = ( n7352 & n7561 ) | ( n7352 & ~n11059 ) | ( n7561 & ~n11059 ) ;
  assign n15353 = ( n3340 & n10444 ) | ( n3340 & ~n11674 ) | ( n10444 & ~n11674 ) ;
  assign n15354 = n1857 ^ n1111 ^ n412 ;
  assign n15355 = ~n319 & n15354 ;
  assign n15356 = n15353 & n15355 ;
  assign n15357 = ( n7988 & n8173 ) | ( n7988 & n15356 ) | ( n8173 & n15356 ) ;
  assign n15359 = n15358 ^ n15357 ^ n671 ;
  assign n15360 = ( ~n1519 & n3441 ) | ( ~n1519 & n7808 ) | ( n3441 & n7808 ) ;
  assign n15361 = n9280 & n15360 ;
  assign n15362 = n11312 & n15361 ;
  assign n15363 = ( n3574 & n10998 ) | ( n3574 & ~n15362 ) | ( n10998 & ~n15362 ) ;
  assign n15364 = n2563 ^ n2034 ^ x166 ;
  assign n15365 = n11688 ^ n2171 ^ 1'b0 ;
  assign n15366 = n11740 & ~n15365 ;
  assign n15367 = ( n9555 & n15364 ) | ( n9555 & n15366 ) | ( n15364 & n15366 ) ;
  assign n15375 = n763 | n10359 ;
  assign n15376 = n15375 ^ n5727 ^ 1'b0 ;
  assign n15370 = n14645 ^ n7563 ^ n5906 ;
  assign n15371 = ( n2971 & ~n13881 ) | ( n2971 & n15370 ) | ( ~n13881 & n15370 ) ;
  assign n15372 = n15371 ^ n4063 ^ 1'b0 ;
  assign n15373 = n7619 & ~n15372 ;
  assign n15368 = n10510 ^ n5580 ^ n5077 ;
  assign n15369 = ( n2280 & ~n14301 ) | ( n2280 & n15368 ) | ( ~n14301 & n15368 ) ;
  assign n15374 = n15373 ^ n15369 ^ n8686 ;
  assign n15377 = n15376 ^ n15374 ^ n6852 ;
  assign n15378 = ( n975 & ~n4273 ) | ( n975 & n4693 ) | ( ~n4273 & n4693 ) ;
  assign n15379 = n15378 ^ n4552 ^ n3354 ;
  assign n15380 = n426 & n15379 ;
  assign n15381 = n15380 ^ n3483 ^ 1'b0 ;
  assign n15382 = n1723 & n8359 ;
  assign n15383 = n15381 & n15382 ;
  assign n15384 = n9849 ^ n3050 ^ n2873 ;
  assign n15385 = n9964 ^ n8923 ^ n6709 ;
  assign n15386 = n6226 ^ n3983 ^ 1'b0 ;
  assign n15387 = ~n13960 & n15386 ;
  assign n15388 = ( n7531 & ~n10932 ) | ( n7531 & n15387 ) | ( ~n10932 & n15387 ) ;
  assign n15389 = ( n3294 & ~n15385 ) | ( n3294 & n15388 ) | ( ~n15385 & n15388 ) ;
  assign n15399 = n2901 ^ n1968 ^ n1852 ;
  assign n15398 = n3899 ^ n3763 ^ 1'b0 ;
  assign n15390 = n5249 | n6993 ;
  assign n15391 = ( n4626 & ~n5463 ) | ( n4626 & n15390 ) | ( ~n5463 & n15390 ) ;
  assign n15392 = n15391 ^ n3096 ^ n2827 ;
  assign n15393 = n6779 ^ n5160 ^ n1916 ;
  assign n15394 = n15393 ^ n12953 ^ n2730 ;
  assign n15395 = n15394 ^ n14662 ^ n2752 ;
  assign n15396 = ( n3617 & n3696 ) | ( n3617 & ~n12539 ) | ( n3696 & ~n12539 ) ;
  assign n15397 = ( ~n15392 & n15395 ) | ( ~n15392 & n15396 ) | ( n15395 & n15396 ) ;
  assign n15400 = n15399 ^ n15398 ^ n15397 ;
  assign n15401 = ( ~n1250 & n2704 ) | ( ~n1250 & n13278 ) | ( n2704 & n13278 ) ;
  assign n15402 = n6625 & ~n7875 ;
  assign n15403 = n15402 ^ n6933 ^ x198 ;
  assign n15404 = n15403 ^ n13452 ^ n7386 ;
  assign n15409 = n7297 ^ n4182 ^ n1704 ;
  assign n15407 = n3964 ^ n3047 ^ n2620 ;
  assign n15406 = ( ~n2858 & n3402 ) | ( ~n2858 & n6232 ) | ( n3402 & n6232 ) ;
  assign n15408 = n15407 ^ n15406 ^ n6021 ;
  assign n15405 = ~n582 & n5175 ;
  assign n15410 = n15409 ^ n15408 ^ n15405 ;
  assign n15411 = ( n452 & n1322 ) | ( n452 & n4120 ) | ( n1322 & n4120 ) ;
  assign n15412 = n15411 ^ n4973 ^ n4209 ;
  assign n15413 = n15412 ^ n10388 ^ n3697 ;
  assign n15414 = n7973 ^ n7880 ^ n1534 ;
  assign n15415 = n11237 & ~n15414 ;
  assign n15416 = n15415 ^ n1717 ^ 1'b0 ;
  assign n15417 = ~n688 & n2437 ;
  assign n15424 = ~n464 & n7000 ;
  assign n15425 = n3210 & n15424 ;
  assign n15423 = ( n3798 & n5373 ) | ( n3798 & n10112 ) | ( n5373 & n10112 ) ;
  assign n15419 = ( n1837 & n1869 ) | ( n1837 & ~n2137 ) | ( n1869 & ~n2137 ) ;
  assign n15420 = n15419 ^ n9341 ^ 1'b0 ;
  assign n15421 = ( ~n7083 & n11724 ) | ( ~n7083 & n15420 ) | ( n11724 & n15420 ) ;
  assign n15418 = n4474 | n13057 ;
  assign n15422 = n15421 ^ n15418 ^ 1'b0 ;
  assign n15426 = n15425 ^ n15423 ^ n15422 ;
  assign n15427 = ( n2397 & n4533 ) | ( n2397 & ~n7431 ) | ( n4533 & ~n7431 ) ;
  assign n15428 = x151 & ~n15427 ;
  assign n15429 = n1669 | n3852 ;
  assign n15430 = n2114 & ~n15429 ;
  assign n15431 = n15430 ^ n9431 ^ n1900 ;
  assign n15432 = ( n8804 & n11964 ) | ( n8804 & ~n14075 ) | ( n11964 & ~n14075 ) ;
  assign n15433 = n15432 ^ n12972 ^ n1630 ;
  assign n15434 = n12594 ^ n3203 ^ x172 ;
  assign n15435 = ( n12984 & ~n13725 ) | ( n12984 & n15434 ) | ( ~n13725 & n15434 ) ;
  assign n15436 = n15435 ^ n15212 ^ n14326 ;
  assign n15437 = ( n15431 & ~n15433 ) | ( n15431 & n15436 ) | ( ~n15433 & n15436 ) ;
  assign n15438 = n2799 | n3207 ;
  assign n15439 = n15438 ^ n2427 ^ 1'b0 ;
  assign n15440 = ( n1709 & n5739 ) | ( n1709 & n15439 ) | ( n5739 & n15439 ) ;
  assign n15441 = n1160 & n15440 ;
  assign n15442 = n1569 & n15441 ;
  assign n15443 = ( n867 & ~n2891 ) | ( n867 & n10301 ) | ( ~n2891 & n10301 ) ;
  assign n15444 = n12516 ^ n5400 ^ x170 ;
  assign n15445 = n15444 ^ n5734 ^ n1953 ;
  assign n15446 = ( n3318 & n15443 ) | ( n3318 & ~n15445 ) | ( n15443 & ~n15445 ) ;
  assign n15447 = ( n6081 & ~n7088 ) | ( n6081 & n15446 ) | ( ~n7088 & n15446 ) ;
  assign n15448 = n6361 ^ n860 ^ x219 ;
  assign n15449 = n7963 | n15448 ;
  assign n15451 = n2525 ^ n2066 ^ n1103 ;
  assign n15450 = n9966 ^ n3826 ^ 1'b0 ;
  assign n15452 = n15451 ^ n15450 ^ 1'b0 ;
  assign n15453 = ( n2197 & n4646 ) | ( n2197 & n4704 ) | ( n4646 & n4704 ) ;
  assign n15454 = ( n763 & n2833 ) | ( n763 & n6038 ) | ( n2833 & n6038 ) ;
  assign n15455 = n15454 ^ n11846 ^ n1928 ;
  assign n15456 = n15455 ^ n13939 ^ n2965 ;
  assign n15457 = n13254 & ~n15456 ;
  assign n15458 = n14861 ^ n4229 ^ n1339 ;
  assign n15459 = n2188 & ~n6058 ;
  assign n15460 = n8565 & n15459 ;
  assign n15461 = n10682 ^ n8215 ^ n4315 ;
  assign n15462 = ( n9453 & n10703 ) | ( n9453 & ~n15461 ) | ( n10703 & ~n15461 ) ;
  assign n15463 = ( n11064 & ~n12354 ) | ( n11064 & n15462 ) | ( ~n12354 & n15462 ) ;
  assign n15464 = ~n15460 & n15463 ;
  assign n15465 = n15464 ^ n11337 ^ 1'b0 ;
  assign n15466 = ~n7232 & n14018 ;
  assign n15467 = ~x88 & n15466 ;
  assign n15468 = n7253 ^ n2896 ^ n1952 ;
  assign n15469 = ( n4670 & ~n5183 ) | ( n4670 & n15468 ) | ( ~n5183 & n15468 ) ;
  assign n15470 = ( ~n4991 & n13839 ) | ( ~n4991 & n15469 ) | ( n13839 & n15469 ) ;
  assign n15471 = n3709 & ~n6689 ;
  assign n15472 = ( ~n1298 & n4699 ) | ( ~n1298 & n6820 ) | ( n4699 & n6820 ) ;
  assign n15483 = n5448 ^ n4562 ^ n665 ;
  assign n15482 = ( n773 & n1945 ) | ( n773 & n8229 ) | ( n1945 & n8229 ) ;
  assign n15481 = ( n1478 & ~n1912 ) | ( n1478 & n13556 ) | ( ~n1912 & n13556 ) ;
  assign n15484 = n15483 ^ n15482 ^ n15481 ;
  assign n15474 = n7842 ^ n4150 ^ n793 ;
  assign n15475 = n15474 ^ n3662 ^ 1'b0 ;
  assign n15476 = ( n7700 & n8973 ) | ( n7700 & ~n15475 ) | ( n8973 & ~n15475 ) ;
  assign n15477 = n9254 | n10417 ;
  assign n15478 = n15477 ^ n882 ^ 1'b0 ;
  assign n15479 = ~n9170 & n15478 ;
  assign n15480 = ( ~n1212 & n15476 ) | ( ~n1212 & n15479 ) | ( n15476 & n15479 ) ;
  assign n15473 = n7796 ^ n2176 ^ 1'b0 ;
  assign n15485 = n15484 ^ n15480 ^ n15473 ;
  assign n15489 = ( n551 & ~n716 ) | ( n551 & n2429 ) | ( ~n716 & n2429 ) ;
  assign n15490 = n658 | n15489 ;
  assign n15491 = n915 | n15490 ;
  assign n15486 = n14322 ^ n6290 ^ 1'b0 ;
  assign n15487 = n2545 | n15486 ;
  assign n15488 = ( n1866 & n13826 ) | ( n1866 & n15487 ) | ( n13826 & n15487 ) ;
  assign n15492 = n15491 ^ n15488 ^ n10779 ;
  assign n15493 = n9381 & n10477 ;
  assign n15494 = n15492 & n15493 ;
  assign n15495 = n15494 ^ n4021 ^ 1'b0 ;
  assign n15496 = n10154 ^ n7963 ^ n1352 ;
  assign n15497 = n15496 ^ n14262 ^ n8245 ;
  assign n15502 = n6803 & ~n7324 ;
  assign n15503 = n15502 ^ n10840 ^ 1'b0 ;
  assign n15499 = n11351 ^ n2458 ^ n1620 ;
  assign n15500 = n10354 ^ n3833 ^ n1446 ;
  assign n15501 = ( ~n6106 & n15499 ) | ( ~n6106 & n15500 ) | ( n15499 & n15500 ) ;
  assign n15498 = ( n11553 & ~n11753 ) | ( n11553 & n13513 ) | ( ~n11753 & n13513 ) ;
  assign n15504 = n15503 ^ n15501 ^ n15498 ;
  assign n15505 = n1551 & n3269 ;
  assign n15506 = n15505 ^ n12578 ^ n8100 ;
  assign n15507 = n15506 ^ n8258 ^ n5679 ;
  assign n15508 = n14353 ^ n7583 ^ 1'b0 ;
  assign n15509 = n15507 & n15508 ;
  assign n15510 = ( ~n6685 & n15504 ) | ( ~n6685 & n15509 ) | ( n15504 & n15509 ) ;
  assign n15511 = n6368 ^ n1698 ^ n1440 ;
  assign n15512 = ( n4590 & n9949 ) | ( n4590 & n15511 ) | ( n9949 & n15511 ) ;
  assign n15513 = ( n5130 & ~n10002 ) | ( n5130 & n15512 ) | ( ~n10002 & n15512 ) ;
  assign n15514 = n14339 ^ n7237 ^ n1481 ;
  assign n15521 = ~n1042 & n4287 ;
  assign n15517 = n9229 ^ n7592 ^ 1'b0 ;
  assign n15518 = n8341 & n15517 ;
  assign n15516 = ( n526 & ~n1731 ) | ( n526 & n5227 ) | ( ~n1731 & n5227 ) ;
  assign n15519 = n15518 ^ n15516 ^ n6578 ;
  assign n15520 = n15519 ^ n9076 ^ x66 ;
  assign n15522 = n15521 ^ n15520 ^ n8107 ;
  assign n15515 = ( n5842 & ~n10918 ) | ( n5842 & n14412 ) | ( ~n10918 & n14412 ) ;
  assign n15523 = n15522 ^ n15515 ^ n2112 ;
  assign n15524 = ( n10401 & n15514 ) | ( n10401 & ~n15523 ) | ( n15514 & ~n15523 ) ;
  assign n15525 = n7557 | n15524 ;
  assign n15526 = ( ~n2726 & n10174 ) | ( ~n2726 & n13344 ) | ( n10174 & n13344 ) ;
  assign n15527 = n15526 ^ n13176 ^ n7178 ;
  assign n15528 = n12721 ^ n11626 ^ n7689 ;
  assign n15529 = n15528 ^ n14681 ^ n9868 ;
  assign n15536 = ( n1010 & n1131 ) | ( n1010 & n4051 ) | ( n1131 & n4051 ) ;
  assign n15530 = n8720 ^ n4222 ^ x124 ;
  assign n15531 = n4085 ^ n1624 ^ 1'b0 ;
  assign n15532 = ~n601 & n15531 ;
  assign n15533 = n15532 ^ n13863 ^ n11277 ;
  assign n15534 = n15533 ^ n2211 ^ 1'b0 ;
  assign n15535 = ( x106 & n15530 ) | ( x106 & n15534 ) | ( n15530 & n15534 ) ;
  assign n15537 = n15536 ^ n15535 ^ n7055 ;
  assign n15538 = n1582 | n2693 ;
  assign n15539 = n6431 | n15538 ;
  assign n15542 = n7454 ^ n3793 ^ x103 ;
  assign n15543 = n15542 ^ n3096 ^ n1651 ;
  assign n15540 = n1077 ^ n615 ^ 1'b0 ;
  assign n15541 = n15540 ^ n9009 ^ n5281 ;
  assign n15544 = n15543 ^ n15541 ^ n8045 ;
  assign n15545 = ( n1811 & n3427 ) | ( n1811 & ~n4753 ) | ( n3427 & ~n4753 ) ;
  assign n15546 = ~n1961 & n2726 ;
  assign n15547 = ~n3543 & n15546 ;
  assign n15548 = n9220 ^ n3533 ^ n1590 ;
  assign n15549 = ~n6946 & n15548 ;
  assign n15550 = n15547 & n15549 ;
  assign n15551 = ( n3247 & ~n15545 ) | ( n3247 & n15550 ) | ( ~n15545 & n15550 ) ;
  assign n15553 = n15072 ^ n9861 ^ n8433 ;
  assign n15556 = n13777 & ~n15355 ;
  assign n15557 = n15556 ^ x224 ^ 1'b0 ;
  assign n15555 = n6914 | n7109 ;
  assign n15558 = n15557 ^ n15555 ^ 1'b0 ;
  assign n15554 = n6535 & ~n10140 ;
  assign n15559 = n15558 ^ n15554 ^ n2440 ;
  assign n15560 = n15553 | n15559 ;
  assign n15552 = ~n3783 & n12267 ;
  assign n15561 = n15560 ^ n15552 ^ 1'b0 ;
  assign n15562 = ( n566 & n5486 ) | ( n566 & ~n9060 ) | ( n5486 & ~n9060 ) ;
  assign n15563 = n13433 | n15562 ;
  assign n15564 = ( n1112 & ~n5278 ) | ( n1112 & n14750 ) | ( ~n5278 & n14750 ) ;
  assign n15565 = ( n4535 & n10922 ) | ( n4535 & ~n15564 ) | ( n10922 & ~n15564 ) ;
  assign n15566 = n15565 ^ n10402 ^ n9608 ;
  assign n15567 = n5409 & ~n15566 ;
  assign n15568 = n5012 ^ n2403 ^ x141 ;
  assign n15569 = ~n1684 & n9567 ;
  assign n15570 = n15569 ^ n1411 ^ 1'b0 ;
  assign n15571 = n15570 ^ n9409 ^ 1'b0 ;
  assign n15572 = n1185 & ~n15571 ;
  assign n15573 = ~n15568 & n15572 ;
  assign n15576 = n3652 ^ n2871 ^ 1'b0 ;
  assign n15575 = n12482 ^ n10985 ^ n7078 ;
  assign n15574 = n9418 ^ n3620 ^ n1708 ;
  assign n15577 = n15576 ^ n15575 ^ n15574 ;
  assign n15578 = n10985 ^ n4664 ^ 1'b0 ;
  assign n15579 = n7986 | n15578 ;
  assign n15580 = ( ~n3622 & n6550 ) | ( ~n3622 & n7770 ) | ( n6550 & n7770 ) ;
  assign n15581 = ( n2143 & ~n4247 ) | ( n2143 & n4906 ) | ( ~n4247 & n4906 ) ;
  assign n15582 = ( ~n2415 & n11232 ) | ( ~n2415 & n15581 ) | ( n11232 & n15581 ) ;
  assign n15583 = ( n13857 & n15580 ) | ( n13857 & n15582 ) | ( n15580 & n15582 ) ;
  assign n15584 = n15583 ^ n2348 ^ 1'b0 ;
  assign n15585 = ~n15579 & n15584 ;
  assign n15586 = n10849 ^ n7109 ^ 1'b0 ;
  assign n15587 = ( n10009 & n12733 ) | ( n10009 & n15586 ) | ( n12733 & n15586 ) ;
  assign n15588 = ( n6817 & ~n8457 ) | ( n6817 & n15587 ) | ( ~n8457 & n15587 ) ;
  assign n15589 = ~n1932 & n15588 ;
  assign n15590 = n15589 ^ n5438 ^ 1'b0 ;
  assign n15591 = n12945 ^ n9017 ^ n2984 ;
  assign n15592 = n4866 | n6711 ;
  assign n15593 = ~x6 & x123 ;
  assign n15594 = ( n990 & n1398 ) | ( n990 & ~n15593 ) | ( n1398 & ~n15593 ) ;
  assign n15595 = n10804 & n15594 ;
  assign n15596 = ~n15592 & n15595 ;
  assign n15597 = n13982 ^ n10617 ^ 1'b0 ;
  assign n15598 = ( n9077 & ~n15596 ) | ( n9077 & n15597 ) | ( ~n15596 & n15597 ) ;
  assign n15599 = n15598 ^ n13132 ^ n9421 ;
  assign n15600 = ( n2257 & ~n7950 ) | ( n2257 & n14518 ) | ( ~n7950 & n14518 ) ;
  assign n15601 = n3064 | n4347 ;
  assign n15602 = n15601 ^ n11169 ^ n9836 ;
  assign n15603 = ( n1595 & n15600 ) | ( n1595 & ~n15602 ) | ( n15600 & ~n15602 ) ;
  assign n15604 = n11517 ^ n9969 ^ n7007 ;
  assign n15605 = n15604 ^ n4321 ^ 1'b0 ;
  assign n15606 = ~n5689 & n15605 ;
  assign n15609 = ~n787 & n10139 ;
  assign n15607 = ( n412 & n1264 ) | ( n412 & ~n7011 ) | ( n1264 & ~n7011 ) ;
  assign n15608 = n15607 ^ n6886 ^ n1755 ;
  assign n15610 = n15609 ^ n15608 ^ n2592 ;
  assign n15613 = n7963 ^ n4995 ^ n2241 ;
  assign n15612 = ( n6746 & ~n7925 ) | ( n6746 & n10783 ) | ( ~n7925 & n10783 ) ;
  assign n15611 = ( n9666 & n10001 ) | ( n9666 & n11828 ) | ( n10001 & n11828 ) ;
  assign n15614 = n15613 ^ n15612 ^ n15611 ;
  assign n15615 = ( ~n2585 & n15610 ) | ( ~n2585 & n15614 ) | ( n15610 & n15614 ) ;
  assign n15616 = ( n11084 & n15606 ) | ( n11084 & ~n15615 ) | ( n15606 & ~n15615 ) ;
  assign n15617 = ( ~x56 & x68 ) | ( ~x56 & n2062 ) | ( x68 & n2062 ) ;
  assign n15618 = ( n3503 & n6813 ) | ( n3503 & n15617 ) | ( n6813 & n15617 ) ;
  assign n15619 = n11111 ^ n331 ^ 1'b0 ;
  assign n15620 = n15619 ^ n3379 ^ n2092 ;
  assign n15621 = ( n7170 & n15618 ) | ( n7170 & n15620 ) | ( n15618 & n15620 ) ;
  assign n15622 = ( n1638 & n1719 ) | ( n1638 & n3982 ) | ( n1719 & n3982 ) ;
  assign n15623 = ( n3419 & n11744 ) | ( n3419 & n15622 ) | ( n11744 & n15622 ) ;
  assign n15624 = n14776 ^ n6984 ^ n2111 ;
  assign n15625 = n15623 & n15624 ;
  assign n15626 = n1726 | n15625 ;
  assign n15627 = n15621 & ~n15626 ;
  assign n15628 = ( n1574 & ~n5645 ) | ( n1574 & n14517 ) | ( ~n5645 & n14517 ) ;
  assign n15629 = n15628 ^ n12037 ^ n7617 ;
  assign n15632 = n13021 ^ n7842 ^ 1'b0 ;
  assign n15630 = n7415 ^ n3813 ^ 1'b0 ;
  assign n15631 = x227 & n15630 ;
  assign n15633 = n15632 ^ n15631 ^ n1223 ;
  assign n15635 = ( n3572 & n3980 ) | ( n3572 & n4607 ) | ( n3980 & n4607 ) ;
  assign n15636 = n15635 ^ n6258 ^ 1'b0 ;
  assign n15634 = ( n685 & n5252 ) | ( n685 & n11684 ) | ( n5252 & n11684 ) ;
  assign n15637 = n15636 ^ n15634 ^ n5739 ;
  assign n15647 = n5465 | n7781 ;
  assign n15648 = n15647 ^ n1835 ^ 1'b0 ;
  assign n15649 = ( ~n312 & n9769 ) | ( ~n312 & n15648 ) | ( n9769 & n15648 ) ;
  assign n15650 = ( ~n3606 & n5700 ) | ( ~n3606 & n15649 ) | ( n5700 & n15649 ) ;
  assign n15638 = n13363 ^ n9407 ^ n7064 ;
  assign n15639 = n1389 | n15638 ;
  assign n15640 = n15639 ^ n7955 ^ 1'b0 ;
  assign n15641 = n4939 & n10584 ;
  assign n15642 = ~n2671 & n15641 ;
  assign n15643 = n15642 ^ n1828 ^ 1'b0 ;
  assign n15644 = ( n1227 & n4049 ) | ( n1227 & ~n15643 ) | ( n4049 & ~n15643 ) ;
  assign n15645 = n15644 ^ n4853 ^ n1405 ;
  assign n15646 = n15640 & n15645 ;
  assign n15651 = n15650 ^ n15646 ^ n14813 ;
  assign n15653 = n5164 ^ n585 ^ 1'b0 ;
  assign n15652 = n13251 ^ n4632 ^ n1008 ;
  assign n15654 = n15653 ^ n15652 ^ n6972 ;
  assign n15657 = n4793 ^ n2309 ^ n473 ;
  assign n15655 = n14525 ^ n6430 ^ n3860 ;
  assign n15656 = ( ~n2911 & n10853 ) | ( ~n2911 & n15655 ) | ( n10853 & n15655 ) ;
  assign n15658 = n15657 ^ n15656 ^ 1'b0 ;
  assign n15659 = n7408 & n15658 ;
  assign n15660 = ( n5691 & ~n9671 ) | ( n5691 & n15659 ) | ( ~n9671 & n15659 ) ;
  assign n15661 = n13997 ^ n12591 ^ n11944 ;
  assign n15662 = n6500 | n9951 ;
  assign n15663 = n15662 ^ n2153 ^ n1738 ;
  assign n15664 = n10219 & n15663 ;
  assign n15665 = ( ~n9332 & n15661 ) | ( ~n9332 & n15664 ) | ( n15661 & n15664 ) ;
  assign n15666 = n3848 ^ n3451 ^ n326 ;
  assign n15667 = ( n2035 & n7012 ) | ( n2035 & ~n13804 ) | ( n7012 & ~n13804 ) ;
  assign n15668 = n15666 & ~n15667 ;
  assign n15669 = n15668 ^ n11270 ^ 1'b0 ;
  assign n15670 = n15669 ^ n6870 ^ x203 ;
  assign n15671 = ( n1951 & ~n11697 ) | ( n1951 & n14253 ) | ( ~n11697 & n14253 ) ;
  assign n15677 = ( n1509 & n2226 ) | ( n1509 & n14007 ) | ( n2226 & n14007 ) ;
  assign n15678 = ( n5886 & n7927 ) | ( n5886 & ~n15677 ) | ( n7927 & ~n15677 ) ;
  assign n15672 = n5188 ^ n3813 ^ 1'b0 ;
  assign n15673 = n4432 & ~n15672 ;
  assign n15674 = ( n1550 & ~n7792 ) | ( n1550 & n15673 ) | ( ~n7792 & n15673 ) ;
  assign n15675 = ( ~n8658 & n13960 ) | ( ~n8658 & n15674 ) | ( n13960 & n15674 ) ;
  assign n15676 = n8346 & ~n15675 ;
  assign n15679 = n15678 ^ n15676 ^ 1'b0 ;
  assign n15680 = n9576 ^ n2572 ^ n2005 ;
  assign n15681 = ( n1479 & ~n9383 ) | ( n1479 & n15680 ) | ( ~n9383 & n15680 ) ;
  assign n15682 = n2418 & ~n11540 ;
  assign n15683 = n12607 & n15682 ;
  assign n15685 = n13952 ^ n1507 ^ n1286 ;
  assign n15684 = n3691 & n7384 ;
  assign n15686 = n15685 ^ n15684 ^ 1'b0 ;
  assign n15687 = ( n2080 & n3989 ) | ( n2080 & ~n7598 ) | ( n3989 & ~n7598 ) ;
  assign n15690 = n7351 ^ n3158 ^ n495 ;
  assign n15691 = n15690 ^ n12716 ^ n6919 ;
  assign n15692 = n8784 | n15691 ;
  assign n15688 = n9281 ^ n4793 ^ 1'b0 ;
  assign n15689 = ~n4143 & n15688 ;
  assign n15693 = n15692 ^ n15689 ^ n8160 ;
  assign n15694 = n9586 ^ n1159 ^ 1'b0 ;
  assign n15695 = ~n15693 & n15694 ;
  assign n15696 = n5602 | n8022 ;
  assign n15697 = n15696 ^ n8148 ^ 1'b0 ;
  assign n15698 = ( n1200 & n5470 ) | ( n1200 & n14494 ) | ( n5470 & n14494 ) ;
  assign n15699 = n13834 & ~n15235 ;
  assign n15700 = n15699 ^ n11645 ^ 1'b0 ;
  assign n15706 = n14840 ^ n5606 ^ n1372 ;
  assign n15707 = n1601 & ~n11784 ;
  assign n15708 = n15706 & n15707 ;
  assign n15703 = ( ~n628 & n5158 ) | ( ~n628 & n12839 ) | ( n5158 & n12839 ) ;
  assign n15702 = n13903 ^ n8365 ^ n5525 ;
  assign n15704 = n15703 ^ n15702 ^ 1'b0 ;
  assign n15701 = ( n12570 & n13494 ) | ( n12570 & ~n13571 ) | ( n13494 & ~n13571 ) ;
  assign n15705 = n15704 ^ n15701 ^ n13971 ;
  assign n15709 = n15708 ^ n15705 ^ n10856 ;
  assign n15720 = n12741 ^ n1383 ^ n608 ;
  assign n15715 = ( n1478 & ~n2446 ) | ( n1478 & n5044 ) | ( ~n2446 & n5044 ) ;
  assign n15716 = n15715 ^ n8013 ^ n7698 ;
  assign n15717 = ( n5807 & n7828 ) | ( n5807 & ~n15716 ) | ( n7828 & ~n15716 ) ;
  assign n15718 = ( n2125 & n8852 ) | ( n2125 & n15717 ) | ( n8852 & n15717 ) ;
  assign n15713 = ( n5314 & n6433 ) | ( n5314 & ~n11517 ) | ( n6433 & ~n11517 ) ;
  assign n15714 = n15713 ^ n4168 ^ 1'b0 ;
  assign n15719 = n15718 ^ n15714 ^ n9430 ;
  assign n15710 = ( n3375 & n4325 ) | ( n3375 & n4784 ) | ( n4325 & n4784 ) ;
  assign n15711 = n15710 ^ n14795 ^ 1'b0 ;
  assign n15712 = n15711 ^ n9782 ^ n5902 ;
  assign n15721 = n15720 ^ n15719 ^ n15712 ;
  assign n15727 = n455 | n4237 ;
  assign n15722 = n3769 | n4618 ;
  assign n15723 = n15722 ^ n3249 ^ 1'b0 ;
  assign n15724 = n15723 ^ n7090 ^ n5265 ;
  assign n15725 = n15724 ^ n4841 ^ n1891 ;
  assign n15726 = n15725 ^ n6636 ^ n4977 ;
  assign n15728 = n15727 ^ n15726 ^ n12032 ;
  assign n15729 = n6031 & ~n12153 ;
  assign n15735 = n853 & n1481 ;
  assign n15736 = n10425 & n15735 ;
  assign n15733 = ( n1186 & n1849 ) | ( n1186 & ~n3434 ) | ( n1849 & ~n3434 ) ;
  assign n15732 = n11497 ^ n983 ^ 1'b0 ;
  assign n15734 = n15733 ^ n15732 ^ n761 ;
  assign n15730 = n1588 | n6328 ;
  assign n15731 = n15730 ^ n6374 ^ 1'b0 ;
  assign n15737 = n15736 ^ n15734 ^ n15731 ;
  assign n15738 = n10316 | n15269 ;
  assign n15739 = n4237 | n15738 ;
  assign n15740 = n15739 ^ n7248 ^ n3681 ;
  assign n15741 = n9566 ^ n8115 ^ n7083 ;
  assign n15742 = ( n7349 & n8369 ) | ( n7349 & n15741 ) | ( n8369 & n15741 ) ;
  assign n15743 = n4566 & n12616 ;
  assign n15744 = ( ~n15740 & n15742 ) | ( ~n15740 & n15743 ) | ( n15742 & n15743 ) ;
  assign n15745 = ( x68 & n3836 ) | ( x68 & ~n13050 ) | ( n3836 & ~n13050 ) ;
  assign n15746 = n15745 ^ n5793 ^ 1'b0 ;
  assign n15747 = n5269 & n15746 ;
  assign n15748 = n11309 ^ n10009 ^ n9401 ;
  assign n15749 = n4224 ^ n2782 ^ n1241 ;
  assign n15750 = n10778 ^ n1056 ^ n492 ;
  assign n15751 = ( n3839 & ~n15749 ) | ( n3839 & n15750 ) | ( ~n15749 & n15750 ) ;
  assign n15752 = n11858 ^ n8854 ^ n3576 ;
  assign n15754 = n5904 ^ n4529 ^ 1'b0 ;
  assign n15755 = n2515 | n15754 ;
  assign n15756 = ( n8845 & n11915 ) | ( n8845 & n15755 ) | ( n11915 & n15755 ) ;
  assign n15753 = ( n1533 & n9584 ) | ( n1533 & ~n11689 ) | ( n9584 & ~n11689 ) ;
  assign n15757 = n15756 ^ n15753 ^ n13461 ;
  assign n15758 = ( n6393 & ~n8618 ) | ( n6393 & n12200 ) | ( ~n8618 & n12200 ) ;
  assign n15759 = n15758 ^ n14799 ^ n7001 ;
  assign n15762 = n5269 ^ n468 ^ 1'b0 ;
  assign n15760 = n8886 ^ n3767 ^ n554 ;
  assign n15761 = n11816 | n15760 ;
  assign n15763 = n15762 ^ n15761 ^ 1'b0 ;
  assign n15764 = n1269 | n6276 ;
  assign n15765 = n15763 | n15764 ;
  assign n15766 = n15765 ^ n10912 ^ n4574 ;
  assign n15767 = ( ~n1541 & n15759 ) | ( ~n1541 & n15766 ) | ( n15759 & n15766 ) ;
  assign n15768 = ( n7216 & n7281 ) | ( n7216 & n12273 ) | ( n7281 & n12273 ) ;
  assign n15769 = n6881 & ~n10935 ;
  assign n15770 = n15769 ^ n7687 ^ 1'b0 ;
  assign n15771 = ~n12256 & n15770 ;
  assign n15781 = n1304 & ~n4151 ;
  assign n15779 = n3506 ^ x128 ^ 1'b0 ;
  assign n15780 = x80 & n15779 ;
  assign n15772 = n3142 ^ n2677 ^ n2217 ;
  assign n15773 = n7396 ^ n2602 ^ x20 ;
  assign n15774 = ( ~n1714 & n15349 ) | ( ~n1714 & n15773 ) | ( n15349 & n15773 ) ;
  assign n15775 = ( n8609 & ~n13752 ) | ( n8609 & n15774 ) | ( ~n13752 & n15774 ) ;
  assign n15776 = n1029 & n15775 ;
  assign n15777 = ( n13857 & n15772 ) | ( n13857 & ~n15776 ) | ( n15772 & ~n15776 ) ;
  assign n15778 = n15777 ^ n12813 ^ n1700 ;
  assign n15782 = n15781 ^ n15780 ^ n15778 ;
  assign n15783 = ( n15768 & ~n15771 ) | ( n15768 & n15782 ) | ( ~n15771 & n15782 ) ;
  assign n15784 = n4566 ^ n2025 ^ 1'b0 ;
  assign n15785 = n15784 ^ n7306 ^ 1'b0 ;
  assign n15786 = n6820 & ~n15785 ;
  assign n15788 = n263 | n10848 ;
  assign n15789 = ( n4063 & ~n4531 ) | ( n4063 & n15788 ) | ( ~n4531 & n15788 ) ;
  assign n15787 = n5066 & n8570 ;
  assign n15790 = n15789 ^ n15787 ^ 1'b0 ;
  assign n15791 = n15790 ^ n1736 ^ 1'b0 ;
  assign n15797 = ( n1396 & ~n7686 ) | ( n1396 & n11685 ) | ( ~n7686 & n11685 ) ;
  assign n15796 = n795 | n10881 ;
  assign n15793 = n1137 & n5929 ;
  assign n15792 = n6857 ^ n4758 ^ n2784 ;
  assign n15794 = n15793 ^ n15792 ^ 1'b0 ;
  assign n15795 = n13150 & ~n15794 ;
  assign n15798 = n15797 ^ n15796 ^ n15795 ;
  assign n15807 = ~n6022 & n15112 ;
  assign n15803 = ( n2068 & ~n3097 ) | ( n2068 & n3318 ) | ( ~n3097 & n3318 ) ;
  assign n15799 = n5332 ^ n682 ^ 1'b0 ;
  assign n15800 = ~n2582 & n15799 ;
  assign n15801 = ~n812 & n15800 ;
  assign n15802 = n15801 ^ n968 ^ 1'b0 ;
  assign n15804 = n15803 ^ n15802 ^ n3040 ;
  assign n15805 = n15804 ^ n11111 ^ 1'b0 ;
  assign n15806 = n2222 | n15805 ;
  assign n15808 = n15807 ^ n15806 ^ 1'b0 ;
  assign n15819 = ( n3780 & ~n10647 ) | ( n3780 & n11027 ) | ( ~n10647 & n11027 ) ;
  assign n15816 = n15356 ^ n5134 ^ 1'b0 ;
  assign n15817 = n5278 & ~n15816 ;
  assign n15809 = n6021 ^ n5131 ^ n4414 ;
  assign n15810 = n13411 ^ n2234 ^ n2025 ;
  assign n15811 = n15810 ^ n4092 ^ n625 ;
  assign n15812 = n15811 ^ n5500 ^ n4428 ;
  assign n15813 = ( n3108 & n7898 ) | ( n3108 & n15812 ) | ( n7898 & n15812 ) ;
  assign n15814 = ( ~n7028 & n12335 ) | ( ~n7028 & n15813 ) | ( n12335 & n15813 ) ;
  assign n15815 = n15809 | n15814 ;
  assign n15818 = n15817 ^ n15815 ^ n9877 ;
  assign n15820 = n15819 ^ n15818 ^ n2970 ;
  assign n15829 = ( n1005 & ~n2369 ) | ( n1005 & n11855 ) | ( ~n2369 & n11855 ) ;
  assign n15830 = n9465 & n15829 ;
  assign n15827 = ( ~n4373 & n10843 ) | ( ~n4373 & n12772 ) | ( n10843 & n12772 ) ;
  assign n15828 = ( ~n7825 & n9387 ) | ( ~n7825 & n15827 ) | ( n9387 & n15827 ) ;
  assign n15821 = ( n347 & ~n5584 ) | ( n347 & n13719 ) | ( ~n5584 & n13719 ) ;
  assign n15822 = ( n4018 & n4427 ) | ( n4018 & ~n15821 ) | ( n4427 & ~n15821 ) ;
  assign n15823 = ( n2410 & n3397 ) | ( n2410 & ~n7489 ) | ( n3397 & ~n7489 ) ;
  assign n15824 = n15823 ^ n8840 ^ n5400 ;
  assign n15825 = n15824 ^ n14246 ^ 1'b0 ;
  assign n15826 = n15822 & ~n15825 ;
  assign n15831 = n15830 ^ n15828 ^ n15826 ;
  assign n15832 = ( n1143 & ~n6123 ) | ( n1143 & n15272 ) | ( ~n6123 & n15272 ) ;
  assign n15833 = n13085 ^ n5587 ^ n4371 ;
  assign n15834 = ( n4960 & n11922 ) | ( n4960 & ~n15833 ) | ( n11922 & ~n15833 ) ;
  assign n15835 = ~n1547 & n15834 ;
  assign n15836 = n15835 ^ n3004 ^ 1'b0 ;
  assign n15837 = ( n6804 & ~n15832 ) | ( n6804 & n15836 ) | ( ~n15832 & n15836 ) ;
  assign n15847 = n12984 ^ n5564 ^ n2976 ;
  assign n15848 = n15847 ^ n9935 ^ n4883 ;
  assign n15849 = n15848 ^ n6351 ^ n2468 ;
  assign n15850 = ( ~n2932 & n13802 ) | ( ~n2932 & n15849 ) | ( n13802 & n15849 ) ;
  assign n15842 = n672 | n10888 ;
  assign n15843 = n15842 ^ n2486 ^ 1'b0 ;
  assign n15844 = n7561 ^ n5209 ^ n4131 ;
  assign n15845 = n15844 ^ n680 ^ x153 ;
  assign n15846 = ~n15843 & n15845 ;
  assign n15838 = ~n2737 & n8116 ;
  assign n15839 = n15838 ^ n7570 ^ 1'b0 ;
  assign n15840 = n15839 ^ n14554 ^ n2609 ;
  assign n15841 = n15840 ^ n1600 ^ 1'b0 ;
  assign n15851 = n15850 ^ n15846 ^ n15841 ;
  assign n15852 = n7554 ^ n1130 ^ n466 ;
  assign n15853 = ( n884 & n6347 ) | ( n884 & ~n15852 ) | ( n6347 & ~n15852 ) ;
  assign n15854 = n15853 ^ n15191 ^ n11726 ;
  assign n15855 = ( n2633 & n11825 ) | ( n2633 & ~n14980 ) | ( n11825 & ~n14980 ) ;
  assign n15856 = ( n7323 & n9553 ) | ( n7323 & ~n12577 ) | ( n9553 & ~n12577 ) ;
  assign n15857 = n13328 ^ n10479 ^ n8736 ;
  assign n15858 = n15857 ^ n4188 ^ 1'b0 ;
  assign n15859 = n13688 & n15858 ;
  assign n15868 = ( ~n8315 & n10484 ) | ( ~n8315 & n11273 ) | ( n10484 & n11273 ) ;
  assign n15860 = n6910 ^ n4310 ^ n1677 ;
  assign n15861 = n15860 ^ n11646 ^ n3977 ;
  assign n15862 = n5927 ^ n4131 ^ 1'b0 ;
  assign n15863 = n6342 | n15862 ;
  assign n15864 = n15863 ^ n4596 ^ 1'b0 ;
  assign n15865 = ( n7457 & n11372 ) | ( n7457 & ~n15864 ) | ( n11372 & ~n15864 ) ;
  assign n15866 = ( x160 & ~n15861 ) | ( x160 & n15865 ) | ( ~n15861 & n15865 ) ;
  assign n15867 = n15866 ^ n9720 ^ 1'b0 ;
  assign n15869 = n15868 ^ n15867 ^ n10082 ;
  assign n15870 = ( n408 & ~n5841 ) | ( n408 & n6345 ) | ( ~n5841 & n6345 ) ;
  assign n15871 = n10835 ^ n7331 ^ n1856 ;
  assign n15872 = n15871 ^ n3995 ^ x45 ;
  assign n15876 = ( n2455 & ~n6223 ) | ( n2455 & n10421 ) | ( ~n6223 & n10421 ) ;
  assign n15873 = n8842 ^ n4590 ^ 1'b0 ;
  assign n15874 = n4659 ^ n4404 ^ 1'b0 ;
  assign n15875 = ( n13685 & n15873 ) | ( n13685 & n15874 ) | ( n15873 & n15874 ) ;
  assign n15877 = n15876 ^ n15875 ^ n5541 ;
  assign n15878 = n4017 ^ n3879 ^ n3190 ;
  assign n15879 = ( n4136 & ~n8268 ) | ( n4136 & n15878 ) | ( ~n8268 & n15878 ) ;
  assign n15880 = ( ~n916 & n5810 ) | ( ~n916 & n10241 ) | ( n5810 & n10241 ) ;
  assign n15881 = n8156 & n15880 ;
  assign n15882 = ( n3610 & ~n15879 ) | ( n3610 & n15881 ) | ( ~n15879 & n15881 ) ;
  assign n15883 = ~n9001 & n15882 ;
  assign n15884 = n15408 ^ n11499 ^ n7573 ;
  assign n15885 = n15884 ^ n9183 ^ n5507 ;
  assign n15886 = ( n3514 & n3988 ) | ( n3514 & n5880 ) | ( n3988 & n5880 ) ;
  assign n15887 = n2381 & ~n15886 ;
  assign n15888 = ( n2119 & ~n3443 ) | ( n2119 & n15887 ) | ( ~n3443 & n15887 ) ;
  assign n15889 = n14759 & ~n14867 ;
  assign n15890 = ( n4218 & n15888 ) | ( n4218 & n15889 ) | ( n15888 & n15889 ) ;
  assign n15891 = ( n4640 & n8708 ) | ( n4640 & ~n10388 ) | ( n8708 & ~n10388 ) ;
  assign n15892 = n5087 ^ n4173 ^ 1'b0 ;
  assign n15893 = ~n3034 & n15892 ;
  assign n15894 = ( n3200 & ~n15891 ) | ( n3200 & n15893 ) | ( ~n15891 & n15893 ) ;
  assign n15895 = n6607 ^ n4378 ^ n3376 ;
  assign n15896 = ( ~n8126 & n9170 ) | ( ~n8126 & n15895 ) | ( n9170 & n15895 ) ;
  assign n15897 = n8082 ^ n6802 ^ n4413 ;
  assign n15898 = ( n2447 & n5755 ) | ( n2447 & ~n15897 ) | ( n5755 & ~n15897 ) ;
  assign n15899 = ( n4684 & n7196 ) | ( n4684 & ~n8092 ) | ( n7196 & ~n8092 ) ;
  assign n15900 = ( n5865 & n15898 ) | ( n5865 & n15899 ) | ( n15898 & n15899 ) ;
  assign n15901 = ( n8637 & n15896 ) | ( n8637 & ~n15900 ) | ( n15896 & ~n15900 ) ;
  assign n15902 = n13161 ^ n9421 ^ n5800 ;
  assign n15903 = n15902 ^ n6472 ^ n1404 ;
  assign n15908 = ( ~n718 & n6540 ) | ( ~n718 & n8048 ) | ( n6540 & n8048 ) ;
  assign n15907 = n12520 ^ n8566 ^ n2171 ;
  assign n15905 = n3950 ^ n2436 ^ n1860 ;
  assign n15904 = n7433 ^ n1736 ^ 1'b0 ;
  assign n15906 = n15905 ^ n15904 ^ n2400 ;
  assign n15909 = n15908 ^ n15907 ^ n15906 ;
  assign n15910 = n15909 ^ n14174 ^ 1'b0 ;
  assign n15911 = n15903 & ~n15910 ;
  assign n15914 = n5683 | n9479 ;
  assign n15915 = n15914 ^ n4520 ^ 1'b0 ;
  assign n15916 = n15915 ^ n4734 ^ 1'b0 ;
  assign n15912 = n10975 ^ n6026 ^ 1'b0 ;
  assign n15913 = n15912 ^ n3676 ^ n3638 ;
  assign n15917 = n15916 ^ n15913 ^ n4340 ;
  assign n15918 = ( n15222 & ~n15911 ) | ( n15222 & n15917 ) | ( ~n15911 & n15917 ) ;
  assign n15919 = ( ~n3404 & n5055 ) | ( ~n3404 & n7384 ) | ( n5055 & n7384 ) ;
  assign n15920 = n15919 ^ n8497 ^ 1'b0 ;
  assign n15921 = ~n15918 & n15920 ;
  assign n15922 = n3848 & n6752 ;
  assign n15923 = n3371 & n15922 ;
  assign n15924 = n6456 ^ n2230 ^ n536 ;
  assign n15925 = ( n4389 & n9097 ) | ( n4389 & n15924 ) | ( n9097 & n15924 ) ;
  assign n15926 = n15925 ^ n8237 ^ 1'b0 ;
  assign n15927 = n15923 | n15926 ;
  assign n15928 = n15927 ^ n14681 ^ n5564 ;
  assign n15929 = ( ~n3630 & n7488 ) | ( ~n3630 & n15928 ) | ( n7488 & n15928 ) ;
  assign n15930 = n7534 & ~n12909 ;
  assign n15931 = n15930 ^ n6616 ^ n990 ;
  assign n15932 = n2828 & n3399 ;
  assign n15933 = ~n13841 & n15932 ;
  assign n15934 = ( n4687 & ~n7257 ) | ( n4687 & n15933 ) | ( ~n7257 & n15933 ) ;
  assign n15935 = n6520 ^ n5200 ^ 1'b0 ;
  assign n15936 = n15935 ^ n11760 ^ n2762 ;
  assign n15937 = n15934 | n15936 ;
  assign n15938 = n15937 ^ n3767 ^ 1'b0 ;
  assign n15947 = ( n1647 & ~n2315 ) | ( n1647 & n11716 ) | ( ~n2315 & n11716 ) ;
  assign n15948 = ( ~n820 & n8941 ) | ( ~n820 & n15947 ) | ( n8941 & n15947 ) ;
  assign n15944 = n7845 ^ n4415 ^ n3011 ;
  assign n15945 = n15944 ^ n1863 ^ 1'b0 ;
  assign n15946 = n9866 | n15945 ;
  assign n15939 = n5784 ^ n2050 ^ 1'b0 ;
  assign n15940 = n13176 & n15939 ;
  assign n15941 = n15940 ^ n8231 ^ n4269 ;
  assign n15942 = n405 & n15941 ;
  assign n15943 = n15942 ^ n3258 ^ 1'b0 ;
  assign n15949 = n15948 ^ n15946 ^ n15943 ;
  assign n15950 = n15949 ^ n6288 ^ 1'b0 ;
  assign n15951 = ( n5467 & n7577 ) | ( n5467 & ~n9662 ) | ( n7577 & ~n9662 ) ;
  assign n15952 = ( ~n9588 & n15325 ) | ( ~n9588 & n15951 ) | ( n15325 & n15951 ) ;
  assign n15953 = n3637 & ~n11755 ;
  assign n15954 = n15953 ^ n1146 ^ 1'b0 ;
  assign n15955 = n7584 ^ n2309 ^ n1487 ;
  assign n15956 = n8678 ^ n1432 ^ 1'b0 ;
  assign n15957 = n15955 | n15956 ;
  assign n15958 = n15774 ^ n1155 ^ 1'b0 ;
  assign n15959 = n15957 | n15958 ;
  assign n15960 = n15878 ^ n4973 ^ n3395 ;
  assign n15961 = n7582 ^ n6143 ^ n2275 ;
  assign n15962 = n15960 & ~n15961 ;
  assign n15963 = n2900 & n15962 ;
  assign n15964 = n15963 ^ n3430 ^ n528 ;
  assign n15965 = n2320 | n6196 ;
  assign n15966 = n15964 & ~n15965 ;
  assign n15967 = n7231 ^ n5694 ^ 1'b0 ;
  assign n15968 = ~n660 & n15967 ;
  assign n15969 = n15968 ^ n10344 ^ n2834 ;
  assign n15970 = n5142 ^ n1104 ^ 1'b0 ;
  assign n15971 = ~n3027 & n15970 ;
  assign n15972 = ( ~n739 & n9068 ) | ( ~n739 & n15971 ) | ( n9068 & n15971 ) ;
  assign n15973 = n15972 ^ n307 ^ 1'b0 ;
  assign n15974 = n9832 ^ n7246 ^ n2700 ;
  assign n15975 = n1648 & n2525 ;
  assign n15976 = ~n378 & n15975 ;
  assign n15977 = n4883 ^ n4712 ^ n2937 ;
  assign n15978 = n3304 | n15977 ;
  assign n15979 = n15976 & ~n15978 ;
  assign n15980 = n4025 ^ n2330 ^ 1'b0 ;
  assign n15981 = n15979 | n15980 ;
  assign n15982 = n15981 ^ n5032 ^ 1'b0 ;
  assign n15983 = ( n6385 & ~n9328 ) | ( n6385 & n15718 ) | ( ~n9328 & n15718 ) ;
  assign n15984 = ( n9730 & n15982 ) | ( n9730 & ~n15983 ) | ( n15982 & ~n15983 ) ;
  assign n15985 = n10082 ^ n318 ^ 1'b0 ;
  assign n15986 = n8210 & ~n15985 ;
  assign n15988 = n1425 & ~n11412 ;
  assign n15989 = ~n1775 & n15988 ;
  assign n15987 = n10122 ^ n5189 ^ 1'b0 ;
  assign n15990 = n15989 ^ n15987 ^ n5511 ;
  assign n15991 = ( ~n4887 & n15986 ) | ( ~n4887 & n15990 ) | ( n15986 & n15990 ) ;
  assign n15992 = n656 ^ n463 ^ 1'b0 ;
  assign n15993 = ( n2418 & ~n4991 ) | ( n2418 & n15992 ) | ( ~n4991 & n15992 ) ;
  assign n15994 = n13531 ^ n457 ^ 1'b0 ;
  assign n15995 = ( ~n3551 & n11993 ) | ( ~n3551 & n13470 ) | ( n11993 & n13470 ) ;
  assign n15996 = n15994 | n15995 ;
  assign n15997 = n14738 | n15996 ;
  assign n15998 = n15997 ^ n15760 ^ n11893 ;
  assign n15999 = n6687 & ~n15998 ;
  assign n16000 = n15999 ^ n3106 ^ 1'b0 ;
  assign n16001 = ( ~n13052 & n15993 ) | ( ~n13052 & n16000 ) | ( n15993 & n16000 ) ;
  assign n16007 = n9760 ^ n3100 ^ 1'b0 ;
  assign n16006 = ( ~n2618 & n3433 ) | ( ~n2618 & n7004 ) | ( n3433 & n7004 ) ;
  assign n16008 = n16007 ^ n16006 ^ n3757 ;
  assign n16002 = n5547 ^ n4324 ^ 1'b0 ;
  assign n16003 = n3134 | n16002 ;
  assign n16004 = ( ~n401 & n2777 ) | ( ~n401 & n16003 ) | ( n2777 & n16003 ) ;
  assign n16005 = n3840 | n16004 ;
  assign n16009 = n16008 ^ n16005 ^ n12074 ;
  assign n16010 = n10903 ^ n5171 ^ 1'b0 ;
  assign n16011 = ( n788 & n4695 ) | ( n788 & ~n6344 ) | ( n4695 & ~n6344 ) ;
  assign n16012 = n9260 & n16011 ;
  assign n16013 = n15266 & n16012 ;
  assign n16014 = ( ~n3177 & n16010 ) | ( ~n3177 & n16013 ) | ( n16010 & n16013 ) ;
  assign n16015 = n15155 ^ n7763 ^ n5867 ;
  assign n16016 = n4500 | n9227 ;
  assign n16018 = ( ~x178 & n1833 ) | ( ~x178 & n8692 ) | ( n1833 & n8692 ) ;
  assign n16017 = ~n3244 & n8573 ;
  assign n16019 = n16018 ^ n16017 ^ n14176 ;
  assign n16020 = ( n16015 & ~n16016 ) | ( n16015 & n16019 ) | ( ~n16016 & n16019 ) ;
  assign n16021 = n16020 ^ n9230 ^ 1'b0 ;
  assign n16022 = ~n1090 & n16021 ;
  assign n16034 = n15896 ^ n7776 ^ n646 ;
  assign n16028 = ( n846 & n3785 ) | ( n846 & ~n4765 ) | ( n3785 & ~n4765 ) ;
  assign n16029 = n16028 ^ n12390 ^ n746 ;
  assign n16030 = n16029 ^ n2948 ^ 1'b0 ;
  assign n16031 = ( n12109 & n13757 ) | ( n12109 & n16030 ) | ( n13757 & n16030 ) ;
  assign n16032 = n16031 ^ n8839 ^ 1'b0 ;
  assign n16023 = n6410 ^ n5727 ^ x174 ;
  assign n16025 = ( n4223 & ~n5684 ) | ( n4223 & n11711 ) | ( ~n5684 & n11711 ) ;
  assign n16024 = ~n1340 & n2565 ;
  assign n16026 = n16025 ^ n16024 ^ n7191 ;
  assign n16027 = ( n14070 & n16023 ) | ( n14070 & ~n16026 ) | ( n16023 & ~n16026 ) ;
  assign n16033 = n16032 ^ n16027 ^ n1045 ;
  assign n16035 = n16034 ^ n16033 ^ n5836 ;
  assign n16036 = n9525 ^ n6293 ^ 1'b0 ;
  assign n16037 = n9041 & ~n16036 ;
  assign n16038 = n4850 ^ n3849 ^ 1'b0 ;
  assign n16039 = ~n11071 & n16038 ;
  assign n16040 = n16039 ^ n10447 ^ x237 ;
  assign n16041 = n12284 & ~n16040 ;
  assign n16043 = ( n6690 & n6948 ) | ( n6690 & n7540 ) | ( n6948 & n7540 ) ;
  assign n16042 = n4176 & ~n5807 ;
  assign n16044 = n16043 ^ n16042 ^ 1'b0 ;
  assign n16045 = ( n9066 & ~n13191 ) | ( n9066 & n16044 ) | ( ~n13191 & n16044 ) ;
  assign n16046 = n16045 ^ n11115 ^ n781 ;
  assign n16047 = ( n7620 & n9930 ) | ( n7620 & ~n10475 ) | ( n9930 & ~n10475 ) ;
  assign n16048 = ( n6288 & n6573 ) | ( n6288 & n16047 ) | ( n6573 & n16047 ) ;
  assign n16049 = n16048 ^ n8391 ^ 1'b0 ;
  assign n16050 = n8539 ^ n6988 ^ n6938 ;
  assign n16051 = n4476 & n5076 ;
  assign n16052 = n16051 ^ n3010 ^ 1'b0 ;
  assign n16053 = n16052 ^ n6975 ^ x200 ;
  assign n16054 = n16031 ^ n10868 ^ 1'b0 ;
  assign n16055 = n16053 & n16054 ;
  assign n16056 = n16050 & n16055 ;
  assign n16057 = n16056 ^ n15068 ^ 1'b0 ;
  assign n16060 = ( n1405 & ~n5108 ) | ( n1405 & n9224 ) | ( ~n5108 & n9224 ) ;
  assign n16058 = ( n3095 & n3224 ) | ( n3095 & n3982 ) | ( n3224 & n3982 ) ;
  assign n16059 = n16058 ^ n7371 ^ n4877 ;
  assign n16061 = n16060 ^ n16059 ^ n6308 ;
  assign n16062 = n15575 ^ n9796 ^ n5672 ;
  assign n16063 = n14846 | n16062 ;
  assign n16064 = n13170 | n16063 ;
  assign n16065 = n6120 & ~n7806 ;
  assign n16066 = n9384 ^ n5184 ^ n2265 ;
  assign n16067 = ( n5901 & n16065 ) | ( n5901 & n16066 ) | ( n16065 & n16066 ) ;
  assign n16071 = n1342 & n4036 ;
  assign n16072 = ( ~n1290 & n15015 ) | ( ~n1290 & n16071 ) | ( n15015 & n16071 ) ;
  assign n16068 = ( ~n7901 & n12394 ) | ( ~n7901 & n15570 ) | ( n12394 & n15570 ) ;
  assign n16069 = n16068 ^ n9804 ^ n4340 ;
  assign n16070 = n2257 & ~n16069 ;
  assign n16073 = n16072 ^ n16070 ^ 1'b0 ;
  assign n16074 = n11681 ^ n6061 ^ 1'b0 ;
  assign n16075 = ~n16073 & n16074 ;
  assign n16076 = n9000 ^ n4934 ^ n439 ;
  assign n16077 = n929 & n16076 ;
  assign n16079 = n836 | n3230 ;
  assign n16080 = n16079 ^ n5457 ^ 1'b0 ;
  assign n16081 = ~n1510 & n16080 ;
  assign n16082 = n4957 ^ n3790 ^ n963 ;
  assign n16083 = n16081 & ~n16082 ;
  assign n16084 = ~n12716 & n16083 ;
  assign n16085 = n16084 ^ n406 ^ 1'b0 ;
  assign n16086 = n5507 & n6698 ;
  assign n16087 = n16086 ^ n1613 ^ 1'b0 ;
  assign n16088 = n4695 & n16087 ;
  assign n16089 = ~n16085 & n16088 ;
  assign n16078 = ( n3249 & n8088 ) | ( n3249 & n12966 ) | ( n8088 & n12966 ) ;
  assign n16090 = n16089 ^ n16078 ^ n11124 ;
  assign n16098 = ( ~n3358 & n5270 ) | ( ~n3358 & n5657 ) | ( n5270 & n5657 ) ;
  assign n16094 = n5648 ^ n4072 ^ n2867 ;
  assign n16095 = n2551 ^ n1103 ^ 1'b0 ;
  assign n16096 = ~n16094 & n16095 ;
  assign n16092 = n10966 ^ n4108 ^ 1'b0 ;
  assign n16093 = n14967 & ~n16092 ;
  assign n16097 = n16096 ^ n16093 ^ n2229 ;
  assign n16091 = ( n2213 & n2350 ) | ( n2213 & ~n9431 ) | ( n2350 & ~n9431 ) ;
  assign n16099 = n16098 ^ n16097 ^ n16091 ;
  assign n16100 = ( ~n525 & n1751 ) | ( ~n525 & n16099 ) | ( n1751 & n16099 ) ;
  assign n16101 = n3554 ^ n2168 ^ 1'b0 ;
  assign n16102 = n12090 ^ n9160 ^ n7070 ;
  assign n16103 = n16102 ^ n5522 ^ n3366 ;
  assign n16104 = n16101 & ~n16103 ;
  assign n16105 = ( n918 & ~n3254 ) | ( n918 & n8684 ) | ( ~n3254 & n8684 ) ;
  assign n16106 = ( n9841 & ~n12970 ) | ( n9841 & n13880 ) | ( ~n12970 & n13880 ) ;
  assign n16107 = ( n13505 & n16105 ) | ( n13505 & ~n16106 ) | ( n16105 & ~n16106 ) ;
  assign n16108 = n8301 ^ n3269 ^ 1'b0 ;
  assign n16109 = ( n1557 & n13679 ) | ( n1557 & ~n16108 ) | ( n13679 & ~n16108 ) ;
  assign n16110 = ~n10075 & n16109 ;
  assign n16111 = n16110 ^ n8279 ^ 1'b0 ;
  assign n16112 = n10603 ^ n6902 ^ n2897 ;
  assign n16113 = n1964 ^ n1709 ^ 1'b0 ;
  assign n16114 = ( n897 & ~n4858 ) | ( n897 & n12758 ) | ( ~n4858 & n12758 ) ;
  assign n16115 = n16114 ^ n12260 ^ n4685 ;
  assign n16117 = n14519 ^ n3599 ^ n2344 ;
  assign n16116 = n10931 ^ n3138 ^ n1456 ;
  assign n16118 = n16117 ^ n16116 ^ n4842 ;
  assign n16119 = ( n16113 & n16115 ) | ( n16113 & ~n16118 ) | ( n16115 & ~n16118 ) ;
  assign n16120 = n7205 ^ n2725 ^ n1020 ;
  assign n16121 = ( n4039 & n5915 ) | ( n4039 & n10164 ) | ( n5915 & n10164 ) ;
  assign n16122 = n16120 & ~n16121 ;
  assign n16123 = n10189 ^ n7371 ^ n877 ;
  assign n16124 = ( n2289 & ~n14577 ) | ( n2289 & n16123 ) | ( ~n14577 & n16123 ) ;
  assign n16125 = n16124 ^ n9887 ^ n5307 ;
  assign n16126 = ( n4783 & n11549 ) | ( n4783 & n16125 ) | ( n11549 & n16125 ) ;
  assign n16127 = ( ~n10820 & n15213 ) | ( ~n10820 & n16126 ) | ( n15213 & n16126 ) ;
  assign n16128 = n15483 ^ n11481 ^ n3778 ;
  assign n16131 = n2983 | n5954 ;
  assign n16129 = ( ~n614 & n4078 ) | ( ~n614 & n10887 ) | ( n4078 & n10887 ) ;
  assign n16130 = x218 & ~n16129 ;
  assign n16132 = n16131 ^ n16130 ^ n4730 ;
  assign n16133 = x171 & ~n2129 ;
  assign n16134 = n16132 & n16133 ;
  assign n16135 = ~n3945 & n8705 ;
  assign n16136 = ( n3326 & n9578 ) | ( n3326 & ~n15427 ) | ( n9578 & ~n15427 ) ;
  assign n16137 = n16136 ^ n13803 ^ n6649 ;
  assign n16138 = ( n1705 & n13800 ) | ( n1705 & ~n14709 ) | ( n13800 & ~n14709 ) ;
  assign n16139 = n16137 | n16138 ;
  assign n16140 = n8503 | n16139 ;
  assign n16141 = n12897 ^ n1940 ^ 1'b0 ;
  assign n16142 = ( n6538 & n13214 ) | ( n6538 & ~n16141 ) | ( n13214 & ~n16141 ) ;
  assign n16143 = n16140 & ~n16142 ;
  assign n16144 = n16143 ^ n15448 ^ 1'b0 ;
  assign n16145 = n11613 ^ n6227 ^ n4131 ;
  assign n16151 = n7442 & ~n8219 ;
  assign n16152 = ~n1092 & n16151 ;
  assign n16147 = n8330 ^ n4850 ^ 1'b0 ;
  assign n16146 = ~n568 & n977 ;
  assign n16148 = n16147 ^ n16146 ^ 1'b0 ;
  assign n16149 = n16148 ^ n3262 ^ n1800 ;
  assign n16150 = n5783 & ~n16149 ;
  assign n16153 = n16152 ^ n16150 ^ 1'b0 ;
  assign n16154 = ( n4678 & n16145 ) | ( n4678 & ~n16153 ) | ( n16145 & ~n16153 ) ;
  assign n16155 = n264 & ~n2200 ;
  assign n16156 = n16155 ^ n14656 ^ n10634 ;
  assign n16157 = n11860 ^ n10822 ^ n288 ;
  assign n16158 = ( n3745 & ~n7596 ) | ( n3745 & n16157 ) | ( ~n7596 & n16157 ) ;
  assign n16159 = ( n2397 & ~n3074 ) | ( n2397 & n3810 ) | ( ~n3074 & n3810 ) ;
  assign n16160 = ~n16158 & n16159 ;
  assign n16161 = n16160 ^ n13987 ^ n10179 ;
  assign n16162 = ( n3548 & n7062 ) | ( n3548 & ~n16161 ) | ( n7062 & ~n16161 ) ;
  assign n16163 = ( n646 & ~n1911 ) | ( n646 & n4433 ) | ( ~n1911 & n4433 ) ;
  assign n16164 = n16163 ^ n14491 ^ n4647 ;
  assign n16165 = ( ~n5015 & n8118 ) | ( ~n5015 & n14843 ) | ( n8118 & n14843 ) ;
  assign n16166 = n16165 ^ n6381 ^ n5065 ;
  assign n16167 = n16164 & ~n16166 ;
  assign n16168 = ( n5031 & n6744 ) | ( n5031 & n10341 ) | ( n6744 & n10341 ) ;
  assign n16169 = ( x251 & ~n2828 ) | ( x251 & n16168 ) | ( ~n2828 & n16168 ) ;
  assign n16170 = ( ~n9210 & n12599 ) | ( ~n9210 & n15134 ) | ( n12599 & n15134 ) ;
  assign n16171 = n16170 ^ n10882 ^ 1'b0 ;
  assign n16172 = n3413 | n16171 ;
  assign n16173 = n10800 & n16172 ;
  assign n16174 = n16173 ^ n1283 ^ 1'b0 ;
  assign n16175 = n4295 & ~n7169 ;
  assign n16176 = ~n9900 & n16175 ;
  assign n16177 = ( ~n3898 & n6922 ) | ( ~n3898 & n16176 ) | ( n6922 & n16176 ) ;
  assign n16178 = ( n729 & ~n2943 ) | ( n729 & n4605 ) | ( ~n2943 & n4605 ) ;
  assign n16179 = n16178 ^ n11539 ^ 1'b0 ;
  assign n16180 = ~n7130 & n16179 ;
  assign n16181 = n16180 ^ n13145 ^ n10081 ;
  assign n16182 = n16181 ^ n15895 ^ n6371 ;
  assign n16183 = ( n721 & n10490 ) | ( n721 & ~n12026 ) | ( n10490 & ~n12026 ) ;
  assign n16184 = n14785 ^ n7141 ^ n813 ;
  assign n16185 = ( n2766 & ~n4481 ) | ( n2766 & n16184 ) | ( ~n4481 & n16184 ) ;
  assign n16186 = n16185 ^ x240 ^ 1'b0 ;
  assign n16187 = n5742 ^ n4573 ^ n4109 ;
  assign n16188 = ( n5204 & n12608 ) | ( n5204 & ~n16187 ) | ( n12608 & ~n16187 ) ;
  assign n16189 = n2500 & ~n16188 ;
  assign n16197 = n414 & ~n11418 ;
  assign n16198 = n16197 ^ n4375 ^ 1'b0 ;
  assign n16194 = n12826 ^ n1568 ^ 1'b0 ;
  assign n16190 = n5006 | n7376 ;
  assign n16191 = n16190 ^ n639 ^ 1'b0 ;
  assign n16192 = n10704 | n16191 ;
  assign n16193 = n16192 ^ n1142 ^ 1'b0 ;
  assign n16195 = n16194 ^ n16193 ^ 1'b0 ;
  assign n16196 = ( n3902 & n10319 ) | ( n3902 & n16195 ) | ( n10319 & n16195 ) ;
  assign n16199 = n16198 ^ n16196 ^ x197 ;
  assign n16200 = ( n6572 & n16189 ) | ( n6572 & n16199 ) | ( n16189 & n16199 ) ;
  assign n16201 = ( n1639 & n4105 ) | ( n1639 & ~n12715 ) | ( n4105 & ~n12715 ) ;
  assign n16202 = ( n2103 & n12825 ) | ( n2103 & ~n13189 ) | ( n12825 & ~n13189 ) ;
  assign n16203 = ( ~n2457 & n10884 ) | ( ~n2457 & n12055 ) | ( n10884 & n12055 ) ;
  assign n16204 = ( n10566 & ~n16202 ) | ( n10566 & n16203 ) | ( ~n16202 & n16203 ) ;
  assign n16209 = ( ~n4632 & n7799 ) | ( ~n4632 & n9431 ) | ( n7799 & n9431 ) ;
  assign n16205 = n4827 ^ n2328 ^ 1'b0 ;
  assign n16206 = n14683 ^ n6118 ^ n5259 ;
  assign n16207 = ~n16205 & n16206 ;
  assign n16208 = n9104 & n16207 ;
  assign n16210 = n16209 ^ n16208 ^ 1'b0 ;
  assign n16211 = n9720 ^ n7917 ^ n319 ;
  assign n16212 = n16211 ^ n11059 ^ 1'b0 ;
  assign n16214 = ( x243 & n4936 ) | ( x243 & ~n9738 ) | ( n4936 & ~n9738 ) ;
  assign n16215 = n16214 ^ n12533 ^ n5310 ;
  assign n16213 = n2594 & n9576 ;
  assign n16216 = n16215 ^ n16213 ^ 1'b0 ;
  assign n16217 = n5772 & n16216 ;
  assign n16218 = n16217 ^ x109 ^ 1'b0 ;
  assign n16219 = n9641 ^ n4382 ^ 1'b0 ;
  assign n16220 = n16219 ^ n6788 ^ x68 ;
  assign n16221 = ( n1408 & n4744 ) | ( n1408 & ~n16220 ) | ( n4744 & ~n16220 ) ;
  assign n16222 = n16221 ^ n14875 ^ n812 ;
  assign n16223 = ( n3208 & n8736 ) | ( n3208 & ~n16222 ) | ( n8736 & ~n16222 ) ;
  assign n16224 = n9144 ^ n5869 ^ n1736 ;
  assign n16225 = n16224 ^ n8663 ^ 1'b0 ;
  assign n16226 = n9478 & ~n16225 ;
  assign n16227 = ~n12390 & n16226 ;
  assign n16228 = n6006 ^ n2697 ^ n1259 ;
  assign n16229 = ( ~n6137 & n9384 ) | ( ~n6137 & n16228 ) | ( n9384 & n16228 ) ;
  assign n16230 = ( n10613 & n15379 ) | ( n10613 & n16229 ) | ( n15379 & n16229 ) ;
  assign n16231 = n12990 ^ n10663 ^ n7108 ;
  assign n16232 = n10927 ^ n2498 ^ 1'b0 ;
  assign n16233 = ~n3541 & n16093 ;
  assign n16234 = n16233 ^ n767 ^ 1'b0 ;
  assign n16237 = n5806 ^ n1937 ^ n1437 ;
  assign n16238 = ( ~n1747 & n5026 ) | ( ~n1747 & n16237 ) | ( n5026 & n16237 ) ;
  assign n16239 = n6023 & n16238 ;
  assign n16240 = n16239 ^ n995 ^ 1'b0 ;
  assign n16235 = ~n5707 & n6025 ;
  assign n16236 = n16235 ^ n1552 ^ 1'b0 ;
  assign n16241 = n16240 ^ n16236 ^ 1'b0 ;
  assign n16242 = ( n1610 & n4151 ) | ( n1610 & n8537 ) | ( n4151 & n8537 ) ;
  assign n16243 = n16242 ^ n8386 ^ n8336 ;
  assign n16249 = ( ~n4097 & n6151 ) | ( ~n4097 & n7396 ) | ( n6151 & n7396 ) ;
  assign n16244 = n3018 & n8391 ;
  assign n16245 = ( ~n3260 & n3584 ) | ( ~n3260 & n16209 ) | ( n3584 & n16209 ) ;
  assign n16246 = n16244 | n16245 ;
  assign n16247 = n16246 ^ n9006 ^ 1'b0 ;
  assign n16248 = ( n2644 & ~n14566 ) | ( n2644 & n16247 ) | ( ~n14566 & n16247 ) ;
  assign n16250 = n16249 ^ n16248 ^ n8476 ;
  assign n16251 = n5691 ^ n4410 ^ n965 ;
  assign n16252 = n5445 & ~n16251 ;
  assign n16253 = n16252 ^ n12386 ^ 1'b0 ;
  assign n16254 = ( n3604 & n6809 ) | ( n3604 & n7750 ) | ( n6809 & n7750 ) ;
  assign n16255 = ~n2092 & n16254 ;
  assign n16256 = ~n16253 & n16255 ;
  assign n16257 = n7096 ^ n284 ^ 1'b0 ;
  assign n16258 = ( n16250 & n16256 ) | ( n16250 & n16257 ) | ( n16256 & n16257 ) ;
  assign n16259 = n10561 ^ n4980 ^ n3397 ;
  assign n16263 = ( ~n2646 & n4414 ) | ( ~n2646 & n9164 ) | ( n4414 & n9164 ) ;
  assign n16264 = n1105 | n16263 ;
  assign n16260 = n6673 ^ n4026 ^ 1'b0 ;
  assign n16261 = n8167 & ~n16260 ;
  assign n16262 = n16261 ^ n12062 ^ n9896 ;
  assign n16265 = n16264 ^ n16262 ^ n11793 ;
  assign n16266 = n10184 ^ n3725 ^ 1'b0 ;
  assign n16267 = ~n3879 & n16266 ;
  assign n16268 = ( ~n884 & n16094 ) | ( ~n884 & n16267 ) | ( n16094 & n16267 ) ;
  assign n16269 = ( n1697 & ~n6450 ) | ( n1697 & n12854 ) | ( ~n6450 & n12854 ) ;
  assign n16270 = ( n3668 & n3820 ) | ( n3668 & n14387 ) | ( n3820 & n14387 ) ;
  assign n16271 = ( n3940 & n16082 ) | ( n3940 & n16270 ) | ( n16082 & n16270 ) ;
  assign n16272 = n16271 ^ n8699 ^ n8561 ;
  assign n16273 = n16272 ^ n10085 ^ n6286 ;
  assign n16274 = ( n16268 & ~n16269 ) | ( n16268 & n16273 ) | ( ~n16269 & n16273 ) ;
  assign n16275 = ( n8291 & n9133 ) | ( n8291 & n13462 ) | ( n9133 & n13462 ) ;
  assign n16276 = ( n4509 & ~n11069 ) | ( n4509 & n15702 ) | ( ~n11069 & n15702 ) ;
  assign n16277 = n16276 ^ n634 ^ n293 ;
  assign n16278 = n5999 ^ n4884 ^ 1'b0 ;
  assign n16279 = n1099 & ~n13348 ;
  assign n16280 = n5494 & n16279 ;
  assign n16281 = n16280 ^ n9952 ^ n4932 ;
  assign n16282 = ( n1455 & n4075 ) | ( n1455 & ~n16281 ) | ( n4075 & ~n16281 ) ;
  assign n16284 = n2977 ^ n1019 ^ 1'b0 ;
  assign n16285 = n4993 & ~n16284 ;
  assign n16286 = ( ~n5547 & n5724 ) | ( ~n5547 & n16285 ) | ( n5724 & n16285 ) ;
  assign n16283 = n13615 ^ n10696 ^ n648 ;
  assign n16287 = n16286 ^ n16283 ^ 1'b0 ;
  assign n16288 = n15331 ^ x177 ^ 1'b0 ;
  assign n16289 = n10091 | n16288 ;
  assign n16290 = n16289 ^ n14307 ^ n5839 ;
  assign n16291 = ( n3957 & n12306 ) | ( n3957 & ~n16290 ) | ( n12306 & ~n16290 ) ;
  assign n16292 = n5251 ^ n4229 ^ 1'b0 ;
  assign n16293 = n8052 ^ n4074 ^ n1678 ;
  assign n16294 = n16293 ^ n1592 ^ 1'b0 ;
  assign n16295 = ~n792 & n16294 ;
  assign n16296 = ~n16292 & n16295 ;
  assign n16297 = n16296 ^ n8107 ^ 1'b0 ;
  assign n16298 = n12692 ^ n8502 ^ 1'b0 ;
  assign n16299 = n1576 & n16298 ;
  assign n16300 = n16299 ^ n7079 ^ n276 ;
  assign n16301 = n8148 ^ n6606 ^ n365 ;
  assign n16302 = n16301 ^ n4791 ^ n1200 ;
  assign n16303 = n16302 ^ n10330 ^ 1'b0 ;
  assign n16304 = ~n16300 & n16303 ;
  assign n16305 = n7990 ^ n4120 ^ n540 ;
  assign n16312 = n9623 ^ n1113 ^ 1'b0 ;
  assign n16313 = n6038 & n16312 ;
  assign n16308 = n15662 ^ n4224 ^ n2782 ;
  assign n16309 = ( ~n590 & n7713 ) | ( ~n590 & n8541 ) | ( n7713 & n8541 ) ;
  assign n16310 = ( ~n15963 & n16308 ) | ( ~n15963 & n16309 ) | ( n16308 & n16309 ) ;
  assign n16306 = n8014 ^ n3648 ^ n3582 ;
  assign n16307 = n363 & n16306 ;
  assign n16311 = n16310 ^ n16307 ^ 1'b0 ;
  assign n16314 = n16313 ^ n16311 ^ n4628 ;
  assign n16316 = n2951 & ~n7194 ;
  assign n16317 = n1328 & n16316 ;
  assign n16318 = ( n3906 & n6172 ) | ( n3906 & ~n16317 ) | ( n6172 & ~n16317 ) ;
  assign n16315 = n9216 ^ n5223 ^ n2245 ;
  assign n16319 = n16318 ^ n16315 ^ n7169 ;
  assign n16320 = n3690 ^ n3073 ^ n468 ;
  assign n16321 = n13295 ^ n8109 ^ n558 ;
  assign n16322 = n16321 ^ n14506 ^ n8372 ;
  assign n16323 = ( n10652 & n16320 ) | ( n10652 & ~n16322 ) | ( n16320 & ~n16322 ) ;
  assign n16324 = ( n2677 & ~n10517 ) | ( n2677 & n15099 ) | ( ~n10517 & n15099 ) ;
  assign n16325 = n4687 | n16324 ;
  assign n16326 = ( ~n1797 & n4743 ) | ( ~n1797 & n7523 ) | ( n4743 & n7523 ) ;
  assign n16327 = ( n6128 & ~n10938 ) | ( n6128 & n16326 ) | ( ~n10938 & n16326 ) ;
  assign n16328 = ( n16323 & n16325 ) | ( n16323 & ~n16327 ) | ( n16325 & ~n16327 ) ;
  assign n16334 = n13261 ^ n3628 ^ 1'b0 ;
  assign n16332 = n13403 ^ n2510 ^ 1'b0 ;
  assign n16331 = n6299 ^ n6105 ^ 1'b0 ;
  assign n16333 = n16332 ^ n16331 ^ n10673 ;
  assign n16329 = n6825 ^ n3563 ^ n1079 ;
  assign n16330 = n16329 ^ n11378 ^ n1069 ;
  assign n16335 = n16334 ^ n16333 ^ n16330 ;
  assign n16336 = n12862 ^ n7534 ^ 1'b0 ;
  assign n16337 = n16336 ^ n15924 ^ n1693 ;
  assign n16341 = n8464 ^ n7042 ^ n602 ;
  assign n16340 = n15992 ^ n6955 ^ n3250 ;
  assign n16342 = n16341 ^ n16340 ^ n15612 ;
  assign n16338 = n12776 ^ x210 ^ 1'b0 ;
  assign n16339 = ( n5590 & n8503 ) | ( n5590 & ~n16338 ) | ( n8503 & ~n16338 ) ;
  assign n16343 = n16342 ^ n16339 ^ n5664 ;
  assign n16344 = n7972 ^ n7331 ^ n1699 ;
  assign n16345 = ( n16236 & ~n16343 ) | ( n16236 & n16344 ) | ( ~n16343 & n16344 ) ;
  assign n16350 = ( n2541 & ~n3320 ) | ( n2541 & n6622 ) | ( ~n3320 & n6622 ) ;
  assign n16351 = n16350 ^ n4625 ^ 1'b0 ;
  assign n16352 = n16351 ^ n9472 ^ n7588 ;
  assign n16346 = n15250 ^ n7897 ^ n292 ;
  assign n16347 = ( ~x179 & n502 ) | ( ~x179 & n16346 ) | ( n502 & n16346 ) ;
  assign n16348 = n9734 ^ n4840 ^ n2296 ;
  assign n16349 = ( n5962 & n16347 ) | ( n5962 & ~n16348 ) | ( n16347 & ~n16348 ) ;
  assign n16353 = n16352 ^ n16349 ^ n4261 ;
  assign n16354 = n1580 ^ n1319 ^ n756 ;
  assign n16358 = n2559 ^ n864 ^ x56 ;
  assign n16355 = n6301 ^ n337 ^ 1'b0 ;
  assign n16356 = n3504 | n7539 ;
  assign n16357 = n16355 | n16356 ;
  assign n16359 = n16358 ^ n16357 ^ n8566 ;
  assign n16360 = ( n4439 & n16354 ) | ( n4439 & ~n16359 ) | ( n16354 & ~n16359 ) ;
  assign n16361 = n5506 & n14123 ;
  assign n16362 = n16361 ^ x200 ^ 1'b0 ;
  assign n16363 = n13091 ^ n4916 ^ n1747 ;
  assign n16364 = ( n2533 & ~n7749 ) | ( n2533 & n16363 ) | ( ~n7749 & n16363 ) ;
  assign n16365 = ( n4099 & n16362 ) | ( n4099 & ~n16364 ) | ( n16362 & ~n16364 ) ;
  assign n16367 = n3833 ^ n3766 ^ n1402 ;
  assign n16366 = n7444 ^ n6790 ^ n6218 ;
  assign n16368 = n16367 ^ n16366 ^ n7067 ;
  assign n16369 = ~n7468 & n8057 ;
  assign n16370 = n439 & ~n9966 ;
  assign n16371 = ~n16369 & n16370 ;
  assign n16372 = ( n4823 & ~n5104 ) | ( n4823 & n5881 ) | ( ~n5104 & n5881 ) ;
  assign n16373 = ( n377 & n2815 ) | ( n377 & ~n6813 ) | ( n2815 & ~n6813 ) ;
  assign n16374 = n16373 ^ n12374 ^ n339 ;
  assign n16375 = n16374 ^ n13574 ^ n3523 ;
  assign n16376 = n15411 & n16375 ;
  assign n16377 = n16376 ^ n1053 ^ 1'b0 ;
  assign n16378 = ~n15199 & n16377 ;
  assign n16381 = n3359 ^ n3001 ^ n2574 ;
  assign n16379 = ( x152 & n2905 ) | ( x152 & ~n3094 ) | ( n2905 & ~n3094 ) ;
  assign n16380 = ( ~n2710 & n11989 ) | ( ~n2710 & n16379 ) | ( n11989 & n16379 ) ;
  assign n16382 = n16381 ^ n16380 ^ 1'b0 ;
  assign n16383 = n11423 ^ n10799 ^ n4229 ;
  assign n16384 = ~n9249 & n16383 ;
  assign n16385 = ~n9419 & n16384 ;
  assign n16386 = n9357 ^ n2886 ^ n2335 ;
  assign n16397 = n4722 ^ n2060 ^ 1'b0 ;
  assign n16398 = n8259 & n16397 ;
  assign n16399 = ( ~n10416 & n10549 ) | ( ~n10416 & n16398 ) | ( n10549 & n16398 ) ;
  assign n16400 = n16399 ^ n8748 ^ n4424 ;
  assign n16387 = n3536 & ~n5500 ;
  assign n16388 = ~n10535 & n16387 ;
  assign n16389 = n16388 ^ n5190 ^ 1'b0 ;
  assign n16390 = n680 | n16389 ;
  assign n16392 = n2629 & n4632 ;
  assign n16393 = n16392 ^ n2615 ^ 1'b0 ;
  assign n16391 = ( n2304 & n5494 ) | ( n2304 & ~n15034 ) | ( n5494 & ~n15034 ) ;
  assign n16394 = n16393 ^ n16391 ^ 1'b0 ;
  assign n16395 = n16390 | n16394 ;
  assign n16396 = n16395 ^ n4513 ^ 1'b0 ;
  assign n16401 = n16400 ^ n16396 ^ n11737 ;
  assign n16402 = n7482 ^ n3962 ^ n1680 ;
  assign n16403 = n16402 ^ n1959 ^ 1'b0 ;
  assign n16404 = ( n1509 & n2800 ) | ( n1509 & n6187 ) | ( n2800 & n6187 ) ;
  assign n16405 = n1558 | n8112 ;
  assign n16406 = n16405 ^ n9578 ^ 1'b0 ;
  assign n16407 = n8190 | n16406 ;
  assign n16408 = n779 & ~n16407 ;
  assign n16409 = n7727 | n16408 ;
  assign n16410 = n16404 & ~n16409 ;
  assign n16411 = n4655 & n7021 ;
  assign n16412 = n16411 ^ n10280 ^ n5166 ;
  assign n16413 = ( n1508 & ~n6172 ) | ( n1508 & n15168 ) | ( ~n6172 & n15168 ) ;
  assign n16414 = n14789 ^ n12936 ^ n308 ;
  assign n16415 = n12840 ^ n6724 ^ 1'b0 ;
  assign n16416 = ( n2646 & n2975 ) | ( n2646 & ~n10877 ) | ( n2975 & ~n10877 ) ;
  assign n16417 = n16381 & ~n16416 ;
  assign n16418 = n8348 ^ n6604 ^ n3535 ;
  assign n16419 = n16418 ^ n16310 ^ n11090 ;
  assign n16420 = n15865 | n16419 ;
  assign n16421 = n5699 | n16420 ;
  assign n16422 = ~n7248 & n16421 ;
  assign n16423 = ~n11740 & n16422 ;
  assign n16424 = ( n2622 & ~n4812 ) | ( n2622 & n16423 ) | ( ~n4812 & n16423 ) ;
  assign n16425 = ( n405 & ~n5803 ) | ( n405 & n13108 ) | ( ~n5803 & n13108 ) ;
  assign n16426 = n12808 & n16425 ;
  assign n16427 = n16426 ^ x84 ^ 1'b0 ;
  assign n16428 = n16427 ^ n13820 ^ 1'b0 ;
  assign n16429 = n6935 ^ n5271 ^ n3416 ;
  assign n16430 = ( n992 & ~n7607 ) | ( n992 & n16429 ) | ( ~n7607 & n16429 ) ;
  assign n16437 = ( n3778 & ~n10055 ) | ( n3778 & n15475 ) | ( ~n10055 & n15475 ) ;
  assign n16438 = n16437 ^ n14495 ^ n10291 ;
  assign n16435 = n11832 ^ n10175 ^ n5073 ;
  assign n16431 = ~n4305 & n15499 ;
  assign n16432 = n16431 ^ n9120 ^ 1'b0 ;
  assign n16433 = ~n5602 & n16432 ;
  assign n16434 = ( n8773 & ~n13561 ) | ( n8773 & n16433 ) | ( ~n13561 & n16433 ) ;
  assign n16436 = n16435 ^ n16434 ^ 1'b0 ;
  assign n16439 = n16438 ^ n16436 ^ n13378 ;
  assign n16440 = ( ~n12673 & n13138 ) | ( ~n12673 & n15940 ) | ( n13138 & n15940 ) ;
  assign n16446 = ( ~x84 & n8220 ) | ( ~x84 & n9143 ) | ( n8220 & n9143 ) ;
  assign n16443 = n4072 ^ n3859 ^ n2605 ;
  assign n16444 = n16443 ^ n13311 ^ n3421 ;
  assign n16445 = n16444 ^ n14147 ^ n10518 ;
  assign n16447 = n16446 ^ n16445 ^ n8885 ;
  assign n16441 = n331 & n9941 ;
  assign n16442 = ~n9301 & n16441 ;
  assign n16448 = n16447 ^ n16442 ^ n5417 ;
  assign n16449 = ( n2303 & ~n16440 ) | ( n2303 & n16448 ) | ( ~n16440 & n16448 ) ;
  assign n16450 = ( n772 & n1075 ) | ( n772 & ~n5022 ) | ( n1075 & ~n5022 ) ;
  assign n16451 = n6099 & ~n16450 ;
  assign n16452 = n16451 ^ n5890 ^ 1'b0 ;
  assign n16459 = n8902 ^ n6544 ^ n2378 ;
  assign n16460 = n16459 ^ n13672 ^ n1828 ;
  assign n16453 = n15042 ^ n4677 ^ n4612 ;
  assign n16454 = n16453 ^ n7830 ^ 1'b0 ;
  assign n16455 = n5130 & ~n10442 ;
  assign n16456 = n1098 | n16455 ;
  assign n16457 = ( n2686 & n14851 ) | ( n2686 & ~n16456 ) | ( n14851 & ~n16456 ) ;
  assign n16458 = ~n16454 & n16457 ;
  assign n16461 = n16460 ^ n16458 ^ 1'b0 ;
  assign n16462 = n16461 ^ n13958 ^ n12760 ;
  assign n16463 = n10925 ^ n6666 ^ n3406 ;
  assign n16464 = n16463 ^ n824 ^ 1'b0 ;
  assign n16465 = n13685 & n16464 ;
  assign n16466 = ( ~x174 & n2473 ) | ( ~x174 & n8972 ) | ( n2473 & n8972 ) ;
  assign n16467 = n16466 ^ n8483 ^ n2176 ;
  assign n16468 = n4813 | n16435 ;
  assign n16469 = n3860 | n16468 ;
  assign n16470 = ( ~n554 & n16467 ) | ( ~n554 & n16469 ) | ( n16467 & n16469 ) ;
  assign n16471 = ( n7273 & n13902 ) | ( n7273 & ~n16470 ) | ( n13902 & ~n16470 ) ;
  assign n16472 = n16471 ^ n15013 ^ n13246 ;
  assign n16473 = ( ~x37 & n1110 ) | ( ~x37 & n2305 ) | ( n1110 & n2305 ) ;
  assign n16474 = n16473 ^ n1233 ^ 1'b0 ;
  assign n16475 = ( ~n4020 & n4362 ) | ( ~n4020 & n16474 ) | ( n4362 & n16474 ) ;
  assign n16476 = n16475 ^ n7927 ^ n7194 ;
  assign n16477 = ( ~n6984 & n16472 ) | ( ~n6984 & n16476 ) | ( n16472 & n16476 ) ;
  assign n16478 = ( n13235 & ~n16465 ) | ( n13235 & n16477 ) | ( ~n16465 & n16477 ) ;
  assign n16479 = ( ~n7378 & n10376 ) | ( ~n7378 & n11755 ) | ( n10376 & n11755 ) ;
  assign n16480 = n16479 ^ n9342 ^ 1'b0 ;
  assign n16481 = ( ~n6213 & n10167 ) | ( ~n6213 & n11300 ) | ( n10167 & n11300 ) ;
  assign n16482 = n14959 ^ n13660 ^ n12159 ;
  assign n16483 = n2737 ^ n1153 ^ 1'b0 ;
  assign n16484 = n12561 & n16483 ;
  assign n16485 = n7787 ^ n5870 ^ 1'b0 ;
  assign n16486 = n6171 & n16485 ;
  assign n16487 = n7852 | n9889 ;
  assign n16488 = n16487 ^ n14557 ^ 1'b0 ;
  assign n16489 = n16486 & n16488 ;
  assign n16490 = ~n16484 & n16489 ;
  assign n16506 = n4465 & n8615 ;
  assign n16507 = ( n2334 & ~n12286 ) | ( n2334 & n16506 ) | ( ~n12286 & n16506 ) ;
  assign n16508 = n1545 | n16507 ;
  assign n16509 = n8728 & ~n16508 ;
  assign n16491 = ( ~n2136 & n6726 ) | ( ~n2136 & n9370 ) | ( n6726 & n9370 ) ;
  assign n16492 = n12813 ^ n4172 ^ n3374 ;
  assign n16493 = n16492 ^ n9517 ^ n5587 ;
  assign n16494 = n5965 & n16493 ;
  assign n16495 = ( ~n1813 & n7334 ) | ( ~n1813 & n16494 ) | ( n7334 & n16494 ) ;
  assign n16496 = n16495 ^ n8133 ^ n6030 ;
  assign n16497 = n3341 ^ n3141 ^ 1'b0 ;
  assign n16498 = n7991 | n16497 ;
  assign n16499 = ( n10716 & ~n14956 ) | ( n10716 & n16498 ) | ( ~n14956 & n16498 ) ;
  assign n16500 = n16499 ^ n9930 ^ n7645 ;
  assign n16501 = n16496 & ~n16500 ;
  assign n16502 = n6914 & n16501 ;
  assign n16503 = ( x86 & ~n6384 ) | ( x86 & n16502 ) | ( ~n6384 & n16502 ) ;
  assign n16504 = ( n10962 & ~n16215 ) | ( n10962 & n16503 ) | ( ~n16215 & n16503 ) ;
  assign n16505 = n16491 & n16504 ;
  assign n16510 = n16509 ^ n16505 ^ 1'b0 ;
  assign n16511 = ( n4211 & ~n5654 ) | ( n4211 & n14509 ) | ( ~n5654 & n14509 ) ;
  assign n16512 = n16511 ^ n8845 ^ 1'b0 ;
  assign n16513 = n4840 & n16512 ;
  assign n16514 = n16513 ^ n10017 ^ n5551 ;
  assign n16515 = n8083 | n16514 ;
  assign n16516 = n10822 ^ n5134 ^ 1'b0 ;
  assign n16517 = n9212 & n16516 ;
  assign n16518 = ( n9283 & n11813 ) | ( n9283 & n16517 ) | ( n11813 & n16517 ) ;
  assign n16519 = n16518 ^ n12531 ^ n4132 ;
  assign n16520 = ~n3517 & n3726 ;
  assign n16521 = ( ~n2565 & n13556 ) | ( ~n2565 & n16520 ) | ( n13556 & n16520 ) ;
  assign n16522 = n727 | n16521 ;
  assign n16523 = n16522 ^ n15469 ^ n5266 ;
  assign n16533 = n9697 ^ n2502 ^ n905 ;
  assign n16534 = n16533 ^ n4411 ^ n1499 ;
  assign n16535 = n4628 & n16534 ;
  assign n16528 = ( n3933 & ~n6298 ) | ( n3933 & n15288 ) | ( ~n6298 & n15288 ) ;
  assign n16529 = n16528 ^ n14136 ^ n4891 ;
  assign n16527 = n12599 ^ n11936 ^ n1698 ;
  assign n16525 = x45 & n6181 ;
  assign n16524 = n11918 ^ n6242 ^ x136 ;
  assign n16526 = n16525 ^ n16524 ^ n9009 ;
  assign n16530 = n16529 ^ n16527 ^ n16526 ;
  assign n16531 = n12852 ^ n5465 ^ 1'b0 ;
  assign n16532 = n16530 & ~n16531 ;
  assign n16536 = n16535 ^ n16532 ^ n8343 ;
  assign n16537 = n3265 | n10277 ;
  assign n16538 = n16537 ^ n494 ^ 1'b0 ;
  assign n16539 = n16538 ^ n9239 ^ n4360 ;
  assign n16546 = n4217 ^ n3293 ^ n2804 ;
  assign n16547 = n16546 ^ n5772 ^ n1656 ;
  assign n16545 = n1127 | n10297 ;
  assign n16548 = n16547 ^ n16545 ^ 1'b0 ;
  assign n16549 = ( n392 & ~n4536 ) | ( n392 & n16548 ) | ( ~n4536 & n16548 ) ;
  assign n16540 = ( n2333 & ~n4222 ) | ( n2333 & n6863 ) | ( ~n4222 & n6863 ) ;
  assign n16541 = n2916 | n16540 ;
  assign n16542 = n2858 | n16541 ;
  assign n16543 = ( n2553 & n14212 ) | ( n2553 & ~n16542 ) | ( n14212 & ~n16542 ) ;
  assign n16544 = ( n1027 & n13322 ) | ( n1027 & n16543 ) | ( n13322 & n16543 ) ;
  assign n16550 = n16549 ^ n16544 ^ n6446 ;
  assign n16551 = n14351 ^ n8692 ^ n965 ;
  assign n16552 = n6328 | n6775 ;
  assign n16553 = n16552 ^ n739 ^ 1'b0 ;
  assign n16554 = n10407 & ~n16553 ;
  assign n16555 = ( ~n14583 & n16551 ) | ( ~n14583 & n16554 ) | ( n16551 & n16554 ) ;
  assign n16556 = n16240 ^ n10001 ^ n5797 ;
  assign n16557 = ~n8685 & n15826 ;
  assign n16558 = n16556 & n16557 ;
  assign n16559 = x41 & ~n16558 ;
  assign n16560 = n16559 ^ n9379 ^ 1'b0 ;
  assign n16562 = n7250 ^ n4162 ^ n3948 ;
  assign n16561 = ( n471 & ~n2496 ) | ( n471 & n8648 ) | ( ~n2496 & n8648 ) ;
  assign n16563 = n16562 ^ n16561 ^ n11136 ;
  assign n16568 = n14198 ^ n2315 ^ 1'b0 ;
  assign n16566 = ( ~n1057 & n8369 ) | ( ~n1057 & n14614 ) | ( n8369 & n14614 ) ;
  assign n16564 = ( n3130 & ~n8554 ) | ( n3130 & n11836 ) | ( ~n8554 & n11836 ) ;
  assign n16565 = ( n7537 & ~n13417 ) | ( n7537 & n16564 ) | ( ~n13417 & n16564 ) ;
  assign n16567 = n16566 ^ n16565 ^ n11050 ;
  assign n16569 = n16568 ^ n16567 ^ 1'b0 ;
  assign n16570 = n13763 & ~n14282 ;
  assign n16571 = ~n13163 & n16570 ;
  assign n16572 = n9545 ^ n7771 ^ n7555 ;
  assign n16573 = n8761 ^ n3387 ^ n1575 ;
  assign n16574 = n16573 ^ n14525 ^ n2706 ;
  assign n16575 = ( n4209 & ~n9551 ) | ( n4209 & n16574 ) | ( ~n9551 & n16574 ) ;
  assign n16578 = n10617 ^ n521 ^ 1'b0 ;
  assign n16579 = ( n868 & ~n16129 ) | ( n868 & n16578 ) | ( ~n16129 & n16578 ) ;
  assign n16580 = n2403 & n16579 ;
  assign n16576 = ~n9441 & n14161 ;
  assign n16577 = ~n14867 & n16576 ;
  assign n16581 = n16580 ^ n16577 ^ 1'b0 ;
  assign n16582 = n4517 & ~n16581 ;
  assign n16583 = ( ~n16572 & n16575 ) | ( ~n16572 & n16582 ) | ( n16575 & n16582 ) ;
  assign n16585 = ( n2078 & n3541 ) | ( n2078 & n7962 ) | ( n3541 & n7962 ) ;
  assign n16584 = n9602 ^ n3168 ^ 1'b0 ;
  assign n16586 = n16585 ^ n16584 ^ n5117 ;
  assign n16592 = n8648 ^ n3462 ^ n2690 ;
  assign n16593 = ( ~x109 & n5157 ) | ( ~x109 & n16592 ) | ( n5157 & n16592 ) ;
  assign n16594 = n3893 & n16593 ;
  assign n16590 = ( x248 & ~n9569 ) | ( x248 & n16158 ) | ( ~n9569 & n16158 ) ;
  assign n16591 = n16590 ^ n15533 ^ n7191 ;
  assign n16587 = ( n1211 & n5645 ) | ( n1211 & n13314 ) | ( n5645 & n13314 ) ;
  assign n16588 = n3167 ^ n1484 ^ 1'b0 ;
  assign n16589 = ~n16587 & n16588 ;
  assign n16595 = n16594 ^ n16591 ^ n16589 ;
  assign n16600 = n6562 ^ n6503 ^ n3947 ;
  assign n16599 = ( n634 & n1531 ) | ( n634 & n10161 ) | ( n1531 & n10161 ) ;
  assign n16596 = n2049 & n11886 ;
  assign n16597 = n16596 ^ n1165 ^ 1'b0 ;
  assign n16598 = n16597 ^ n14697 ^ n12721 ;
  assign n16601 = n16600 ^ n16599 ^ n16598 ;
  assign n16606 = ( n1987 & n2851 ) | ( n1987 & ~n12853 ) | ( n2851 & ~n12853 ) ;
  assign n16607 = n16606 ^ n5021 ^ n1983 ;
  assign n16602 = ( ~n1896 & n4258 ) | ( ~n1896 & n5918 ) | ( n4258 & n5918 ) ;
  assign n16603 = n16602 ^ n4364 ^ n2684 ;
  assign n16604 = ( n2112 & n13935 ) | ( n2112 & n16603 ) | ( n13935 & n16603 ) ;
  assign n16605 = n16604 ^ n14719 ^ n6733 ;
  assign n16608 = n16607 ^ n16605 ^ 1'b0 ;
  assign n16609 = n2444 ^ n2126 ^ n1293 ;
  assign n16610 = n6585 ^ n2815 ^ 1'b0 ;
  assign n16611 = ( n10334 & ~n16609 ) | ( n10334 & n16610 ) | ( ~n16609 & n16610 ) ;
  assign n16612 = n14640 ^ n417 ^ 1'b0 ;
  assign n16613 = n16611 & ~n16612 ;
  assign n16616 = n9917 ^ n6392 ^ 1'b0 ;
  assign n16614 = n6413 ^ n3605 ^ x83 ;
  assign n16615 = ( ~n1713 & n10911 ) | ( ~n1713 & n16614 ) | ( n10911 & n16614 ) ;
  assign n16617 = n16616 ^ n16615 ^ n2700 ;
  assign n16618 = n16617 ^ n10496 ^ 1'b0 ;
  assign n16619 = n16613 & n16618 ;
  assign n16620 = n15827 ^ n9361 ^ n7619 ;
  assign n16621 = n1511 & n2698 ;
  assign n16622 = n16621 ^ n9750 ^ n7636 ;
  assign n16623 = n16622 ^ n8318 ^ 1'b0 ;
  assign n16624 = n16623 ^ n9131 ^ 1'b0 ;
  assign n16626 = n8127 ^ n7364 ^ n6353 ;
  assign n16625 = n305 | n6113 ;
  assign n16627 = n16626 ^ n16625 ^ 1'b0 ;
  assign n16628 = n6936 ^ n6694 ^ n1550 ;
  assign n16629 = n16628 ^ n9591 ^ x188 ;
  assign n16630 = ~n16627 & n16629 ;
  assign n16631 = n16630 ^ n3374 ^ 1'b0 ;
  assign n16632 = n9359 ^ n5655 ^ 1'b0 ;
  assign n16633 = n4998 & n16632 ;
  assign n16637 = ( n495 & n4693 ) | ( n495 & ~n15623 ) | ( n4693 & ~n15623 ) ;
  assign n16635 = ( n379 & n538 ) | ( n379 & ~n5442 ) | ( n538 & ~n5442 ) ;
  assign n16634 = ( n5131 & n6134 ) | ( n5131 & ~n8903 ) | ( n6134 & ~n8903 ) ;
  assign n16636 = n16635 ^ n16634 ^ n3701 ;
  assign n16638 = n16637 ^ n16636 ^ n8316 ;
  assign n16639 = ( n799 & ~n7656 ) | ( n799 & n9059 ) | ( ~n7656 & n9059 ) ;
  assign n16640 = ~n2211 & n12282 ;
  assign n16644 = n10475 ^ n2197 ^ n526 ;
  assign n16643 = ( n9532 & n10390 ) | ( n9532 & ~n15511 ) | ( n10390 & ~n15511 ) ;
  assign n16641 = ( n2081 & n2824 ) | ( n2081 & n9382 ) | ( n2824 & n9382 ) ;
  assign n16642 = n16641 ^ n9950 ^ n2308 ;
  assign n16645 = n16644 ^ n16643 ^ n16642 ;
  assign n16646 = n16375 ^ n12185 ^ n4223 ;
  assign n16647 = ( n4571 & ~n5138 ) | ( n4571 & n15866 ) | ( ~n5138 & n15866 ) ;
  assign n16648 = n13823 ^ n3359 ^ 1'b0 ;
  assign n16649 = n7532 | n16648 ;
  assign n16650 = n16354 ^ n5483 ^ n1420 ;
  assign n16651 = ( n6412 & n16649 ) | ( n6412 & n16650 ) | ( n16649 & n16650 ) ;
  assign n16652 = n16651 ^ n7209 ^ n5673 ;
  assign n16657 = n9062 ^ n6185 ^ n3027 ;
  assign n16653 = x88 & ~n14217 ;
  assign n16654 = n14217 & n16653 ;
  assign n16655 = ( ~n5061 & n14675 ) | ( ~n5061 & n16654 ) | ( n14675 & n16654 ) ;
  assign n16656 = n1590 & ~n16655 ;
  assign n16658 = n16657 ^ n16656 ^ 1'b0 ;
  assign n16659 = ( n6684 & n10551 ) | ( n6684 & ~n11034 ) | ( n10551 & ~n11034 ) ;
  assign n16660 = n287 & n3737 ;
  assign n16661 = n16660 ^ n13645 ^ n316 ;
  assign n16662 = n3580 ^ n2826 ^ 1'b0 ;
  assign n16663 = ( ~n3892 & n5132 ) | ( ~n3892 & n16662 ) | ( n5132 & n16662 ) ;
  assign n16664 = ( n1149 & n3360 ) | ( n1149 & ~n5291 ) | ( n3360 & ~n5291 ) ;
  assign n16665 = n16664 ^ n14145 ^ n1094 ;
  assign n16667 = n5806 ^ n2225 ^ 1'b0 ;
  assign n16668 = n11099 ^ n5684 ^ 1'b0 ;
  assign n16669 = ( ~n8895 & n16667 ) | ( ~n8895 & n16668 ) | ( n16667 & n16668 ) ;
  assign n16666 = n5591 | n10845 ;
  assign n16670 = n16669 ^ n16666 ^ 1'b0 ;
  assign n16671 = ( n3298 & n6502 ) | ( n3298 & n9411 ) | ( n6502 & n9411 ) ;
  assign n16672 = ( n7507 & n14137 ) | ( n7507 & n16671 ) | ( n14137 & n16671 ) ;
  assign n16673 = n16672 ^ n9627 ^ 1'b0 ;
  assign n16674 = n12453 ^ n5829 ^ n1868 ;
  assign n16675 = ~n9331 & n11946 ;
  assign n16676 = n15881 ^ n9372 ^ n3565 ;
  assign n16677 = n13708 ^ n12320 ^ n1344 ;
  assign n16678 = ( n7348 & ~n16676 ) | ( n7348 & n16677 ) | ( ~n16676 & n16677 ) ;
  assign n16679 = ( n2594 & n4034 ) | ( n2594 & n6265 ) | ( n4034 & n6265 ) ;
  assign n16685 = n8577 ^ n2968 ^ n2152 ;
  assign n16686 = n16685 ^ n14949 ^ n2343 ;
  assign n16683 = n4436 ^ n3866 ^ n3573 ;
  assign n16680 = n5155 ^ n3463 ^ 1'b0 ;
  assign n16681 = n4257 & n16680 ;
  assign n16682 = n16681 ^ n15998 ^ n1872 ;
  assign n16684 = n16683 ^ n16682 ^ n13205 ;
  assign n16687 = n16686 ^ n16684 ^ n1483 ;
  assign n16688 = n11202 ^ n6693 ^ n757 ;
  assign n16689 = n8210 ^ n3334 ^ n2509 ;
  assign n16690 = ~n16309 & n16689 ;
  assign n16691 = n11806 ^ n11141 ^ n6113 ;
  assign n16692 = n4752 ^ n3326 ^ n2931 ;
  assign n16693 = ( n16690 & n16691 ) | ( n16690 & ~n16692 ) | ( n16691 & ~n16692 ) ;
  assign n16694 = ( ~n2665 & n16688 ) | ( ~n2665 & n16693 ) | ( n16688 & n16693 ) ;
  assign n16695 = n1083 & ~n2539 ;
  assign n16696 = n16219 & n16695 ;
  assign n16697 = ~n16694 & n16696 ;
  assign n16698 = n2950 & ~n5893 ;
  assign n16699 = n16698 ^ n1135 ^ 1'b0 ;
  assign n16700 = n12312 ^ n6031 ^ n4466 ;
  assign n16701 = ~n3904 & n7066 ;
  assign n16702 = n16701 ^ n10956 ^ n1233 ;
  assign n16703 = n6278 | n14683 ;
  assign n16704 = n10931 | n16703 ;
  assign n16705 = ( n7719 & n16702 ) | ( n7719 & ~n16704 ) | ( n16702 & ~n16704 ) ;
  assign n16706 = ( n16699 & n16700 ) | ( n16699 & ~n16705 ) | ( n16700 & ~n16705 ) ;
  assign n16707 = n7787 | n8036 ;
  assign n16708 = n12760 ^ n4724 ^ n845 ;
  assign n16709 = ( n2033 & ~n2265 ) | ( n2033 & n4663 ) | ( ~n2265 & n4663 ) ;
  assign n16710 = n16709 ^ n3671 ^ 1'b0 ;
  assign n16711 = n16708 & ~n16710 ;
  assign n16712 = n16707 & n16711 ;
  assign n16713 = ( x216 & ~n5031 ) | ( x216 & n7672 ) | ( ~n5031 & n7672 ) ;
  assign n16714 = n411 | n2927 ;
  assign n16715 = ( n4989 & ~n11106 ) | ( n4989 & n16714 ) | ( ~n11106 & n16714 ) ;
  assign n16716 = n9292 & n16715 ;
  assign n16717 = ~n16713 & n16716 ;
  assign n16718 = ~n482 & n7694 ;
  assign n16719 = n16718 ^ n15817 ^ 1'b0 ;
  assign n16720 = n6281 & ~n16719 ;
  assign n16721 = ( n9822 & n16717 ) | ( n9822 & ~n16720 ) | ( n16717 & ~n16720 ) ;
  assign n16722 = x251 & n1268 ;
  assign n16723 = ~n1745 & n16722 ;
  assign n16724 = n6616 | n16723 ;
  assign n16725 = n16724 ^ n12884 ^ 1'b0 ;
  assign n16726 = ( ~n10624 & n11314 ) | ( ~n10624 & n12284 ) | ( n11314 & n12284 ) ;
  assign n16727 = n16725 | n16726 ;
  assign n16728 = n4725 & ~n16727 ;
  assign n16729 = n13878 ^ n6665 ^ 1'b0 ;
  assign n16730 = n5324 | n10278 ;
  assign n16731 = ( n595 & n1862 ) | ( n595 & ~n4064 ) | ( n1862 & ~n4064 ) ;
  assign n16732 = ~n1130 & n11674 ;
  assign n16733 = ( n2560 & ~n16731 ) | ( n2560 & n16732 ) | ( ~n16731 & n16732 ) ;
  assign n16734 = ( n2993 & n6776 ) | ( n2993 & ~n16733 ) | ( n6776 & ~n16733 ) ;
  assign n16735 = ~n15430 & n16734 ;
  assign n16736 = n2875 | n16735 ;
  assign n16737 = n8804 ^ n2323 ^ n1482 ;
  assign n16738 = ( x71 & ~n9559 ) | ( x71 & n16737 ) | ( ~n9559 & n16737 ) ;
  assign n16739 = n16738 ^ n5736 ^ 1'b0 ;
  assign n16740 = n4203 | n14364 ;
  assign n16741 = ( ~n13637 & n15099 ) | ( ~n13637 & n16740 ) | ( n15099 & n16740 ) ;
  assign n16742 = n2223 | n7867 ;
  assign n16743 = n11995 | n16742 ;
  assign n16744 = n1476 | n8055 ;
  assign n16745 = n5963 & ~n8698 ;
  assign n16746 = ( n2146 & n13686 ) | ( n2146 & n16745 ) | ( n13686 & n16745 ) ;
  assign n16747 = n16746 ^ n5270 ^ 1'b0 ;
  assign n16748 = n9254 | n16747 ;
  assign n16749 = ( n1169 & n13100 ) | ( n1169 & n16748 ) | ( n13100 & n16748 ) ;
  assign n16750 = ( n1367 & ~n7445 ) | ( n1367 & n9828 ) | ( ~n7445 & n9828 ) ;
  assign n16751 = ~n3972 & n7432 ;
  assign n16752 = ( n1959 & n16750 ) | ( n1959 & n16751 ) | ( n16750 & n16751 ) ;
  assign n16756 = n10595 ^ n5073 ^ n4366 ;
  assign n16757 = ( ~n366 & n1071 ) | ( ~n366 & n2231 ) | ( n1071 & n2231 ) ;
  assign n16758 = n15760 ^ n4552 ^ n1533 ;
  assign n16759 = ( n9610 & n16757 ) | ( n9610 & n16758 ) | ( n16757 & n16758 ) ;
  assign n16760 = ( n4922 & n16756 ) | ( n4922 & n16759 ) | ( n16756 & n16759 ) ;
  assign n16753 = n5090 ^ n4247 ^ 1'b0 ;
  assign n16754 = n16753 ^ n884 ^ 1'b0 ;
  assign n16755 = n1824 & ~n16754 ;
  assign n16761 = n16760 ^ n16755 ^ n15108 ;
  assign n16762 = n6675 ^ n5071 ^ n844 ;
  assign n16763 = n8299 ^ n5157 ^ n1960 ;
  assign n16764 = n16763 ^ n4551 ^ n1905 ;
  assign n16768 = n3685 ^ n2527 ^ 1'b0 ;
  assign n16766 = ~n7796 & n15643 ;
  assign n16767 = n16766 ^ x144 ^ 1'b0 ;
  assign n16765 = ( n5258 & ~n5474 ) | ( n5258 & n8532 ) | ( ~n5474 & n8532 ) ;
  assign n16769 = n16768 ^ n16767 ^ n16765 ;
  assign n16770 = n7037 & n16769 ;
  assign n16771 = n16764 | n16770 ;
  assign n16772 = n16762 & ~n16771 ;
  assign n16773 = n12448 ^ n4285 ^ x240 ;
  assign n16774 = ( ~n522 & n3173 ) | ( ~n522 & n16773 ) | ( n3173 & n16773 ) ;
  assign n16775 = n9542 & ~n16381 ;
  assign n16776 = ~n3921 & n16775 ;
  assign n16777 = n8595 ^ n2854 ^ 1'b0 ;
  assign n16778 = n16776 | n16777 ;
  assign n16779 = ( ~n13440 & n16774 ) | ( ~n13440 & n16778 ) | ( n16774 & n16778 ) ;
  assign n16780 = ( n5774 & ~n6857 ) | ( n5774 & n13083 ) | ( ~n6857 & n13083 ) ;
  assign n16781 = n8692 ^ n3985 ^ 1'b0 ;
  assign n16782 = ( n2385 & n10800 ) | ( n2385 & ~n16781 ) | ( n10800 & ~n16781 ) ;
  assign n16783 = ( n6389 & n16780 ) | ( n6389 & n16782 ) | ( n16780 & n16782 ) ;
  assign n16784 = ( n3846 & n4836 ) | ( n3846 & n8017 ) | ( n4836 & n8017 ) ;
  assign n16785 = n16784 ^ n4607 ^ n2794 ;
  assign n16786 = n16785 ^ n15662 ^ n2572 ;
  assign n16787 = ( ~n4755 & n6396 ) | ( ~n4755 & n11140 ) | ( n6396 & n11140 ) ;
  assign n16788 = n16787 ^ n9116 ^ n5697 ;
  assign n16789 = n16788 ^ n4029 ^ n286 ;
  assign n16790 = n16789 ^ n6732 ^ n4749 ;
  assign n16791 = n7767 ^ n4934 ^ n4565 ;
  assign n16792 = n10673 ^ n9418 ^ n2530 ;
  assign n16793 = n16792 ^ n7040 ^ 1'b0 ;
  assign n16794 = ( n4311 & n16791 ) | ( n4311 & n16793 ) | ( n16791 & n16793 ) ;
  assign n16795 = n16794 ^ n12718 ^ 1'b0 ;
  assign n16796 = ~n16790 & n16795 ;
  assign n16797 = n16796 ^ n661 ^ 1'b0 ;
  assign n16798 = n3404 ^ n698 ^ 1'b0 ;
  assign n16799 = n1960 | n16798 ;
  assign n16800 = ( n6010 & n12023 ) | ( n6010 & n16799 ) | ( n12023 & n16799 ) ;
  assign n16801 = n16800 ^ n9041 ^ n5154 ;
  assign n16802 = n16801 ^ n13018 ^ 1'b0 ;
  assign n16803 = ~n16797 & n16802 ;
  assign n16804 = n12663 & n12742 ;
  assign n16805 = ~n2460 & n16804 ;
  assign n16806 = n13403 ^ n13150 ^ n4208 ;
  assign n16807 = ( n7297 & n14608 ) | ( n7297 & n16806 ) | ( n14608 & n16806 ) ;
  assign n16808 = ~n2263 & n16807 ;
  assign n16809 = n16805 & n16808 ;
  assign n16810 = n13461 ^ n10514 ^ n10256 ;
  assign n16811 = n12516 ^ n11862 ^ 1'b0 ;
  assign n16812 = n16811 ^ n8289 ^ 1'b0 ;
  assign n16813 = n2594 & n16812 ;
  assign n16814 = n11758 & n12422 ;
  assign n16815 = ~n6067 & n16814 ;
  assign n16816 = ( ~n2234 & n13615 ) | ( ~n2234 & n16815 ) | ( n13615 & n16815 ) ;
  assign n16817 = n1469 & n5376 ;
  assign n16818 = n16817 ^ n12881 ^ 1'b0 ;
  assign n16819 = n10638 & ~n16818 ;
  assign n16820 = n16819 ^ n9960 ^ 1'b0 ;
  assign n16821 = n16820 ^ n16718 ^ 1'b0 ;
  assign n16822 = ~n3866 & n16231 ;
  assign n16823 = ~n888 & n15173 ;
  assign n16824 = n12053 ^ n9277 ^ n4294 ;
  assign n16825 = x103 & n5457 ;
  assign n16826 = ~n1756 & n16825 ;
  assign n16827 = n16568 | n16826 ;
  assign n16828 = n16827 ^ n1785 ^ n1238 ;
  assign n16829 = x130 | n3991 ;
  assign n16830 = ( ~n12667 & n16828 ) | ( ~n12667 & n16829 ) | ( n16828 & n16829 ) ;
  assign n16833 = ( n1133 & n2711 ) | ( n1133 & ~n6797 ) | ( n2711 & ~n6797 ) ;
  assign n16831 = ( n5258 & n7039 ) | ( n5258 & n11078 ) | ( n7039 & n11078 ) ;
  assign n16832 = n14536 & ~n16831 ;
  assign n16834 = n16833 ^ n16832 ^ 1'b0 ;
  assign n16840 = n4631 | n13136 ;
  assign n16841 = n16840 ^ n11494 ^ 1'b0 ;
  assign n16835 = n1055 | n11845 ;
  assign n16836 = n2896 | n16835 ;
  assign n16837 = n5573 & n16836 ;
  assign n16838 = n16837 ^ n6094 ^ 1'b0 ;
  assign n16839 = ( n2833 & n16714 ) | ( n2833 & ~n16838 ) | ( n16714 & ~n16838 ) ;
  assign n16842 = n16841 ^ n16839 ^ n2251 ;
  assign n16843 = n16842 ^ n6627 ^ n2697 ;
  assign n16844 = ( n16830 & n16834 ) | ( n16830 & n16843 ) | ( n16834 & n16843 ) ;
  assign n16863 = ( x214 & ~n1082 ) | ( x214 & n14252 ) | ( ~n1082 & n14252 ) ;
  assign n16860 = ( n5053 & n6146 ) | ( n5053 & n7192 ) | ( n6146 & n7192 ) ;
  assign n16861 = n16860 ^ n5917 ^ 1'b0 ;
  assign n16862 = n8610 | n16861 ;
  assign n16845 = ( ~n304 & n1112 ) | ( ~n304 & n3480 ) | ( n1112 & n3480 ) ;
  assign n16846 = n2385 & n14569 ;
  assign n16847 = ( ~n7304 & n10711 ) | ( ~n7304 & n16846 ) | ( n10711 & n16846 ) ;
  assign n16848 = n16847 ^ n8332 ^ n3173 ;
  assign n16849 = n16848 ^ n8451 ^ 1'b0 ;
  assign n16850 = ( n3814 & n4804 ) | ( n3814 & ~n16849 ) | ( n4804 & ~n16849 ) ;
  assign n16851 = n16845 & n16850 ;
  assign n16852 = n16851 ^ n4525 ^ 1'b0 ;
  assign n16853 = ~n9159 & n16203 ;
  assign n16854 = n16852 & n16853 ;
  assign n16855 = ( n4324 & n5656 ) | ( n4324 & ~n11345 ) | ( n5656 & ~n11345 ) ;
  assign n16856 = n7830 & ~n12238 ;
  assign n16857 = ~n16855 & n16856 ;
  assign n16858 = ( n1768 & n7339 ) | ( n1768 & n16857 ) | ( n7339 & n16857 ) ;
  assign n16859 = ( ~n8688 & n16854 ) | ( ~n8688 & n16858 ) | ( n16854 & n16858 ) ;
  assign n16864 = n16863 ^ n16862 ^ n16859 ;
  assign n16872 = ( n5887 & n9807 ) | ( n5887 & ~n13014 ) | ( n9807 & ~n13014 ) ;
  assign n16868 = n11474 ^ n1996 ^ 1'b0 ;
  assign n16869 = n16868 ^ n8052 ^ n4829 ;
  assign n16865 = n8325 ^ n4658 ^ n4619 ;
  assign n16866 = ( n4479 & n8537 ) | ( n4479 & n16865 ) | ( n8537 & n16865 ) ;
  assign n16867 = ( n9809 & ~n13563 ) | ( n9809 & n16866 ) | ( ~n13563 & n16866 ) ;
  assign n16870 = n16869 ^ n16867 ^ n6357 ;
  assign n16871 = n12265 & n16870 ;
  assign n16873 = n16872 ^ n16871 ^ 1'b0 ;
  assign n16874 = n2976 & n6979 ;
  assign n16875 = n633 & ~n10966 ;
  assign n16876 = n13888 ^ n9589 ^ n6740 ;
  assign n16878 = ~n5262 & n6212 ;
  assign n16879 = n16878 ^ n434 ^ 1'b0 ;
  assign n16880 = ~n16242 & n16879 ;
  assign n16881 = n16880 ^ n5783 ^ 1'b0 ;
  assign n16882 = ( n7064 & ~n9837 ) | ( n7064 & n16881 ) | ( ~n9837 & n16881 ) ;
  assign n16883 = ( n1360 & ~n3077 ) | ( n1360 & n4890 ) | ( ~n3077 & n4890 ) ;
  assign n16884 = ( n2462 & ~n16882 ) | ( n2462 & n16883 ) | ( ~n16882 & n16883 ) ;
  assign n16877 = n16318 ^ x174 ^ x73 ;
  assign n16885 = n16884 ^ n16877 ^ n15311 ;
  assign n16890 = ( n2616 & n8684 ) | ( n2616 & ~n11922 ) | ( n8684 & ~n11922 ) ;
  assign n16886 = ( ~n4369 & n7078 ) | ( ~n4369 & n14286 ) | ( n7078 & n14286 ) ;
  assign n16887 = ( n286 & n5656 ) | ( n286 & n9272 ) | ( n5656 & n9272 ) ;
  assign n16888 = n16887 ^ n13178 ^ 1'b0 ;
  assign n16889 = ~n16886 & n16888 ;
  assign n16891 = n16890 ^ n16889 ^ n3320 ;
  assign n16892 = n8330 ^ n4816 ^ n4007 ;
  assign n16893 = n16402 ^ n4559 ^ 1'b0 ;
  assign n16894 = n557 & n16893 ;
  assign n16895 = n16894 ^ n3250 ^ n2626 ;
  assign n16896 = ( n10746 & n16892 ) | ( n10746 & n16895 ) | ( n16892 & n16895 ) ;
  assign n16897 = n15768 ^ n6308 ^ n5550 ;
  assign n16898 = n16897 ^ n11678 ^ n11291 ;
  assign n16899 = n16898 ^ n16819 ^ n15488 ;
  assign n16900 = ~n860 & n6661 ;
  assign n16901 = n7760 & n16900 ;
  assign n16902 = n1902 | n16901 ;
  assign n16903 = n16902 ^ n7917 ^ 1'b0 ;
  assign n16904 = ( ~n3177 & n16899 ) | ( ~n3177 & n16903 ) | ( n16899 & n16903 ) ;
  assign n16905 = ( ~n5625 & n5771 ) | ( ~n5625 & n10435 ) | ( n5771 & n10435 ) ;
  assign n16906 = ~n2016 & n15902 ;
  assign n16907 = n16905 & n16906 ;
  assign n16908 = n16907 ^ n10775 ^ n7911 ;
  assign n16912 = ( n1825 & n14111 ) | ( n1825 & n14281 ) | ( n14111 & n14281 ) ;
  assign n16911 = n12372 ^ n1427 ^ n370 ;
  assign n16909 = ( n3902 & n5479 ) | ( n3902 & ~n13538 ) | ( n5479 & ~n13538 ) ;
  assign n16910 = ( n5294 & ~n5573 ) | ( n5294 & n16909 ) | ( ~n5573 & n16909 ) ;
  assign n16913 = n16912 ^ n16911 ^ n16910 ;
  assign n16914 = ~n8378 & n16336 ;
  assign n16915 = n16914 ^ n14791 ^ 1'b0 ;
  assign n16916 = n4015 & ~n13213 ;
  assign n16917 = n16916 ^ n13877 ^ 1'b0 ;
  assign n16918 = n16917 ^ n6830 ^ n1136 ;
  assign n16919 = n8706 ^ n7013 ^ 1'b0 ;
  assign n16921 = n5933 ^ n3771 ^ 1'b0 ;
  assign n16922 = ~n779 & n16921 ;
  assign n16920 = ( ~n2146 & n2895 ) | ( ~n2146 & n11176 ) | ( n2895 & n11176 ) ;
  assign n16923 = n16922 ^ n16920 ^ n3266 ;
  assign n16924 = ( n13741 & n16919 ) | ( n13741 & ~n16923 ) | ( n16919 & ~n16923 ) ;
  assign n16926 = ( n3008 & n3248 ) | ( n3008 & ~n9624 ) | ( n3248 & ~n9624 ) ;
  assign n16925 = ( n2731 & n4841 ) | ( n2731 & n12417 ) | ( n4841 & n12417 ) ;
  assign n16927 = n16926 ^ n16925 ^ n6027 ;
  assign n16928 = n2546 ^ n838 ^ 1'b0 ;
  assign n16929 = ( n5218 & ~n16927 ) | ( n5218 & n16928 ) | ( ~n16927 & n16928 ) ;
  assign n16930 = n10029 ^ n3834 ^ 1'b0 ;
  assign n16931 = n8963 | n15227 ;
  assign n16932 = n6295 & n9904 ;
  assign n16933 = n16932 ^ n16379 ^ 1'b0 ;
  assign n16934 = ( n799 & n6550 ) | ( n799 & n16933 ) | ( n6550 & n16933 ) ;
  assign n16935 = n16934 ^ n8027 ^ n3564 ;
  assign n16936 = n13507 ^ n8977 ^ n3397 ;
  assign n16937 = ~n7455 & n16936 ;
  assign n16938 = ( n10678 & n16935 ) | ( n10678 & n16937 ) | ( n16935 & n16937 ) ;
  assign n16939 = n9634 ^ n8254 ^ n6288 ;
  assign n16940 = ( n4208 & ~n7871 ) | ( n4208 & n11281 ) | ( ~n7871 & n11281 ) ;
  assign n16942 = ( n2172 & ~n6897 ) | ( n2172 & n8506 ) | ( ~n6897 & n8506 ) ;
  assign n16941 = n6620 | n10018 ;
  assign n16943 = n16942 ^ n16941 ^ 1'b0 ;
  assign n16944 = n16943 ^ n12731 ^ n897 ;
  assign n16945 = n16944 ^ n15181 ^ n12714 ;
  assign n16946 = ( ~n6630 & n16940 ) | ( ~n6630 & n16945 ) | ( n16940 & n16945 ) ;
  assign n16947 = n7054 ^ n5087 ^ n3614 ;
  assign n16948 = n16947 ^ x1 ^ 1'b0 ;
  assign n16949 = n16948 ^ n16379 ^ n4792 ;
  assign n16950 = n12984 ^ n4496 ^ n777 ;
  assign n16951 = n16950 ^ n4623 ^ 1'b0 ;
  assign n16953 = ( ~n363 & n1960 ) | ( ~n363 & n2483 ) | ( n1960 & n2483 ) ;
  assign n16952 = n11075 ^ n9248 ^ 1'b0 ;
  assign n16954 = n16953 ^ n16952 ^ n11612 ;
  assign n16955 = n16954 ^ n13437 ^ n12808 ;
  assign n16957 = n9668 ^ n1908 ^ n1117 ;
  assign n16956 = ( ~n2717 & n5703 ) | ( ~n2717 & n10017 ) | ( n5703 & n10017 ) ;
  assign n16958 = n16957 ^ n16956 ^ n3471 ;
  assign n16959 = ( n16951 & n16955 ) | ( n16951 & ~n16958 ) | ( n16955 & ~n16958 ) ;
  assign n16960 = n3542 & n4454 ;
  assign n16961 = n16960 ^ n5003 ^ x43 ;
  assign n16962 = n6017 ^ n2178 ^ 1'b0 ;
  assign n16963 = n7052 & ~n16962 ;
  assign n16964 = n7067 ^ n2647 ^ 1'b0 ;
  assign n16965 = n1581 & ~n16964 ;
  assign n16968 = n13630 | n15136 ;
  assign n16966 = n13532 ^ n6152 ^ 1'b0 ;
  assign n16967 = n16966 ^ n5650 ^ n5343 ;
  assign n16969 = n16968 ^ n16967 ^ n12572 ;
  assign n16970 = ( n4535 & n6018 ) | ( n4535 & ~n10183 ) | ( n6018 & ~n10183 ) ;
  assign n16971 = n16970 ^ n6746 ^ n4504 ;
  assign n16972 = ( n5021 & n11969 ) | ( n5021 & ~n16971 ) | ( n11969 & ~n16971 ) ;
  assign n16973 = n7510 | n15706 ;
  assign n16974 = n4414 | n16973 ;
  assign n16975 = n4916 ^ n968 ^ 1'b0 ;
  assign n16976 = n16975 ^ n13101 ^ n1302 ;
  assign n16977 = ( n4327 & n11295 ) | ( n4327 & ~n16976 ) | ( n11295 & ~n16976 ) ;
  assign n16978 = n8104 ^ n4939 ^ n821 ;
  assign n16979 = ( n644 & n5077 ) | ( n644 & n6958 ) | ( n5077 & n6958 ) ;
  assign n16980 = n4788 ^ n3058 ^ 1'b0 ;
  assign n16981 = n16980 ^ n9846 ^ n7026 ;
  assign n16982 = ( ~n262 & n5719 ) | ( ~n262 & n6250 ) | ( n5719 & n6250 ) ;
  assign n16983 = ( n16979 & n16981 ) | ( n16979 & ~n16982 ) | ( n16981 & ~n16982 ) ;
  assign n16984 = n11277 ^ n11002 ^ n6606 ;
  assign n16985 = ( n5032 & n7061 ) | ( n5032 & ~n16984 ) | ( n7061 & ~n16984 ) ;
  assign n16986 = n14237 ^ n7011 ^ n5948 ;
  assign n16987 = ( n9343 & ~n12115 ) | ( n9343 & n16986 ) | ( ~n12115 & n16986 ) ;
  assign n16988 = n12533 ^ n6078 ^ n641 ;
  assign n16989 = ~n12856 & n16988 ;
  assign n16990 = ~n16987 & n16989 ;
  assign n16991 = n16985 | n16990 ;
  assign n16995 = ( n365 & n5734 ) | ( n365 & ~n10296 ) | ( n5734 & ~n10296 ) ;
  assign n16992 = n14042 ^ n9038 ^ n3637 ;
  assign n16993 = n7796 ^ n6878 ^ n1157 ;
  assign n16994 = ~n16992 & n16993 ;
  assign n16996 = n16995 ^ n16994 ^ 1'b0 ;
  assign n16997 = n2037 ^ n1009 ^ 1'b0 ;
  assign n16998 = n16997 ^ n8227 ^ n4304 ;
  assign n16999 = ~n850 & n6157 ;
  assign n17000 = ~n16998 & n16999 ;
  assign n17001 = n6429 & n17000 ;
  assign n17002 = n17001 ^ n12824 ^ n6454 ;
  assign n17003 = ( n621 & ~n6712 ) | ( n621 & n7432 ) | ( ~n6712 & n7432 ) ;
  assign n17004 = n17003 ^ n7027 ^ 1'b0 ;
  assign n17005 = n17002 & ~n17004 ;
  assign n17009 = n7792 ^ n6988 ^ n2427 ;
  assign n17006 = n1831 ^ n1397 ^ 1'b0 ;
  assign n17007 = n10838 ^ n6076 ^ n439 ;
  assign n17008 = ( x158 & n17006 ) | ( x158 & ~n17007 ) | ( n17006 & ~n17007 ) ;
  assign n17010 = n17009 ^ n17008 ^ n1416 ;
  assign n17011 = n1024 ^ n796 ^ 1'b0 ;
  assign n17012 = ~n7525 & n17011 ;
  assign n17013 = ( n2433 & ~n4748 ) | ( n2433 & n17012 ) | ( ~n4748 & n17012 ) ;
  assign n17015 = n2221 ^ n297 ^ 1'b0 ;
  assign n17016 = n1597 | n17015 ;
  assign n17014 = n8254 ^ n4652 ^ 1'b0 ;
  assign n17017 = n17016 ^ n17014 ^ n3658 ;
  assign n17018 = n10214 ^ n4087 ^ n2337 ;
  assign n17019 = n17018 ^ n6042 ^ n1736 ;
  assign n17022 = ( n1827 & ~n7253 ) | ( n1827 & n12544 ) | ( ~n7253 & n12544 ) ;
  assign n17020 = ~n6904 & n10765 ;
  assign n17021 = ~n13681 & n17020 ;
  assign n17023 = n17022 ^ n17021 ^ 1'b0 ;
  assign n17024 = n17019 & ~n17023 ;
  assign n17025 = n14465 ^ n14372 ^ n9469 ;
  assign n17026 = n9207 | n17025 ;
  assign n17027 = n2498 & ~n3560 ;
  assign n17028 = n3954 & n17027 ;
  assign n17029 = n13348 | n17028 ;
  assign n17030 = n10704 ^ n3925 ^ n385 ;
  assign n17031 = n1676 | n17030 ;
  assign n17032 = n13647 & ~n17031 ;
  assign n17033 = n1324 & ~n1807 ;
  assign n17034 = n17033 ^ n7299 ^ 1'b0 ;
  assign n17035 = ~n2421 & n17034 ;
  assign n17036 = ( n17029 & ~n17032 ) | ( n17029 & n17035 ) | ( ~n17032 & n17035 ) ;
  assign n17037 = ( n901 & ~n6303 ) | ( n901 & n8785 ) | ( ~n6303 & n8785 ) ;
  assign n17038 = n4025 ^ n437 ^ 1'b0 ;
  assign n17039 = ( n4319 & n17037 ) | ( n4319 & ~n17038 ) | ( n17037 & ~n17038 ) ;
  assign n17040 = n3520 ^ n3116 ^ 1'b0 ;
  assign n17041 = n9455 ^ n5429 ^ n2700 ;
  assign n17042 = ( ~n17016 & n17040 ) | ( ~n17016 & n17041 ) | ( n17040 & n17041 ) ;
  assign n17043 = n17042 ^ n2568 ^ 1'b0 ;
  assign n17044 = n1645 & ~n17043 ;
  assign n17045 = n17044 ^ n4063 ^ n3848 ;
  assign n17046 = x144 & ~n17045 ;
  assign n17047 = ~n17039 & n17046 ;
  assign n17049 = n7432 & ~n8112 ;
  assign n17050 = ~x190 & n17049 ;
  assign n17048 = ( ~n11007 & n13312 ) | ( ~n11007 & n15144 ) | ( n13312 & n15144 ) ;
  assign n17051 = n17050 ^ n17048 ^ n7294 ;
  assign n17056 = n12803 ^ n2494 ^ x216 ;
  assign n17052 = ( x152 & n1646 ) | ( x152 & ~n8603 ) | ( n1646 & ~n8603 ) ;
  assign n17053 = n17052 ^ n4530 ^ 1'b0 ;
  assign n17054 = n986 & n17053 ;
  assign n17055 = ( n7560 & n9457 ) | ( n7560 & ~n17054 ) | ( n9457 & ~n17054 ) ;
  assign n17057 = n17056 ^ n17055 ^ n7063 ;
  assign n17058 = n5671 ^ n1839 ^ n669 ;
  assign n17059 = n10540 ^ n8537 ^ n3519 ;
  assign n17060 = n17059 ^ n10844 ^ n8637 ;
  assign n17061 = ( n6430 & ~n11858 ) | ( n6430 & n17060 ) | ( ~n11858 & n17060 ) ;
  assign n17062 = ( n6166 & ~n6177 ) | ( n6166 & n6292 ) | ( ~n6177 & n6292 ) ;
  assign n17063 = ( n5838 & n7159 ) | ( n5838 & n10099 ) | ( n7159 & n10099 ) ;
  assign n17064 = n17063 ^ n10657 ^ n6866 ;
  assign n17065 = ( ~n4504 & n7554 ) | ( ~n4504 & n17064 ) | ( n7554 & n17064 ) ;
  assign n17066 = n13427 ^ n11923 ^ n7415 ;
  assign n17067 = ( n5903 & n12775 ) | ( n5903 & ~n17066 ) | ( n12775 & ~n17066 ) ;
  assign n17068 = ~n9703 & n15637 ;
  assign n17069 = ( n6860 & n6906 ) | ( n6860 & ~n11566 ) | ( n6906 & ~n11566 ) ;
  assign n17070 = ( n3543 & ~n5843 ) | ( n3543 & n17069 ) | ( ~n5843 & n17069 ) ;
  assign n17071 = n17070 ^ n2514 ^ n359 ;
  assign n17072 = n436 ^ n323 ^ 1'b0 ;
  assign n17073 = n716 & n17072 ;
  assign n17074 = ( n1535 & n4293 ) | ( n1535 & n17073 ) | ( n4293 & n17073 ) ;
  assign n17075 = n11151 ^ n2856 ^ 1'b0 ;
  assign n17076 = ( n1519 & ~n17074 ) | ( n1519 & n17075 ) | ( ~n17074 & n17075 ) ;
  assign n17077 = ( n3292 & n4700 ) | ( n3292 & n8126 ) | ( n4700 & n8126 ) ;
  assign n17078 = ( n1691 & ~n4437 ) | ( n1691 & n6366 ) | ( ~n4437 & n6366 ) ;
  assign n17079 = ( ~n6594 & n8965 ) | ( ~n6594 & n17078 ) | ( n8965 & n17078 ) ;
  assign n17080 = ( ~n12578 & n17077 ) | ( ~n12578 & n17079 ) | ( n17077 & n17079 ) ;
  assign n17081 = ( n4479 & n7971 ) | ( n4479 & n9831 ) | ( n7971 & n9831 ) ;
  assign n17082 = n7363 ^ n6285 ^ n3289 ;
  assign n17083 = n17081 & n17082 ;
  assign n17084 = ~n5909 & n17083 ;
  assign n17087 = n5090 ^ n4628 ^ n3230 ;
  assign n17085 = n11818 ^ n5056 ^ n1614 ;
  assign n17086 = n17085 ^ n4188 ^ n2870 ;
  assign n17088 = n17087 ^ n17086 ^ 1'b0 ;
  assign n17089 = ( n17080 & n17084 ) | ( n17080 & ~n17088 ) | ( n17084 & ~n17088 ) ;
  assign n17090 = n15886 ^ n12134 ^ n12093 ;
  assign n17091 = x17 & n1809 ;
  assign n17092 = n17091 ^ n3605 ^ 1'b0 ;
  assign n17093 = ~n16731 & n17092 ;
  assign n17094 = n17093 ^ n1646 ^ 1'b0 ;
  assign n17096 = n13305 ^ n10618 ^ n2465 ;
  assign n17097 = n17096 ^ n15713 ^ n10787 ;
  assign n17095 = ( n4254 & n12446 ) | ( n4254 & ~n13166 ) | ( n12446 & ~n13166 ) ;
  assign n17098 = n17097 ^ n17095 ^ n9697 ;
  assign n17104 = ( ~n734 & n1185 ) | ( ~n734 & n13173 ) | ( n1185 & n13173 ) ;
  assign n17105 = n8268 | n17104 ;
  assign n17106 = n12042 & ~n17105 ;
  assign n17101 = n1869 & ~n8135 ;
  assign n17102 = ~n7436 & n17101 ;
  assign n17103 = n17102 ^ n3380 ^ 1'b0 ;
  assign n17099 = n10557 ^ n9029 ^ n3765 ;
  assign n17100 = ( n3461 & n12904 ) | ( n3461 & n17099 ) | ( n12904 & n17099 ) ;
  assign n17107 = n17106 ^ n17103 ^ n17100 ;
  assign n17108 = ~n857 & n8259 ;
  assign n17109 = ( n4381 & n15334 ) | ( n4381 & n17108 ) | ( n15334 & n17108 ) ;
  assign n17116 = n10607 ^ n7614 ^ 1'b0 ;
  assign n17117 = n5330 & ~n17116 ;
  assign n17118 = n17117 ^ n9309 ^ 1'b0 ;
  assign n17119 = n5203 & n17118 ;
  assign n17114 = n13750 ^ n9521 ^ n3097 ;
  assign n17115 = n11772 & n17114 ;
  assign n17120 = n17119 ^ n17115 ^ 1'b0 ;
  assign n17110 = n6957 ^ n6835 ^ x199 ;
  assign n17111 = n9402 & ~n9492 ;
  assign n17112 = ~n5854 & n17111 ;
  assign n17113 = ( n16102 & n17110 ) | ( n16102 & n17112 ) | ( n17110 & n17112 ) ;
  assign n17121 = n17120 ^ n17113 ^ n9243 ;
  assign n17122 = ( n16827 & n17109 ) | ( n16827 & n17121 ) | ( n17109 & n17121 ) ;
  assign n17123 = ( ~n3731 & n6508 ) | ( ~n3731 & n6984 ) | ( n6508 & n6984 ) ;
  assign n17124 = n17123 ^ n6029 ^ 1'b0 ;
  assign n17125 = n11645 & n17124 ;
  assign n17126 = n17125 ^ n15306 ^ 1'b0 ;
  assign n17127 = ( n4436 & n6464 ) | ( n4436 & ~n17126 ) | ( n6464 & ~n17126 ) ;
  assign n17128 = n15331 ^ n10359 ^ n1228 ;
  assign n17129 = ( n12573 & n16830 ) | ( n12573 & n17128 ) | ( n16830 & n17128 ) ;
  assign n17131 = ( n5609 & n8590 ) | ( n5609 & n8996 ) | ( n8590 & n8996 ) ;
  assign n17132 = ( n5731 & n8237 ) | ( n5731 & n17131 ) | ( n8237 & n17131 ) ;
  assign n17133 = n1221 & ~n4478 ;
  assign n17134 = n2104 & n17133 ;
  assign n17135 = ( n12531 & ~n17132 ) | ( n12531 & n17134 ) | ( ~n17132 & n17134 ) ;
  assign n17130 = n6540 | n8679 ;
  assign n17136 = n17135 ^ n17130 ^ 1'b0 ;
  assign n17144 = n12031 ^ n5160 ^ n3920 ;
  assign n17141 = ~n4151 & n10608 ;
  assign n17142 = n17141 ^ n1714 ^ 1'b0 ;
  assign n17139 = n4785 ^ n4077 ^ n1606 ;
  assign n17137 = n1024 & ~n11429 ;
  assign n17138 = n17137 ^ n13505 ^ n11855 ;
  assign n17140 = n17139 ^ n17138 ^ n2932 ;
  assign n17143 = n17142 ^ n17140 ^ n2688 ;
  assign n17145 = n17144 ^ n17143 ^ n7191 ;
  assign n17146 = ( n3610 & n11182 ) | ( n3610 & ~n16066 ) | ( n11182 & ~n16066 ) ;
  assign n17147 = n9913 ^ n3181 ^ 1'b0 ;
  assign n17148 = n17146 & n17147 ;
  assign n17149 = n7557 ^ n5196 ^ n2170 ;
  assign n17150 = n17149 ^ n16745 ^ 1'b0 ;
  assign n17151 = ~n3785 & n17150 ;
  assign n17152 = n17151 ^ n8390 ^ n3661 ;
  assign n17159 = x185 & ~n10111 ;
  assign n17160 = n17159 ^ n7584 ^ n4897 ;
  assign n17155 = n13147 ^ n3932 ^ n1939 ;
  assign n17156 = n9106 ^ n8617 ^ n5725 ;
  assign n17157 = n17156 ^ n12171 ^ 1'b0 ;
  assign n17158 = ( n2492 & n17155 ) | ( n2492 & n17157 ) | ( n17155 & n17157 ) ;
  assign n17153 = ( n948 & n1053 ) | ( n948 & n10467 ) | ( n1053 & n10467 ) ;
  assign n17154 = n17153 ^ n6824 ^ 1'b0 ;
  assign n17161 = n17160 ^ n17158 ^ n17154 ;
  assign n17167 = n14586 ^ n2363 ^ 1'b0 ;
  assign n17168 = ~n1822 & n17167 ;
  assign n17162 = n8056 ^ n5041 ^ n4093 ;
  assign n17163 = n5506 & ~n17162 ;
  assign n17164 = n10833 & n17163 ;
  assign n17165 = n17164 ^ n6832 ^ n5776 ;
  assign n17166 = n8981 & ~n17165 ;
  assign n17169 = n17168 ^ n17166 ^ n17045 ;
  assign n17170 = n516 | n3431 ;
  assign n17171 = n12005 | n17170 ;
  assign n17172 = n5306 & ~n8364 ;
  assign n17173 = n17172 ^ n9889 ^ 1'b0 ;
  assign n17174 = n14468 ^ n13988 ^ 1'b0 ;
  assign n17175 = n2906 & n17174 ;
  assign n17176 = n17173 & n17175 ;
  assign n17177 = ~n17171 & n17176 ;
  assign n17178 = n15279 ^ n10420 ^ 1'b0 ;
  assign n17179 = ~n2444 & n17178 ;
  assign n17180 = n545 & ~n3491 ;
  assign n17181 = n6811 & ~n17180 ;
  assign n17182 = ( ~n2800 & n15038 ) | ( ~n2800 & n17181 ) | ( n15038 & n17181 ) ;
  assign n17183 = n8652 ^ n4101 ^ n478 ;
  assign n17184 = n8464 ^ n2491 ^ 1'b0 ;
  assign n17185 = n14961 ^ n4032 ^ x253 ;
  assign n17186 = ( ~n11395 & n14087 ) | ( ~n11395 & n17185 ) | ( n14087 & n17185 ) ;
  assign n17187 = ( n8197 & n9485 ) | ( n8197 & ~n17186 ) | ( n9485 & ~n17186 ) ;
  assign n17188 = ( n17183 & ~n17184 ) | ( n17183 & n17187 ) | ( ~n17184 & n17187 ) ;
  assign n17189 = ( n4312 & ~n16710 ) | ( n4312 & n17188 ) | ( ~n16710 & n17188 ) ;
  assign n17193 = ( n9772 & ~n10896 ) | ( n9772 & n12984 ) | ( ~n10896 & n12984 ) ;
  assign n17190 = ( n1629 & ~n4671 ) | ( n1629 & n11747 ) | ( ~n4671 & n11747 ) ;
  assign n17191 = ( n1147 & n6940 ) | ( n1147 & n17190 ) | ( n6940 & n17190 ) ;
  assign n17192 = n9896 & ~n17191 ;
  assign n17194 = n17193 ^ n17192 ^ 1'b0 ;
  assign n17195 = n4652 ^ n3526 ^ 1'b0 ;
  assign n17196 = n2637 & ~n17195 ;
  assign n17197 = n17196 ^ n15742 ^ 1'b0 ;
  assign n17198 = n5804 ^ n2399 ^ 1'b0 ;
  assign n17199 = n10006 & ~n17198 ;
  assign n17200 = ( n9579 & n12193 ) | ( n9579 & n17199 ) | ( n12193 & n17199 ) ;
  assign n17201 = ( n4833 & ~n5871 ) | ( n4833 & n7791 ) | ( ~n5871 & n7791 ) ;
  assign n17202 = n17201 ^ n7521 ^ n977 ;
  assign n17211 = n10243 ^ n6182 ^ 1'b0 ;
  assign n17203 = ~n6609 & n12960 ;
  assign n17204 = ( n2896 & n4847 ) | ( n2896 & n15262 ) | ( n4847 & n15262 ) ;
  assign n17205 = n17204 ^ n5591 ^ 1'b0 ;
  assign n17206 = n17203 | n17205 ;
  assign n17207 = n10861 | n17206 ;
  assign n17208 = ( n2570 & n5436 ) | ( n2570 & ~n10977 ) | ( n5436 & ~n10977 ) ;
  assign n17209 = ~n4011 & n17208 ;
  assign n17210 = ~n17207 & n17209 ;
  assign n17212 = n17211 ^ n17210 ^ n13550 ;
  assign n17213 = n5283 ^ n1185 ^ 1'b0 ;
  assign n17214 = n17213 ^ n3689 ^ n799 ;
  assign n17215 = n17214 ^ n10521 ^ 1'b0 ;
  assign n17216 = ( ~n7619 & n16437 ) | ( ~n7619 & n17215 ) | ( n16437 & n17215 ) ;
  assign n17220 = n6339 ^ n2853 ^ n2050 ;
  assign n17221 = n17220 ^ n5173 ^ 1'b0 ;
  assign n17218 = ( n2267 & ~n9199 ) | ( n2267 & n16060 ) | ( ~n9199 & n16060 ) ;
  assign n17217 = n11481 ^ n10711 ^ 1'b0 ;
  assign n17219 = n17218 ^ n17217 ^ n13040 ;
  assign n17222 = n17221 ^ n17219 ^ n10335 ;
  assign n17224 = ( ~n2619 & n2901 ) | ( ~n2619 & n4229 ) | ( n2901 & n4229 ) ;
  assign n17223 = n6404 ^ n4705 ^ n2371 ;
  assign n17225 = n17224 ^ n17223 ^ n1689 ;
  assign n17228 = n8804 ^ x242 ^ 1'b0 ;
  assign n17229 = n5625 & n17228 ;
  assign n17230 = n4970 ^ n2799 ^ 1'b0 ;
  assign n17231 = n17229 & n17230 ;
  assign n17232 = n17231 ^ n13902 ^ n7694 ;
  assign n17226 = n2440 ^ n1706 ^ 1'b0 ;
  assign n17227 = n17226 ^ n4540 ^ n2339 ;
  assign n17233 = n17232 ^ n17227 ^ n582 ;
  assign n17234 = n17233 ^ n7016 ^ n4432 ;
  assign n17235 = n3565 ^ n1616 ^ 1'b0 ;
  assign n17236 = ( n850 & n4643 ) | ( n850 & n16453 ) | ( n4643 & n16453 ) ;
  assign n17237 = ( n14510 & ~n17235 ) | ( n14510 & n17236 ) | ( ~n17235 & n17236 ) ;
  assign n17238 = n3879 ^ n2145 ^ 1'b0 ;
  assign n17239 = ( ~n4288 & n5068 ) | ( ~n4288 & n15781 ) | ( n5068 & n15781 ) ;
  assign n17242 = n1876 ^ n891 ^ n287 ;
  assign n17240 = n3718 & ~n12890 ;
  assign n17241 = n9341 & n17240 ;
  assign n17243 = n17242 ^ n17241 ^ n3012 ;
  assign n17244 = ( n2510 & n9739 ) | ( n2510 & ~n17243 ) | ( n9739 & ~n17243 ) ;
  assign n17245 = n16276 ^ n9342 ^ 1'b0 ;
  assign n17246 = ( n3505 & n5875 ) | ( n3505 & ~n10536 ) | ( n5875 & ~n10536 ) ;
  assign n17247 = n17246 ^ n9379 ^ n3172 ;
  assign n17248 = n4752 & ~n16466 ;
  assign n17249 = ( n8209 & n10892 ) | ( n8209 & ~n17248 ) | ( n10892 & ~n17248 ) ;
  assign n17250 = ( n2919 & ~n9274 ) | ( n2919 & n17249 ) | ( ~n9274 & n17249 ) ;
  assign n17253 = ( n1359 & n6699 ) | ( n1359 & ~n16676 ) | ( n6699 & ~n16676 ) ;
  assign n17251 = n3584 ^ n3178 ^ n3093 ;
  assign n17252 = n3494 | n17251 ;
  assign n17254 = n17253 ^ n17252 ^ 1'b0 ;
  assign n17255 = ~n774 & n4063 ;
  assign n17256 = ~n14843 & n17255 ;
  assign n17261 = ( ~n5590 & n7576 ) | ( ~n5590 & n10513 ) | ( n7576 & n10513 ) ;
  assign n17257 = n6595 ^ n1475 ^ 1'b0 ;
  assign n17258 = ( ~n2894 & n6103 ) | ( ~n2894 & n17257 ) | ( n6103 & n17257 ) ;
  assign n17259 = n16292 ^ n6987 ^ 1'b0 ;
  assign n17260 = n17258 & n17259 ;
  assign n17262 = n17261 ^ n17260 ^ 1'b0 ;
  assign n17263 = n17262 ^ n829 ^ 1'b0 ;
  assign n17264 = ~n17256 & n17263 ;
  assign n17265 = ( n7048 & n14976 ) | ( n7048 & ~n17264 ) | ( n14976 & ~n17264 ) ;
  assign n17266 = n9214 ^ n5446 ^ n794 ;
  assign n17267 = n11424 ^ n7693 ^ 1'b0 ;
  assign n17268 = ( x107 & n2631 ) | ( x107 & ~n6314 ) | ( n2631 & ~n6314 ) ;
  assign n17269 = n17268 ^ n4183 ^ n3547 ;
  assign n17276 = ( n5424 & n10256 ) | ( n5424 & ~n15036 ) | ( n10256 & ~n15036 ) ;
  assign n17275 = ( n5304 & n9625 ) | ( n5304 & n9635 ) | ( n9625 & n9635 ) ;
  assign n17270 = ( n6048 & ~n7666 ) | ( n6048 & n14679 ) | ( ~n7666 & n14679 ) ;
  assign n17271 = ( n3112 & n13634 ) | ( n3112 & ~n17270 ) | ( n13634 & ~n17270 ) ;
  assign n17272 = ( x67 & x208 ) | ( x67 & ~n10592 ) | ( x208 & ~n10592 ) ;
  assign n17273 = n17271 & n17272 ;
  assign n17274 = n7211 & n17273 ;
  assign n17277 = n17276 ^ n17275 ^ n17274 ;
  assign n17278 = n3408 ^ n3308 ^ n1709 ;
  assign n17283 = ( ~n3981 & n4907 ) | ( ~n3981 & n15015 ) | ( n4907 & n15015 ) ;
  assign n17284 = n17283 ^ n6127 ^ n697 ;
  assign n17279 = ~n2555 & n6501 ;
  assign n17280 = n9327 & n17279 ;
  assign n17281 = n5988 | n17280 ;
  assign n17282 = n17281 ^ n9461 ^ 1'b0 ;
  assign n17285 = n17284 ^ n17282 ^ n8147 ;
  assign n17286 = ( ~n7380 & n17278 ) | ( ~n7380 & n17285 ) | ( n17278 & n17285 ) ;
  assign n17287 = ( n4156 & n8471 ) | ( n4156 & ~n13717 ) | ( n8471 & ~n13717 ) ;
  assign n17288 = ( ~n7055 & n8612 ) | ( ~n7055 & n17287 ) | ( n8612 & n17287 ) ;
  assign n17289 = n9435 ^ n2530 ^ 1'b0 ;
  assign n17290 = n11789 ^ n11301 ^ n1541 ;
  assign n17291 = ( n12147 & ~n17289 ) | ( n12147 & n17290 ) | ( ~n17289 & n17290 ) ;
  assign n17292 = ( n9537 & n11647 ) | ( n9537 & n17291 ) | ( n11647 & n17291 ) ;
  assign n17294 = ( n1611 & n6873 ) | ( n1611 & n16082 ) | ( n6873 & n16082 ) ;
  assign n17293 = n10917 | n11211 ;
  assign n17295 = n17294 ^ n17293 ^ 1'b0 ;
  assign n17296 = n13967 & n17295 ;
  assign n17297 = n10860 & n17296 ;
  assign n17298 = n5189 | n8845 ;
  assign n17299 = n13526 & ~n17298 ;
  assign n17300 = ( n5504 & ~n11010 ) | ( n5504 & n17299 ) | ( ~n11010 & n17299 ) ;
  assign n17301 = n2502 | n4586 ;
  assign n17302 = ~n14208 & n17301 ;
  assign n17308 = n5472 ^ n4253 ^ 1'b0 ;
  assign n17304 = n16228 ^ n1132 ^ n871 ;
  assign n17305 = n17304 ^ n9753 ^ n4090 ;
  assign n17306 = n7096 | n17305 ;
  assign n17303 = n1073 & ~n10936 ;
  assign n17307 = n17306 ^ n17303 ^ 1'b0 ;
  assign n17309 = n17308 ^ n17307 ^ n9723 ;
  assign n17310 = ( n16130 & n17302 ) | ( n16130 & ~n17309 ) | ( n17302 & ~n17309 ) ;
  assign n17311 = n3470 & ~n11408 ;
  assign n17312 = n17311 ^ n14256 ^ n3503 ;
  assign n17313 = n7330 ^ n2519 ^ x96 ;
  assign n17314 = n17313 ^ n3958 ^ 1'b0 ;
  assign n17315 = n13672 | n17314 ;
  assign n17316 = ( ~n4533 & n9040 ) | ( ~n4533 & n12034 ) | ( n9040 & n12034 ) ;
  assign n17317 = n11441 & n17316 ;
  assign n17318 = n17315 & n17317 ;
  assign n17319 = n17318 ^ n8547 ^ 1'b0 ;
  assign n17320 = n5267 ^ n5213 ^ n3339 ;
  assign n17321 = n9433 & n17320 ;
  assign n17322 = ( n3790 & n11615 ) | ( n3790 & n13340 ) | ( n11615 & n13340 ) ;
  assign n17323 = n17322 ^ n17045 ^ n7319 ;
  assign n17324 = n13084 ^ n10383 ^ 1'b0 ;
  assign n17325 = ~n8547 & n17324 ;
  assign n17326 = n12118 ^ n3181 ^ 1'b0 ;
  assign n17327 = n1889 & n8963 ;
  assign n17328 = n9975 & n17327 ;
  assign n17329 = n6929 ^ n4823 ^ n2516 ;
  assign n17330 = n6774 | n17329 ;
  assign n17331 = n11373 & ~n17330 ;
  assign n17332 = n7742 & ~n17331 ;
  assign n17333 = n17332 ^ n3808 ^ 1'b0 ;
  assign n17334 = ( ~n1760 & n2615 ) | ( ~n1760 & n9097 ) | ( n2615 & n9097 ) ;
  assign n17335 = n17334 ^ n10084 ^ n2808 ;
  assign n17336 = n7871 ^ n4571 ^ n3874 ;
  assign n17337 = ( x48 & ~n1723 ) | ( x48 & n17336 ) | ( ~n1723 & n17336 ) ;
  assign n17338 = ( n1962 & n17335 ) | ( n1962 & ~n17337 ) | ( n17335 & ~n17337 ) ;
  assign n17339 = n17159 ^ n6759 ^ n1626 ;
  assign n17340 = ( n1200 & ~n10269 ) | ( n1200 & n17339 ) | ( ~n10269 & n17339 ) ;
  assign n17341 = n13914 ^ n4804 ^ 1'b0 ;
  assign n17342 = ( ~n10873 & n17340 ) | ( ~n10873 & n17341 ) | ( n17340 & n17341 ) ;
  assign n17343 = ( n5108 & ~n17338 ) | ( n5108 & n17342 ) | ( ~n17338 & n17342 ) ;
  assign n17344 = n16619 ^ n16589 ^ n870 ;
  assign n17345 = n14807 ^ n9361 ^ n5006 ;
  assign n17346 = n17345 ^ n9672 ^ 1'b0 ;
  assign n17347 = n12728 | n17346 ;
  assign n17348 = ( n1787 & n3766 ) | ( n1787 & n11211 ) | ( n3766 & n11211 ) ;
  assign n17349 = n12378 | n17348 ;
  assign n17350 = n17349 ^ n3885 ^ 1'b0 ;
  assign n17356 = ( ~n5450 & n8745 ) | ( ~n5450 & n11750 ) | ( n8745 & n11750 ) ;
  assign n17353 = n6632 | n8333 ;
  assign n17354 = n17353 ^ n8528 ^ 1'b0 ;
  assign n17355 = n17354 ^ n7168 ^ n3625 ;
  assign n17351 = ( n862 & n1446 ) | ( n862 & ~n16369 ) | ( n1446 & ~n16369 ) ;
  assign n17352 = n17351 ^ n15666 ^ n9916 ;
  assign n17357 = n17356 ^ n17355 ^ n17352 ;
  assign n17363 = n8368 ^ n4837 ^ x69 ;
  assign n17361 = ( n3116 & ~n9566 ) | ( n3116 & n13404 ) | ( ~n9566 & n13404 ) ;
  assign n17362 = n17361 ^ n6914 ^ 1'b0 ;
  assign n17364 = n17363 ^ n17362 ^ n5836 ;
  assign n17358 = n861 & ~n16406 ;
  assign n17359 = n17358 ^ n1142 ^ 1'b0 ;
  assign n17360 = ( n1231 & ~n12685 ) | ( n1231 & n17359 ) | ( ~n12685 & n17359 ) ;
  assign n17365 = n17364 ^ n17360 ^ n3774 ;
  assign n17366 = n364 & ~n4981 ;
  assign n17367 = n10300 & ~n10938 ;
  assign n17368 = n10212 & n17367 ;
  assign n17369 = ( ~n355 & n7564 ) | ( ~n355 & n9799 ) | ( n7564 & n9799 ) ;
  assign n17370 = ( n17366 & ~n17368 ) | ( n17366 & n17369 ) | ( ~n17368 & n17369 ) ;
  assign n17371 = n3767 ^ n3375 ^ n2544 ;
  assign n17372 = ( n2344 & n6194 ) | ( n2344 & n17371 ) | ( n6194 & n17371 ) ;
  assign n17373 = ( n4113 & n15523 ) | ( n4113 & n17372 ) | ( n15523 & n17372 ) ;
  assign n17374 = ( n1554 & n3366 ) | ( n1554 & n13375 ) | ( n3366 & n13375 ) ;
  assign n17375 = n10433 ^ n9042 ^ n2643 ;
  assign n17376 = n8797 ^ n6901 ^ n5584 ;
  assign n17377 = ( ~n6114 & n9572 ) | ( ~n6114 & n11284 ) | ( n9572 & n11284 ) ;
  assign n17378 = ( ~n4741 & n6893 ) | ( ~n4741 & n7329 ) | ( n6893 & n7329 ) ;
  assign n17379 = ( n17376 & n17377 ) | ( n17376 & ~n17378 ) | ( n17377 & ~n17378 ) ;
  assign n17380 = n17379 ^ n5977 ^ n1644 ;
  assign n17381 = n17380 ^ n16731 ^ n15848 ;
  assign n17382 = n13117 ^ n7873 ^ x226 ;
  assign n17383 = ( n742 & ~n11828 ) | ( n742 & n17382 ) | ( ~n11828 & n17382 ) ;
  assign n17384 = n17383 ^ n16671 ^ 1'b0 ;
  assign n17385 = ( n988 & ~n7563 ) | ( n988 & n17384 ) | ( ~n7563 & n17384 ) ;
  assign n17386 = n318 | n7192 ;
  assign n17387 = n9236 & n17386 ;
  assign n17388 = ( n7563 & ~n13114 ) | ( n7563 & n13470 ) | ( ~n13114 & n13470 ) ;
  assign n17389 = ( n4982 & ~n15010 ) | ( n4982 & n17388 ) | ( ~n15010 & n17388 ) ;
  assign n17390 = n17389 ^ n8457 ^ n4049 ;
  assign n17391 = n3395 ^ n2726 ^ n2598 ;
  assign n17392 = ( ~n3286 & n5208 ) | ( ~n3286 & n17391 ) | ( n5208 & n17391 ) ;
  assign n17393 = n15034 ^ n6866 ^ n770 ;
  assign n17394 = n17392 & ~n17393 ;
  assign n17395 = ~n6195 & n17394 ;
  assign n17409 = ( n286 & n1459 ) | ( n286 & ~n5250 ) | ( n1459 & ~n5250 ) ;
  assign n17403 = n568 | n2208 ;
  assign n17404 = n10082 & ~n17403 ;
  assign n17405 = n2943 & ~n3132 ;
  assign n17406 = ~n17404 & n17405 ;
  assign n17396 = n7090 & ~n15354 ;
  assign n17397 = n10787 ^ n9545 ^ n295 ;
  assign n17398 = n17397 ^ n12960 ^ n5396 ;
  assign n17399 = n16950 ^ n2528 ^ n2041 ;
  assign n17400 = ( ~n7019 & n10341 ) | ( ~n7019 & n17399 ) | ( n10341 & n17399 ) ;
  assign n17401 = ( ~n8773 & n14034 ) | ( ~n8773 & n17400 ) | ( n14034 & n17400 ) ;
  assign n17402 = ( n17396 & n17398 ) | ( n17396 & ~n17401 ) | ( n17398 & ~n17401 ) ;
  assign n17407 = n17406 ^ n17402 ^ n16363 ;
  assign n17408 = ( n409 & n6432 ) | ( n409 & n17407 ) | ( n6432 & n17407 ) ;
  assign n17410 = n17409 ^ n17408 ^ n1398 ;
  assign n17412 = n17034 ^ n10607 ^ n3984 ;
  assign n17413 = n17412 ^ n11717 ^ 1'b0 ;
  assign n17411 = ~n5326 & n14150 ;
  assign n17414 = n17413 ^ n17411 ^ 1'b0 ;
  assign n17415 = ( n1566 & ~n8036 ) | ( n1566 & n8591 ) | ( ~n8036 & n8591 ) ;
  assign n17416 = n1034 | n8272 ;
  assign n17417 = n17415 | n17416 ;
  assign n17418 = ( n4329 & ~n8511 ) | ( n4329 & n10358 ) | ( ~n8511 & n10358 ) ;
  assign n17419 = ( ~n671 & n9370 ) | ( ~n671 & n17418 ) | ( n9370 & n17418 ) ;
  assign n17420 = n13175 ^ n10887 ^ n9933 ;
  assign n17421 = n10344 ^ n7719 ^ n2307 ;
  assign n17422 = n17421 ^ n12031 ^ n7439 ;
  assign n17423 = n17422 ^ n7448 ^ n1306 ;
  assign n17424 = ( n1477 & n2799 ) | ( n1477 & ~n5838 ) | ( n2799 & ~n5838 ) ;
  assign n17425 = ( ~n3053 & n13712 ) | ( ~n3053 & n17424 ) | ( n13712 & n17424 ) ;
  assign n17426 = n17425 ^ n13630 ^ x34 ;
  assign n17427 = n17426 ^ n10534 ^ n10009 ;
  assign n17428 = ~n17423 & n17427 ;
  assign n17429 = ( n14328 & n17420 ) | ( n14328 & ~n17428 ) | ( n17420 & ~n17428 ) ;
  assign n17430 = n1062 ^ n1001 ^ 1'b0 ;
  assign n17431 = ~n2278 & n17430 ;
  assign n17432 = ~n1939 & n17431 ;
  assign n17433 = n9354 ^ n3604 ^ 1'b0 ;
  assign n17434 = ~n388 & n17433 ;
  assign n17435 = ( n4757 & n17432 ) | ( n4757 & ~n17434 ) | ( n17432 & ~n17434 ) ;
  assign n17436 = n10934 ^ n10447 ^ n8104 ;
  assign n17437 = ( n8755 & ~n11647 ) | ( n8755 & n17436 ) | ( ~n11647 & n17436 ) ;
  assign n17438 = n17437 ^ n8024 ^ 1'b0 ;
  assign n17439 = ( ~n5125 & n8197 ) | ( ~n5125 & n17438 ) | ( n8197 & n17438 ) ;
  assign n17440 = n11043 ^ n2385 ^ 1'b0 ;
  assign n17442 = ( n2006 & n2215 ) | ( n2006 & ~n7444 ) | ( n2215 & ~n7444 ) ;
  assign n17443 = ( ~n14378 & n16157 ) | ( ~n14378 & n17442 ) | ( n16157 & n17442 ) ;
  assign n17441 = n15025 ^ n8905 ^ n1395 ;
  assign n17444 = n17443 ^ n17441 ^ 1'b0 ;
  assign n17445 = n14050 & n17444 ;
  assign n17446 = n9962 ^ n4494 ^ n1748 ;
  assign n17447 = ( ~n11411 & n12271 ) | ( ~n11411 & n17446 ) | ( n12271 & n17446 ) ;
  assign n17448 = ( n3644 & n10744 ) | ( n3644 & n12707 ) | ( n10744 & n12707 ) ;
  assign n17450 = n9189 ^ n7146 ^ n2341 ;
  assign n17449 = ( ~n6113 & n7538 ) | ( ~n6113 & n8240 ) | ( n7538 & n8240 ) ;
  assign n17451 = n17450 ^ n17449 ^ n6431 ;
  assign n17452 = ( n733 & ~n17448 ) | ( n733 & n17451 ) | ( ~n17448 & n17451 ) ;
  assign n17453 = ~n5337 & n17452 ;
  assign n17454 = ( n3258 & n3784 ) | ( n3258 & n11957 ) | ( n3784 & n11957 ) ;
  assign n17455 = n17454 ^ n4620 ^ 1'b0 ;
  assign n17456 = n10567 ^ n3488 ^ 1'b0 ;
  assign n17457 = n7492 & ~n10458 ;
  assign n17458 = ~n4239 & n17457 ;
  assign n17459 = ( x136 & n1636 ) | ( x136 & ~n2416 ) | ( n1636 & ~n2416 ) ;
  assign n17460 = ( ~n910 & n5581 ) | ( ~n910 & n17459 ) | ( n5581 & n17459 ) ;
  assign n17461 = ( ~n10132 & n17458 ) | ( ~n10132 & n17460 ) | ( n17458 & n17460 ) ;
  assign n17462 = ( n10358 & n15027 ) | ( n10358 & n17461 ) | ( n15027 & n17461 ) ;
  assign n17467 = n9108 ^ n2731 ^ n1553 ;
  assign n17468 = ( n6776 & ~n16109 ) | ( n6776 & n17467 ) | ( ~n16109 & n17467 ) ;
  assign n17463 = ~n9149 & n10240 ;
  assign n17464 = ( n5245 & n10663 ) | ( n5245 & ~n17463 ) | ( n10663 & ~n17463 ) ;
  assign n17465 = ( n815 & ~n2565 ) | ( n815 & n17464 ) | ( ~n2565 & n17464 ) ;
  assign n17466 = n17465 ^ n13041 ^ n7544 ;
  assign n17469 = n17468 ^ n17466 ^ 1'b0 ;
  assign n17471 = n10950 ^ n4216 ^ 1'b0 ;
  assign n17470 = ( x126 & n6330 ) | ( x126 & ~n9958 ) | ( n6330 & ~n9958 ) ;
  assign n17472 = n17471 ^ n17470 ^ n2710 ;
  assign n17473 = ( n3865 & n12622 ) | ( n3865 & n17472 ) | ( n12622 & n17472 ) ;
  assign n17474 = n16184 ^ n6250 ^ n954 ;
  assign n17475 = n15607 ^ n2631 ^ 1'b0 ;
  assign n17476 = n12146 & n17475 ;
  assign n17478 = n7048 ^ n5531 ^ n1564 ;
  assign n17477 = ( n3680 & ~n3683 ) | ( n3680 & n4256 ) | ( ~n3683 & n4256 ) ;
  assign n17479 = n17478 ^ n17477 ^ n14206 ;
  assign n17480 = ( n15955 & n17476 ) | ( n15955 & n17479 ) | ( n17476 & n17479 ) ;
  assign n17481 = ( n12635 & n17474 ) | ( n12635 & n17480 ) | ( n17474 & n17480 ) ;
  assign n17482 = n5811 ^ n3756 ^ 1'b0 ;
  assign n17483 = n592 | n17482 ;
  assign n17484 = ~n8606 & n12073 ;
  assign n17485 = n17484 ^ n8126 ^ 1'b0 ;
  assign n17486 = n4724 ^ n3494 ^ 1'b0 ;
  assign n17487 = n10169 | n17486 ;
  assign n17488 = ( ~n1501 & n5600 ) | ( ~n1501 & n6154 ) | ( n5600 & n6154 ) ;
  assign n17489 = ( ~n2762 & n17487 ) | ( ~n2762 & n17488 ) | ( n17487 & n17488 ) ;
  assign n17490 = ( n1816 & ~n17485 ) | ( n1816 & n17489 ) | ( ~n17485 & n17489 ) ;
  assign n17491 = ( n7044 & n7324 ) | ( n7044 & n12892 ) | ( n7324 & n12892 ) ;
  assign n17492 = n15823 ^ n7757 ^ x75 ;
  assign n17493 = ( ~n1443 & n9577 ) | ( ~n1443 & n14896 ) | ( n9577 & n14896 ) ;
  assign n17494 = ( n12282 & n17492 ) | ( n12282 & n17493 ) | ( n17492 & n17493 ) ;
  assign n17495 = ( n10914 & n17491 ) | ( n10914 & n17494 ) | ( n17491 & n17494 ) ;
  assign n17496 = n6364 ^ n5072 ^ n336 ;
  assign n17497 = n4759 ^ n2970 ^ 1'b0 ;
  assign n17498 = n17496 & n17497 ;
  assign n17499 = ~n7898 & n17498 ;
  assign n17505 = n15139 ^ n8032 ^ n3987 ;
  assign n17501 = ( x162 & n4670 ) | ( x162 & n5270 ) | ( n4670 & n5270 ) ;
  assign n17502 = n2827 & ~n5602 ;
  assign n17503 = n17502 ^ n14862 ^ 1'b0 ;
  assign n17504 = ( n15951 & ~n17501 ) | ( n15951 & n17503 ) | ( ~n17501 & n17503 ) ;
  assign n17500 = ( n6559 & ~n9727 ) | ( n6559 & n14351 ) | ( ~n9727 & n14351 ) ;
  assign n17506 = n17505 ^ n17504 ^ n17500 ;
  assign n17507 = ~n326 & n6870 ;
  assign n17508 = n17507 ^ n16866 ^ n8610 ;
  assign n17509 = n17508 ^ n12162 ^ n6503 ;
  assign n17510 = ~n13928 & n16168 ;
  assign n17511 = n14227 & n17510 ;
  assign n17516 = ( n846 & ~n3042 ) | ( n846 & n4115 ) | ( ~n3042 & n4115 ) ;
  assign n17512 = n10849 ^ n7975 ^ n468 ;
  assign n17513 = n9600 ^ n6065 ^ n903 ;
  assign n17514 = n17513 ^ n9874 ^ 1'b0 ;
  assign n17515 = ( n519 & n17512 ) | ( n519 & ~n17514 ) | ( n17512 & ~n17514 ) ;
  assign n17517 = n17516 ^ n17515 ^ n15080 ;
  assign n17518 = ( ~n5074 & n7923 ) | ( ~n5074 & n9111 ) | ( n7923 & n9111 ) ;
  assign n17519 = ~n9921 & n17518 ;
  assign n17520 = ( n5838 & n6579 ) | ( n5838 & ~n17519 ) | ( n6579 & ~n17519 ) ;
  assign n17521 = ( n9235 & ~n11951 ) | ( n9235 & n15048 ) | ( ~n11951 & n15048 ) ;
  assign n17522 = n12302 ^ n5372 ^ n3630 ;
  assign n17523 = ( n1387 & n3718 ) | ( n1387 & n4681 ) | ( n3718 & n4681 ) ;
  assign n17524 = ( n5671 & n17522 ) | ( n5671 & n17523 ) | ( n17522 & n17523 ) ;
  assign n17525 = n16886 ^ n12354 ^ n8382 ;
  assign n17526 = n7290 ^ n1317 ^ 1'b0 ;
  assign n17527 = n1595 | n17526 ;
  assign n17528 = n17527 ^ n12340 ^ n6919 ;
  assign n17529 = n17528 ^ n8461 ^ n692 ;
  assign n17530 = ( n855 & n1897 ) | ( n855 & n3119 ) | ( n1897 & n3119 ) ;
  assign n17531 = ( n3084 & n9761 ) | ( n3084 & n17530 ) | ( n9761 & n17530 ) ;
  assign n17532 = ( n7357 & n9597 ) | ( n7357 & ~n17531 ) | ( n9597 & ~n17531 ) ;
  assign n17533 = n6669 & ~n10252 ;
  assign n17534 = ( n2937 & n11396 ) | ( n2937 & ~n13231 ) | ( n11396 & ~n13231 ) ;
  assign n17535 = ( n4972 & n8823 ) | ( n4972 & n17534 ) | ( n8823 & n17534 ) ;
  assign n17536 = n14706 ^ n13510 ^ 1'b0 ;
  assign n17537 = n10084 ^ n7141 ^ n5289 ;
  assign n17538 = ~n2327 & n17537 ;
  assign n17539 = ~n17536 & n17538 ;
  assign n17540 = ( n1689 & n14493 ) | ( n1689 & n15356 ) | ( n14493 & n15356 ) ;
  assign n17541 = ( ~n7061 & n8728 ) | ( ~n7061 & n15185 ) | ( n8728 & n15185 ) ;
  assign n17542 = n4465 ^ n1767 ^ 1'b0 ;
  assign n17543 = n2096 & n17542 ;
  assign n17544 = n17543 ^ n4448 ^ n1876 ;
  assign n17545 = ( x11 & x200 ) | ( x11 & n3987 ) | ( x200 & n3987 ) ;
  assign n17546 = n17545 ^ n4900 ^ 1'b0 ;
  assign n17547 = n17544 & ~n17546 ;
  assign n17548 = n14121 ^ n739 ^ n448 ;
  assign n17549 = ~n4948 & n17548 ;
  assign n17550 = ( n5244 & n17356 ) | ( n5244 & n17549 ) | ( n17356 & n17549 ) ;
  assign n17551 = n17550 ^ n10767 ^ 1'b0 ;
  assign n17552 = ( n15610 & n17547 ) | ( n15610 & ~n17551 ) | ( n17547 & ~n17551 ) ;
  assign n17553 = ( n1523 & n3560 ) | ( n1523 & ~n8241 ) | ( n3560 & ~n8241 ) ;
  assign n17554 = n1215 & ~n17553 ;
  assign n17557 = n7691 ^ n1296 ^ x79 ;
  assign n17558 = ~n1500 & n7150 ;
  assign n17559 = ~n17557 & n17558 ;
  assign n17555 = n4972 & n9311 ;
  assign n17556 = n12666 | n17555 ;
  assign n17560 = n17559 ^ n17556 ^ n10950 ;
  assign n17561 = ~n1296 & n5195 ;
  assign n17562 = n17561 ^ n3380 ^ 1'b0 ;
  assign n17563 = ( n6177 & ~n7760 ) | ( n6177 & n8503 ) | ( ~n7760 & n8503 ) ;
  assign n17564 = ( ~n9970 & n10704 ) | ( ~n9970 & n16614 ) | ( n10704 & n16614 ) ;
  assign n17565 = n8833 ^ x137 ^ 1'b0 ;
  assign n17566 = ~n17564 & n17565 ;
  assign n17567 = ( n17562 & n17563 ) | ( n17562 & ~n17566 ) | ( n17563 & ~n17566 ) ;
  assign n17568 = n9148 ^ n7609 ^ n2248 ;
  assign n17569 = n13301 & n17568 ;
  assign n17571 = ( n6919 & ~n11094 ) | ( n6919 & n14903 ) | ( ~n11094 & n14903 ) ;
  assign n17570 = ( ~n2927 & n2954 ) | ( ~n2927 & n11377 ) | ( n2954 & n11377 ) ;
  assign n17572 = n17571 ^ n17570 ^ n2120 ;
  assign n17574 = n5178 ^ n1411 ^ 1'b0 ;
  assign n17575 = n9624 ^ n3570 ^ 1'b0 ;
  assign n17576 = n17574 | n17575 ;
  assign n17577 = ( x33 & n6443 ) | ( x33 & n17576 ) | ( n6443 & n17576 ) ;
  assign n17578 = n17577 ^ n12743 ^ n1824 ;
  assign n17573 = n11395 ^ n3978 ^ n3872 ;
  assign n17579 = n17578 ^ n17573 ^ n3058 ;
  assign n17580 = n17579 ^ n6739 ^ 1'b0 ;
  assign n17581 = n13175 ^ n8038 ^ 1'b0 ;
  assign n17582 = n9361 & n14166 ;
  assign n17583 = n17582 ^ n8770 ^ n6349 ;
  assign n17584 = ~n5310 & n17583 ;
  assign n17585 = ~n17322 & n17584 ;
  assign n17586 = n9841 & n14500 ;
  assign n17587 = n17586 ^ n16704 ^ n15963 ;
  assign n17588 = n4051 ^ n1034 ^ 1'b0 ;
  assign n17589 = n9224 | n17588 ;
  assign n17590 = n10271 & ~n17589 ;
  assign n17591 = ( n1050 & ~n1180 ) | ( n1050 & n1419 ) | ( ~n1180 & n1419 ) ;
  assign n17592 = n17591 ^ n8784 ^ n1986 ;
  assign n17593 = ( n3498 & n5217 ) | ( n3498 & ~n17592 ) | ( n5217 & ~n17592 ) ;
  assign n17594 = n9501 ^ n3629 ^ x16 ;
  assign n17595 = ( n9206 & n12701 ) | ( n9206 & ~n17594 ) | ( n12701 & ~n17594 ) ;
  assign n17596 = n10777 ^ n1428 ^ x1 ;
  assign n17597 = n6197 & ~n17042 ;
  assign n17598 = ~n12814 & n17597 ;
  assign n17599 = n17596 & n17598 ;
  assign n17600 = n4670 & ~n16770 ;
  assign n17601 = n17600 ^ n2975 ^ 1'b0 ;
  assign n17602 = ( n5205 & n6751 ) | ( n5205 & ~n17601 ) | ( n6751 & ~n17601 ) ;
  assign n17604 = n9995 ^ n3174 ^ n1599 ;
  assign n17603 = ~n965 & n4391 ;
  assign n17605 = n17604 ^ n17603 ^ 1'b0 ;
  assign n17607 = n9900 ^ n9091 ^ n8794 ;
  assign n17606 = n7727 & ~n12332 ;
  assign n17608 = n17607 ^ n17606 ^ n1500 ;
  assign n17611 = n16094 ^ n8716 ^ n2299 ;
  assign n17612 = n13069 & n17611 ;
  assign n17610 = n898 & n2335 ;
  assign n17613 = n17612 ^ n17610 ^ 1'b0 ;
  assign n17614 = n17613 ^ n9680 ^ n5406 ;
  assign n17609 = ( n2613 & n12792 ) | ( n2613 & n15503 ) | ( n12792 & n15503 ) ;
  assign n17615 = n17614 ^ n17609 ^ 1'b0 ;
  assign n17616 = n17608 & ~n17615 ;
  assign n17624 = n12989 ^ n7593 ^ 1'b0 ;
  assign n17621 = ( ~n1001 & n5855 ) | ( ~n1001 & n12648 ) | ( n5855 & n12648 ) ;
  assign n17622 = n1528 | n17621 ;
  assign n17620 = ( n651 & n1223 ) | ( n651 & ~n6287 ) | ( n1223 & ~n6287 ) ;
  assign n17619 = n9568 ^ n6043 ^ n4098 ;
  assign n17623 = n17622 ^ n17620 ^ n17619 ;
  assign n17617 = n7319 & ~n9834 ;
  assign n17618 = ( n4511 & ~n7135 ) | ( n4511 & n17617 ) | ( ~n7135 & n17617 ) ;
  assign n17625 = n17624 ^ n17623 ^ n17618 ;
  assign n17626 = n17625 ^ n12778 ^ n4839 ;
  assign n17627 = ( ~n2404 & n10837 ) | ( ~n2404 & n11091 ) | ( n10837 & n11091 ) ;
  assign n17628 = n17627 ^ n8459 ^ n8439 ;
  assign n17629 = n16300 ^ n6038 ^ n1226 ;
  assign n17630 = ( n14364 & ~n16733 ) | ( n14364 & n17629 ) | ( ~n16733 & n17629 ) ;
  assign n17631 = n9925 | n17630 ;
  assign n17632 = n14021 & ~n15058 ;
  assign n17633 = n17632 ^ n431 ^ 1'b0 ;
  assign n17634 = ( ~n4724 & n17631 ) | ( ~n4724 & n17633 ) | ( n17631 & n17633 ) ;
  assign n17635 = n13826 ^ n4441 ^ 1'b0 ;
  assign n17638 = n10267 ^ n5841 ^ n589 ;
  assign n17636 = n9995 ^ n7964 ^ 1'b0 ;
  assign n17637 = n17636 ^ n9762 ^ n9613 ;
  assign n17639 = n17638 ^ n17637 ^ n7341 ;
  assign n17640 = n17040 ^ n9937 ^ n362 ;
  assign n17641 = ( n6778 & ~n9857 ) | ( n6778 & n17640 ) | ( ~n9857 & n17640 ) ;
  assign n17642 = n17641 ^ n17386 ^ n3272 ;
  assign n17643 = n11467 & ~n17642 ;
  assign n17644 = ~n17639 & n17643 ;
  assign n17645 = n12368 ^ n7082 ^ 1'b0 ;
  assign n17646 = ~n12827 & n17645 ;
  assign n17647 = ~n15701 & n17646 ;
  assign n17648 = n10187 ^ n8225 ^ n4956 ;
  assign n17649 = ( n6600 & ~n16733 ) | ( n6600 & n17648 ) | ( ~n16733 & n17648 ) ;
  assign n17650 = n868 ^ n795 ^ 1'b0 ;
  assign n17651 = n14007 ^ n4591 ^ n3710 ;
  assign n17652 = n17651 ^ n4082 ^ 1'b0 ;
  assign n17653 = ( n12716 & ~n17650 ) | ( n12716 & n17652 ) | ( ~n17650 & n17652 ) ;
  assign n17654 = n17653 ^ n11417 ^ n3755 ;
  assign n17655 = n16689 ^ n8777 ^ n5093 ;
  assign n17656 = ~n6718 & n17655 ;
  assign n17657 = n17654 & n17656 ;
  assign n17658 = n8002 ^ n5355 ^ 1'b0 ;
  assign n17659 = ~n1419 & n17658 ;
  assign n17660 = n17659 ^ n3293 ^ n442 ;
  assign n17661 = n1427 & ~n2182 ;
  assign n17662 = n17661 ^ n5924 ^ 1'b0 ;
  assign n17663 = ( n5486 & n9081 ) | ( n5486 & ~n17662 ) | ( n9081 & ~n17662 ) ;
  assign n17664 = n8111 ^ n3113 ^ 1'b0 ;
  assign n17665 = ( n17660 & n17663 ) | ( n17660 & ~n17664 ) | ( n17663 & ~n17664 ) ;
  assign n17668 = n10664 ^ n9153 ^ n3328 ;
  assign n17666 = ( ~n1691 & n2268 ) | ( ~n1691 & n5737 ) | ( n2268 & n5737 ) ;
  assign n17667 = ( n5831 & n11770 ) | ( n5831 & ~n17666 ) | ( n11770 & ~n17666 ) ;
  assign n17669 = n17668 ^ n17667 ^ 1'b0 ;
  assign n17670 = ( ~n5474 & n5757 ) | ( ~n5474 & n17553 ) | ( n5757 & n17553 ) ;
  assign n17678 = n11141 ^ n4362 ^ n1445 ;
  assign n17677 = n10045 ^ n5185 ^ 1'b0 ;
  assign n17671 = n2722 ^ n1804 ^ 1'b0 ;
  assign n17672 = n2278 | n17671 ;
  assign n17673 = n5899 | n17672 ;
  assign n17674 = n17673 ^ n7717 ^ 1'b0 ;
  assign n17675 = ( n764 & n4935 ) | ( n764 & ~n17674 ) | ( n4935 & ~n17674 ) ;
  assign n17676 = ( n9551 & ~n12416 ) | ( n9551 & n17675 ) | ( ~n12416 & n17675 ) ;
  assign n17679 = n17678 ^ n17677 ^ n17676 ;
  assign n17680 = n16023 ^ n4194 ^ 1'b0 ;
  assign n17681 = n6749 & n17680 ;
  assign n17682 = n4165 ^ n2935 ^ n1139 ;
  assign n17683 = ( ~n10458 & n13586 ) | ( ~n10458 & n17682 ) | ( n13586 & n17682 ) ;
  assign n17684 = ( n6429 & n6562 ) | ( n6429 & n9129 ) | ( n6562 & n9129 ) ;
  assign n17685 = ( n5347 & ~n6278 ) | ( n5347 & n17684 ) | ( ~n6278 & n17684 ) ;
  assign n17686 = ( n267 & n17683 ) | ( n267 & n17685 ) | ( n17683 & n17685 ) ;
  assign n17687 = ( n7910 & n17681 ) | ( n7910 & n17686 ) | ( n17681 & n17686 ) ;
  assign n17688 = ( ~n10830 & n15001 ) | ( ~n10830 & n17687 ) | ( n15001 & n17687 ) ;
  assign n17689 = n7562 ^ n6937 ^ n3392 ;
  assign n17690 = ~n2773 & n5445 ;
  assign n17691 = n6223 & n17690 ;
  assign n17692 = n17691 ^ n1157 ^ n292 ;
  assign n17693 = ( ~n8528 & n17689 ) | ( ~n8528 & n17692 ) | ( n17689 & n17692 ) ;
  assign n17694 = n2176 ^ n448 ^ 1'b0 ;
  assign n17695 = n17693 | n17694 ;
  assign n17696 = n7265 ^ n2783 ^ 1'b0 ;
  assign n17697 = n8020 | n17696 ;
  assign n17698 = n2233 | n17697 ;
  assign n17699 = ( n578 & n2963 ) | ( n578 & ~n6777 ) | ( n2963 & ~n6777 ) ;
  assign n17700 = n17699 ^ n13070 ^ 1'b0 ;
  assign n17701 = n13573 ^ n10385 ^ n4040 ;
  assign n17702 = ( x50 & ~n12596 ) | ( x50 & n17701 ) | ( ~n12596 & n17701 ) ;
  assign n17703 = ( n4000 & n4443 ) | ( n4000 & ~n12266 ) | ( n4443 & ~n12266 ) ;
  assign n17704 = ( n2724 & ~n17702 ) | ( n2724 & n17703 ) | ( ~n17702 & n17703 ) ;
  assign n17707 = n17000 ^ x193 ^ 1'b0 ;
  assign n17708 = n17707 ^ n11999 ^ n2490 ;
  assign n17705 = n15278 ^ n8099 ^ 1'b0 ;
  assign n17706 = n6297 & n17705 ;
  assign n17709 = n17708 ^ n17706 ^ n10792 ;
  assign n17710 = ~n12566 & n17709 ;
  assign n17711 = n17710 ^ n14451 ^ 1'b0 ;
  assign n17712 = n8147 ^ n7419 ^ n1499 ;
  assign n17713 = ( n5117 & ~n8832 ) | ( n5117 & n17712 ) | ( ~n8832 & n17712 ) ;
  assign n17716 = ( n1372 & n4905 ) | ( n1372 & n9210 ) | ( n4905 & n9210 ) ;
  assign n17717 = ( n10725 & n13378 ) | ( n10725 & n17716 ) | ( n13378 & n17716 ) ;
  assign n17718 = ~n3560 & n17717 ;
  assign n17719 = n7464 & n17718 ;
  assign n17714 = ( n487 & n3916 ) | ( n487 & ~n4534 ) | ( n3916 & ~n4534 ) ;
  assign n17715 = ( n2704 & ~n17553 ) | ( n2704 & n17714 ) | ( ~n17553 & n17714 ) ;
  assign n17720 = n17719 ^ n17715 ^ n1129 ;
  assign n17721 = n3948 | n4170 ;
  assign n17723 = n3983 ^ n3318 ^ n2920 ;
  assign n17722 = n10140 ^ n4355 ^ n781 ;
  assign n17724 = n17723 ^ n17722 ^ 1'b0 ;
  assign n17725 = n5436 & ~n17724 ;
  assign n17726 = ~n11188 & n17725 ;
  assign n17727 = n17726 ^ n377 ^ 1'b0 ;
  assign n17728 = n17727 ^ n16538 ^ 1'b0 ;
  assign n17729 = n17728 ^ n9082 ^ n1407 ;
  assign n17730 = ( ~n4705 & n17721 ) | ( ~n4705 & n17729 ) | ( n17721 & n17729 ) ;
  assign n17731 = n2528 ^ n2250 ^ n809 ;
  assign n17732 = n17731 ^ n5961 ^ 1'b0 ;
  assign n17733 = n16850 ^ n12374 ^ 1'b0 ;
  assign n17734 = n9376 & n17733 ;
  assign n17735 = ( ~n5213 & n8410 ) | ( ~n5213 & n17734 ) | ( n8410 & n17734 ) ;
  assign n17736 = ( n6238 & n11570 ) | ( n6238 & ~n16258 ) | ( n11570 & ~n16258 ) ;
  assign n17737 = ( n8750 & n9249 ) | ( n8750 & ~n11696 ) | ( n9249 & ~n11696 ) ;
  assign n17738 = ( n10191 & n13147 ) | ( n10191 & ~n13994 ) | ( n13147 & ~n13994 ) ;
  assign n17739 = ( n6554 & ~n11457 ) | ( n6554 & n17738 ) | ( ~n11457 & n17738 ) ;
  assign n17740 = n14666 ^ n8769 ^ 1'b0 ;
  assign n17741 = ~x227 & n16670 ;
  assign n17742 = ( n3022 & n4607 ) | ( n3022 & ~n12125 ) | ( n4607 & ~n12125 ) ;
  assign n17743 = ~n6621 & n10888 ;
  assign n17744 = n17743 ^ n1636 ^ 1'b0 ;
  assign n17745 = n10274 & ~n17744 ;
  assign n17746 = ~n9441 & n17745 ;
  assign n17747 = n17742 & n17746 ;
  assign n17748 = n4006 | n17747 ;
  assign n17749 = n7843 ^ n7517 ^ n3580 ;
  assign n17750 = ( n594 & n2660 ) | ( n594 & ~n17749 ) | ( n2660 & ~n17749 ) ;
  assign n17751 = ( n4643 & n6610 ) | ( n4643 & ~n17750 ) | ( n6610 & ~n17750 ) ;
  assign n17752 = n697 | n12828 ;
  assign n17753 = ( n2018 & ~n12223 ) | ( n2018 & n15961 ) | ( ~n12223 & n15961 ) ;
  assign n17754 = n17753 ^ n8398 ^ 1'b0 ;
  assign n17755 = n15058 ^ n7574 ^ 1'b0 ;
  assign n17756 = n17754 & ~n17755 ;
  assign n17757 = n17756 ^ n12232 ^ n11225 ;
  assign n17758 = ( n6926 & n17752 ) | ( n6926 & ~n17757 ) | ( n17752 & ~n17757 ) ;
  assign n17759 = ( n4466 & n17751 ) | ( n4466 & ~n17758 ) | ( n17751 & ~n17758 ) ;
  assign n17760 = ~n4426 & n6943 ;
  assign n17761 = n11337 ^ n6690 ^ n6486 ;
  assign n17762 = n12828 ^ n8075 ^ n2112 ;
  assign n17763 = ( ~n8955 & n17761 ) | ( ~n8955 & n17762 ) | ( n17761 & n17762 ) ;
  assign n17764 = n11385 & n15507 ;
  assign n17765 = ( n17760 & n17763 ) | ( n17760 & n17764 ) | ( n17763 & n17764 ) ;
  assign n17766 = n14412 ^ n12715 ^ 1'b0 ;
  assign n17767 = n5456 & ~n17766 ;
  assign n17773 = ~n4687 & n12344 ;
  assign n17774 = ~n4780 & n17773 ;
  assign n17775 = ( n2024 & n16432 ) | ( n2024 & n17774 ) | ( n16432 & n17774 ) ;
  assign n17768 = ( n885 & n4241 ) | ( n885 & n14570 ) | ( n4241 & n14570 ) ;
  assign n17769 = n17768 ^ n3605 ^ 1'b0 ;
  assign n17770 = n17248 ^ n8738 ^ 1'b0 ;
  assign n17771 = ~n17769 & n17770 ;
  assign n17772 = n17262 & n17771 ;
  assign n17776 = n17775 ^ n17772 ^ 1'b0 ;
  assign n17784 = ( ~n535 & n4005 ) | ( ~n535 & n14371 ) | ( n4005 & n14371 ) ;
  assign n17780 = n1285 | n3279 ;
  assign n17781 = n5273 & ~n17780 ;
  assign n17782 = ( n5328 & ~n7747 ) | ( n5328 & n17781 ) | ( ~n7747 & n17781 ) ;
  assign n17779 = ( x104 & n8051 ) | ( x104 & ~n12685 ) | ( n8051 & ~n12685 ) ;
  assign n17777 = ( n8261 & n8765 ) | ( n8261 & n11466 ) | ( n8765 & n11466 ) ;
  assign n17778 = n17777 ^ n8876 ^ n511 ;
  assign n17783 = n17782 ^ n17779 ^ n17778 ;
  assign n17785 = n17784 ^ n17783 ^ 1'b0 ;
  assign n17786 = ( n312 & n6408 ) | ( n312 & n13667 ) | ( n6408 & n13667 ) ;
  assign n17787 = n9395 ^ n4792 ^ n3785 ;
  assign n17788 = n17787 ^ n12349 ^ 1'b0 ;
  assign n17789 = n7681 & ~n17788 ;
  assign n17791 = n15891 ^ n13014 ^ n5689 ;
  assign n17790 = ( ~n733 & n4109 ) | ( ~n733 & n11390 ) | ( n4109 & n11390 ) ;
  assign n17792 = n17791 ^ n17790 ^ n5840 ;
  assign n17803 = n8900 ^ n4100 ^ n683 ;
  assign n17804 = n17803 ^ n1733 ^ n518 ;
  assign n17805 = ( n4996 & ~n15518 ) | ( n4996 & n17804 ) | ( ~n15518 & n17804 ) ;
  assign n17806 = n17805 ^ n9616 ^ 1'b0 ;
  assign n17800 = n14840 ^ n7594 ^ 1'b0 ;
  assign n17801 = n12496 & ~n17800 ;
  assign n17798 = ( x25 & ~n889 ) | ( x25 & n1868 ) | ( ~n889 & n1868 ) ;
  assign n17799 = n3478 & n17798 ;
  assign n17802 = n17801 ^ n17799 ^ 1'b0 ;
  assign n17807 = n17806 ^ n17802 ^ n12456 ;
  assign n17793 = x227 ^ x87 ^ 1'b0 ;
  assign n17794 = ~n16621 & n17793 ;
  assign n17795 = ( ~x143 & n7764 ) | ( ~x143 & n17794 ) | ( n7764 & n17794 ) ;
  assign n17796 = ( n3149 & n7686 ) | ( n3149 & ~n17795 ) | ( n7686 & ~n17795 ) ;
  assign n17797 = n17796 ^ n8943 ^ n8747 ;
  assign n17808 = n17807 ^ n17797 ^ n11779 ;
  assign n17809 = ( ~n8582 & n10425 ) | ( ~n8582 & n17808 ) | ( n10425 & n17808 ) ;
  assign n17811 = n6798 & ~n11302 ;
  assign n17812 = n3079 & n17811 ;
  assign n17810 = n16236 ^ n13594 ^ n8455 ;
  assign n17813 = n17812 ^ n17810 ^ n2224 ;
  assign n17814 = n16081 ^ n14945 ^ n6414 ;
  assign n17815 = n17814 ^ n6491 ^ n4209 ;
  assign n17816 = ( n2439 & n8006 ) | ( n2439 & ~n10328 ) | ( n8006 & ~n10328 ) ;
  assign n17817 = ( n774 & ~n3347 ) | ( n774 & n17816 ) | ( ~n3347 & n17816 ) ;
  assign n17818 = n4725 | n13860 ;
  assign n17819 = n17818 ^ n5637 ^ 1'b0 ;
  assign n17820 = ( n4212 & n4847 ) | ( n4212 & n15904 ) | ( n4847 & n15904 ) ;
  assign n17821 = n17820 ^ n9628 ^ n4980 ;
  assign n17822 = n1749 ^ n1623 ^ 1'b0 ;
  assign n17823 = ~n903 & n17822 ;
  assign n17824 = ( x161 & n4222 ) | ( x161 & n17823 ) | ( n4222 & n17823 ) ;
  assign n17825 = ( ~n17819 & n17821 ) | ( ~n17819 & n17824 ) | ( n17821 & n17824 ) ;
  assign n17826 = n17825 ^ n5640 ^ 1'b0 ;
  assign n17827 = ~n17817 & n17826 ;
  assign n17828 = n8777 ^ n7070 ^ 1'b0 ;
  assign n17829 = n2846 & ~n17828 ;
  assign n17830 = n5504 ^ n1390 ^ 1'b0 ;
  assign n17831 = n3553 & n17830 ;
  assign n17832 = ~n8269 & n17831 ;
  assign n17833 = n11918 & n17832 ;
  assign n17834 = n8760 ^ n5204 ^ 1'b0 ;
  assign n17835 = n511 | n17834 ;
  assign n17836 = n17660 & n17835 ;
  assign n17837 = n17833 & n17836 ;
  assign n17838 = ( n599 & n793 ) | ( n599 & n15878 ) | ( n793 & n15878 ) ;
  assign n17839 = ( n12610 & ~n13718 ) | ( n12610 & n17838 ) | ( ~n13718 & n17838 ) ;
  assign n17840 = n13594 ^ n12667 ^ 1'b0 ;
  assign n17841 = n5242 & n17840 ;
  assign n17842 = n1753 | n6030 ;
  assign n17843 = n17842 ^ n3823 ^ 1'b0 ;
  assign n17844 = ( n7882 & n11212 ) | ( n7882 & ~n17843 ) | ( n11212 & ~n17843 ) ;
  assign n17845 = ( n3791 & n17841 ) | ( n3791 & n17844 ) | ( n17841 & n17844 ) ;
  assign n17846 = ( n952 & ~n1896 ) | ( n952 & n8145 ) | ( ~n1896 & n8145 ) ;
  assign n17847 = n12742 ^ n5780 ^ n1140 ;
  assign n17848 = n17847 ^ n9788 ^ n9532 ;
  assign n17849 = ( n3870 & ~n11789 ) | ( n3870 & n13759 ) | ( ~n11789 & n13759 ) ;
  assign n17850 = ( ~n841 & n13114 ) | ( ~n841 & n17849 ) | ( n13114 & n17849 ) ;
  assign n17851 = n10598 ^ n9507 ^ n8937 ;
  assign n17852 = ~n2983 & n17851 ;
  assign n17853 = ( n9681 & n11697 ) | ( n9681 & ~n12245 ) | ( n11697 & ~n12245 ) ;
  assign n17854 = n17853 ^ n16767 ^ n8121 ;
  assign n17855 = ( n840 & n17386 ) | ( n840 & n17854 ) | ( n17386 & n17854 ) ;
  assign n17856 = n1323 ^ n1071 ^ 1'b0 ;
  assign n17857 = n17856 ^ n7013 ^ 1'b0 ;
  assign n17858 = ~n13342 & n16774 ;
  assign n17859 = n17858 ^ n12173 ^ 1'b0 ;
  assign n17866 = n12479 ^ n5643 ^ 1'b0 ;
  assign n17867 = n8737 | n17866 ;
  assign n17868 = n15880 & ~n17867 ;
  assign n17869 = n8884 & n17868 ;
  assign n17863 = n5253 | n7942 ;
  assign n17864 = ( n4105 & n5314 ) | ( n4105 & n17863 ) | ( n5314 & n17863 ) ;
  assign n17865 = x21 & n17864 ;
  assign n17870 = n17869 ^ n17865 ^ n2168 ;
  assign n17860 = n5142 ^ n4626 ^ n3116 ;
  assign n17861 = ~n3469 & n17860 ;
  assign n17862 = ( n771 & n17348 ) | ( n771 & n17861 ) | ( n17348 & n17861 ) ;
  assign n17871 = n17870 ^ n17862 ^ n15706 ;
  assign n17872 = n7504 ^ n1954 ^ 1'b0 ;
  assign n17873 = n13053 & n17872 ;
  assign n17874 = ( n852 & n1321 ) | ( n852 & n12838 ) | ( n1321 & n12838 ) ;
  assign n17878 = n10984 ^ n3753 ^ n926 ;
  assign n17879 = ( n8154 & n13293 ) | ( n8154 & ~n17878 ) | ( n13293 & ~n17878 ) ;
  assign n17875 = n2870 ^ n417 ^ 1'b0 ;
  assign n17876 = ( n8412 & n12142 ) | ( n8412 & n17875 ) | ( n12142 & n17875 ) ;
  assign n17877 = n17876 ^ n14588 ^ n443 ;
  assign n17880 = n17879 ^ n17877 ^ n8293 ;
  assign n17881 = ( n3429 & ~n17874 ) | ( n3429 & n17880 ) | ( ~n17874 & n17880 ) ;
  assign n17882 = ( n4257 & ~n17873 ) | ( n4257 & n17881 ) | ( ~n17873 & n17881 ) ;
  assign n17883 = n1690 ^ n893 ^ x248 ;
  assign n17886 = ( n528 & n4546 ) | ( n528 & n6190 ) | ( n4546 & n6190 ) ;
  assign n17884 = n9892 ^ n5778 ^ n5702 ;
  assign n17885 = n9339 | n17884 ;
  assign n17887 = n17886 ^ n17885 ^ n9421 ;
  assign n17888 = ( ~x183 & n17883 ) | ( ~x183 & n17887 ) | ( n17883 & n17887 ) ;
  assign n17898 = ( ~n887 & n5872 ) | ( ~n887 & n14214 ) | ( n5872 & n14214 ) ;
  assign n17895 = ( n3120 & n6950 ) | ( n3120 & n7346 ) | ( n6950 & n7346 ) ;
  assign n17896 = n9013 ^ n5811 ^ 1'b0 ;
  assign n17897 = ( n11785 & n17895 ) | ( n11785 & n17896 ) | ( n17895 & n17896 ) ;
  assign n17889 = ( n2876 & n3267 ) | ( n2876 & n11134 ) | ( n3267 & n11134 ) ;
  assign n17890 = ( n1175 & n9699 ) | ( n1175 & n17889 ) | ( n9699 & n17889 ) ;
  assign n17891 = ( n3073 & n8256 ) | ( n3073 & ~n17890 ) | ( n8256 & ~n17890 ) ;
  assign n17892 = n6865 ^ n2711 ^ 1'b0 ;
  assign n17893 = n17891 | n17892 ;
  assign n17894 = n17893 ^ n11225 ^ 1'b0 ;
  assign n17899 = n17898 ^ n17897 ^ n17894 ;
  assign n17901 = n13670 & n15519 ;
  assign n17900 = ( n2628 & n4458 ) | ( n2628 & ~n5728 ) | ( n4458 & ~n5728 ) ;
  assign n17902 = n17901 ^ n17900 ^ n11381 ;
  assign n17903 = n12389 ^ n1042 ^ 1'b0 ;
  assign n17911 = n15924 ^ n3872 ^ 1'b0 ;
  assign n17912 = ~n11195 & n17911 ;
  assign n17904 = n16286 ^ n9940 ^ n7872 ;
  assign n17906 = n2399 ^ n558 ^ 1'b0 ;
  assign n17907 = n4569 & ~n17906 ;
  assign n17905 = ( ~n2091 & n5409 ) | ( ~n2091 & n17576 ) | ( n5409 & n17576 ) ;
  assign n17908 = n17907 ^ n17905 ^ n4877 ;
  assign n17909 = ( ~n5590 & n6141 ) | ( ~n5590 & n17908 ) | ( n6141 & n17908 ) ;
  assign n17910 = ~n17904 & n17909 ;
  assign n17913 = n17912 ^ n17910 ^ n8585 ;
  assign n17915 = n9503 & n10895 ;
  assign n17916 = n17915 ^ n2386 ^ 1'b0 ;
  assign n17917 = n17916 ^ n17399 ^ n16587 ;
  assign n17914 = ~n4897 & n8241 ;
  assign n17918 = n17917 ^ n17914 ^ 1'b0 ;
  assign n17919 = ~n2211 & n17918 ;
  assign n17920 = ( n5078 & n17913 ) | ( n5078 & n17919 ) | ( n17913 & n17919 ) ;
  assign n17921 = ( n15433 & ~n17903 ) | ( n15433 & n17920 ) | ( ~n17903 & n17920 ) ;
  assign n17922 = ( n4759 & n7646 ) | ( n4759 & n10660 ) | ( n7646 & n10660 ) ;
  assign n17923 = ( n11417 & ~n14729 ) | ( n11417 & n17922 ) | ( ~n14729 & n17922 ) ;
  assign n17924 = ( x200 & ~n5654 ) | ( x200 & n17264 ) | ( ~n5654 & n17264 ) ;
  assign n17925 = n17221 ^ n1123 ^ 1'b0 ;
  assign n17926 = n5308 | n17925 ;
  assign n17927 = ( n5999 & n6906 ) | ( n5999 & ~n17926 ) | ( n6906 & ~n17926 ) ;
  assign n17928 = n9227 ^ n468 ^ 1'b0 ;
  assign n17929 = n8296 & n17928 ;
  assign n17930 = n17929 ^ n11980 ^ n5735 ;
  assign n17933 = n5215 ^ n1629 ^ 1'b0 ;
  assign n17934 = n12996 & ~n17933 ;
  assign n17931 = n16578 ^ n2791 ^ n2131 ;
  assign n17932 = n17931 ^ n12862 ^ n9630 ;
  assign n17935 = n17934 ^ n17932 ^ n6126 ;
  assign n17936 = ( n7557 & n17930 ) | ( n7557 & n17935 ) | ( n17930 & n17935 ) ;
  assign n17937 = ( ~n1162 & n17927 ) | ( ~n1162 & n17936 ) | ( n17927 & n17936 ) ;
  assign n17938 = n6436 ^ n4209 ^ 1'b0 ;
  assign n17939 = n15493 & n17938 ;
  assign n17940 = ~n15306 & n17939 ;
  assign n17941 = n13823 ^ n7332 ^ 1'b0 ;
  assign n17942 = n1959 | n17941 ;
  assign n17948 = n1908 ^ n1777 ^ n1303 ;
  assign n17943 = ( n525 & ~n1443 ) | ( n525 & n7209 ) | ( ~n1443 & n7209 ) ;
  assign n17944 = n10439 ^ n4637 ^ n1310 ;
  assign n17945 = ( ~n13620 & n17943 ) | ( ~n13620 & n17944 ) | ( n17943 & n17944 ) ;
  assign n17946 = n17945 ^ n6935 ^ n3359 ;
  assign n17947 = n17946 ^ n10361 ^ n4718 ;
  assign n17949 = n17948 ^ n17947 ^ n8606 ;
  assign n17950 = n17949 ^ n16607 ^ n6696 ;
  assign n17951 = n16342 ^ n14613 ^ n11912 ;
  assign n17952 = n17951 ^ n3060 ^ n1746 ;
  assign n17953 = n2996 ^ n2768 ^ 1'b0 ;
  assign n17954 = ( ~n3993 & n5813 ) | ( ~n3993 & n15393 ) | ( n5813 & n15393 ) ;
  assign n17955 = ( n16457 & n17114 ) | ( n16457 & n17954 ) | ( n17114 & n17954 ) ;
  assign n17956 = n2780 ^ n1087 ^ n844 ;
  assign n17957 = ( n1927 & n3470 ) | ( n1927 & ~n10875 ) | ( n3470 & ~n10875 ) ;
  assign n17958 = n17957 ^ n7055 ^ n5894 ;
  assign n17959 = n971 & ~n17958 ;
  assign n17960 = ~n17956 & n17959 ;
  assign n17961 = n812 | n17960 ;
  assign n17962 = n17955 | n17961 ;
  assign n17963 = n4919 ^ n1253 ^ 1'b0 ;
  assign n17964 = n3744 & ~n6591 ;
  assign n17965 = ~n3707 & n17964 ;
  assign n17966 = n6441 ^ n5828 ^ n682 ;
  assign n17967 = ( n5852 & ~n14761 ) | ( n5852 & n17966 ) | ( ~n14761 & n17966 ) ;
  assign n17968 = n8267 & n17967 ;
  assign n17969 = n17968 ^ n8782 ^ 1'b0 ;
  assign n17970 = ( n17963 & n17965 ) | ( n17963 & n17969 ) | ( n17965 & n17969 ) ;
  assign n17971 = ( n3031 & ~n17740 ) | ( n3031 & n17970 ) | ( ~n17740 & n17970 ) ;
  assign n17972 = n13735 ^ x212 ^ 1'b0 ;
  assign n17973 = n2838 & n17972 ;
  assign n17975 = ( ~n1877 & n6330 ) | ( ~n1877 & n15152 ) | ( n6330 & n15152 ) ;
  assign n17974 = ( n831 & n1471 ) | ( n831 & n2877 ) | ( n1471 & n2877 ) ;
  assign n17976 = n17975 ^ n17974 ^ n7371 ;
  assign n17977 = ( n8822 & n17973 ) | ( n8822 & ~n17976 ) | ( n17973 & ~n17976 ) ;
  assign n17983 = n4714 ^ n3604 ^ 1'b0 ;
  assign n17984 = ~n15642 & n17983 ;
  assign n17985 = ~n4453 & n12588 ;
  assign n17986 = ( n6376 & n13559 ) | ( n6376 & ~n17985 ) | ( n13559 & ~n17985 ) ;
  assign n17987 = n17984 & n17986 ;
  assign n17988 = ( n6901 & n8427 ) | ( n6901 & ~n17987 ) | ( n8427 & ~n17987 ) ;
  assign n17982 = n1816 & n4749 ;
  assign n17989 = n17988 ^ n17982 ^ 1'b0 ;
  assign n17981 = n7185 & ~n9608 ;
  assign n17990 = n17989 ^ n17981 ^ 1'b0 ;
  assign n17978 = n1558 ^ x241 ^ 1'b0 ;
  assign n17979 = n10047 & ~n17978 ;
  assign n17980 = ( n2408 & ~n3525 ) | ( n2408 & n17979 ) | ( ~n3525 & n17979 ) ;
  assign n17991 = n17990 ^ n17980 ^ n6789 ;
  assign n17992 = n6240 ^ n1321 ^ n600 ;
  assign n17993 = n17992 ^ n9276 ^ n3027 ;
  assign n17994 = n4362 | n17993 ;
  assign n17995 = n14046 | n17994 ;
  assign n17996 = ( n12668 & ~n17991 ) | ( n12668 & n17995 ) | ( ~n17991 & n17995 ) ;
  assign n17997 = n10699 ^ n860 ^ 1'b0 ;
  assign n17998 = n17428 & n17997 ;
  assign n18001 = ( n3042 & n6923 ) | ( n3042 & n13471 ) | ( n6923 & n13471 ) ;
  assign n18000 = ( n1522 & n2243 ) | ( n1522 & ~n12221 ) | ( n2243 & ~n12221 ) ;
  assign n17999 = ( x190 & n12018 ) | ( x190 & n16079 ) | ( n12018 & n16079 ) ;
  assign n18002 = n18001 ^ n18000 ^ n17999 ;
  assign n18003 = n1908 & n11801 ;
  assign n18004 = n18003 ^ n13108 ^ 1'b0 ;
  assign n18005 = ( n6782 & ~n11828 ) | ( n6782 & n13877 ) | ( ~n11828 & n13877 ) ;
  assign n18006 = n18005 ^ n17117 ^ n16758 ;
  assign n18007 = n18006 ^ n4224 ^ 1'b0 ;
  assign n18008 = n16572 & n18007 ;
  assign n18009 = ( n15232 & n18004 ) | ( n15232 & n18008 ) | ( n18004 & n18008 ) ;
  assign n18014 = n2494 | n9964 ;
  assign n18015 = n16425 | n18014 ;
  assign n18010 = n4877 ^ n766 ^ 1'b0 ;
  assign n18011 = ( n8095 & n8536 ) | ( n8095 & n18010 ) | ( n8536 & n18010 ) ;
  assign n18012 = ( n763 & ~n7880 ) | ( n763 & n18011 ) | ( ~n7880 & n18011 ) ;
  assign n18013 = n18012 ^ n13529 ^ n7693 ;
  assign n18016 = n18015 ^ n18013 ^ n5641 ;
  assign n18017 = n16263 ^ n2190 ^ n296 ;
  assign n18018 = n12817 ^ n6718 ^ n4478 ;
  assign n18019 = ( n10335 & ~n12185 ) | ( n10335 & n18018 ) | ( ~n12185 & n18018 ) ;
  assign n18020 = n16842 ^ n11305 ^ 1'b0 ;
  assign n18021 = n3512 | n18020 ;
  assign n18022 = n1641 | n3012 ;
  assign n18023 = n3836 & ~n18022 ;
  assign n18024 = n18023 ^ n10626 ^ n2804 ;
  assign n18025 = n15673 ^ n9185 ^ 1'b0 ;
  assign n18026 = n18025 ^ n8720 ^ n4341 ;
  assign n18027 = n18026 ^ n8034 ^ n998 ;
  assign n18028 = ( ~n16585 & n18024 ) | ( ~n16585 & n18027 ) | ( n18024 & n18027 ) ;
  assign n18029 = ( n1314 & n1608 ) | ( n1314 & n2327 ) | ( n1608 & n2327 ) ;
  assign n18030 = n7828 ^ n6922 ^ 1'b0 ;
  assign n18031 = n10694 | n18030 ;
  assign n18032 = ( n5923 & n18029 ) | ( n5923 & ~n18031 ) | ( n18029 & ~n18031 ) ;
  assign n18033 = ( n3231 & ~n6989 ) | ( n3231 & n9625 ) | ( ~n6989 & n9625 ) ;
  assign n18034 = n18033 ^ n11868 ^ 1'b0 ;
  assign n18035 = n6312 | n18034 ;
  assign n18036 = n14351 ^ n3341 ^ n682 ;
  assign n18037 = n15731 ^ n12853 ^ n11534 ;
  assign n18038 = ( n5179 & ~n6354 ) | ( n5179 & n16622 ) | ( ~n6354 & n16622 ) ;
  assign n18039 = n18038 ^ n13464 ^ x236 ;
  assign n18040 = ( n12470 & n15228 ) | ( n12470 & n18039 ) | ( n15228 & n18039 ) ;
  assign n18041 = ( ~n11429 & n18037 ) | ( ~n11429 & n18040 ) | ( n18037 & n18040 ) ;
  assign n18042 = ( ~n8233 & n18036 ) | ( ~n8233 & n18041 ) | ( n18036 & n18041 ) ;
  assign n18043 = n16867 ^ n5003 ^ 1'b0 ;
  assign n18044 = ( n6772 & n6963 ) | ( n6772 & ~n11405 ) | ( n6963 & ~n11405 ) ;
  assign n18045 = n9911 | n11978 ;
  assign n18046 = n18044 & ~n18045 ;
  assign n18047 = ( n3497 & n17397 ) | ( n3497 & ~n18046 ) | ( n17397 & ~n18046 ) ;
  assign n18048 = n8261 & n12205 ;
  assign n18049 = n5811 | n18048 ;
  assign n18050 = ( x194 & n5382 ) | ( x194 & ~n14840 ) | ( n5382 & ~n14840 ) ;
  assign n18051 = n10932 ^ n7485 ^ x16 ;
  assign n18052 = ( n3236 & ~n13857 ) | ( n3236 & n18051 ) | ( ~n13857 & n18051 ) ;
  assign n18053 = ( n4097 & n8395 ) | ( n4097 & ~n8806 ) | ( n8395 & ~n8806 ) ;
  assign n18054 = n18053 ^ n1143 ^ n301 ;
  assign n18055 = n1450 & n4536 ;
  assign n18056 = n3925 & n4521 ;
  assign n18057 = n18056 ^ n5152 ^ 1'b0 ;
  assign n18058 = x182 & n18057 ;
  assign n18059 = n18058 ^ n12244 ^ 1'b0 ;
  assign n18060 = n18059 ^ n11742 ^ n10232 ;
  assign n18061 = ( n7997 & n18055 ) | ( n7997 & n18060 ) | ( n18055 & n18060 ) ;
  assign n18062 = ( n4372 & ~n6584 ) | ( n4372 & n6679 ) | ( ~n6584 & n6679 ) ;
  assign n18063 = n18062 ^ n15168 ^ n11268 ;
  assign n18064 = ( n1535 & ~n2706 ) | ( n1535 & n4015 ) | ( ~n2706 & n4015 ) ;
  assign n18065 = ( n3679 & n4109 ) | ( n3679 & n5988 ) | ( n4109 & n5988 ) ;
  assign n18066 = ( n7011 & n9713 ) | ( n7011 & n14845 ) | ( n9713 & n14845 ) ;
  assign n18067 = ( n18064 & ~n18065 ) | ( n18064 & n18066 ) | ( ~n18065 & n18066 ) ;
  assign n18068 = ( ~n12233 & n14382 ) | ( ~n12233 & n18067 ) | ( n14382 & n18067 ) ;
  assign n18069 = ~n16453 & n17073 ;
  assign n18071 = n7374 ^ n5807 ^ n4963 ;
  assign n18072 = n18071 ^ n15622 ^ n13344 ;
  assign n18073 = n6351 ^ n4208 ^ n2763 ;
  assign n18074 = n18073 ^ n7748 ^ n637 ;
  assign n18075 = ( n7882 & n18072 ) | ( n7882 & ~n18074 ) | ( n18072 & ~n18074 ) ;
  assign n18076 = ( ~n8796 & n14472 ) | ( ~n8796 & n18075 ) | ( n14472 & n18075 ) ;
  assign n18070 = n11516 & ~n13223 ;
  assign n18077 = n18076 ^ n18070 ^ 1'b0 ;
  assign n18078 = ~n7325 & n8661 ;
  assign n18079 = n18078 ^ n12529 ^ 1'b0 ;
  assign n18080 = n18079 ^ n12898 ^ n12162 ;
  assign n18087 = ( n2228 & ~n5779 ) | ( n2228 & n13235 ) | ( ~n5779 & n13235 ) ;
  assign n18088 = n9550 | n18087 ;
  assign n18081 = n514 & n2741 ;
  assign n18082 = n13339 & n17295 ;
  assign n18083 = n18081 & n18082 ;
  assign n18084 = n18083 ^ n15936 ^ n5330 ;
  assign n18085 = n18084 ^ n1419 ^ 1'b0 ;
  assign n18086 = ~n17371 & n18085 ;
  assign n18089 = n18088 ^ n18086 ^ n16455 ;
  assign n18090 = n2571 | n8695 ;
  assign n18091 = ( n5929 & n10636 ) | ( n5929 & ~n14999 ) | ( n10636 & ~n14999 ) ;
  assign n18092 = n12710 ^ n9756 ^ n1157 ;
  assign n18095 = ( ~n424 & n1544 ) | ( ~n424 & n1710 ) | ( n1544 & n1710 ) ;
  assign n18093 = ( n5196 & n10692 ) | ( n5196 & n12449 ) | ( n10692 & n12449 ) ;
  assign n18094 = n1961 | n18093 ;
  assign n18096 = n18095 ^ n18094 ^ 1'b0 ;
  assign n18097 = n16117 ^ n11919 ^ n1048 ;
  assign n18098 = ~n13304 & n18097 ;
  assign n18099 = ~n18096 & n18098 ;
  assign n18100 = ( n4689 & ~n7395 ) | ( n4689 & n7796 ) | ( ~n7395 & n7796 ) ;
  assign n18101 = n16429 ^ n4227 ^ 1'b0 ;
  assign n18102 = n9354 & n18101 ;
  assign n18103 = n12730 ^ n9209 ^ n6425 ;
  assign n18104 = ( n7387 & n9200 ) | ( n7387 & n18103 ) | ( n9200 & n18103 ) ;
  assign n18105 = ( n6597 & n18102 ) | ( n6597 & n18104 ) | ( n18102 & n18104 ) ;
  assign n18106 = ( n14860 & n18100 ) | ( n14860 & n18105 ) | ( n18100 & n18105 ) ;
  assign n18107 = ( n7402 & ~n8101 ) | ( n7402 & n8494 ) | ( ~n8101 & n8494 ) ;
  assign n18108 = n6212 & n8736 ;
  assign n18109 = n18108 ^ n4127 ^ 1'b0 ;
  assign n18110 = n11143 & n18109 ;
  assign n18111 = n18110 ^ n4678 ^ n912 ;
  assign n18112 = ( ~n4702 & n18107 ) | ( ~n4702 & n18111 ) | ( n18107 & n18111 ) ;
  assign n18114 = n7411 ^ n6492 ^ n2605 ;
  assign n18113 = ( n434 & n3629 ) | ( n434 & n13875 ) | ( n3629 & n13875 ) ;
  assign n18115 = n18114 ^ n18113 ^ n1807 ;
  assign n18123 = ( n2100 & ~n2192 ) | ( n2100 & n6881 ) | ( ~n2192 & n6881 ) ;
  assign n18124 = ( n7925 & n8020 ) | ( n7925 & n18123 ) | ( n8020 & n18123 ) ;
  assign n18116 = n10865 ^ n3176 ^ n464 ;
  assign n18117 = n18116 ^ n8301 ^ n3477 ;
  assign n18118 = n6844 & n12720 ;
  assign n18119 = ~n7492 & n18118 ;
  assign n18120 = ( n2895 & n5843 ) | ( n2895 & n18119 ) | ( n5843 & n18119 ) ;
  assign n18121 = n5834 & ~n18120 ;
  assign n18122 = ~n18117 & n18121 ;
  assign n18125 = n18124 ^ n18122 ^ n823 ;
  assign n18126 = ( n5279 & n13564 ) | ( n5279 & n17422 ) | ( n13564 & n17422 ) ;
  assign n18127 = n16189 ^ n2948 ^ 1'b0 ;
  assign n18128 = n5839 & ~n18127 ;
  assign n18129 = ( n4213 & n10310 ) | ( n4213 & n18128 ) | ( n10310 & n18128 ) ;
  assign n18130 = ( n5380 & ~n8891 ) | ( n5380 & n18129 ) | ( ~n8891 & n18129 ) ;
  assign n18131 = n2757 ^ n882 ^ 1'b0 ;
  assign n18132 = n1279 | n18131 ;
  assign n18133 = n18132 ^ n5237 ^ 1'b0 ;
  assign n18134 = n15949 & n18133 ;
  assign n18135 = n4647 & n15133 ;
  assign n18136 = ( n4192 & n4978 ) | ( n4192 & ~n18135 ) | ( n4978 & ~n18135 ) ;
  assign n18137 = ( n17199 & n18134 ) | ( n17199 & ~n18136 ) | ( n18134 & ~n18136 ) ;
  assign n18138 = n6549 ^ n5134 ^ n3813 ;
  assign n18139 = n18138 ^ n14488 ^ 1'b0 ;
  assign n18140 = n4375 ^ n3652 ^ 1'b0 ;
  assign n18141 = n3176 & n18140 ;
  assign n18145 = n2012 & ~n2920 ;
  assign n18146 = n11887 | n18145 ;
  assign n18147 = n6739 | n18146 ;
  assign n18148 = ( ~n2275 & n7168 ) | ( ~n2275 & n18147 ) | ( n7168 & n18147 ) ;
  assign n18142 = n1699 & ~n3764 ;
  assign n18143 = n8100 & n18142 ;
  assign n18144 = n18143 ^ n12551 ^ n2641 ;
  assign n18149 = n18148 ^ n18144 ^ 1'b0 ;
  assign n18150 = ~n16233 & n16522 ;
  assign n18151 = n18150 ^ n5689 ^ n4616 ;
  assign n18152 = n14727 ^ n10184 ^ n5723 ;
  assign n18153 = ( n5030 & ~n6756 ) | ( n5030 & n18152 ) | ( ~n6756 & n18152 ) ;
  assign n18154 = ( n10119 & ~n12148 ) | ( n10119 & n12629 ) | ( ~n12148 & n12629 ) ;
  assign n18155 = n2812 ^ x26 ^ 1'b0 ;
  assign n18156 = n2856 & ~n15336 ;
  assign n18157 = n8994 & ~n18156 ;
  assign n18158 = n18157 ^ x66 ^ 1'b0 ;
  assign n18159 = ( n16263 & ~n18155 ) | ( n16263 & n18158 ) | ( ~n18155 & n18158 ) ;
  assign n18160 = ( n928 & ~n6287 ) | ( n928 & n7386 ) | ( ~n6287 & n7386 ) ;
  assign n18161 = ( ~n1596 & n7974 ) | ( ~n1596 & n18160 ) | ( n7974 & n18160 ) ;
  assign n18162 = n18161 ^ n3626 ^ n445 ;
  assign n18163 = ( n2863 & n2974 ) | ( n2863 & n7870 ) | ( n2974 & n7870 ) ;
  assign n18164 = n15770 | n18163 ;
  assign n18165 = n18164 ^ n4802 ^ 1'b0 ;
  assign n18166 = ~n14938 & n18165 ;
  assign n18167 = n7389 & n15616 ;
  assign n18168 = ~n7279 & n18167 ;
  assign n18169 = ~n10187 & n13777 ;
  assign n18170 = n18169 ^ n6179 ^ 1'b0 ;
  assign n18177 = n1864 ^ n1087 ^ n725 ;
  assign n18178 = ( ~n10870 & n15060 ) | ( ~n10870 & n18177 ) | ( n15060 & n18177 ) ;
  assign n18176 = x205 & n3936 ;
  assign n18179 = n18178 ^ n18176 ^ 1'b0 ;
  assign n18172 = n7513 ^ n6161 ^ 1'b0 ;
  assign n18173 = n18172 ^ n14444 ^ n3176 ;
  assign n18171 = n15814 ^ n13815 ^ 1'b0 ;
  assign n18174 = n18173 ^ n18171 ^ n5041 ;
  assign n18175 = n18174 ^ n16863 ^ n4938 ;
  assign n18180 = n18179 ^ n18175 ^ n15030 ;
  assign n18181 = n10405 | n18180 ;
  assign n18182 = n9060 & ~n18181 ;
  assign n18183 = n18182 ^ n592 ^ 1'b0 ;
  assign n18184 = ( n1125 & n6328 ) | ( n1125 & n10737 ) | ( n6328 & n10737 ) ;
  assign n18185 = ( ~n2512 & n7082 ) | ( ~n2512 & n18184 ) | ( n7082 & n18184 ) ;
  assign n18186 = ( ~n4503 & n5745 ) | ( ~n4503 & n18185 ) | ( n5745 & n18185 ) ;
  assign n18187 = n15254 ^ n2251 ^ 1'b0 ;
  assign n18188 = n2896 & ~n18187 ;
  assign n18190 = ~n377 & n5339 ;
  assign n18189 = n7298 ^ n4132 ^ n2988 ;
  assign n18191 = n18190 ^ n18189 ^ n6911 ;
  assign n18195 = ( n3377 & n3772 ) | ( n3377 & ~n9475 ) | ( n3772 & ~n9475 ) ;
  assign n18192 = n3936 & ~n6022 ;
  assign n18193 = n12404 & ~n18192 ;
  assign n18194 = ( n9749 & n11631 ) | ( n9749 & n18193 ) | ( n11631 & n18193 ) ;
  assign n18196 = n18195 ^ n18194 ^ 1'b0 ;
  assign n18197 = n17537 ^ n12688 ^ n2217 ;
  assign n18200 = n5952 ^ n3138 ^ n466 ;
  assign n18198 = n15256 ^ n7088 ^ n6654 ;
  assign n18199 = n13413 | n18198 ;
  assign n18201 = n18200 ^ n18199 ^ 1'b0 ;
  assign n18203 = n11180 ^ n4981 ^ n870 ;
  assign n18202 = n5962 | n10499 ;
  assign n18204 = n18203 ^ n18202 ^ 1'b0 ;
  assign n18205 = n17881 & ~n18204 ;
  assign n18206 = n18205 ^ n8618 ^ 1'b0 ;
  assign n18207 = n13563 ^ n9550 ^ n7936 ;
  assign n18208 = ( n583 & ~n5660 ) | ( n583 & n6854 ) | ( ~n5660 & n6854 ) ;
  assign n18209 = n18208 ^ n9018 ^ n6555 ;
  assign n18210 = ( n4662 & ~n18207 ) | ( n4662 & n18209 ) | ( ~n18207 & n18209 ) ;
  assign n18211 = n15498 ^ n10635 ^ n4554 ;
  assign n18212 = ( ~n1322 & n1914 ) | ( ~n1322 & n14510 ) | ( n1914 & n14510 ) ;
  assign n18213 = n14045 | n17781 ;
  assign n18214 = n12490 | n18213 ;
  assign n18215 = n8624 ^ n4403 ^ n4313 ;
  assign n18216 = n18215 ^ n14198 ^ 1'b0 ;
  assign n18217 = n18214 & ~n18216 ;
  assign n18218 = ~n18212 & n18217 ;
  assign n18219 = ~n1574 & n18218 ;
  assign n18220 = n18211 & ~n18219 ;
  assign n18221 = ~n18210 & n18220 ;
  assign n18222 = ~n606 & n17001 ;
  assign n18223 = n18222 ^ x164 ^ 1'b0 ;
  assign n18224 = n18223 ^ n14880 ^ n13031 ;
  assign n18225 = n5288 ^ n3546 ^ x198 ;
  assign n18226 = ( n6765 & n10582 ) | ( n6765 & n18225 ) | ( n10582 & n18225 ) ;
  assign n18227 = n4412 | n18226 ;
  assign n18228 = ( n3671 & ~n8902 ) | ( n3671 & n11197 ) | ( ~n8902 & n11197 ) ;
  assign n18229 = n18228 ^ n17986 ^ n13079 ;
  assign n18230 = ( n4988 & n11416 ) | ( n4988 & n16976 ) | ( n11416 & n16976 ) ;
  assign n18231 = n13442 | n18230 ;
  assign n18232 = n7803 ^ n1851 ^ 1'b0 ;
  assign n18233 = ( n7013 & n8254 ) | ( n7013 & n11375 ) | ( n8254 & n11375 ) ;
  assign n18234 = n16874 & ~n18233 ;
  assign n18235 = n18234 ^ n13869 ^ 1'b0 ;
  assign n18236 = n5517 ^ n2762 ^ 1'b0 ;
  assign n18237 = ( n556 & n6063 ) | ( n556 & n12384 ) | ( n6063 & n12384 ) ;
  assign n18238 = n18237 ^ n10543 ^ 1'b0 ;
  assign n18239 = ~n18236 & n18238 ;
  assign n18240 = n18239 ^ n10792 ^ n7514 ;
  assign n18241 = n9510 ^ n4849 ^ n3147 ;
  assign n18242 = n16866 & ~n18241 ;
  assign n18243 = n5308 & n18242 ;
  assign n18244 = ( n1057 & n6038 ) | ( n1057 & ~n9357 ) | ( n6038 & ~n9357 ) ;
  assign n18245 = ( n10656 & n13856 ) | ( n10656 & n18244 ) | ( n13856 & n18244 ) ;
  assign n18246 = ( n716 & ~n18243 ) | ( n716 & n18245 ) | ( ~n18243 & n18245 ) ;
  assign n18247 = n15898 ^ n13009 ^ n5014 ;
  assign n18248 = n9913 ^ n6787 ^ 1'b0 ;
  assign n18249 = ( ~n2039 & n6231 ) | ( ~n2039 & n18248 ) | ( n6231 & n18248 ) ;
  assign n18251 = n11170 ^ n3106 ^ n952 ;
  assign n18250 = n15547 ^ n14430 ^ n11302 ;
  assign n18252 = n18251 ^ n18250 ^ n9907 ;
  assign n18253 = ( n9794 & n13863 ) | ( n9794 & ~n16895 ) | ( n13863 & ~n16895 ) ;
  assign n18254 = ( n8573 & n9176 ) | ( n8573 & n18253 ) | ( n9176 & n18253 ) ;
  assign n18256 = n2403 ^ n2056 ^ n1572 ;
  assign n18255 = n7796 ^ n2255 ^ 1'b0 ;
  assign n18257 = n18256 ^ n18255 ^ n2627 ;
  assign n18258 = n5453 ^ n5253 ^ n4647 ;
  assign n18259 = ~n7178 & n18258 ;
  assign n18260 = ~n2766 & n18259 ;
  assign n18261 = ( n6354 & n18257 ) | ( n6354 & n18260 ) | ( n18257 & n18260 ) ;
  assign n18263 = n13856 ^ n11645 ^ n334 ;
  assign n18264 = x169 & n18263 ;
  assign n18262 = n3819 ^ n3512 ^ x244 ;
  assign n18265 = n18264 ^ n18262 ^ x152 ;
  assign n18266 = n8960 & ~n18265 ;
  assign n18267 = n18261 & n18266 ;
  assign n18268 = n2672 & n13364 ;
  assign n18269 = n18268 ^ n16163 ^ 1'b0 ;
  assign n18270 = n12150 & ~n12869 ;
  assign n18271 = n18270 ^ n9791 ^ 1'b0 ;
  assign n18272 = n18271 ^ x240 ^ 1'b0 ;
  assign n18273 = n17898 ^ n13703 ^ n7602 ;
  assign n18274 = n3037 ^ n485 ^ x50 ;
  assign n18275 = n8019 ^ n5506 ^ n4876 ;
  assign n18276 = n18275 ^ n1920 ^ n1432 ;
  assign n18277 = ( n1266 & n3565 ) | ( n1266 & ~n18276 ) | ( n3565 & ~n18276 ) ;
  assign n18278 = n18274 | n18277 ;
  assign n18282 = n4901 & n9162 ;
  assign n18279 = n6430 & ~n7236 ;
  assign n18280 = n18279 ^ n463 ^ 1'b0 ;
  assign n18281 = n18280 ^ n17613 ^ n4474 ;
  assign n18283 = n18282 ^ n18281 ^ n9781 ;
  assign n18284 = n13965 ^ n9688 ^ n2187 ;
  assign n18285 = n18284 ^ n9833 ^ n6628 ;
  assign n18286 = ( ~n3634 & n3855 ) | ( ~n3634 & n18285 ) | ( n3855 & n18285 ) ;
  assign n18287 = n10252 & ~n18286 ;
  assign n18288 = n18287 ^ n6999 ^ 1'b0 ;
  assign n18289 = ~n1045 & n18288 ;
  assign n18290 = n18283 & n18289 ;
  assign n18292 = ( n4359 & n5593 ) | ( n4359 & n9958 ) | ( n5593 & n9958 ) ;
  assign n18291 = ( n2278 & ~n5080 ) | ( n2278 & n11929 ) | ( ~n5080 & n11929 ) ;
  assign n18293 = n18292 ^ n18291 ^ 1'b0 ;
  assign n18294 = n18290 | n18293 ;
  assign n18295 = ~n748 & n3979 ;
  assign n18296 = n1197 & n18295 ;
  assign n18297 = n3576 & n8325 ;
  assign n18298 = ~n14290 & n18297 ;
  assign n18299 = n18298 ^ n10286 ^ n8320 ;
  assign n18300 = ( n17121 & ~n18296 ) | ( n17121 & n18299 ) | ( ~n18296 & n18299 ) ;
  assign n18302 = n4405 ^ n2477 ^ n2387 ;
  assign n18303 = ~n788 & n18302 ;
  assign n18304 = ~n1631 & n18303 ;
  assign n18301 = n7873 & n10244 ;
  assign n18305 = n18304 ^ n18301 ^ n9639 ;
  assign n18306 = ( n2400 & ~n10359 ) | ( n2400 & n18305 ) | ( ~n10359 & n18305 ) ;
  assign n18307 = n18306 ^ n3049 ^ 1'b0 ;
  assign n18308 = n12274 ^ n3715 ^ n3093 ;
  assign n18309 = n18308 ^ n6796 ^ n4809 ;
  assign n18319 = ( n1930 & n4158 ) | ( n1930 & n5699 ) | ( n4158 & n5699 ) ;
  assign n18316 = ~n1205 & n1411 ;
  assign n18317 = n18316 ^ n7205 ^ n1308 ;
  assign n18318 = ( n6081 & n9295 ) | ( n6081 & n18317 ) | ( n9295 & n18317 ) ;
  assign n18320 = n18319 ^ n18318 ^ n13833 ;
  assign n18321 = n18320 ^ n10383 ^ 1'b0 ;
  assign n18322 = ~n4812 & n18321 ;
  assign n18312 = n9574 ^ n5880 ^ n4318 ;
  assign n18313 = n4749 & n18312 ;
  assign n18314 = n17893 & n18313 ;
  assign n18310 = n2873 & n4700 ;
  assign n18311 = n18310 ^ n3209 ^ 1'b0 ;
  assign n18315 = n18314 ^ n18311 ^ 1'b0 ;
  assign n18323 = n18322 ^ n18315 ^ n9749 ;
  assign n18334 = ( ~n2213 & n3618 ) | ( ~n2213 & n5150 ) | ( n3618 & n5150 ) ;
  assign n18324 = n9041 ^ n585 ^ 1'b0 ;
  assign n18325 = ( n2285 & ~n5389 ) | ( n2285 & n18324 ) | ( ~n5389 & n18324 ) ;
  assign n18326 = ( n14345 & n16805 ) | ( n14345 & n18325 ) | ( n16805 & n18325 ) ;
  assign n18327 = n16214 ^ n6936 ^ n2750 ;
  assign n18328 = n3023 ^ n1004 ^ x91 ;
  assign n18329 = ( n1259 & n1919 ) | ( n1259 & ~n3129 ) | ( n1919 & ~n3129 ) ;
  assign n18330 = ( ~n1807 & n7679 ) | ( ~n1807 & n18329 ) | ( n7679 & n18329 ) ;
  assign n18331 = ( n3073 & n18328 ) | ( n3073 & ~n18330 ) | ( n18328 & ~n18330 ) ;
  assign n18332 = ( n4420 & ~n18327 ) | ( n4420 & n18331 ) | ( ~n18327 & n18331 ) ;
  assign n18333 = ~n18326 & n18332 ;
  assign n18335 = n18334 ^ n18333 ^ 1'b0 ;
  assign n18336 = n11404 ^ n3315 ^ n2204 ;
  assign n18337 = n4669 & n10579 ;
  assign n18338 = n18337 ^ n18214 ^ 1'b0 ;
  assign n18339 = n9237 & ~n18338 ;
  assign n18340 = n18336 & n18339 ;
  assign n18341 = n18257 ^ n6351 ^ x36 ;
  assign n18342 = n13498 ^ n6990 ^ n1099 ;
  assign n18343 = n4487 | n8173 ;
  assign n18344 = n18342 & ~n18343 ;
  assign n18345 = n18344 ^ n2680 ^ 1'b0 ;
  assign n18346 = n6810 & n18345 ;
  assign n18347 = ( n6007 & n8201 ) | ( n6007 & n8267 ) | ( n8201 & n8267 ) ;
  assign n18348 = n18347 ^ n2374 ^ 1'b0 ;
  assign n18349 = n4212 ^ n1932 ^ n980 ;
  assign n18350 = ~n3526 & n18349 ;
  assign n18351 = ( n6355 & ~n17215 ) | ( n6355 & n18350 ) | ( ~n17215 & n18350 ) ;
  assign n18352 = n5946 ^ n3525 ^ n1483 ;
  assign n18353 = n10207 | n18352 ;
  assign n18354 = ( n1586 & n18351 ) | ( n1586 & n18353 ) | ( n18351 & n18353 ) ;
  assign n18355 = n2237 | n4354 ;
  assign n18356 = n2471 | n18355 ;
  assign n18357 = n18356 ^ n15406 ^ n12213 ;
  assign n18358 = ~n10511 & n18357 ;
  assign n18359 = ~n3431 & n4789 ;
  assign n18360 = n16805 ^ n3197 ^ 1'b0 ;
  assign n18361 = ~n18359 & n18360 ;
  assign n18362 = ( n2136 & n5647 ) | ( n2136 & ~n8605 ) | ( n5647 & ~n8605 ) ;
  assign n18363 = n12862 ^ n5223 ^ n3769 ;
  assign n18364 = ( n2226 & n15176 ) | ( n2226 & n18363 ) | ( n15176 & n18363 ) ;
  assign n18365 = ( n5693 & n11111 ) | ( n5693 & n11547 ) | ( n11111 & n11547 ) ;
  assign n18366 = n5937 & n18365 ;
  assign n18367 = n18364 & n18366 ;
  assign n18368 = n18367 ^ n4745 ^ 1'b0 ;
  assign n18369 = n6059 | n12856 ;
  assign n18370 = n18369 ^ n4317 ^ 1'b0 ;
  assign n18371 = ( ~n3498 & n5620 ) | ( ~n3498 & n16380 ) | ( n5620 & n16380 ) ;
  assign n18372 = n18370 & ~n18371 ;
  assign n18374 = ( n3633 & ~n4101 ) | ( n3633 & n5278 ) | ( ~n4101 & n5278 ) ;
  assign n18375 = ~n9372 & n15507 ;
  assign n18376 = ~n6118 & n18375 ;
  assign n18377 = n18376 ^ n4405 ^ n3707 ;
  assign n18378 = ( ~n11301 & n18374 ) | ( ~n11301 & n18377 ) | ( n18374 & n18377 ) ;
  assign n18373 = ( n2979 & ~n13296 ) | ( n2979 & n15512 ) | ( ~n13296 & n15512 ) ;
  assign n18379 = n18378 ^ n18373 ^ n6184 ;
  assign n18380 = n18379 ^ n2609 ^ 1'b0 ;
  assign n18381 = ( n439 & ~n11679 ) | ( n439 & n14632 ) | ( ~n11679 & n14632 ) ;
  assign n18382 = n13536 | n18381 ;
  assign n18383 = n1985 & n6581 ;
  assign n18384 = n18383 ^ n8783 ^ n4458 ;
  assign n18385 = ( ~n6073 & n6913 ) | ( ~n6073 & n10365 ) | ( n6913 & n10365 ) ;
  assign n18386 = n18385 ^ n10023 ^ 1'b0 ;
  assign n18387 = n10902 & n18386 ;
  assign n18388 = ( n557 & n2500 ) | ( n557 & ~n13322 ) | ( n2500 & ~n13322 ) ;
  assign n18389 = n5926 ^ n1461 ^ n1243 ;
  assign n18390 = ( n3610 & n5838 ) | ( n3610 & n18389 ) | ( n5838 & n18389 ) ;
  assign n18391 = ( n2418 & n8250 ) | ( n2418 & ~n12921 ) | ( n8250 & ~n12921 ) ;
  assign n18392 = n18391 ^ n5467 ^ n1722 ;
  assign n18393 = ( n2247 & ~n18390 ) | ( n2247 & n18392 ) | ( ~n18390 & n18392 ) ;
  assign n18394 = n18025 ^ n1963 ^ n810 ;
  assign n18395 = ( ~n927 & n4525 ) | ( ~n927 & n8178 ) | ( n4525 & n8178 ) ;
  assign n18402 = n10091 | n12002 ;
  assign n18397 = n9021 ^ n2773 ^ n1801 ;
  assign n18398 = ( n7888 & n17449 ) | ( n7888 & n18397 ) | ( n17449 & n18397 ) ;
  assign n18399 = n6940 & ~n11094 ;
  assign n18400 = ~n18398 & n18399 ;
  assign n18396 = n13767 ^ n13543 ^ n3277 ;
  assign n18401 = n18400 ^ n18396 ^ n15339 ;
  assign n18403 = n18402 ^ n18401 ^ n16863 ;
  assign n18404 = ( n18394 & n18395 ) | ( n18394 & n18403 ) | ( n18395 & n18403 ) ;
  assign n18405 = ( ~n18388 & n18393 ) | ( ~n18388 & n18404 ) | ( n18393 & n18404 ) ;
  assign n18406 = n8719 & n16934 ;
  assign n18407 = n17168 & n18406 ;
  assign n18408 = n18407 ^ n13063 ^ 1'b0 ;
  assign n18409 = ( ~n1809 & n5994 ) | ( ~n1809 & n9060 ) | ( n5994 & n9060 ) ;
  assign n18410 = n15082 ^ n5555 ^ n283 ;
  assign n18411 = n18410 ^ n16776 ^ 1'b0 ;
  assign n18412 = n18409 | n18411 ;
  assign n18413 = ( ~n5188 & n14734 ) | ( ~n5188 & n18412 ) | ( n14734 & n18412 ) ;
  assign n18414 = ( n4638 & n9367 ) | ( n4638 & ~n11877 ) | ( n9367 & ~n11877 ) ;
  assign n18415 = n2713 | n4289 ;
  assign n18418 = ( ~n3707 & n4761 ) | ( ~n3707 & n8155 ) | ( n4761 & n8155 ) ;
  assign n18419 = n18418 ^ n17208 ^ n5812 ;
  assign n18416 = n16221 ^ n4325 ^ 1'b0 ;
  assign n18417 = n7701 & ~n18416 ;
  assign n18420 = n18419 ^ n18417 ^ n8025 ;
  assign n18421 = ( n9309 & n18415 ) | ( n9309 & ~n18420 ) | ( n18415 & ~n18420 ) ;
  assign n18422 = ~n6410 & n7433 ;
  assign n18426 = ( n1329 & ~n6508 ) | ( n1329 & n7194 ) | ( ~n6508 & n7194 ) ;
  assign n18423 = n4954 ^ n2400 ^ 1'b0 ;
  assign n18424 = ( n11670 & ~n17138 ) | ( n11670 & n18423 ) | ( ~n17138 & n18423 ) ;
  assign n18425 = n1769 | n18424 ;
  assign n18427 = n18426 ^ n18425 ^ 1'b0 ;
  assign n18428 = n15087 ^ n14330 ^ n7131 ;
  assign n18429 = n9857 ^ n7094 ^ n5493 ;
  assign n18430 = n3582 | n18429 ;
  assign n18431 = n18430 ^ n2533 ^ 1'b0 ;
  assign n18432 = n18431 ^ n6331 ^ n728 ;
  assign n18433 = n14112 ^ n11491 ^ n10692 ;
  assign n18435 = n1474 & n6010 ;
  assign n18436 = n13400 ^ n3063 ^ 1'b0 ;
  assign n18437 = n18435 | n18436 ;
  assign n18438 = n18437 ^ n7872 ^ n1245 ;
  assign n18439 = n18438 ^ n16668 ^ n2539 ;
  assign n18441 = n5843 & ~n14961 ;
  assign n18440 = n5708 ^ n2042 ^ 1'b0 ;
  assign n18442 = n18441 ^ n18440 ^ n15101 ;
  assign n18443 = n18439 & n18442 ;
  assign n18444 = n18443 ^ n6472 ^ 1'b0 ;
  assign n18445 = n17270 | n18444 ;
  assign n18434 = n15334 & ~n15615 ;
  assign n18446 = n18445 ^ n18434 ^ 1'b0 ;
  assign n18447 = ( ~n2494 & n9399 ) | ( ~n2494 & n13692 ) | ( n9399 & n13692 ) ;
  assign n18448 = n18447 ^ n5814 ^ n1575 ;
  assign n18449 = ( n1518 & n6989 ) | ( n1518 & n7548 ) | ( n6989 & n7548 ) ;
  assign n18450 = n18449 ^ n13363 ^ n8909 ;
  assign n18451 = n11046 ^ n4959 ^ n1007 ;
  assign n18452 = ( n3633 & ~n5858 ) | ( n3633 & n18451 ) | ( ~n5858 & n18451 ) ;
  assign n18453 = n15923 ^ n13387 ^ n592 ;
  assign n18454 = ~n13361 & n18453 ;
  assign n18455 = n18454 ^ n4211 ^ 1'b0 ;
  assign n18456 = n18452 & ~n18455 ;
  assign n18459 = n3791 | n12034 ;
  assign n18460 = n16467 | n18459 ;
  assign n18461 = ( ~n949 & n5235 ) | ( ~n949 & n18460 ) | ( n5235 & n18460 ) ;
  assign n18457 = n11188 ^ n4958 ^ n2429 ;
  assign n18458 = n15951 & ~n18457 ;
  assign n18462 = n18461 ^ n18458 ^ 1'b0 ;
  assign n18463 = n6280 | n10982 ;
  assign n18464 = n522 | n18463 ;
  assign n18477 = ( x241 & n1499 ) | ( x241 & ~n6614 ) | ( n1499 & ~n6614 ) ;
  assign n18471 = n7104 ^ n952 ^ x152 ;
  assign n18472 = ( n652 & n9616 ) | ( n652 & ~n16826 ) | ( n9616 & ~n16826 ) ;
  assign n18473 = n13735 & ~n14637 ;
  assign n18474 = ~n18472 & n18473 ;
  assign n18475 = n18471 & n18474 ;
  assign n18468 = n5453 ^ n1999 ^ 1'b0 ;
  assign n18465 = n8980 ^ n2141 ^ 1'b0 ;
  assign n18466 = n3186 & n18465 ;
  assign n18467 = n18466 ^ n11152 ^ n290 ;
  assign n18469 = n18468 ^ n18467 ^ n6227 ;
  assign n18470 = n18469 ^ n15257 ^ n1372 ;
  assign n18476 = n18475 ^ n18470 ^ n9756 ;
  assign n18478 = n18477 ^ n18476 ^ 1'b0 ;
  assign n18479 = n9782 ^ n2855 ^ n2496 ;
  assign n18480 = ( x91 & ~n1774 ) | ( x91 & n7235 ) | ( ~n1774 & n7235 ) ;
  assign n18481 = n18480 ^ n9258 ^ 1'b0 ;
  assign n18485 = ( n1656 & n5873 ) | ( n1656 & ~n8459 ) | ( n5873 & ~n8459 ) ;
  assign n18486 = ( n11227 & n17391 ) | ( n11227 & ~n18485 ) | ( n17391 & ~n18485 ) ;
  assign n18482 = ~n1784 & n11026 ;
  assign n18483 = n18482 ^ n6454 ^ 1'b0 ;
  assign n18484 = n18483 ^ n3456 ^ n2594 ;
  assign n18487 = n18486 ^ n18484 ^ n15756 ;
  assign n18488 = ( ~n278 & n7325 ) | ( ~n278 & n15116 ) | ( n7325 & n15116 ) ;
  assign n18489 = ( n3421 & ~n6868 ) | ( n3421 & n17459 ) | ( ~n6868 & n17459 ) ;
  assign n18490 = n7161 ^ n4754 ^ n1398 ;
  assign n18491 = ( n2686 & n18489 ) | ( n2686 & n18490 ) | ( n18489 & n18490 ) ;
  assign n18492 = ( n282 & n1411 ) | ( n282 & n18491 ) | ( n1411 & n18491 ) ;
  assign n18493 = ( n2091 & n6919 ) | ( n2091 & n10219 ) | ( n6919 & n10219 ) ;
  assign n18497 = ( n2459 & n2586 ) | ( n2459 & n3290 ) | ( n2586 & n3290 ) ;
  assign n18498 = n18497 ^ n2564 ^ n1055 ;
  assign n18499 = n9090 & n18498 ;
  assign n18494 = n1962 ^ x174 ^ 1'b0 ;
  assign n18495 = n18494 ^ n6688 ^ n5717 ;
  assign n18496 = ( n1730 & n5831 ) | ( n1730 & ~n18495 ) | ( n5831 & ~n18495 ) ;
  assign n18500 = n18499 ^ n18496 ^ 1'b0 ;
  assign n18501 = n18493 | n18500 ;
  assign n18502 = ( ~n7108 & n11508 ) | ( ~n7108 & n17500 ) | ( n11508 & n17500 ) ;
  assign n18503 = n10407 ^ n8471 ^ n5403 ;
  assign n18504 = n18503 ^ n9076 ^ 1'b0 ;
  assign n18505 = ~n4704 & n18504 ;
  assign n18506 = n8471 ^ n6243 ^ 1'b0 ;
  assign n18507 = n18505 & ~n18506 ;
  assign n18508 = ( ~n4701 & n9144 ) | ( ~n4701 & n18507 ) | ( n9144 & n18507 ) ;
  assign n18509 = ( n3345 & ~n4011 ) | ( n3345 & n18508 ) | ( ~n4011 & n18508 ) ;
  assign n18512 = n9551 ^ n649 ^ 1'b0 ;
  assign n18513 = n12737 | n18512 ;
  assign n18510 = n16947 ^ n11375 ^ 1'b0 ;
  assign n18511 = ( n1457 & n4867 ) | ( n1457 & ~n18510 ) | ( n4867 & ~n18510 ) ;
  assign n18514 = n18513 ^ n18511 ^ 1'b0 ;
  assign n18515 = ( ~n7470 & n9375 ) | ( ~n7470 & n18363 ) | ( n9375 & n18363 ) ;
  assign n18516 = ( ~n7595 & n12929 ) | ( ~n7595 & n15195 ) | ( n12929 & n15195 ) ;
  assign n18517 = n18516 ^ n7971 ^ n6031 ;
  assign n18518 = n3940 & ~n18517 ;
  assign n18519 = n18515 & n18518 ;
  assign n18520 = ~n1136 & n5756 ;
  assign n18521 = n18520 ^ n8837 ^ 1'b0 ;
  assign n18528 = ~n4094 & n16562 ;
  assign n18529 = n18528 ^ x172 ^ 1'b0 ;
  assign n18522 = n15812 ^ n12487 ^ 1'b0 ;
  assign n18523 = n14374 | n18522 ;
  assign n18524 = n10829 | n18523 ;
  assign n18525 = ( n5409 & n15609 ) | ( n5409 & ~n18524 ) | ( n15609 & ~n18524 ) ;
  assign n18526 = ~n9307 & n18525 ;
  assign n18527 = n18526 ^ n7819 ^ 1'b0 ;
  assign n18530 = n18529 ^ n18527 ^ n11470 ;
  assign n18531 = n8470 ^ n1528 ^ 1'b0 ;
  assign n18532 = n18530 & n18531 ;
  assign n18533 = n18532 ^ n16244 ^ n10252 ;
  assign n18534 = ( n3625 & n5400 ) | ( n3625 & ~n15608 ) | ( n5400 & ~n15608 ) ;
  assign n18535 = n11502 & n18534 ;
  assign n18536 = n18535 ^ n7289 ^ n5903 ;
  assign n18537 = ~n597 & n7229 ;
  assign n18538 = n3732 & n18537 ;
  assign n18539 = n11858 ^ n1404 ^ 1'b0 ;
  assign n18540 = n11174 & ~n11204 ;
  assign n18541 = ~n1290 & n18540 ;
  assign n18542 = ( n16548 & n18539 ) | ( n16548 & ~n18541 ) | ( n18539 & ~n18541 ) ;
  assign n18546 = n12261 & n18177 ;
  assign n18547 = ~n8259 & n18546 ;
  assign n18543 = n7504 ^ n7425 ^ n3187 ;
  assign n18544 = n18543 ^ n6760 ^ n4772 ;
  assign n18545 = n16258 | n18544 ;
  assign n18548 = n18547 ^ n18545 ^ 1'b0 ;
  assign n18549 = ( n445 & ~n4863 ) | ( n445 & n17855 ) | ( ~n4863 & n17855 ) ;
  assign n18550 = n7505 ^ n997 ^ 1'b0 ;
  assign n18551 = n4668 | n18550 ;
  assign n18552 = n1402 & n18551 ;
  assign n18553 = ( n3264 & n5638 ) | ( n3264 & n18552 ) | ( n5638 & n18552 ) ;
  assign n18554 = n18553 ^ n15167 ^ n4612 ;
  assign n18555 = n14861 ^ n10949 ^ n1275 ;
  assign n18556 = n5689 | n5845 ;
  assign n18557 = n4808 | n18556 ;
  assign n18558 = ( n8903 & n14879 ) | ( n8903 & ~n18557 ) | ( n14879 & ~n18557 ) ;
  assign n18559 = n18558 ^ n3295 ^ 1'b0 ;
  assign n18560 = n18559 ^ n6422 ^ n2362 ;
  assign n18561 = n18560 ^ n13346 ^ n11098 ;
  assign n18562 = n2899 ^ n1536 ^ 1'b0 ;
  assign n18563 = n10861 & n18562 ;
  assign n18564 = ( n2010 & n7646 ) | ( n2010 & n14759 ) | ( n7646 & n14759 ) ;
  assign n18565 = n18564 ^ n16553 ^ 1'b0 ;
  assign n18566 = ( ~n14410 & n18563 ) | ( ~n14410 & n18565 ) | ( n18563 & n18565 ) ;
  assign n18567 = n6773 | n7693 ;
  assign n18568 = n9409 | n18567 ;
  assign n18569 = ( ~n1107 & n1543 ) | ( ~n1107 & n5700 ) | ( n1543 & n5700 ) ;
  assign n18570 = ~n18568 & n18569 ;
  assign n18571 = n12300 ^ n12188 ^ n778 ;
  assign n18572 = n6864 & n7594 ;
  assign n18573 = n18572 ^ n18439 ^ n10897 ;
  assign n18574 = ( n4340 & ~n13960 ) | ( n4340 & n17283 ) | ( ~n13960 & n17283 ) ;
  assign n18575 = ( ~n5323 & n7634 ) | ( ~n5323 & n18574 ) | ( n7634 & n18574 ) ;
  assign n18576 = n18575 ^ n1846 ^ 1'b0 ;
  assign n18577 = ~n15278 & n18576 ;
  assign n18578 = ~n16758 & n18577 ;
  assign n18579 = ( n1303 & ~n1378 ) | ( n1303 & n8850 ) | ( ~n1378 & n8850 ) ;
  assign n18580 = n5755 ^ n3807 ^ n2396 ;
  assign n18581 = n18580 ^ n17086 ^ 1'b0 ;
  assign n18582 = n14680 ^ n5461 ^ n4563 ;
  assign n18583 = n18582 ^ n6396 ^ n5346 ;
  assign n18584 = n18583 ^ n5107 ^ n1455 ;
  assign n18585 = n8517 & ~n10004 ;
  assign n18586 = ( n1739 & n6199 ) | ( n1739 & n18585 ) | ( n6199 & n18585 ) ;
  assign n18587 = n4795 | n18586 ;
  assign n18588 = n4075 & ~n18587 ;
  assign n18589 = ( n6002 & n9501 ) | ( n6002 & n18588 ) | ( n9501 & n18588 ) ;
  assign n18590 = n5168 & n17009 ;
  assign n18591 = n18589 | n18590 ;
  assign n18592 = n2531 ^ n2193 ^ n1142 ;
  assign n18593 = ( n2672 & ~n17221 ) | ( n2672 & n18592 ) | ( ~n17221 & n18592 ) ;
  assign n18594 = n5028 | n18593 ;
  assign n18595 = n18594 ^ n10955 ^ n10441 ;
  assign n18596 = n10269 ^ n9155 ^ n611 ;
  assign n18597 = ~n18595 & n18596 ;
  assign n18601 = n9720 | n13439 ;
  assign n18602 = n8747 | n18601 ;
  assign n18598 = ( n5456 & n6745 ) | ( n5456 & ~n6868 ) | ( n6745 & ~n6868 ) ;
  assign n18599 = n18598 ^ n13372 ^ n12257 ;
  assign n18600 = n5833 & ~n18599 ;
  assign n18603 = n18602 ^ n18600 ^ 1'b0 ;
  assign n18604 = n16321 ^ n15898 ^ n9844 ;
  assign n18605 = ( ~n1430 & n7658 ) | ( ~n1430 & n18604 ) | ( n7658 & n18604 ) ;
  assign n18606 = n14481 ^ n6752 ^ n2729 ;
  assign n18607 = n3588 & ~n12238 ;
  assign n18608 = ~n6346 & n18607 ;
  assign n18609 = n18608 ^ n3204 ^ 1'b0 ;
  assign n18610 = n18609 ^ n9871 ^ n7860 ;
  assign n18611 = ( n8816 & n13454 ) | ( n8816 & ~n18610 ) | ( n13454 & ~n18610 ) ;
  assign n18612 = n983 | n18611 ;
  assign n18613 = n7225 | n18612 ;
  assign n18614 = n2983 ^ n2626 ^ 1'b0 ;
  assign n18615 = n2989 & ~n7211 ;
  assign n18616 = n18615 ^ n1308 ^ 1'b0 ;
  assign n18617 = ~n3352 & n3739 ;
  assign n18618 = n1097 & n18617 ;
  assign n18619 = ( n346 & n18616 ) | ( n346 & n18618 ) | ( n18616 & n18618 ) ;
  assign n18620 = n18619 ^ n18616 ^ 1'b0 ;
  assign n18621 = ~n2562 & n9509 ;
  assign n18622 = ( n3004 & n3942 ) | ( n3004 & ~n18621 ) | ( n3942 & ~n18621 ) ;
  assign n18623 = n14141 ^ n11417 ^ n6027 ;
  assign n18624 = n5071 ^ n2998 ^ n2782 ;
  assign n18625 = n6448 ^ n5910 ^ n894 ;
  assign n18626 = ( n14720 & n18624 ) | ( n14720 & ~n18625 ) | ( n18624 & ~n18625 ) ;
  assign n18627 = n7542 ^ n661 ^ 1'b0 ;
  assign n18628 = n18627 ^ n4403 ^ n1207 ;
  assign n18629 = n362 & n13563 ;
  assign n18630 = n3640 & n18629 ;
  assign n18631 = ( n10796 & n10904 ) | ( n10796 & ~n12186 ) | ( n10904 & ~n12186 ) ;
  assign n18632 = n5171 & n18631 ;
  assign n18633 = n18632 ^ n5595 ^ 1'b0 ;
  assign n18634 = ( x9 & n5161 ) | ( x9 & n15051 ) | ( n5161 & n15051 ) ;
  assign n18635 = ( n14949 & ~n15540 ) | ( n14949 & n18634 ) | ( ~n15540 & n18634 ) ;
  assign n18636 = n6540 | n16689 ;
  assign n18637 = n18636 ^ n4970 ^ 1'b0 ;
  assign n18638 = ( n2082 & n7159 ) | ( n2082 & n18637 ) | ( n7159 & n18637 ) ;
  assign n18639 = ( n10298 & ~n16699 ) | ( n10298 & n18638 ) | ( ~n16699 & n18638 ) ;
  assign n18640 = ( n12600 & n18635 ) | ( n12600 & n18639 ) | ( n18635 & n18639 ) ;
  assign n18641 = ( n740 & n4868 ) | ( n740 & n11682 ) | ( n4868 & n11682 ) ;
  assign n18642 = n18641 ^ n16425 ^ n3056 ;
  assign n18643 = n15634 ^ n7815 ^ 1'b0 ;
  assign n18644 = n18643 ^ n11589 ^ n810 ;
  assign n18645 = n18644 ^ n11532 ^ n4987 ;
  assign n18646 = n9569 ^ n5106 ^ n2440 ;
  assign n18647 = n1923 | n18646 ;
  assign n18648 = ( n3106 & n5918 ) | ( n3106 & n10200 ) | ( n5918 & n10200 ) ;
  assign n18649 = n4110 & ~n10012 ;
  assign n18650 = n15979 & n18649 ;
  assign n18651 = n7292 | n9653 ;
  assign n18652 = n18651 ^ n6930 ^ 1'b0 ;
  assign n18653 = ( ~n18648 & n18650 ) | ( ~n18648 & n18652 ) | ( n18650 & n18652 ) ;
  assign n18654 = ( n2814 & n6866 ) | ( n2814 & ~n15662 ) | ( n6866 & ~n15662 ) ;
  assign n18655 = n2248 & ~n4574 ;
  assign n18656 = ( ~x244 & n580 ) | ( ~x244 & n18655 ) | ( n580 & n18655 ) ;
  assign n18661 = n6317 ^ n752 ^ n308 ;
  assign n18659 = n12212 ^ n3746 ^ x233 ;
  assign n18657 = n8502 ^ n6323 ^ n391 ;
  assign n18658 = n18657 ^ n9979 ^ n4270 ;
  assign n18660 = n18659 ^ n18658 ^ n3467 ;
  assign n18662 = n18661 ^ n18660 ^ 1'b0 ;
  assign n18663 = ( ~n18654 & n18656 ) | ( ~n18654 & n18662 ) | ( n18656 & n18662 ) ;
  assign n18664 = ~n5238 & n9848 ;
  assign n18665 = ( n5840 & n13369 ) | ( n5840 & n18664 ) | ( n13369 & n18664 ) ;
  assign n18666 = n7229 ^ n6059 ^ 1'b0 ;
  assign n18667 = n13282 | n18666 ;
  assign n18668 = n18667 ^ n13049 ^ n2546 ;
  assign n18669 = n6599 ^ n2935 ^ n330 ;
  assign n18670 = ( n4489 & ~n9549 ) | ( n4489 & n18669 ) | ( ~n9549 & n18669 ) ;
  assign n18671 = n13499 ^ x159 ^ 1'b0 ;
  assign n18672 = ( n1993 & n8750 ) | ( n1993 & ~n18671 ) | ( n8750 & ~n18671 ) ;
  assign n18673 = ( n14926 & ~n17366 ) | ( n14926 & n18672 ) | ( ~n17366 & n18672 ) ;
  assign n18674 = ( x102 & n13045 ) | ( x102 & ~n18673 ) | ( n13045 & ~n18673 ) ;
  assign n18675 = ( n18668 & n18670 ) | ( n18668 & ~n18674 ) | ( n18670 & ~n18674 ) ;
  assign n18676 = ~n12972 & n13528 ;
  assign n18677 = n16292 ^ n13182 ^ 1'b0 ;
  assign n18678 = n4809 | n18677 ;
  assign n18679 = n18678 ^ n8873 ^ n1754 ;
  assign n18680 = ( n1825 & n16793 ) | ( n1825 & n17617 ) | ( n16793 & n17617 ) ;
  assign n18681 = ~n2183 & n18680 ;
  assign n18683 = n1317 & n3375 ;
  assign n18684 = n9636 ^ n2978 ^ 1'b0 ;
  assign n18685 = n18683 & n18684 ;
  assign n18682 = n1406 | n17040 ;
  assign n18686 = n18685 ^ n18682 ^ 1'b0 ;
  assign n18687 = n13152 ^ n6815 ^ n4191 ;
  assign n18689 = n3047 & ~n4304 ;
  assign n18688 = ( n2401 & n7722 ) | ( n2401 & ~n18160 ) | ( n7722 & ~n18160 ) ;
  assign n18690 = n18689 ^ n18688 ^ n9640 ;
  assign n18691 = ~n18055 & n18690 ;
  assign n18693 = n16427 ^ n8665 ^ n6839 ;
  assign n18692 = n17738 ^ n12966 ^ n5000 ;
  assign n18694 = n18693 ^ n18692 ^ n16954 ;
  assign n18696 = n6027 ^ n4732 ^ n4554 ;
  assign n18697 = x71 & ~n18696 ;
  assign n18695 = ( n7523 & n10867 ) | ( n7523 & ~n13569 ) | ( n10867 & ~n13569 ) ;
  assign n18698 = n18697 ^ n18695 ^ n3215 ;
  assign n18699 = n13200 ^ n9853 ^ 1'b0 ;
  assign n18700 = n18699 ^ n11146 ^ 1'b0 ;
  assign n18701 = n18698 & n18700 ;
  assign n18705 = ( n3860 & n5567 ) | ( n3860 & ~n6506 ) | ( n5567 & ~n6506 ) ;
  assign n18706 = n18705 ^ n9311 ^ n2480 ;
  assign n18702 = n2725 & ~n14235 ;
  assign n18703 = n18702 ^ n2907 ^ 1'b0 ;
  assign n18704 = n18703 ^ n14960 ^ n12013 ;
  assign n18707 = n18706 ^ n18704 ^ n8356 ;
  assign n18708 = ( n1143 & n7775 ) | ( n1143 & ~n18707 ) | ( n7775 & ~n18707 ) ;
  assign n18709 = n18708 ^ n10247 ^ 1'b0 ;
  assign n18710 = ~n15961 & n18709 ;
  assign n18711 = n18710 ^ n6603 ^ n3189 ;
  assign n18721 = ~n7570 & n12273 ;
  assign n18716 = n5829 & n8150 ;
  assign n18717 = ( n697 & n3560 ) | ( n697 & n8747 ) | ( n3560 & n8747 ) ;
  assign n18718 = ( n3427 & n18716 ) | ( n3427 & n18717 ) | ( n18716 & n18717 ) ;
  assign n18719 = ( n11299 & n14198 ) | ( n11299 & ~n18718 ) | ( n14198 & ~n18718 ) ;
  assign n18713 = n6218 ^ n4164 ^ n3703 ;
  assign n18712 = n3066 ^ n2537 ^ n1489 ;
  assign n18714 = n18713 ^ n18712 ^ n7591 ;
  assign n18715 = n18714 ^ n3570 ^ 1'b0 ;
  assign n18720 = n18719 ^ n18715 ^ n12367 ;
  assign n18722 = n18721 ^ n18720 ^ n4849 ;
  assign n18723 = n4418 & ~n17000 ;
  assign n18724 = n6972 ^ n2809 ^ 1'b0 ;
  assign n18725 = n4489 ^ n3227 ^ n2297 ;
  assign n18726 = n12286 & n18725 ;
  assign n18727 = n18726 ^ n2594 ^ 1'b0 ;
  assign n18728 = ( ~n7995 & n18724 ) | ( ~n7995 & n18727 ) | ( n18724 & n18727 ) ;
  assign n18729 = n18728 ^ n12536 ^ n1562 ;
  assign n18730 = n12930 ^ n4453 ^ n530 ;
  assign n18731 = n18730 ^ n14693 ^ n2633 ;
  assign n18732 = n18731 ^ n5418 ^ n5165 ;
  assign n18733 = n1351 | n8093 ;
  assign n18734 = n18733 ^ n2519 ^ 1'b0 ;
  assign n18735 = ( ~n1157 & n4876 ) | ( ~n1157 & n14231 ) | ( n4876 & n14231 ) ;
  assign n18736 = ( n1173 & ~n10820 ) | ( n1173 & n18735 ) | ( ~n10820 & n18735 ) ;
  assign n18737 = n18736 ^ n9353 ^ 1'b0 ;
  assign n18738 = n8178 | n15468 ;
  assign n18739 = ( ~n6383 & n7388 ) | ( ~n6383 & n18738 ) | ( n7388 & n18738 ) ;
  assign n18740 = ( n3783 & n12388 ) | ( n3783 & n18739 ) | ( n12388 & n18739 ) ;
  assign n18741 = n18740 ^ n6934 ^ n2848 ;
  assign n18742 = ( ~n6285 & n8251 ) | ( ~n6285 & n18741 ) | ( n8251 & n18741 ) ;
  assign n18743 = n631 & n8019 ;
  assign n18744 = ( n4082 & n5415 ) | ( n4082 & n10184 ) | ( n5415 & n10184 ) ;
  assign n18745 = n10459 ^ n6626 ^ 1'b0 ;
  assign n18746 = n10430 | n18745 ;
  assign n18747 = n18744 & ~n18746 ;
  assign n18748 = n18747 ^ n6464 ^ 1'b0 ;
  assign n18749 = ( n5393 & n18743 ) | ( n5393 & ~n18748 ) | ( n18743 & ~n18748 ) ;
  assign n18750 = ( n4071 & n18742 ) | ( n4071 & n18749 ) | ( n18742 & n18749 ) ;
  assign n18754 = ( ~n2479 & n5389 ) | ( ~n2479 & n16699 ) | ( n5389 & n16699 ) ;
  assign n18751 = ~n1937 & n16588 ;
  assign n18752 = ~n9419 & n18751 ;
  assign n18753 = ( n9297 & ~n18145 ) | ( n9297 & n18752 ) | ( ~n18145 & n18752 ) ;
  assign n18755 = n18754 ^ n18753 ^ n7299 ;
  assign n18756 = n12930 ^ n5805 ^ 1'b0 ;
  assign n18757 = n18756 ^ n8950 ^ n1898 ;
  assign n18758 = n5307 ^ n4130 ^ 1'b0 ;
  assign n18759 = n18758 ^ n14018 ^ n13214 ;
  assign n18760 = n8758 ^ n2525 ^ n264 ;
  assign n18761 = n11199 ^ n3287 ^ n2483 ;
  assign n18762 = ( n9851 & n18760 ) | ( n9851 & n18761 ) | ( n18760 & n18761 ) ;
  assign n18763 = ( n14824 & n18688 ) | ( n14824 & ~n18762 ) | ( n18688 & ~n18762 ) ;
  assign n18764 = ( n3700 & n5205 ) | ( n3700 & ~n11473 ) | ( n5205 & ~n11473 ) ;
  assign n18765 = n18764 ^ n3422 ^ 1'b0 ;
  assign n18766 = n3783 | n4743 ;
  assign n18767 = ~n18765 & n18766 ;
  assign n18768 = n16003 ^ n13664 ^ n2835 ;
  assign n18769 = n18768 ^ n14106 ^ n6971 ;
  assign n18771 = ( n16882 & n17518 ) | ( n16882 & ~n18572 ) | ( n17518 & ~n18572 ) ;
  assign n18772 = n18771 ^ n1927 ^ 1'b0 ;
  assign n18770 = ( n1004 & n8962 ) | ( n1004 & ~n15239 ) | ( n8962 & ~n15239 ) ;
  assign n18773 = n18772 ^ n18770 ^ 1'b0 ;
  assign n18782 = n8183 & n14097 ;
  assign n18775 = n1342 | n5333 ;
  assign n18776 = n11993 | n18775 ;
  assign n18779 = ( ~n3363 & n12525 ) | ( ~n3363 & n15106 ) | ( n12525 & n15106 ) ;
  assign n18777 = n12254 ^ n2617 ^ n2541 ;
  assign n18778 = n9292 & n18777 ;
  assign n18780 = n18779 ^ n18778 ^ 1'b0 ;
  assign n18781 = n18776 & ~n18780 ;
  assign n18774 = ( ~n3703 & n4353 ) | ( ~n3703 & n4936 ) | ( n4353 & n4936 ) ;
  assign n18783 = n18782 ^ n18781 ^ n18774 ;
  assign n18784 = ( ~x140 & n3255 ) | ( ~x140 & n18064 ) | ( n3255 & n18064 ) ;
  assign n18785 = n4741 & ~n18784 ;
  assign n18786 = ( n3015 & n3873 ) | ( n3015 & n18785 ) | ( n3873 & n18785 ) ;
  assign n18790 = n1800 & ~n12398 ;
  assign n18788 = n17804 ^ n9705 ^ n8050 ;
  assign n18787 = ( n4415 & n8711 ) | ( n4415 & ~n11103 ) | ( n8711 & ~n11103 ) ;
  assign n18789 = n18788 ^ n18787 ^ n1047 ;
  assign n18791 = n18790 ^ n18789 ^ n5268 ;
  assign n18792 = n10879 & n18791 ;
  assign n18793 = ~n15648 & n18792 ;
  assign n18794 = n4128 ^ n3545 ^ n2119 ;
  assign n18795 = n6206 | n18794 ;
  assign n18796 = n18795 ^ n12439 ^ 1'b0 ;
  assign n18797 = ( ~n11487 & n14979 ) | ( ~n11487 & n18373 ) | ( n14979 & n18373 ) ;
  assign n18798 = n4474 & ~n18797 ;
  assign n18799 = ~n18796 & n18798 ;
  assign n18800 = n10908 & ~n11965 ;
  assign n18803 = ( n771 & n4207 ) | ( n771 & n14449 ) | ( n4207 & n14449 ) ;
  assign n18801 = ~n1571 & n7026 ;
  assign n18802 = n18801 ^ n13112 ^ n2932 ;
  assign n18804 = n18803 ^ n18802 ^ n1387 ;
  assign n18805 = n9349 ^ n7020 ^ n4945 ;
  assign n18806 = n10728 ^ n9523 ^ n5576 ;
  assign n18807 = ( n6494 & ~n18805 ) | ( n6494 & n18806 ) | ( ~n18805 & n18806 ) ;
  assign n18808 = n6080 & ~n14078 ;
  assign n18809 = n5074 & n18808 ;
  assign n18810 = n4773 ^ n3247 ^ n1642 ;
  assign n18811 = n16350 ^ n11883 ^ n2936 ;
  assign n18812 = n18811 ^ n4714 ^ n2971 ;
  assign n18813 = n3948 ^ n1936 ^ n1896 ;
  assign n18814 = n18813 ^ n6585 ^ n963 ;
  assign n18815 = ( n9343 & n18812 ) | ( n9343 & n18814 ) | ( n18812 & n18814 ) ;
  assign n18816 = n8315 ^ n427 ^ 1'b0 ;
  assign n18817 = n7294 & n18816 ;
  assign n18818 = n18817 ^ n2828 ^ n1486 ;
  assign n18819 = ~n778 & n18818 ;
  assign n18820 = n1419 & n18819 ;
  assign n18822 = ( ~n366 & n9986 ) | ( ~n366 & n13081 ) | ( n9986 & n13081 ) ;
  assign n18821 = n278 | n7192 ;
  assign n18823 = n18822 ^ n18821 ^ 1'b0 ;
  assign n18824 = n16969 ^ n10541 ^ n5725 ;
  assign n18825 = ( n3507 & ~n5302 ) | ( n3507 & n8806 ) | ( ~n5302 & n8806 ) ;
  assign n18826 = n11070 & n18825 ;
  assign n18827 = n12369 ^ n11750 ^ n9263 ;
  assign n18831 = n1879 ^ x171 ^ x36 ;
  assign n18828 = n15749 ^ n4276 ^ x85 ;
  assign n18829 = n18828 ^ n11650 ^ n10147 ;
  assign n18830 = x220 & ~n18829 ;
  assign n18832 = n18831 ^ n18830 ^ 1'b0 ;
  assign n18833 = n18832 ^ n5010 ^ n3458 ;
  assign n18834 = n12020 ^ n10168 ^ 1'b0 ;
  assign n18835 = n1476 & ~n18834 ;
  assign n18836 = ( ~n4849 & n17522 ) | ( ~n4849 & n18835 ) | ( n17522 & n18835 ) ;
  assign n18837 = n7156 ^ n5871 ^ n5301 ;
  assign n18838 = n18837 ^ n6925 ^ 1'b0 ;
  assign n18839 = ~n18836 & n18838 ;
  assign n18840 = ( n571 & ~n1767 ) | ( n571 & n5278 ) | ( ~n1767 & n5278 ) ;
  assign n18841 = n18840 ^ n15708 ^ n12720 ;
  assign n18842 = ( n4938 & ~n6357 ) | ( n4938 & n7510 ) | ( ~n6357 & n7510 ) ;
  assign n18843 = ( ~n1616 & n2106 ) | ( ~n1616 & n8707 ) | ( n2106 & n8707 ) ;
  assign n18844 = ( ~n7816 & n18842 ) | ( ~n7816 & n18843 ) | ( n18842 & n18843 ) ;
  assign n18845 = n18844 ^ n16912 ^ 1'b0 ;
  assign n18846 = ( ~n5787 & n18841 ) | ( ~n5787 & n18845 ) | ( n18841 & n18845 ) ;
  assign n18850 = ( ~n2610 & n6825 ) | ( ~n2610 & n13457 ) | ( n6825 & n13457 ) ;
  assign n18848 = ( n1802 & ~n4899 ) | ( n1802 & n10319 ) | ( ~n4899 & n10319 ) ;
  assign n18849 = n18848 ^ n18147 ^ n10266 ;
  assign n18847 = ( n4509 & n9244 ) | ( n4509 & ~n15273 ) | ( n9244 & ~n15273 ) ;
  assign n18851 = n18850 ^ n18849 ^ n18847 ;
  assign n18853 = ( ~x193 & n327 ) | ( ~x193 & n5733 ) | ( n327 & n5733 ) ;
  assign n18852 = n8700 ^ n7648 ^ 1'b0 ;
  assign n18854 = n18853 ^ n18852 ^ 1'b0 ;
  assign n18855 = n2344 ^ n2002 ^ 1'b0 ;
  assign n18856 = n7209 & n18855 ;
  assign n18857 = n7050 | n9012 ;
  assign n18858 = ( ~n3120 & n3887 ) | ( ~n3120 & n18857 ) | ( n3887 & n18857 ) ;
  assign n18859 = n18858 ^ n3861 ^ 1'b0 ;
  assign n18860 = ( n17063 & ~n18856 ) | ( n17063 & n18859 ) | ( ~n18856 & n18859 ) ;
  assign n18861 = n18860 ^ n1382 ^ n814 ;
  assign n18862 = n5493 ^ n1849 ^ 1'b0 ;
  assign n18863 = n1999 | n18862 ;
  assign n18864 = ( n5530 & n7691 ) | ( n5530 & n18863 ) | ( n7691 & n18863 ) ;
  assign n18865 = n18864 ^ n6984 ^ n3756 ;
  assign n18866 = n14338 ^ n3242 ^ n2846 ;
  assign n18867 = n18866 ^ n15263 ^ n4452 ;
  assign n18868 = ( n11341 & ~n16352 ) | ( n11341 & n18867 ) | ( ~n16352 & n18867 ) ;
  assign n18869 = ( n13781 & ~n18865 ) | ( n13781 & n18868 ) | ( ~n18865 & n18868 ) ;
  assign n18870 = n10320 ^ n9501 ^ 1'b0 ;
  assign n18871 = ~n17183 & n18870 ;
  assign n18872 = n18871 ^ n17458 ^ 1'b0 ;
  assign n18873 = n18610 ^ n15755 ^ 1'b0 ;
  assign n18874 = ( ~n6014 & n8943 ) | ( ~n6014 & n13400 ) | ( n8943 & n13400 ) ;
  assign n18875 = n18874 ^ n16658 ^ 1'b0 ;
  assign n18876 = n18873 & n18875 ;
  assign n18877 = ~n1155 & n16995 ;
  assign n18878 = n18877 ^ n18145 ^ n4977 ;
  assign n18879 = ( ~n4623 & n13285 ) | ( ~n4623 & n14099 ) | ( n13285 & n14099 ) ;
  assign n18880 = ( n1301 & ~n18878 ) | ( n1301 & n18879 ) | ( ~n18878 & n18879 ) ;
  assign n18881 = ( n948 & ~n9822 ) | ( n948 & n10365 ) | ( ~n9822 & n10365 ) ;
  assign n18882 = n748 | n3631 ;
  assign n18883 = ~n18881 & n18882 ;
  assign n18884 = n18883 ^ n16872 ^ 1'b0 ;
  assign n18885 = n11909 ^ n7124 ^ n2068 ;
  assign n18886 = n11014 ^ n10858 ^ n1028 ;
  assign n18887 = n659 & n18886 ;
  assign n18888 = n17210 & n18887 ;
  assign n18897 = ( n2486 & ~n3464 ) | ( n2486 & n9009 ) | ( ~n3464 & n9009 ) ;
  assign n18898 = ( ~n5767 & n17929 ) | ( ~n5767 & n18897 ) | ( n17929 & n18897 ) ;
  assign n18895 = n10247 | n18113 ;
  assign n18893 = ( ~n806 & n6226 ) | ( ~n806 & n8205 ) | ( n6226 & n8205 ) ;
  assign n18891 = ( ~n4306 & n6063 ) | ( ~n4306 & n12019 ) | ( n6063 & n12019 ) ;
  assign n18892 = n18891 ^ n10908 ^ n10049 ;
  assign n18894 = n18893 ^ n18892 ^ n5777 ;
  assign n18896 = n18895 ^ n18894 ^ n8310 ;
  assign n18889 = n18568 ^ n7070 ^ 1'b0 ;
  assign n18890 = n8622 & n18889 ;
  assign n18899 = n18898 ^ n18896 ^ n18890 ;
  assign n18900 = n868 | n2590 ;
  assign n18901 = n18900 ^ n5328 ^ 1'b0 ;
  assign n18902 = n18901 ^ n14252 ^ n3950 ;
  assign n18903 = n10367 ^ n6601 ^ n465 ;
  assign n18904 = ( ~n11281 & n18902 ) | ( ~n11281 & n18903 ) | ( n18902 & n18903 ) ;
  assign n18905 = ( n3852 & n10115 ) | ( n3852 & ~n13613 ) | ( n10115 & ~n13613 ) ;
  assign n18906 = n3879 ^ n1323 ^ n641 ;
  assign n18907 = ( ~n3705 & n7359 ) | ( ~n3705 & n18906 ) | ( n7359 & n18906 ) ;
  assign n18908 = ~n2881 & n15661 ;
  assign n18909 = ( n18905 & n18907 ) | ( n18905 & n18908 ) | ( n18907 & n18908 ) ;
  assign n18915 = n1954 & n5549 ;
  assign n18910 = ( ~n2375 & n6497 ) | ( ~n2375 & n8438 ) | ( n6497 & n8438 ) ;
  assign n18911 = ( x141 & n14240 ) | ( x141 & ~n18910 ) | ( n14240 & ~n18910 ) ;
  assign n18912 = n18911 ^ n9393 ^ n1680 ;
  assign n18913 = ( n1620 & ~n2478 ) | ( n1620 & n18912 ) | ( ~n2478 & n18912 ) ;
  assign n18914 = n5149 & ~n18913 ;
  assign n18916 = n18915 ^ n18914 ^ 1'b0 ;
  assign n18923 = n4744 ^ n1863 ^ 1'b0 ;
  assign n18924 = n4557 & n18923 ;
  assign n18921 = ( n3433 & ~n5697 ) | ( n3433 & n11146 ) | ( ~n5697 & n11146 ) ;
  assign n18922 = ( n2036 & ~n10762 ) | ( n2036 & n18921 ) | ( ~n10762 & n18921 ) ;
  assign n18917 = ( ~n6639 & n10022 ) | ( ~n6639 & n11381 ) | ( n10022 & n11381 ) ;
  assign n18918 = n7926 | n18917 ;
  assign n18919 = n18918 ^ n18107 ^ 1'b0 ;
  assign n18920 = n14193 & n18919 ;
  assign n18925 = n18924 ^ n18922 ^ n18920 ;
  assign n18926 = n884 | n5377 ;
  assign n18927 = ( ~n10191 & n11413 ) | ( ~n10191 & n15097 ) | ( n11413 & n15097 ) ;
  assign n18928 = ( n3794 & n6888 ) | ( n3794 & n10914 ) | ( n6888 & n10914 ) ;
  assign n18929 = n18928 ^ n7285 ^ n1208 ;
  assign n18933 = n8980 ^ n5793 ^ n3845 ;
  assign n18934 = n17496 & n18933 ;
  assign n18935 = n18934 ^ n11799 ^ 1'b0 ;
  assign n18936 = n18935 ^ n1946 ^ n1125 ;
  assign n18932 = ( n6707 & n7905 ) | ( n6707 & n12805 ) | ( n7905 & n12805 ) ;
  assign n18930 = n8160 ^ n407 ^ 1'b0 ;
  assign n18931 = ( n1963 & n8489 ) | ( n1963 & ~n18930 ) | ( n8489 & ~n18930 ) ;
  assign n18937 = n18936 ^ n18932 ^ n18931 ;
  assign n18938 = n18937 ^ n18046 ^ n6991 ;
  assign n18939 = n16662 ^ n16271 ^ 1'b0 ;
  assign n18940 = ( x142 & n1588 ) | ( x142 & ~n18893 ) | ( n1588 & ~n18893 ) ;
  assign n18941 = ( ~n4267 & n5831 ) | ( ~n4267 & n18940 ) | ( n5831 & n18940 ) ;
  assign n18942 = n10679 | n18941 ;
  assign n18943 = ( n7229 & ~n11870 ) | ( n7229 & n18942 ) | ( ~n11870 & n18942 ) ;
  assign n18944 = n18943 ^ n14161 ^ n8282 ;
  assign n18945 = n10054 ^ n6102 ^ 1'b0 ;
  assign n18946 = n14463 & ~n18945 ;
  assign n18947 = n18946 ^ n6841 ^ n5571 ;
  assign n18948 = x6 & ~n18947 ;
  assign n18949 = n18948 ^ n13781 ^ 1'b0 ;
  assign n18950 = ( n424 & ~n10297 ) | ( n424 & n16685 ) | ( ~n10297 & n16685 ) ;
  assign n18954 = n2644 & ~n4908 ;
  assign n18955 = n18954 ^ n5584 ^ 1'b0 ;
  assign n18951 = n12745 ^ n8430 ^ 1'b0 ;
  assign n18952 = ( n8674 & n16542 ) | ( n8674 & n18951 ) | ( n16542 & n18951 ) ;
  assign n18953 = ( n3142 & ~n11508 ) | ( n3142 & n18952 ) | ( ~n11508 & n18952 ) ;
  assign n18956 = n18955 ^ n18953 ^ 1'b0 ;
  assign n18957 = n2468 ^ x245 ^ 1'b0 ;
  assign n18958 = n18957 ^ n3467 ^ 1'b0 ;
  assign n18959 = ( n15250 & n18483 ) | ( n15250 & n18958 ) | ( n18483 & n18958 ) ;
  assign n18960 = n18959 ^ n15855 ^ 1'b0 ;
  assign n18961 = ( ~n2103 & n3553 ) | ( ~n2103 & n10123 ) | ( n3553 & n10123 ) ;
  assign n18962 = n18961 ^ n15638 ^ n7660 ;
  assign n18963 = x148 & ~n9054 ;
  assign n18964 = ( n3640 & ~n9841 ) | ( n3640 & n18963 ) | ( ~n9841 & n18963 ) ;
  assign n18965 = n6802 & ~n18964 ;
  assign n18966 = ( n7698 & n18962 ) | ( n7698 & n18965 ) | ( n18962 & n18965 ) ;
  assign n18967 = n18966 ^ n16651 ^ n2296 ;
  assign n18968 = ( n4877 & n5189 ) | ( n4877 & n8481 ) | ( n5189 & n8481 ) ;
  assign n18969 = ( n1170 & n1614 ) | ( n1170 & ~n18968 ) | ( n1614 & ~n18968 ) ;
  assign n18970 = n18969 ^ n12168 ^ n6574 ;
  assign n18971 = ~n2129 & n5059 ;
  assign n18972 = n15179 & n18971 ;
  assign n18973 = n4023 ^ n1815 ^ x65 ;
  assign n18974 = n18973 ^ n10268 ^ n2687 ;
  assign n18975 = ( n17087 & n18972 ) | ( n17087 & n18974 ) | ( n18972 & n18974 ) ;
  assign n18976 = n18975 ^ n1281 ^ 1'b0 ;
  assign n18977 = n2799 | n6221 ;
  assign n18978 = n18977 ^ n17339 ^ 1'b0 ;
  assign n18979 = n18978 ^ n2620 ^ 1'b0 ;
  assign n18980 = n5870 | n18979 ;
  assign n18981 = n18896 ^ n17691 ^ 1'b0 ;
  assign n18982 = n13974 ^ n7883 ^ n3215 ;
  assign n18983 = n16621 ^ n10043 ^ n7217 ;
  assign n18984 = ( n12343 & n17333 ) | ( n12343 & n18983 ) | ( n17333 & n18983 ) ;
  assign n18985 = ( n10053 & ~n18982 ) | ( n10053 & n18984 ) | ( ~n18982 & n18984 ) ;
  assign n18986 = ~n1310 & n14010 ;
  assign n18987 = n18986 ^ n9831 ^ 1'b0 ;
  assign n18988 = n18987 ^ n15014 ^ n7300 ;
  assign n18989 = n6733 & n14490 ;
  assign n18990 = n18989 ^ n6699 ^ 1'b0 ;
  assign n18991 = n4984 & n14519 ;
  assign n18992 = n18990 & n18991 ;
  assign n18996 = n7075 ^ n4708 ^ n2157 ;
  assign n18995 = ( n722 & ~n3422 ) | ( n722 & n14307 ) | ( ~n3422 & n14307 ) ;
  assign n18997 = n18996 ^ n18995 ^ n1006 ;
  assign n18993 = n16696 ^ n8197 ^ n7325 ;
  assign n18994 = n5767 & n18993 ;
  assign n18998 = n18997 ^ n18994 ^ 1'b0 ;
  assign n18999 = ~n12332 & n15153 ;
  assign n19000 = n10559 & ~n18999 ;
  assign n19001 = n19000 ^ n6841 ^ n3915 ;
  assign n19002 = ( n436 & n4338 ) | ( n436 & n5237 ) | ( n4338 & n5237 ) ;
  assign n19003 = ( n1965 & ~n14612 ) | ( n1965 & n19002 ) | ( ~n14612 & n19002 ) ;
  assign n19004 = n19003 ^ n11638 ^ 1'b0 ;
  assign n19013 = ( ~n12377 & n16806 ) | ( ~n12377 & n17073 ) | ( n16806 & n17073 ) ;
  assign n19012 = n6801 ^ n5722 ^ n5230 ;
  assign n19005 = n14501 ^ n5990 ^ 1'b0 ;
  assign n19006 = n697 | n19005 ;
  assign n19007 = n10657 ^ n6240 ^ n1656 ;
  assign n19008 = n19007 ^ n11373 ^ n8036 ;
  assign n19009 = ( ~n13439 & n19006 ) | ( ~n13439 & n19008 ) | ( n19006 & n19008 ) ;
  assign n19010 = n13778 & ~n19009 ;
  assign n19011 = n4823 & n19010 ;
  assign n19014 = n19013 ^ n19012 ^ n19011 ;
  assign n19015 = n19014 ^ n7371 ^ n852 ;
  assign n19021 = n3421 | n8708 ;
  assign n19016 = ( n5039 & n8584 ) | ( n5039 & ~n15010 ) | ( n8584 & ~n15010 ) ;
  assign n19017 = ( n1560 & n5246 ) | ( n1560 & ~n19016 ) | ( n5246 & ~n19016 ) ;
  assign n19018 = n13122 ^ n2741 ^ 1'b0 ;
  assign n19019 = n19017 & ~n19018 ;
  assign n19020 = n19019 ^ n9271 ^ n7000 ;
  assign n19022 = n19021 ^ n19020 ^ n7955 ;
  assign n19024 = ( n10177 & n11876 ) | ( n10177 & n13029 ) | ( n11876 & n13029 ) ;
  assign n19023 = n4978 ^ n1793 ^ n1436 ;
  assign n19025 = n19024 ^ n19023 ^ n8419 ;
  assign n19026 = n10130 ^ n9623 ^ n4247 ;
  assign n19027 = ( n4724 & n12172 ) | ( n4724 & ~n19026 ) | ( n12172 & ~n19026 ) ;
  assign n19028 = n11652 ^ n5193 ^ n2841 ;
  assign n19031 = ( n2979 & ~n4109 ) | ( n2979 & n6196 ) | ( ~n4109 & n6196 ) ;
  assign n19029 = ~n7494 & n9497 ;
  assign n19030 = n17679 & ~n19029 ;
  assign n19032 = n19031 ^ n19030 ^ 1'b0 ;
  assign n19033 = n7395 ^ n3685 ^ n623 ;
  assign n19034 = ( ~n1882 & n8197 ) | ( ~n1882 & n18802 ) | ( n8197 & n18802 ) ;
  assign n19036 = ( n5394 & n9880 ) | ( n5394 & ~n12030 ) | ( n9880 & ~n12030 ) ;
  assign n19035 = ( n635 & ~n5390 ) | ( n635 & n12062 ) | ( ~n5390 & n12062 ) ;
  assign n19037 = n19036 ^ n19035 ^ n498 ;
  assign n19038 = n8211 ^ n2362 ^ 1'b0 ;
  assign n19039 = n19037 & ~n19038 ;
  assign n19040 = n768 & ~n6980 ;
  assign n19041 = ~n19039 & n19040 ;
  assign n19042 = ( n19033 & n19034 ) | ( n19033 & n19041 ) | ( n19034 & n19041 ) ;
  assign n19043 = n18426 ^ n15846 ^ n4538 ;
  assign n19044 = n19043 ^ n8447 ^ n7212 ;
  assign n19046 = ( ~n462 & n5198 ) | ( ~n462 & n7316 ) | ( n5198 & n7316 ) ;
  assign n19045 = n18654 ^ n13794 ^ 1'b0 ;
  assign n19047 = n19046 ^ n19045 ^ n15828 ;
  assign n19048 = n19047 ^ n12524 ^ 1'b0 ;
  assign n19049 = n10298 & ~n19048 ;
  assign n19050 = n14491 ^ n7517 ^ n6297 ;
  assign n19051 = n19050 ^ n17814 ^ n4382 ;
  assign n19052 = n6430 & ~n10172 ;
  assign n19053 = n19052 ^ n1826 ^ 1'b0 ;
  assign n19054 = n19053 ^ n17910 ^ 1'b0 ;
  assign n19055 = n3732 & ~n19054 ;
  assign n19057 = ( ~x240 & n2898 ) | ( ~x240 & n4431 ) | ( n2898 & n4431 ) ;
  assign n19056 = ( n3699 & ~n9883 ) | ( n3699 & n13471 ) | ( ~n9883 & n13471 ) ;
  assign n19058 = n19057 ^ n19056 ^ n16509 ;
  assign n19059 = n19058 ^ n7268 ^ n2928 ;
  assign n19060 = ( ~n4141 & n18400 ) | ( ~n4141 & n18446 ) | ( n18400 & n18446 ) ;
  assign n19062 = n8186 ^ n2467 ^ x239 ;
  assign n19061 = n6798 & ~n13083 ;
  assign n19063 = n19062 ^ n19061 ^ n10424 ;
  assign n19064 = n18046 ^ n10490 ^ n8431 ;
  assign n19065 = n12053 & ~n19064 ;
  assign n19066 = n19065 ^ n6399 ^ 1'b0 ;
  assign n19067 = ( n2342 & n6237 ) | ( n2342 & ~n11461 ) | ( n6237 & ~n11461 ) ;
  assign n19068 = n1207 & ~n12523 ;
  assign n19069 = n19068 ^ n13730 ^ 1'b0 ;
  assign n19070 = n19069 ^ n10177 ^ n6951 ;
  assign n19071 = n15810 ^ n8398 ^ 1'b0 ;
  assign n19072 = ( ~n4966 & n7565 ) | ( ~n4966 & n19071 ) | ( n7565 & n19071 ) ;
  assign n19073 = n12850 & n19072 ;
  assign n19074 = n12321 & n19073 ;
  assign n19075 = n12942 ^ n8344 ^ n4641 ;
  assign n19076 = ( n5100 & ~n14062 ) | ( n5100 & n19075 ) | ( ~n14062 & n19075 ) ;
  assign n19077 = ~n3512 & n5445 ;
  assign n19078 = n19077 ^ n12614 ^ n3365 ;
  assign n19079 = ( ~n5967 & n10461 ) | ( ~n5967 & n19078 ) | ( n10461 & n19078 ) ;
  assign n19080 = n2528 & ~n6026 ;
  assign n19081 = n19080 ^ n8487 ^ n5000 ;
  assign n19082 = n17689 & ~n19081 ;
  assign n19083 = n17079 ^ n15406 ^ 1'b0 ;
  assign n19084 = n11370 | n15904 ;
  assign n19085 = n19083 & ~n19084 ;
  assign n19086 = n4812 & ~n19085 ;
  assign n19087 = n8497 ^ n4191 ^ n724 ;
  assign n19088 = n522 | n4431 ;
  assign n19089 = ( n2052 & n19087 ) | ( n2052 & n19088 ) | ( n19087 & n19088 ) ;
  assign n19090 = ( n8438 & n8697 ) | ( n8438 & ~n14420 ) | ( n8697 & ~n14420 ) ;
  assign n19091 = ( n11071 & ~n19089 ) | ( n11071 & n19090 ) | ( ~n19089 & n19090 ) ;
  assign n19092 = n10249 ^ n7893 ^ n7070 ;
  assign n19093 = n10636 ^ n2278 ^ n1408 ;
  assign n19094 = n19093 ^ n3863 ^ 1'b0 ;
  assign n19095 = n3264 & ~n19094 ;
  assign n19096 = n19095 ^ n8294 ^ n7381 ;
  assign n19097 = n5991 ^ n4298 ^ 1'b0 ;
  assign n19098 = n9347 | n19097 ;
  assign n19099 = n6955 & ~n19098 ;
  assign n19100 = n13320 ^ n7308 ^ 1'b0 ;
  assign n19102 = n6070 ^ n5601 ^ n718 ;
  assign n19101 = ( ~n590 & n2974 ) | ( ~n590 & n15747 ) | ( n2974 & n15747 ) ;
  assign n19103 = n19102 ^ n19101 ^ n4359 ;
  assign n19104 = n16211 ^ n6480 ^ n3342 ;
  assign n19105 = n17571 ^ n7313 ^ x99 ;
  assign n19106 = n19105 ^ n17974 ^ n6772 ;
  assign n19111 = n11573 ^ n10100 ^ n2275 ;
  assign n19109 = ( n4972 & n10787 ) | ( n4972 & n10932 ) | ( n10787 & n10932 ) ;
  assign n19110 = n19109 ^ n4553 ^ n831 ;
  assign n19107 = ( x200 & ~n3120 ) | ( x200 & n7235 ) | ( ~n3120 & n7235 ) ;
  assign n19108 = ( n5200 & n15282 ) | ( n5200 & ~n19107 ) | ( n15282 & ~n19107 ) ;
  assign n19112 = n19111 ^ n19110 ^ n19108 ;
  assign n19113 = ( n2565 & n11998 ) | ( n2565 & ~n19112 ) | ( n11998 & ~n19112 ) ;
  assign n19114 = ( n1112 & ~n7884 ) | ( n1112 & n16886 ) | ( ~n7884 & n16886 ) ;
  assign n19115 = n5861 & n6632 ;
  assign n19116 = ( n3265 & n19114 ) | ( n3265 & n19115 ) | ( n19114 & n19115 ) ;
  assign n19117 = n6560 ^ n4732 ^ n4173 ;
  assign n19118 = n4544 ^ n4099 ^ n1034 ;
  assign n19119 = n5831 | n7394 ;
  assign n19120 = n19119 ^ n2967 ^ 1'b0 ;
  assign n19121 = n19120 ^ n16905 ^ n453 ;
  assign n19122 = n12439 ^ n7455 ^ 1'b0 ;
  assign n19123 = n19121 | n19122 ;
  assign n19124 = ( ~n2807 & n10002 ) | ( ~n2807 & n19123 ) | ( n10002 & n19123 ) ;
  assign n19125 = ~n19118 & n19124 ;
  assign n19126 = ~n19117 & n19125 ;
  assign n19127 = n11963 ^ n4745 ^ 1'b0 ;
  assign n19128 = n19127 ^ n16744 ^ n3137 ;
  assign n19129 = n7839 ^ n3018 ^ n2023 ;
  assign n19130 = ~n2937 & n19129 ;
  assign n19131 = n19130 ^ n2291 ^ 1'b0 ;
  assign n19132 = n12151 ^ n2453 ^ 1'b0 ;
  assign n19133 = ~n12403 & n19132 ;
  assign n19134 = n2087 & n14295 ;
  assign n19135 = n19134 ^ n964 ^ 1'b0 ;
  assign n19136 = ( ~n3845 & n10147 ) | ( ~n3845 & n19135 ) | ( n10147 & n19135 ) ;
  assign n19137 = n11424 ^ n6586 ^ n303 ;
  assign n19138 = n4205 & ~n14314 ;
  assign n19139 = n19138 ^ n11372 ^ 1'b0 ;
  assign n19140 = n19139 ^ n14850 ^ 1'b0 ;
  assign n19141 = n673 & n19140 ;
  assign n19142 = n4141 & ~n11532 ;
  assign n19143 = ( n932 & ~n19141 ) | ( n932 & n19142 ) | ( ~n19141 & n19142 ) ;
  assign n19144 = ( n5260 & ~n18478 ) | ( n5260 & n19143 ) | ( ~n18478 & n19143 ) ;
  assign n19145 = n9368 ^ n9320 ^ n8110 ;
  assign n19146 = n10073 ^ n6491 ^ n1641 ;
  assign n19147 = ( n4458 & n8590 ) | ( n4458 & ~n19146 ) | ( n8590 & ~n19146 ) ;
  assign n19148 = n14501 ^ n3444 ^ n1470 ;
  assign n19149 = n6258 ^ n3964 ^ n1597 ;
  assign n19150 = ( n8127 & ~n8436 ) | ( n8127 & n19149 ) | ( ~n8436 & n19149 ) ;
  assign n19151 = n19150 ^ n18065 ^ n9352 ;
  assign n19152 = ( ~n1065 & n11952 ) | ( ~n1065 & n19151 ) | ( n11952 & n19151 ) ;
  assign n19153 = ( n4281 & ~n6566 ) | ( n4281 & n19152 ) | ( ~n6566 & n19152 ) ;
  assign n19154 = ( n18957 & n19148 ) | ( n18957 & n19153 ) | ( n19148 & n19153 ) ;
  assign n19155 = ( n7798 & ~n10397 ) | ( n7798 & n12795 ) | ( ~n10397 & n12795 ) ;
  assign n19156 = n19155 ^ n7799 ^ n2782 ;
  assign n19159 = n14124 ^ n6993 ^ x184 ;
  assign n19158 = n2867 | n18263 ;
  assign n19157 = n12194 ^ n7052 ^ x60 ;
  assign n19160 = n19159 ^ n19158 ^ n19157 ;
  assign n19161 = n19156 & ~n19160 ;
  assign n19162 = n19161 ^ n15995 ^ 1'b0 ;
  assign n19163 = n9317 ^ n9310 ^ n4718 ;
  assign n19168 = ~n5181 & n6870 ;
  assign n19169 = n10558 & n19168 ;
  assign n19170 = ( ~n9691 & n11900 ) | ( ~n9691 & n19169 ) | ( n11900 & n19169 ) ;
  assign n19164 = ( n2909 & n3097 ) | ( n2909 & ~n5108 ) | ( n3097 & ~n5108 ) ;
  assign n19165 = ( n5073 & n6287 ) | ( n5073 & ~n11588 ) | ( n6287 & ~n11588 ) ;
  assign n19166 = n19165 ^ n8225 ^ 1'b0 ;
  assign n19167 = n19164 & n19166 ;
  assign n19171 = n19170 ^ n19167 ^ 1'b0 ;
  assign n19172 = n14494 ^ n2247 ^ 1'b0 ;
  assign n19173 = n19172 ^ n8854 ^ n6680 ;
  assign n19174 = ( n6061 & n7828 ) | ( n6061 & ~n11519 ) | ( n7828 & ~n11519 ) ;
  assign n19182 = ( ~n1691 & n2386 ) | ( ~n1691 & n6024 ) | ( n2386 & n6024 ) ;
  assign n19180 = ( ~n1221 & n2261 ) | ( ~n1221 & n10828 ) | ( n2261 & n10828 ) ;
  assign n19181 = ( n4234 & n9264 ) | ( n4234 & ~n19180 ) | ( n9264 & ~n19180 ) ;
  assign n19183 = n19182 ^ n19181 ^ n12059 ;
  assign n19184 = n19183 ^ n6973 ^ n4741 ;
  assign n19185 = n19184 ^ n1360 ^ 1'b0 ;
  assign n19176 = n6903 | n16767 ;
  assign n19177 = n2315 | n19176 ;
  assign n19175 = ~n2681 & n11564 ;
  assign n19178 = n19177 ^ n19175 ^ 1'b0 ;
  assign n19179 = n11687 & ~n19178 ;
  assign n19186 = n19185 ^ n19179 ^ n14659 ;
  assign n19187 = ( n7594 & n19174 ) | ( n7594 & ~n19186 ) | ( n19174 & ~n19186 ) ;
  assign n19188 = ( ~n12338 & n13006 ) | ( ~n12338 & n13468 ) | ( n13006 & n13468 ) ;
  assign n19189 = n8166 ^ n997 ^ n617 ;
  assign n19190 = ( n16700 & n19188 ) | ( n16700 & ~n19189 ) | ( n19188 & ~n19189 ) ;
  assign n19191 = ( n9737 & n11734 ) | ( n9737 & ~n13186 ) | ( n11734 & ~n13186 ) ;
  assign n19192 = n6137 | n15749 ;
  assign n19193 = n19192 ^ n13213 ^ n10067 ;
  assign n19194 = n19191 & ~n19193 ;
  assign n19195 = ~n1714 & n19194 ;
  assign n19196 = n1339 & ~n19195 ;
  assign n19197 = n19190 & n19196 ;
  assign n19198 = ( n1609 & n2378 ) | ( n1609 & ~n9564 ) | ( n2378 & ~n9564 ) ;
  assign n19199 = n19198 ^ n4710 ^ n667 ;
  assign n19200 = n19199 ^ n18351 ^ 1'b0 ;
  assign n19201 = n15288 ^ n9455 ^ n7370 ;
  assign n19202 = n19200 | n19201 ;
  assign n19207 = n15225 ^ n10809 ^ n278 ;
  assign n19208 = ( n1886 & n14301 ) | ( n1886 & n19207 ) | ( n14301 & n19207 ) ;
  assign n19209 = ~n16451 & n19208 ;
  assign n19203 = n15749 ^ n10339 ^ n960 ;
  assign n19204 = ~n16507 & n19203 ;
  assign n19205 = ~n4775 & n19204 ;
  assign n19206 = n16927 & ~n19205 ;
  assign n19210 = n19209 ^ n19206 ^ 1'b0 ;
  assign n19211 = n8308 ^ n2258 ^ n1908 ;
  assign n19212 = n19211 ^ n16882 ^ n12012 ;
  assign n19213 = ( ~n11067 & n12743 ) | ( ~n11067 & n13329 ) | ( n12743 & n13329 ) ;
  assign n19214 = n7364 ^ n3315 ^ n2555 ;
  assign n19215 = n3108 & n14201 ;
  assign n19216 = n19215 ^ n3467 ^ n2630 ;
  assign n19217 = ( n19213 & n19214 ) | ( n19213 & ~n19216 ) | ( n19214 & ~n19216 ) ;
  assign n19218 = ~n7904 & n17819 ;
  assign n19219 = n19218 ^ n5215 ^ 1'b0 ;
  assign n19220 = ~n1525 & n6020 ;
  assign n19221 = n19220 ^ n10711 ^ 1'b0 ;
  assign n19222 = n19221 ^ n7874 ^ n2842 ;
  assign n19229 = n15390 ^ n3717 ^ 1'b0 ;
  assign n19223 = ~n8565 & n13569 ;
  assign n19224 = n10709 & ~n12343 ;
  assign n19225 = n19223 & n19224 ;
  assign n19226 = n2583 ^ n1847 ^ n733 ;
  assign n19227 = ( n11295 & n15426 ) | ( n11295 & ~n19226 ) | ( n15426 & ~n19226 ) ;
  assign n19228 = ~n19225 & n19227 ;
  assign n19230 = n19229 ^ n19228 ^ 1'b0 ;
  assign n19231 = ( n19219 & n19222 ) | ( n19219 & ~n19230 ) | ( n19222 & ~n19230 ) ;
  assign n19232 = n4517 ^ n3082 ^ n2115 ;
  assign n19233 = n14551 ^ n14088 ^ n6111 ;
  assign n19234 = n19232 & ~n19233 ;
  assign n19235 = n19234 ^ n17448 ^ 1'b0 ;
  assign n19236 = ( n3616 & n9200 ) | ( n3616 & ~n19235 ) | ( n9200 & ~n19235 ) ;
  assign n19237 = n19236 ^ n18061 ^ n16524 ;
  assign n19247 = n12996 ^ n7053 ^ n1462 ;
  assign n19238 = n1707 & ~n2451 ;
  assign n19239 = n19238 ^ n5244 ^ 1'b0 ;
  assign n19243 = n3206 & ~n9911 ;
  assign n19241 = ( n3645 & n8542 ) | ( n3645 & ~n17843 ) | ( n8542 & ~n17843 ) ;
  assign n19240 = n6212 ^ n3037 ^ n2610 ;
  assign n19242 = n19241 ^ n19240 ^ n5551 ;
  assign n19244 = n19243 ^ n19242 ^ n8407 ;
  assign n19245 = ~n19239 & n19244 ;
  assign n19246 = ~x187 & n19245 ;
  assign n19248 = n19247 ^ n19246 ^ n7181 ;
  assign n19249 = ( n1342 & ~n1996 ) | ( n1342 & n4596 ) | ( ~n1996 & n4596 ) ;
  assign n19250 = n19249 ^ n5888 ^ n4466 ;
  assign n19251 = n19250 ^ n11042 ^ n7852 ;
  assign n19252 = n19251 ^ n18397 ^ n1280 ;
  assign n19253 = n2209 & n18001 ;
  assign n19254 = n2903 & n19253 ;
  assign n19257 = n15843 ^ n15169 ^ 1'b0 ;
  assign n19258 = n3847 & ~n19257 ;
  assign n19259 = n19258 ^ n7911 ^ n5900 ;
  assign n19255 = n4866 ^ n2706 ^ n728 ;
  assign n19256 = n19255 ^ n2825 ^ n1645 ;
  assign n19260 = n19259 ^ n19256 ^ n11142 ;
  assign n19266 = ( n10417 & n12372 ) | ( n10417 & ~n17543 ) | ( n12372 & ~n17543 ) ;
  assign n19267 = ( n914 & n1659 ) | ( n914 & ~n6158 ) | ( n1659 & ~n6158 ) ;
  assign n19268 = ( n553 & n3214 ) | ( n553 & ~n19267 ) | ( n3214 & ~n19267 ) ;
  assign n19269 = n6358 & ~n19268 ;
  assign n19270 = n5020 | n9329 ;
  assign n19271 = ( n3791 & n3975 ) | ( n3791 & ~n15570 ) | ( n3975 & ~n15570 ) ;
  assign n19272 = ~n19270 & n19271 ;
  assign n19273 = n19269 & n19272 ;
  assign n19274 = n19273 ^ n9616 ^ n6260 ;
  assign n19275 = ( n4853 & n19266 ) | ( n4853 & ~n19274 ) | ( n19266 & ~n19274 ) ;
  assign n19261 = n1779 ^ n457 ^ 1'b0 ;
  assign n19262 = ~n5698 & n19261 ;
  assign n19263 = ( ~n812 & n11685 ) | ( ~n812 & n19262 ) | ( n11685 & n19262 ) ;
  assign n19264 = n19263 ^ n4903 ^ n3379 ;
  assign n19265 = n16955 & n19264 ;
  assign n19276 = n19275 ^ n19265 ^ n6689 ;
  assign n19277 = n1525 | n19276 ;
  assign n19278 = n4639 | n19277 ;
  assign n19279 = n18468 ^ n13526 ^ n1396 ;
  assign n19280 = n7476 ^ n2332 ^ n1736 ;
  assign n19281 = n19280 ^ n14500 ^ n12050 ;
  assign n19282 = n17974 ^ n3796 ^ 1'b0 ;
  assign n19283 = n19281 & ~n19282 ;
  assign n19284 = n1411 & ~n6441 ;
  assign n19285 = ~n3608 & n19284 ;
  assign n19286 = n10628 ^ n1634 ^ n1012 ;
  assign n19287 = ( n17903 & n19285 ) | ( n17903 & ~n19286 ) | ( n19285 & ~n19286 ) ;
  assign n19288 = n11942 ^ n11150 ^ n6035 ;
  assign n19289 = n9030 ^ n2527 ^ n2146 ;
  assign n19290 = n19289 ^ n13493 ^ n5681 ;
  assign n19291 = n12658 & ~n19290 ;
  assign n19292 = n19288 & n19291 ;
  assign n19293 = n12488 ^ n11966 ^ n5399 ;
  assign n19294 = n2037 & ~n8295 ;
  assign n19295 = n19294 ^ n13450 ^ n12640 ;
  assign n19301 = n18610 ^ n16290 ^ n5149 ;
  assign n19296 = ( n682 & n7190 ) | ( n682 & n11579 ) | ( n7190 & n11579 ) ;
  assign n19297 = ( ~n2979 & n4773 ) | ( ~n2979 & n19296 ) | ( n4773 & n19296 ) ;
  assign n19298 = n19297 ^ n3519 ^ 1'b0 ;
  assign n19299 = n17424 & n19298 ;
  assign n19300 = n19299 ^ n13442 ^ n11801 ;
  assign n19302 = n19301 ^ n19300 ^ n5219 ;
  assign n19303 = ( n4289 & n19295 ) | ( n4289 & n19302 ) | ( n19295 & n19302 ) ;
  assign n19305 = n3725 | n10763 ;
  assign n19306 = n19305 ^ n17348 ^ n7774 ;
  assign n19304 = ~n18852 & n19152 ;
  assign n19307 = n19306 ^ n19304 ^ 1'b0 ;
  assign n19308 = n18593 ^ n11601 ^ n9966 ;
  assign n19309 = ( ~n10189 & n11746 ) | ( ~n10189 & n19308 ) | ( n11746 & n19308 ) ;
  assign n19310 = n9963 ^ n2117 ^ n1068 ;
  assign n19311 = ( n9012 & n12785 ) | ( n9012 & n13237 ) | ( n12785 & n13237 ) ;
  assign n19312 = ( ~n9053 & n19310 ) | ( ~n9053 & n19311 ) | ( n19310 & n19311 ) ;
  assign n19317 = x68 & ~n10014 ;
  assign n19313 = ( n3605 & n4690 ) | ( n3605 & n8295 ) | ( n4690 & n8295 ) ;
  assign n19314 = ( n949 & ~n3205 ) | ( n949 & n14722 ) | ( ~n3205 & n14722 ) ;
  assign n19315 = ( n10086 & n11273 ) | ( n10086 & ~n14018 ) | ( n11273 & ~n14018 ) ;
  assign n19316 = ( n19313 & ~n19314 ) | ( n19313 & n19315 ) | ( ~n19314 & n19315 ) ;
  assign n19318 = n19317 ^ n19316 ^ 1'b0 ;
  assign n19319 = n8896 & n19318 ;
  assign n19320 = n5677 ^ n1478 ^ 1'b0 ;
  assign n19321 = n13317 & ~n19320 ;
  assign n19324 = n1138 & n9899 ;
  assign n19325 = n19324 ^ n11732 ^ 1'b0 ;
  assign n19326 = n9199 & ~n19325 ;
  assign n19322 = ( ~x149 & n1549 ) | ( ~x149 & n5647 ) | ( n1549 & n5647 ) ;
  assign n19323 = n19322 ^ n9831 ^ n6371 ;
  assign n19327 = n19326 ^ n19323 ^ n6673 ;
  assign n19328 = n19327 ^ n16667 ^ 1'b0 ;
  assign n19329 = n19321 & ~n19328 ;
  assign n19330 = ( n3927 & ~n5379 ) | ( n3927 & n6589 ) | ( ~n5379 & n6589 ) ;
  assign n19333 = n7807 ^ n1050 ^ 1'b0 ;
  assign n19331 = n4529 & n15169 ;
  assign n19332 = n19331 ^ n14318 ^ 1'b0 ;
  assign n19334 = n19333 ^ n19332 ^ n9732 ;
  assign n19335 = ( n19314 & ~n19330 ) | ( n19314 & n19334 ) | ( ~n19330 & n19334 ) ;
  assign n19336 = n2157 | n4186 ;
  assign n19337 = ( ~n2623 & n14463 ) | ( ~n2623 & n19336 ) | ( n14463 & n19336 ) ;
  assign n19340 = n11591 ^ n2856 ^ n2035 ;
  assign n19338 = n10158 ^ n395 ^ 1'b0 ;
  assign n19339 = ( n5930 & n7505 ) | ( n5930 & n19338 ) | ( n7505 & n19338 ) ;
  assign n19341 = n19340 ^ n19339 ^ 1'b0 ;
  assign n19342 = n4795 | n19341 ;
  assign n19343 = n19342 ^ n17528 ^ n5211 ;
  assign n19344 = ( ~n14395 & n19337 ) | ( ~n14395 & n19343 ) | ( n19337 & n19343 ) ;
  assign n19345 = n19344 ^ n4378 ^ n3355 ;
  assign n19346 = ( n1159 & n10326 ) | ( n1159 & n18296 ) | ( n10326 & n18296 ) ;
  assign n19347 = ( ~n4638 & n14003 ) | ( ~n4638 & n19346 ) | ( n14003 & n19346 ) ;
  assign n19348 = n2487 | n18510 ;
  assign n19349 = ~n4245 & n19348 ;
  assign n19350 = n19347 & n19349 ;
  assign n19351 = ( n4082 & n5813 ) | ( n4082 & ~n19350 ) | ( n5813 & ~n19350 ) ;
  assign n19352 = n19351 ^ n14160 ^ n7458 ;
  assign n19353 = ( n5154 & ~n5815 ) | ( n5154 & n7167 ) | ( ~n5815 & n7167 ) ;
  assign n19354 = ( ~n4763 & n6862 ) | ( ~n4763 & n19353 ) | ( n6862 & n19353 ) ;
  assign n19355 = n6443 ^ n5185 ^ n3433 ;
  assign n19356 = n1319 | n6123 ;
  assign n19357 = ( n7585 & n19355 ) | ( n7585 & ~n19356 ) | ( n19355 & ~n19356 ) ;
  assign n19358 = n19357 ^ n17378 ^ n8227 ;
  assign n19359 = n9283 ^ n7734 ^ n3202 ;
  assign n19360 = ( n4574 & ~n6154 ) | ( n4574 & n19359 ) | ( ~n6154 & n19359 ) ;
  assign n19361 = n19360 ^ n8309 ^ n1454 ;
  assign n19362 = ( n4825 & n7776 ) | ( n4825 & n7791 ) | ( n7776 & n7791 ) ;
  assign n19363 = n10934 | n19362 ;
  assign n19364 = n3481 & ~n19363 ;
  assign n19367 = x130 & ~n1610 ;
  assign n19368 = ~n9407 & n19367 ;
  assign n19369 = n5917 & n19368 ;
  assign n19365 = n2337 | n12861 ;
  assign n19366 = ~n17867 & n19365 ;
  assign n19370 = n19369 ^ n19366 ^ 1'b0 ;
  assign n19371 = ( n8509 & n11951 ) | ( n8509 & n19370 ) | ( n11951 & n19370 ) ;
  assign n19372 = n8045 ^ n5489 ^ 1'b0 ;
  assign n19373 = n7509 | n19372 ;
  assign n19374 = n19371 & ~n19373 ;
  assign n19375 = n15902 ^ n1846 ^ n1574 ;
  assign n19376 = n19375 ^ n18314 ^ n2134 ;
  assign n19377 = n19376 ^ n10084 ^ n2877 ;
  assign n19378 = n16406 ^ n13624 ^ x2 ;
  assign n19379 = n4798 & n19378 ;
  assign n19380 = ~n887 & n7433 ;
  assign n19381 = n19380 ^ n12397 ^ n1916 ;
  assign n19382 = n19381 ^ n16561 ^ n15243 ;
  assign n19385 = n7006 & ~n13235 ;
  assign n19386 = n10469 & n19385 ;
  assign n19383 = n4599 ^ n1565 ^ x169 ;
  assign n19384 = ( ~n1269 & n5090 ) | ( ~n1269 & n19383 ) | ( n5090 & n19383 ) ;
  assign n19387 = n19386 ^ n19384 ^ 1'b0 ;
  assign n19388 = n19382 | n19387 ;
  assign n19389 = ( ~n10129 & n14458 ) | ( ~n10129 & n19388 ) | ( n14458 & n19388 ) ;
  assign n19390 = ~n2080 & n6772 ;
  assign n19391 = n2941 & ~n13719 ;
  assign n19392 = ( n5341 & n10932 ) | ( n5341 & ~n19391 ) | ( n10932 & ~n19391 ) ;
  assign n19393 = n2424 & n3721 ;
  assign n19394 = n1219 | n7047 ;
  assign n19395 = ( ~n5191 & n19393 ) | ( ~n5191 & n19394 ) | ( n19393 & n19394 ) ;
  assign n19396 = ( n3454 & n19392 ) | ( n3454 & n19395 ) | ( n19392 & n19395 ) ;
  assign n19397 = ( n12809 & n19390 ) | ( n12809 & n19396 ) | ( n19390 & n19396 ) ;
  assign n19412 = n297 & n7019 ;
  assign n19413 = n19412 ^ n18706 ^ n6429 ;
  assign n19401 = n4159 ^ n3471 ^ 1'b0 ;
  assign n19402 = n9415 & n19401 ;
  assign n19403 = ( n8161 & n14546 ) | ( n8161 & ~n19402 ) | ( n14546 & ~n19402 ) ;
  assign n19404 = n6066 ^ n5286 ^ 1'b0 ;
  assign n19405 = ( n1985 & n19317 ) | ( n1985 & ~n19404 ) | ( n19317 & ~n19404 ) ;
  assign n19406 = n19403 & ~n19405 ;
  assign n19407 = n19406 ^ n16098 ^ 1'b0 ;
  assign n19398 = ~n4368 & n13976 ;
  assign n19399 = n19398 ^ n5150 ^ 1'b0 ;
  assign n19400 = n19399 ^ n15609 ^ n2609 ;
  assign n19408 = n19407 ^ n19400 ^ n18357 ;
  assign n19409 = n14022 ^ n6429 ^ n2224 ;
  assign n19410 = ( n10760 & ~n19408 ) | ( n10760 & n19409 ) | ( ~n19408 & n19409 ) ;
  assign n19411 = n3770 & ~n19410 ;
  assign n19414 = n19413 ^ n19411 ^ 1'b0 ;
  assign n19419 = x149 & ~n8635 ;
  assign n19420 = n19419 ^ n12214 ^ 1'b0 ;
  assign n19418 = n13280 ^ n8975 ^ x202 ;
  assign n19415 = n6827 ^ n6459 ^ n2022 ;
  assign n19416 = n8481 | n19415 ;
  assign n19417 = n19416 ^ n12940 ^ 1'b0 ;
  assign n19421 = n19420 ^ n19418 ^ n19417 ;
  assign n19422 = ( ~n2733 & n10558 ) | ( ~n2733 & n13499 ) | ( n10558 & n13499 ) ;
  assign n19423 = n1199 & n4016 ;
  assign n19424 = n1082 & n19423 ;
  assign n19425 = n15638 ^ n14174 ^ 1'b0 ;
  assign n19426 = n19425 ^ n5565 ^ 1'b0 ;
  assign n19427 = ( n16691 & ~n19424 ) | ( n16691 & n19426 ) | ( ~n19424 & n19426 ) ;
  assign n19428 = ( x2 & ~x72 ) | ( x2 & n1149 ) | ( ~x72 & n1149 ) ;
  assign n19429 = n7170 & n19428 ;
  assign n19430 = n6986 ^ n5031 ^ n2049 ;
  assign n19431 = n19430 ^ n13995 ^ n1629 ;
  assign n19432 = n19431 ^ n7839 ^ n4049 ;
  assign n19433 = ( n7178 & n19429 ) | ( n7178 & n19432 ) | ( n19429 & n19432 ) ;
  assign n19434 = ( n2478 & n4371 ) | ( n2478 & ~n4821 ) | ( n4371 & ~n4821 ) ;
  assign n19435 = ( n3998 & ~n7034 ) | ( n3998 & n7090 ) | ( ~n7034 & n7090 ) ;
  assign n19436 = ~n3172 & n9748 ;
  assign n19437 = ( n19434 & ~n19435 ) | ( n19434 & n19436 ) | ( ~n19435 & n19436 ) ;
  assign n19438 = n457 & n551 ;
  assign n19439 = n19438 ^ n16433 ^ n4990 ;
  assign n19440 = n19439 ^ n8039 ^ n5909 ;
  assign n19441 = ( n13119 & ~n18418 ) | ( n13119 & n19251 ) | ( ~n18418 & n19251 ) ;
  assign n19442 = ( n8934 & n13818 ) | ( n8934 & n16696 ) | ( n13818 & n16696 ) ;
  assign n19443 = n19442 ^ n13480 ^ n4294 ;
  assign n19444 = n16020 ^ n1724 ^ 1'b0 ;
  assign n19445 = n2265 & n19444 ;
  assign n19446 = n14349 ^ n5147 ^ x202 ;
  assign n19447 = n19446 ^ n18953 ^ n15215 ;
  assign n19451 = ~n3170 & n6834 ;
  assign n19452 = n4937 & ~n19451 ;
  assign n19448 = ( n5742 & n6394 ) | ( n5742 & ~n8742 ) | ( n6394 & ~n8742 ) ;
  assign n19449 = n11356 ^ n1669 ^ 1'b0 ;
  assign n19450 = ( n3967 & n19448 ) | ( n3967 & ~n19449 ) | ( n19448 & ~n19449 ) ;
  assign n19453 = n19452 ^ n19450 ^ n6532 ;
  assign n19454 = n13544 ^ n12949 ^ n8912 ;
  assign n19455 = n19454 ^ n8688 ^ 1'b0 ;
  assign n19464 = ( n411 & n1552 ) | ( n411 & n12770 ) | ( n1552 & n12770 ) ;
  assign n19462 = ~n5417 & n13175 ;
  assign n19463 = n19462 ^ n4669 ^ n1834 ;
  assign n19465 = n19464 ^ n19463 ^ n9040 ;
  assign n19456 = n16593 ^ n3998 ^ 1'b0 ;
  assign n19457 = n5784 | n19456 ;
  assign n19458 = n12584 ^ n2805 ^ 1'b0 ;
  assign n19459 = n19457 | n19458 ;
  assign n19460 = ( n1405 & ~n9738 ) | ( n1405 & n19459 ) | ( ~n9738 & n19459 ) ;
  assign n19461 = n19460 ^ n11355 ^ n10430 ;
  assign n19466 = n19465 ^ n19461 ^ n12856 ;
  assign n19467 = n19455 & ~n19466 ;
  assign n19468 = n2716 | n10428 ;
  assign n19469 = n19468 ^ n3579 ^ 1'b0 ;
  assign n19470 = ( n792 & ~n12324 ) | ( n792 & n12858 ) | ( ~n12324 & n12858 ) ;
  assign n19471 = n19469 | n19470 ;
  assign n19472 = ( ~n12546 & n12645 ) | ( ~n12546 & n19471 ) | ( n12645 & n19471 ) ;
  assign n19473 = n6797 ^ n3585 ^ 1'b0 ;
  assign n19474 = n18688 | n19473 ;
  assign n19476 = ( n901 & n12758 ) | ( n901 & ~n14466 ) | ( n12758 & ~n14466 ) ;
  assign n19475 = ~n2797 & n4404 ;
  assign n19477 = n19476 ^ n19475 ^ n12525 ;
  assign n19478 = ( n9269 & ~n12515 ) | ( n9269 & n19477 ) | ( ~n12515 & n19477 ) ;
  assign n19479 = n16075 ^ n15622 ^ 1'b0 ;
  assign n19480 = ~n7729 & n19479 ;
  assign n19481 = n18753 ^ n13662 ^ n12185 ;
  assign n19482 = ( n8612 & ~n8848 ) | ( n8612 & n9395 ) | ( ~n8848 & n9395 ) ;
  assign n19488 = n9205 ^ n8177 ^ 1'b0 ;
  assign n19483 = n1773 & ~n5275 ;
  assign n19484 = n19483 ^ n16249 ^ 1'b0 ;
  assign n19485 = x14 & n6866 ;
  assign n19486 = n19485 ^ n11361 ^ 1'b0 ;
  assign n19487 = n19484 & n19486 ;
  assign n19489 = n19488 ^ n19487 ^ 1'b0 ;
  assign n19490 = n15072 ^ n11408 ^ n3264 ;
  assign n19491 = ( n11371 & ~n16184 ) | ( n11371 & n19490 ) | ( ~n16184 & n19490 ) ;
  assign n19492 = n12708 ^ n9930 ^ n6287 ;
  assign n19493 = n19492 ^ n6613 ^ n1611 ;
  assign n19494 = ( n3925 & n8890 ) | ( n3925 & n19493 ) | ( n8890 & n19493 ) ;
  assign n19495 = ( n6834 & n19491 ) | ( n6834 & ~n19494 ) | ( n19491 & ~n19494 ) ;
  assign n19496 = n2907 | n17723 ;
  assign n19497 = ( ~n1064 & n12665 ) | ( ~n1064 & n19496 ) | ( n12665 & n19496 ) ;
  assign n19498 = n3109 | n7085 ;
  assign n19499 = n4892 ^ n1063 ^ 1'b0 ;
  assign n19500 = n19498 & n19499 ;
  assign n19502 = n10117 ^ n2108 ^ n1623 ;
  assign n19501 = n10367 ^ n4614 ^ n2803 ;
  assign n19503 = n19502 ^ n19501 ^ n8860 ;
  assign n19504 = ( n2757 & n5813 ) | ( n2757 & n15255 ) | ( n5813 & n15255 ) ;
  assign n19505 = ( n7271 & n8061 ) | ( n7271 & ~n9279 ) | ( n8061 & ~n9279 ) ;
  assign n19506 = n9771 ^ n3729 ^ n1050 ;
  assign n19507 = ( ~n388 & n15823 ) | ( ~n388 & n15997 ) | ( n15823 & n15997 ) ;
  assign n19508 = ( ~n4692 & n19506 ) | ( ~n4692 & n19507 ) | ( n19506 & n19507 ) ;
  assign n19509 = n14190 ^ n6729 ^ 1'b0 ;
  assign n19510 = ( ~x149 & n447 ) | ( ~x149 & n3031 ) | ( n447 & n3031 ) ;
  assign n19511 = n3913 & ~n19510 ;
  assign n19512 = n19511 ^ n11452 ^ 1'b0 ;
  assign n19513 = n10219 ^ n2597 ^ n2122 ;
  assign n19514 = ( n3968 & n11351 ) | ( n3968 & ~n15373 ) | ( n11351 & ~n15373 ) ;
  assign n19515 = ( n1047 & n8545 ) | ( n1047 & n19514 ) | ( n8545 & n19514 ) ;
  assign n19516 = ( ~n4900 & n7668 ) | ( ~n4900 & n7923 ) | ( n7668 & n7923 ) ;
  assign n19518 = ( n333 & ~n1278 ) | ( n333 & n2242 ) | ( ~n1278 & n2242 ) ;
  assign n19517 = n17275 ^ n7088 ^ x207 ;
  assign n19519 = n19518 ^ n19517 ^ n2474 ;
  assign n19520 = n19516 & ~n19519 ;
  assign n19521 = n19515 & n19520 ;
  assign n19522 = ( n4037 & ~n19513 ) | ( n4037 & n19521 ) | ( ~n19513 & n19521 ) ;
  assign n19523 = ( n2408 & n3183 ) | ( n2408 & ~n10473 ) | ( n3183 & ~n10473 ) ;
  assign n19524 = n19523 ^ n11048 ^ n8440 ;
  assign n19525 = ( n2583 & ~n7322 ) | ( n2583 & n13189 ) | ( ~n7322 & n13189 ) ;
  assign n19526 = n19525 ^ n13351 ^ n2484 ;
  assign n19527 = ( ~n1963 & n3642 ) | ( ~n1963 & n12278 ) | ( n3642 & n12278 ) ;
  assign n19528 = n17651 ^ n15112 ^ n1049 ;
  assign n19529 = ( n15697 & n19527 ) | ( n15697 & ~n19528 ) | ( n19527 & ~n19528 ) ;
  assign n19530 = n14560 ^ n1588 ^ n410 ;
  assign n19531 = n7733 ^ n7491 ^ n6189 ;
  assign n19532 = ( n724 & n12306 ) | ( n724 & n19531 ) | ( n12306 & n19531 ) ;
  assign n19533 = ( n8050 & n18609 ) | ( n8050 & n19532 ) | ( n18609 & n19532 ) ;
  assign n19534 = ~n19530 & n19533 ;
  assign n19535 = n18277 ^ n14417 ^ n11895 ;
  assign n19536 = n19535 ^ n3987 ^ 1'b0 ;
  assign n19537 = ~n5904 & n19536 ;
  assign n19538 = n2873 & ~n12409 ;
  assign n19539 = n19538 ^ n19403 ^ 1'b0 ;
  assign n19540 = ( n2036 & n10804 ) | ( n2036 & n19539 ) | ( n10804 & n19539 ) ;
  assign n19548 = n7352 & ~n19078 ;
  assign n19549 = n19548 ^ n4771 ^ n3116 ;
  assign n19541 = ( n503 & n5893 ) | ( n503 & n6872 ) | ( n5893 & n6872 ) ;
  assign n19542 = n7954 & ~n19541 ;
  assign n19543 = n15099 & n19542 ;
  assign n19544 = n7759 ^ n3900 ^ n2138 ;
  assign n19545 = ( n3162 & n8523 ) | ( n3162 & n19544 ) | ( n8523 & n19544 ) ;
  assign n19546 = ( n7949 & n19543 ) | ( n7949 & ~n19545 ) | ( n19543 & ~n19545 ) ;
  assign n19547 = n8934 & n19546 ;
  assign n19550 = n19549 ^ n19547 ^ 1'b0 ;
  assign n19551 = n11592 ^ n6447 ^ n5422 ;
  assign n19552 = n7468 ^ n2226 ^ 1'b0 ;
  assign n19553 = ( x16 & n5504 ) | ( x16 & ~n19552 ) | ( n5504 & ~n19552 ) ;
  assign n19554 = ( n15392 & ~n19551 ) | ( n15392 & n19553 ) | ( ~n19551 & n19553 ) ;
  assign n19555 = ( n813 & n1456 ) | ( n813 & n2664 ) | ( n1456 & n2664 ) ;
  assign n19556 = ~n5346 & n8213 ;
  assign n19557 = n4026 & n19556 ;
  assign n19558 = ( x206 & n647 ) | ( x206 & n7425 ) | ( n647 & n7425 ) ;
  assign n19559 = ( n19555 & n19557 ) | ( n19555 & ~n19558 ) | ( n19557 & ~n19558 ) ;
  assign n19560 = n19559 ^ n12809 ^ 1'b0 ;
  assign n19561 = ( n5994 & n19554 ) | ( n5994 & ~n19560 ) | ( n19554 & ~n19560 ) ;
  assign n19564 = n4310 ^ x246 ^ 1'b0 ;
  assign n19562 = n8780 ^ x91 ^ 1'b0 ;
  assign n19563 = n9227 | n19562 ;
  assign n19565 = n19564 ^ n19563 ^ 1'b0 ;
  assign n19566 = n15657 | n18353 ;
  assign n19567 = n16520 ^ n7248 ^ 1'b0 ;
  assign n19568 = n19567 ^ n1819 ^ 1'b0 ;
  assign n19569 = n19566 & ~n19568 ;
  assign n19570 = x191 & ~n14343 ;
  assign n19571 = ( n4512 & ~n6213 ) | ( n4512 & n9601 ) | ( ~n6213 & n9601 ) ;
  assign n19572 = n915 & ~n19571 ;
  assign n19573 = n19572 ^ n2982 ^ 1'b0 ;
  assign n19574 = ( ~n3487 & n5704 ) | ( ~n3487 & n17096 ) | ( n5704 & n17096 ) ;
  assign n19575 = n19574 ^ n12842 ^ n8710 ;
  assign n19576 = n5391 & ~n14107 ;
  assign n19577 = ( ~n3303 & n11818 ) | ( ~n3303 & n19576 ) | ( n11818 & n19576 ) ;
  assign n19578 = ( ~n9003 & n13474 ) | ( ~n9003 & n19577 ) | ( n13474 & n19577 ) ;
  assign n19579 = ( ~n2291 & n11971 ) | ( ~n2291 & n17468 ) | ( n11971 & n17468 ) ;
  assign n19580 = ( n9243 & n9826 ) | ( n9243 & ~n13110 ) | ( n9826 & ~n13110 ) ;
  assign n19581 = ( ~n1988 & n4920 ) | ( ~n1988 & n12723 ) | ( n4920 & n12723 ) ;
  assign n19582 = ( n17135 & n18403 ) | ( n17135 & ~n19581 ) | ( n18403 & ~n19581 ) ;
  assign n19583 = ( n8841 & ~n19580 ) | ( n8841 & n19582 ) | ( ~n19580 & n19582 ) ;
  assign n19584 = n12560 ^ n3693 ^ 1'b0 ;
  assign n19585 = n13144 ^ n11257 ^ 1'b0 ;
  assign n19586 = n19584 | n19585 ;
  assign n19587 = ( ~n5840 & n6745 ) | ( ~n5840 & n10260 ) | ( n6745 & n10260 ) ;
  assign n19588 = ( n3011 & n10465 ) | ( n3011 & ~n14588 ) | ( n10465 & ~n14588 ) ;
  assign n19589 = n19588 ^ n19108 ^ n5142 ;
  assign n19590 = n13298 ^ n7995 ^ 1'b0 ;
  assign n19591 = n18029 ^ n11714 ^ n4630 ;
  assign n19592 = ( n2320 & ~n3789 ) | ( n2320 & n4375 ) | ( ~n3789 & n4375 ) ;
  assign n19593 = ( n3316 & n12670 ) | ( n3316 & n15715 ) | ( n12670 & n15715 ) ;
  assign n19594 = n19593 ^ n9160 ^ n6802 ;
  assign n19595 = ( ~n14379 & n19592 ) | ( ~n14379 & n19594 ) | ( n19592 & n19594 ) ;
  assign n19596 = ( n9545 & n14271 ) | ( n9545 & ~n19595 ) | ( n14271 & ~n19595 ) ;
  assign n19597 = ( n345 & ~n19591 ) | ( n345 & n19596 ) | ( ~n19591 & n19596 ) ;
  assign n19598 = ( ~n1511 & n2700 ) | ( ~n1511 & n9616 ) | ( n2700 & n9616 ) ;
  assign n19599 = n19598 ^ n10045 ^ n2691 ;
  assign n19600 = n1875 | n2073 ;
  assign n19601 = n19599 | n19600 ;
  assign n19602 = n7539 ^ n5233 ^ n4706 ;
  assign n19603 = n19602 ^ n4131 ^ 1'b0 ;
  assign n19604 = ~n9537 & n19603 ;
  assign n19605 = ( ~n7427 & n9459 ) | ( ~n7427 & n11181 ) | ( n9459 & n11181 ) ;
  assign n19606 = ( n4368 & ~n13637 ) | ( n4368 & n19605 ) | ( ~n13637 & n19605 ) ;
  assign n19607 = ( ~n4943 & n19604 ) | ( ~n4943 & n19606 ) | ( n19604 & n19606 ) ;
  assign n19608 = n19607 ^ n17885 ^ n1993 ;
  assign n19609 = n11165 ^ n2324 ^ 1'b0 ;
  assign n19610 = n19609 ^ n18670 ^ n10894 ;
  assign n19611 = n13347 ^ n2562 ^ n2216 ;
  assign n19612 = ( n776 & n3074 ) | ( n776 & n19611 ) | ( n3074 & n19611 ) ;
  assign n19613 = n19612 ^ n14895 ^ 1'b0 ;
  assign n19614 = n5552 ^ n1608 ^ 1'b0 ;
  assign n19615 = ~n9274 & n19614 ;
  assign n19616 = ~n1669 & n19615 ;
  assign n19617 = n19616 ^ n9381 ^ 1'b0 ;
  assign n19618 = ( n10382 & ~n19613 ) | ( n10382 & n19617 ) | ( ~n19613 & n19617 ) ;
  assign n19619 = n14523 ^ n8397 ^ 1'b0 ;
  assign n19620 = ~n8983 & n19619 ;
  assign n19621 = n14282 | n19620 ;
  assign n19622 = ( n4748 & n9079 ) | ( n4748 & ~n14164 ) | ( n9079 & ~n14164 ) ;
  assign n19623 = ( n8377 & n15570 ) | ( n8377 & n17132 ) | ( n15570 & n17132 ) ;
  assign n19624 = ( n2921 & n14443 ) | ( n2921 & ~n19623 ) | ( n14443 & ~n19623 ) ;
  assign n19625 = ( n4683 & n11083 ) | ( n4683 & n16699 ) | ( n11083 & n16699 ) ;
  assign n19626 = n19625 ^ n11672 ^ n10650 ;
  assign n19627 = n1962 | n8472 ;
  assign n19628 = n19626 | n19627 ;
  assign n19629 = n7455 & n19628 ;
  assign n19630 = n19034 ^ n16905 ^ 1'b0 ;
  assign n19631 = n5602 | n19630 ;
  assign n19632 = n15725 ^ n1481 ^ 1'b0 ;
  assign n19633 = ( n4915 & ~n6090 ) | ( n4915 & n7027 ) | ( ~n6090 & n7027 ) ;
  assign n19634 = ( n14661 & n14951 ) | ( n14661 & n18415 ) | ( n14951 & n18415 ) ;
  assign n19635 = ~n5505 & n19634 ;
  assign n19636 = n19633 & n19635 ;
  assign n19637 = n19636 ^ n7672 ^ n1673 ;
  assign n19638 = n1212 | n3347 ;
  assign n19639 = n3397 ^ x186 ^ 1'b0 ;
  assign n19640 = n14591 & n19639 ;
  assign n19641 = n19640 ^ n2794 ^ n2368 ;
  assign n19642 = n19641 ^ n8545 ^ n3044 ;
  assign n19643 = ( n5836 & ~n11152 ) | ( n5836 & n15951 ) | ( ~n11152 & n15951 ) ;
  assign n19644 = n16519 ^ n11005 ^ 1'b0 ;
  assign n19652 = n4948 ^ n4294 ^ n3800 ;
  assign n19650 = n1430 & ~n10687 ;
  assign n19651 = n8794 & n19650 ;
  assign n19653 = n19652 ^ n19651 ^ n5071 ;
  assign n19646 = ( ~n6888 & n8937 ) | ( ~n6888 & n16271 ) | ( n8937 & n16271 ) ;
  assign n19647 = ( ~n1393 & n5479 ) | ( ~n1393 & n19646 ) | ( n5479 & n19646 ) ;
  assign n19648 = ( ~n1137 & n10138 ) | ( ~n1137 & n19647 ) | ( n10138 & n19647 ) ;
  assign n19649 = n1289 & ~n19648 ;
  assign n19654 = n19653 ^ n19649 ^ 1'b0 ;
  assign n19645 = ~n6977 & n9037 ;
  assign n19655 = n19654 ^ n19645 ^ 1'b0 ;
  assign n19658 = ( ~n1958 & n4283 ) | ( ~n1958 & n6452 ) | ( n4283 & n6452 ) ;
  assign n19659 = n5019 & n8523 ;
  assign n19660 = ( ~n15489 & n19658 ) | ( ~n15489 & n19659 ) | ( n19658 & n19659 ) ;
  assign n19656 = n7084 ^ n281 ^ 1'b0 ;
  assign n19657 = ( ~n9981 & n15025 ) | ( ~n9981 & n19656 ) | ( n15025 & n19656 ) ;
  assign n19661 = n19660 ^ n19657 ^ n10612 ;
  assign n19662 = ( n3535 & n19548 ) | ( n3535 & n19661 ) | ( n19548 & n19661 ) ;
  assign n19663 = n17388 ^ n7693 ^ n4015 ;
  assign n19664 = n19663 ^ n5969 ^ n2942 ;
  assign n19665 = n19664 ^ n11167 ^ 1'b0 ;
  assign n19666 = ( x94 & n2553 ) | ( x94 & n17692 ) | ( n2553 & n17692 ) ;
  assign n19667 = ( n6744 & n10442 ) | ( n6744 & n19666 ) | ( n10442 & n19666 ) ;
  assign n19668 = n11650 | n15039 ;
  assign n19669 = n19668 ^ n3833 ^ 1'b0 ;
  assign n19670 = ( n3702 & n9161 ) | ( n3702 & ~n19669 ) | ( n9161 & ~n19669 ) ;
  assign n19671 = n19670 ^ n13265 ^ 1'b0 ;
  assign n19672 = n19671 ^ n9636 ^ 1'b0 ;
  assign n19673 = n14893 & n19672 ;
  assign n19674 = ( n5496 & n7765 ) | ( n5496 & ~n19673 ) | ( n7765 & ~n19673 ) ;
  assign n19675 = n13337 ^ n9576 ^ n5983 ;
  assign n19676 = n5223 & ~n19675 ;
  assign n19679 = n13838 ^ n7562 ^ n1779 ;
  assign n19677 = n6749 & ~n9206 ;
  assign n19678 = n16478 | n19677 ;
  assign n19680 = n19679 ^ n19678 ^ 1'b0 ;
  assign n19683 = n19656 ^ n16547 ^ n727 ;
  assign n19681 = n1427 & n3109 ;
  assign n19682 = n19681 ^ n18396 ^ 1'b0 ;
  assign n19684 = n19683 ^ n19682 ^ n16610 ;
  assign n19685 = n19684 ^ n9698 ^ n3789 ;
  assign n19686 = ( n3725 & n12792 ) | ( n3725 & ~n17659 ) | ( n12792 & ~n17659 ) ;
  assign n19687 = n19686 ^ n6502 ^ n2454 ;
  assign n19691 = n2900 ^ n1118 ^ n283 ;
  assign n19688 = n15607 ^ n7567 ^ n2586 ;
  assign n19689 = ~n9637 & n19688 ;
  assign n19690 = n19689 ^ n15594 ^ n7371 ;
  assign n19692 = n19691 ^ n19690 ^ n8263 ;
  assign n19693 = n1362 & n16072 ;
  assign n19694 = n19693 ^ n8123 ^ 1'b0 ;
  assign n19695 = ( ~n12787 & n19692 ) | ( ~n12787 & n19694 ) | ( n19692 & n19694 ) ;
  assign n19696 = ~n11921 & n12287 ;
  assign n19697 = n19696 ^ n5795 ^ 1'b0 ;
  assign n19698 = n16979 ^ n2381 ^ 1'b0 ;
  assign n19699 = n15880 & ~n19698 ;
  assign n19700 = ( ~n19626 & n19697 ) | ( ~n19626 & n19699 ) | ( n19697 & n19699 ) ;
  assign n19701 = ( x170 & n18031 ) | ( x170 & n19226 ) | ( n18031 & n19226 ) ;
  assign n19702 = n19701 ^ n14838 ^ n5558 ;
  assign n19703 = ( ~n7162 & n9788 ) | ( ~n7162 & n18280 ) | ( n9788 & n18280 ) ;
  assign n19704 = n18611 ^ n11353 ^ n8102 ;
  assign n19705 = n7414 ^ n1122 ^ 1'b0 ;
  assign n19706 = n11641 & n19705 ;
  assign n19707 = ~n11961 & n19706 ;
  assign n19708 = n19707 ^ n16161 ^ 1'b0 ;
  assign n19709 = ( n2146 & ~n5937 ) | ( n2146 & n9901 ) | ( ~n5937 & n9901 ) ;
  assign n19710 = ( n4942 & ~n9385 ) | ( n4942 & n10380 ) | ( ~n9385 & n10380 ) ;
  assign n19711 = n13624 ^ n8969 ^ n4607 ;
  assign n19712 = n19711 ^ n1979 ^ 1'b0 ;
  assign n19713 = n19710 & ~n19712 ;
  assign n19714 = n19709 & n19713 ;
  assign n19715 = n3394 & n19714 ;
  assign n19716 = n5676 ^ n4559 ^ 1'b0 ;
  assign n19717 = n4206 | n19716 ;
  assign n19718 = n2656 & ~n3743 ;
  assign n19719 = n19718 ^ n6864 ^ 1'b0 ;
  assign n19720 = ( ~n8052 & n19717 ) | ( ~n8052 & n19719 ) | ( n19717 & n19719 ) ;
  assign n19721 = n19720 ^ n18637 ^ n5398 ;
  assign n19722 = n2563 & ~n18283 ;
  assign n19723 = n19721 & n19722 ;
  assign n19724 = n14762 ^ n5471 ^ n5089 ;
  assign n19725 = n19724 ^ n4841 ^ n937 ;
  assign n19726 = n3601 & ~n19725 ;
  assign n19727 = n19726 ^ n19269 ^ n628 ;
  assign n19735 = ( n944 & ~n3983 ) | ( n944 & n12774 ) | ( ~n3983 & n12774 ) ;
  assign n19736 = n19735 ^ n1033 ^ 1'b0 ;
  assign n19737 = n3538 & ~n19736 ;
  assign n19738 = n17805 & n19737 ;
  assign n19739 = n19738 ^ n2567 ^ 1'b0 ;
  assign n19732 = ( ~n4315 & n8419 ) | ( ~n4315 & n12219 ) | ( n8419 & n12219 ) ;
  assign n19728 = n12831 ^ n12592 ^ n5178 ;
  assign n19729 = n19728 ^ n8694 ^ n3497 ;
  assign n19730 = n19729 ^ n9428 ^ 1'b0 ;
  assign n19731 = n6937 | n19730 ;
  assign n19733 = n19732 ^ n19731 ^ 1'b0 ;
  assign n19734 = n5030 & ~n19733 ;
  assign n19740 = n19739 ^ n19734 ^ n747 ;
  assign n19741 = n6187 & n7570 ;
  assign n19742 = n19741 ^ n8405 ^ n8008 ;
  assign n19743 = n9647 ^ n3395 ^ 1'b0 ;
  assign n19744 = ~n14728 & n19743 ;
  assign n19745 = ( ~n7232 & n7384 ) | ( ~n7232 & n8902 ) | ( n7384 & n8902 ) ;
  assign n19746 = ( n9828 & n15898 ) | ( n9828 & n19745 ) | ( n15898 & n19745 ) ;
  assign n19747 = ( n2231 & n2821 ) | ( n2231 & ~n14111 ) | ( n2821 & ~n14111 ) ;
  assign n19748 = n19747 ^ n19266 ^ n14136 ;
  assign n19749 = ( n18564 & n19746 ) | ( n18564 & ~n19748 ) | ( n19746 & ~n19748 ) ;
  assign n19750 = n13884 ^ n5370 ^ n4903 ;
  assign n19751 = n7952 ^ n5187 ^ n1686 ;
  assign n19752 = n19751 ^ n13380 ^ 1'b0 ;
  assign n19753 = n19574 ^ n11541 ^ n1951 ;
  assign n19754 = ( n19750 & n19752 ) | ( n19750 & ~n19753 ) | ( n19752 & ~n19753 ) ;
  assign n19755 = n15887 ^ n13170 ^ 1'b0 ;
  assign n19756 = n16059 & ~n19755 ;
  assign n19757 = n3675 ^ n3035 ^ n1742 ;
  assign n19758 = ( n1594 & n3044 ) | ( n1594 & n3281 ) | ( n3044 & n3281 ) ;
  assign n19759 = n19757 | n19758 ;
  assign n19760 = n3142 | n19759 ;
  assign n19761 = ( n5413 & n19756 ) | ( n5413 & ~n19760 ) | ( n19756 & ~n19760 ) ;
  assign n19762 = ( n1005 & n2602 ) | ( n1005 & ~n7273 ) | ( n2602 & ~n7273 ) ;
  assign n19763 = ( n2002 & n4644 ) | ( n2002 & n19762 ) | ( n4644 & n19762 ) ;
  assign n19764 = n19763 ^ n16437 ^ 1'b0 ;
  assign n19765 = n8951 ^ n6357 ^ n3608 ;
  assign n19767 = n18864 ^ n15809 ^ n7352 ;
  assign n19768 = n5243 & ~n19767 ;
  assign n19769 = n19768 ^ n15917 ^ n14736 ;
  assign n19766 = n346 & n8710 ;
  assign n19770 = n19769 ^ n19766 ^ 1'b0 ;
  assign n19771 = ( ~n2570 & n4654 ) | ( ~n2570 & n5660 ) | ( n4654 & n5660 ) ;
  assign n19772 = ( n1411 & ~n6829 ) | ( n1411 & n19771 ) | ( ~n6829 & n19771 ) ;
  assign n19773 = ( ~n278 & n3294 ) | ( ~n278 & n3544 ) | ( n3294 & n3544 ) ;
  assign n19774 = n19773 ^ n14410 ^ n13623 ;
  assign n19775 = n19774 ^ n13216 ^ x72 ;
  assign n19776 = n11482 ^ n7969 ^ n1411 ;
  assign n19777 = ( n516 & n1569 ) | ( n516 & ~n12856 ) | ( n1569 & ~n12856 ) ;
  assign n19778 = ( n6431 & n19776 ) | ( n6431 & n19777 ) | ( n19776 & n19777 ) ;
  assign n19779 = n6040 ^ n5325 ^ n5319 ;
  assign n19780 = ( n9503 & n17923 ) | ( n9503 & n19779 ) | ( n17923 & n19779 ) ;
  assign n19785 = n5296 | n17625 ;
  assign n19786 = n17743 & ~n19785 ;
  assign n19783 = n3756 ^ n3181 ^ 1'b0 ;
  assign n19784 = n19783 ^ n6572 ^ n3109 ;
  assign n19781 = n6445 & ~n7902 ;
  assign n19782 = n19781 ^ n8130 ^ 1'b0 ;
  assign n19787 = n19786 ^ n19784 ^ n19782 ;
  assign n19788 = ( ~n5422 & n5684 ) | ( ~n5422 & n17769 ) | ( n5684 & n17769 ) ;
  assign n19789 = ( n5851 & n8019 ) | ( n5851 & ~n19788 ) | ( n8019 & ~n19788 ) ;
  assign n19790 = n11502 ^ n4391 ^ n3899 ;
  assign n19791 = n7124 ^ n6228 ^ n5087 ;
  assign n19792 = n11016 | n19791 ;
  assign n19793 = ( ~n6054 & n19790 ) | ( ~n6054 & n19792 ) | ( n19790 & n19792 ) ;
  assign n19796 = n1310 | n6387 ;
  assign n19797 = n19796 ^ n12374 ^ 1'b0 ;
  assign n19798 = n19797 ^ n8188 ^ n6786 ;
  assign n19799 = n19798 ^ n5014 ^ x207 ;
  assign n19794 = n7795 & ~n13282 ;
  assign n19795 = n1444 & n19794 ;
  assign n19800 = n19799 ^ n19795 ^ 1'b0 ;
  assign n19801 = ( ~n2974 & n8377 ) | ( ~n2974 & n19800 ) | ( n8377 & n19800 ) ;
  assign n19802 = n19801 ^ n8718 ^ n1464 ;
  assign n19803 = n17185 ^ n5566 ^ 1'b0 ;
  assign n19804 = n1694 & ~n19803 ;
  assign n19805 = ~n10704 & n17753 ;
  assign n19806 = ~n1833 & n19805 ;
  assign n19807 = n19806 ^ n18120 ^ 1'b0 ;
  assign n19808 = ( n2197 & n3304 ) | ( n2197 & ~n3451 ) | ( n3304 & ~n3451 ) ;
  assign n19809 = n6616 ^ n649 ^ 1'b0 ;
  assign n19810 = n9414 & ~n19809 ;
  assign n19811 = ( n1172 & n19808 ) | ( n1172 & n19810 ) | ( n19808 & n19810 ) ;
  assign n19812 = ( n1561 & ~n10062 ) | ( n1561 & n19811 ) | ( ~n10062 & n19811 ) ;
  assign n19813 = n17073 ^ n4673 ^ n2246 ;
  assign n19814 = n19139 & n19813 ;
  assign n19815 = ~n2292 & n19814 ;
  assign n19816 = n19815 ^ n13408 ^ n8033 ;
  assign n19817 = n16447 ^ n4932 ^ 1'b0 ;
  assign n19818 = n19817 ^ n7397 ^ 1'b0 ;
  assign n19819 = n19818 ^ n10600 ^ 1'b0 ;
  assign n19820 = n19819 ^ n3693 ^ x219 ;
  assign n19821 = ( n6346 & n8258 ) | ( n6346 & ~n10779 ) | ( n8258 & ~n10779 ) ;
  assign n19822 = ( n2499 & n7317 ) | ( n2499 & n19821 ) | ( n7317 & n19821 ) ;
  assign n19823 = ( n2965 & n10217 ) | ( n2965 & ~n19822 ) | ( n10217 & ~n19822 ) ;
  assign n19824 = ( n1107 & ~n11180 ) | ( n1107 & n15199 ) | ( ~n11180 & n15199 ) ;
  assign n19825 = n19824 ^ n7496 ^ 1'b0 ;
  assign n19826 = n19823 & ~n19825 ;
  assign n19827 = n19826 ^ n13663 ^ n10079 ;
  assign n19829 = ( ~n2932 & n7162 ) | ( ~n2932 & n15811 ) | ( n7162 & n15811 ) ;
  assign n19828 = n6803 ^ n1690 ^ 1'b0 ;
  assign n19830 = n19829 ^ n19828 ^ 1'b0 ;
  assign n19831 = ~n1868 & n6275 ;
  assign n19832 = ~n17398 & n19831 ;
  assign n19833 = n11626 ^ n7786 ^ n6355 ;
  assign n19834 = ( n464 & n18968 ) | ( n464 & ~n19833 ) | ( n18968 & ~n19833 ) ;
  assign n19835 = n19834 ^ n3155 ^ n1569 ;
  assign n19836 = ( n3855 & ~n19832 ) | ( n3855 & n19835 ) | ( ~n19832 & n19835 ) ;
  assign n19839 = ( n1807 & n8815 ) | ( n1807 & ~n18262 ) | ( n8815 & ~n18262 ) ;
  assign n19840 = n19839 ^ n4946 ^ n4718 ;
  assign n19837 = n19671 ^ n5230 ^ 1'b0 ;
  assign n19838 = n4903 & ~n19837 ;
  assign n19841 = n19840 ^ n19838 ^ n2029 ;
  assign n19842 = n7901 | n18503 ;
  assign n19843 = n19842 ^ n8103 ^ 1'b0 ;
  assign n19844 = n18378 & ~n19843 ;
  assign n19845 = n6968 & ~n12825 ;
  assign n19846 = n14820 ^ n13360 ^ 1'b0 ;
  assign n19847 = n19845 & ~n19846 ;
  assign n19848 = ( ~n3165 & n3281 ) | ( ~n3165 & n10547 ) | ( n3281 & n10547 ) ;
  assign n19849 = ( n1739 & n13463 ) | ( n1739 & n19848 ) | ( n13463 & n19848 ) ;
  assign n19850 = ( ~n3819 & n11617 ) | ( ~n3819 & n19849 ) | ( n11617 & n19849 ) ;
  assign n19851 = ( n9805 & ~n9817 ) | ( n9805 & n13069 ) | ( ~n9817 & n13069 ) ;
  assign n19852 = n15173 ^ n5779 ^ n1336 ;
  assign n19853 = n19852 ^ n803 ^ 1'b0 ;
  assign n19854 = n1842 & n19853 ;
  assign n19855 = ( n3488 & n19851 ) | ( n3488 & n19854 ) | ( n19851 & n19854 ) ;
  assign n19856 = ( ~x182 & n6525 ) | ( ~x182 & n19855 ) | ( n6525 & n19855 ) ;
  assign n19857 = ( n693 & n11630 ) | ( n693 & ~n12634 ) | ( n11630 & ~n12634 ) ;
  assign n19858 = n19857 ^ n11603 ^ n264 ;
  assign n19859 = n19858 ^ n17307 ^ n13318 ;
  assign n19860 = ( n4528 & ~n14176 ) | ( n4528 & n19859 ) | ( ~n14176 & n19859 ) ;
  assign n19866 = n13787 ^ n3520 ^ 1'b0 ;
  assign n19867 = n4724 & ~n19866 ;
  assign n19861 = ~n1677 & n3429 ;
  assign n19862 = n6809 & n19861 ;
  assign n19863 = n15311 ^ n10140 ^ n1649 ;
  assign n19864 = ( n578 & ~n19862 ) | ( n578 & n19863 ) | ( ~n19862 & n19863 ) ;
  assign n19865 = n19864 ^ n16982 ^ n5108 ;
  assign n19868 = n19867 ^ n19865 ^ n1416 ;
  assign n19869 = ( ~n9040 & n14468 ) | ( ~n9040 & n18529 ) | ( n14468 & n18529 ) ;
  assign n19870 = ( n15649 & n17660 ) | ( n15649 & n19869 ) | ( n17660 & n19869 ) ;
  assign n19871 = n561 | n10006 ;
  assign n19872 = n19871 ^ n8653 ^ 1'b0 ;
  assign n19873 = ~n3207 & n19872 ;
  assign n19874 = n19873 ^ n13233 ^ n2625 ;
  assign n19875 = n19078 ^ n7881 ^ n4999 ;
  assign n19876 = ( ~n739 & n7544 ) | ( ~n739 & n8147 ) | ( n7544 & n8147 ) ;
  assign n19877 = ( n535 & n12526 ) | ( n535 & ~n19876 ) | ( n12526 & ~n19876 ) ;
  assign n19878 = ( n12730 & n19875 ) | ( n12730 & n19877 ) | ( n19875 & n19877 ) ;
  assign n19887 = n10048 ^ n4241 ^ n2517 ;
  assign n19888 = n19887 ^ n5118 ^ n2217 ;
  assign n19879 = n13573 ^ n10873 ^ n5848 ;
  assign n19880 = n12037 ^ n5084 ^ n1767 ;
  assign n19881 = n10698 & ~n19880 ;
  assign n19882 = n19881 ^ n8559 ^ n8531 ;
  assign n19883 = n19882 ^ n19033 ^ n3976 ;
  assign n19884 = n11829 & ~n17315 ;
  assign n19885 = n19883 & n19884 ;
  assign n19886 = ( n1278 & n19879 ) | ( n1278 & n19885 ) | ( n19879 & n19885 ) ;
  assign n19889 = n19888 ^ n19886 ^ n12897 ;
  assign n19890 = ( n451 & ~n3270 ) | ( n451 & n13782 ) | ( ~n3270 & n13782 ) ;
  assign n19891 = n6330 ^ n851 ^ 1'b0 ;
  assign n19892 = ~n8485 & n19891 ;
  assign n19893 = n5906 & n9074 ;
  assign n19896 = ~n3108 & n3534 ;
  assign n19897 = n19896 ^ n14513 ^ n7281 ;
  assign n19894 = n11589 ^ n3167 ^ n2477 ;
  assign n19895 = n19894 ^ n1599 ^ n903 ;
  assign n19898 = n19897 ^ n19895 ^ n17355 ;
  assign n19905 = ( n1829 & n7399 ) | ( n1829 & ~n15206 ) | ( n7399 & ~n15206 ) ;
  assign n19902 = ( n2812 & ~n9786 ) | ( n2812 & n12183 ) | ( ~n9786 & n12183 ) ;
  assign n19903 = n19902 ^ n15198 ^ n2551 ;
  assign n19900 = n297 & ~n16451 ;
  assign n19901 = n1282 & n19900 ;
  assign n19904 = n19903 ^ n19901 ^ n14025 ;
  assign n19906 = n19905 ^ n19904 ^ n15039 ;
  assign n19899 = n8985 ^ n8486 ^ n1019 ;
  assign n19907 = n19906 ^ n19899 ^ n7828 ;
  assign n19908 = ( n2289 & n4344 ) | ( n2289 & ~n6866 ) | ( n4344 & ~n6866 ) ;
  assign n19909 = n19908 ^ n1795 ^ 1'b0 ;
  assign n19910 = ( n1997 & ~n3367 ) | ( n1997 & n8996 ) | ( ~n3367 & n8996 ) ;
  assign n19911 = ( ~n3429 & n13887 ) | ( ~n3429 & n19910 ) | ( n13887 & n19910 ) ;
  assign n19912 = n8708 ^ n8221 ^ n7034 ;
  assign n19914 = ( n1627 & n4394 ) | ( n1627 & ~n4664 ) | ( n4394 & ~n4664 ) ;
  assign n19915 = ( ~n6512 & n13378 ) | ( ~n6512 & n19914 ) | ( n13378 & n19914 ) ;
  assign n19913 = n12045 & n16365 ;
  assign n19916 = n19915 ^ n19913 ^ 1'b0 ;
  assign n19919 = n16363 ^ n5572 ^ n3049 ;
  assign n19917 = ( n962 & n5979 ) | ( n962 & n17870 ) | ( n5979 & n17870 ) ;
  assign n19918 = ( n16741 & ~n17768 ) | ( n16741 & n19917 ) | ( ~n17768 & n19917 ) ;
  assign n19920 = n19919 ^ n19918 ^ n6647 ;
  assign n19923 = n18917 ^ n539 ^ 1'b0 ;
  assign n19921 = ( n7468 & n10209 ) | ( n7468 & n13088 ) | ( n10209 & n13088 ) ;
  assign n19922 = n19921 ^ n12811 ^ n10258 ;
  assign n19924 = n19923 ^ n19922 ^ n7822 ;
  assign n19925 = n18474 ^ n15164 ^ 1'b0 ;
  assign n19926 = n10673 ^ n8076 ^ n2064 ;
  assign n19927 = n7344 ^ n3669 ^ n1806 ;
  assign n19933 = n9958 ^ n8737 ^ n308 ;
  assign n19928 = n7795 & n8689 ;
  assign n19929 = n6527 & n19928 ;
  assign n19930 = ( ~n1423 & n4920 ) | ( ~n1423 & n19929 ) | ( n4920 & n19929 ) ;
  assign n19931 = n19930 ^ n4560 ^ 1'b0 ;
  assign n19932 = ~n544 & n19931 ;
  assign n19934 = n19933 ^ n19932 ^ n15680 ;
  assign n19935 = n19927 | n19934 ;
  assign n19936 = n19368 ^ n15706 ^ n11131 ;
  assign n19937 = ( n1465 & n11980 ) | ( n1465 & n18695 ) | ( n11980 & n18695 ) ;
  assign n19938 = ( n595 & n19936 ) | ( n595 & n19937 ) | ( n19936 & n19937 ) ;
  assign n19939 = n3076 & ~n15657 ;
  assign n19940 = n17491 | n19939 ;
  assign n19941 = n3266 ^ n1373 ^ x241 ;
  assign n19942 = ( n13959 & n14229 ) | ( n13959 & n19941 ) | ( n14229 & n19941 ) ;
  assign n19943 = n17322 & ~n19942 ;
  assign n19944 = n11463 & n19943 ;
  assign n19945 = ( n13090 & n14594 ) | ( n13090 & n15254 ) | ( n14594 & n15254 ) ;
  assign n19946 = ~n11281 & n19945 ;
  assign n19947 = n19946 ^ n457 ^ 1'b0 ;
  assign n19948 = n13090 ^ n2898 ^ 1'b0 ;
  assign n19949 = ( n5135 & n16030 ) | ( n5135 & n17261 ) | ( n16030 & n17261 ) ;
  assign n19950 = ( n4213 & n19948 ) | ( n4213 & ~n19949 ) | ( n19948 & ~n19949 ) ;
  assign n19951 = n5325 | n18683 ;
  assign n19952 = n19951 ^ n7178 ^ n427 ;
  assign n19953 = n19952 ^ n5003 ^ n4676 ;
  assign n19954 = n19953 ^ n2292 ^ n1366 ;
  assign n19956 = n5791 ^ n4729 ^ n493 ;
  assign n19955 = n12599 ^ n2224 ^ n764 ;
  assign n19957 = n19956 ^ n19955 ^ n1587 ;
  assign n19961 = n6432 & ~n7149 ;
  assign n19962 = n19961 ^ n9870 ^ n4596 ;
  assign n19958 = n9780 & ~n18828 ;
  assign n19959 = ~n11760 & n19958 ;
  assign n19960 = n19959 ^ n13889 ^ n771 ;
  assign n19963 = n19962 ^ n19960 ^ n9669 ;
  assign n19964 = n3096 ^ n2235 ^ 1'b0 ;
  assign n19965 = n10977 & ~n19964 ;
  assign n19966 = ( n2991 & ~n19336 ) | ( n2991 & n19965 ) | ( ~n19336 & n19965 ) ;
  assign n19967 = n19966 ^ n17399 ^ n2659 ;
  assign n19968 = ~n11418 & n19967 ;
  assign n19969 = n15946 & n19968 ;
  assign n19973 = ~n2331 & n3637 ;
  assign n19974 = n7624 & n19973 ;
  assign n19972 = ~n3947 & n12146 ;
  assign n19975 = n19974 ^ n19972 ^ 1'b0 ;
  assign n19970 = n19102 ^ n11392 ^ 1'b0 ;
  assign n19971 = n19970 ^ n5010 ^ x215 ;
  assign n19976 = n19975 ^ n19971 ^ n7232 ;
  assign n19977 = ( n2094 & n5270 ) | ( n2094 & ~n5456 ) | ( n5270 & ~n5456 ) ;
  assign n19978 = n19977 ^ n5782 ^ n5777 ;
  assign n19979 = ( ~n3514 & n3715 ) | ( ~n3514 & n19978 ) | ( n3715 & n19978 ) ;
  assign n19980 = n12564 ^ n4255 ^ 1'b0 ;
  assign n19981 = n9874 & ~n19980 ;
  assign n19982 = n1554 & ~n3311 ;
  assign n19983 = n19982 ^ n1766 ^ 1'b0 ;
  assign n19984 = n7792 ^ n6376 ^ n2325 ;
  assign n19985 = ( n4547 & ~n14308 ) | ( n4547 & n19984 ) | ( ~n14308 & n19984 ) ;
  assign n19986 = n19985 ^ n7317 ^ 1'b0 ;
  assign n19987 = ( n5224 & ~n19983 ) | ( n5224 & n19986 ) | ( ~n19983 & n19986 ) ;
  assign n19988 = n18761 ^ n7382 ^ n1438 ;
  assign n19989 = ( n5551 & n11076 ) | ( n5551 & ~n19988 ) | ( n11076 & ~n19988 ) ;
  assign n19990 = n14137 ^ n9809 ^ n996 ;
  assign n19998 = n6661 ^ n6325 ^ n1220 ;
  assign n19999 = ( n530 & ~n7046 ) | ( n530 & n19998 ) | ( ~n7046 & n19998 ) ;
  assign n19995 = ( n1231 & n4590 ) | ( n1231 & n6595 ) | ( n4590 & n6595 ) ;
  assign n19991 = ~n8777 & n16546 ;
  assign n19992 = n15896 & n19991 ;
  assign n19993 = ( n1507 & n4481 ) | ( n1507 & ~n14252 ) | ( n4481 & ~n14252 ) ;
  assign n19994 = ( n12697 & n19992 ) | ( n12697 & n19993 ) | ( n19992 & n19993 ) ;
  assign n19996 = n19995 ^ n19994 ^ n15602 ;
  assign n19997 = n12660 & n19996 ;
  assign n20000 = n19999 ^ n19997 ^ n14405 ;
  assign n20002 = n11993 ^ n11005 ^ n4107 ;
  assign n20001 = n10672 ^ n6974 ^ 1'b0 ;
  assign n20003 = n20002 ^ n20001 ^ n17541 ;
  assign n20005 = n5344 ^ n4781 ^ n2399 ;
  assign n20004 = n2520 & ~n6269 ;
  assign n20006 = n20005 ^ n20004 ^ n14845 ;
  assign n20007 = n3507 & n20006 ;
  assign n20019 = ( n412 & n4761 ) | ( n412 & n8773 ) | ( n4761 & n8773 ) ;
  assign n20015 = n15516 ^ n12609 ^ n4168 ;
  assign n20016 = n20015 ^ n770 ^ 1'b0 ;
  assign n20017 = ~n7078 & n20016 ;
  assign n20018 = n20017 ^ n6241 ^ 1'b0 ;
  assign n20010 = n5279 ^ n2885 ^ n2526 ;
  assign n20011 = n20010 ^ n6113 ^ 1'b0 ;
  assign n20012 = n5408 & n20011 ;
  assign n20013 = n20012 ^ n6969 ^ n5172 ;
  assign n20008 = ( ~n3534 & n5250 ) | ( ~n3534 & n5361 ) | ( n5250 & n5361 ) ;
  assign n20009 = ( n10673 & ~n14273 ) | ( n10673 & n20008 ) | ( ~n14273 & n20008 ) ;
  assign n20014 = n20013 ^ n20009 ^ n16902 ;
  assign n20020 = n20019 ^ n20018 ^ n20014 ;
  assign n20021 = ( n8846 & n9532 ) | ( n8846 & ~n16240 ) | ( n9532 & ~n16240 ) ;
  assign n20022 = n20021 ^ n14761 ^ 1'b0 ;
  assign n20023 = n20022 ^ n14317 ^ 1'b0 ;
  assign n20024 = ( ~n1390 & n5886 ) | ( ~n1390 & n6833 ) | ( n5886 & n6833 ) ;
  assign n20025 = n11621 ^ n7100 ^ n3961 ;
  assign n20026 = n10416 ^ n1242 ^ n1134 ;
  assign n20027 = n11497 & ~n12104 ;
  assign n20028 = ~n10431 & n20027 ;
  assign n20029 = ( n690 & n1712 ) | ( n690 & n6740 ) | ( n1712 & n6740 ) ;
  assign n20030 = ( n10165 & n10673 ) | ( n10165 & n20029 ) | ( n10673 & n20029 ) ;
  assign n20031 = n8517 ^ n8016 ^ n6745 ;
  assign n20032 = n20031 ^ n15414 ^ n11221 ;
  assign n20033 = ( n12519 & ~n20030 ) | ( n12519 & n20032 ) | ( ~n20030 & n20032 ) ;
  assign n20034 = ( ~n2171 & n20028 ) | ( ~n2171 & n20033 ) | ( n20028 & n20033 ) ;
  assign n20035 = ( ~n8099 & n20026 ) | ( ~n8099 & n20034 ) | ( n20026 & n20034 ) ;
  assign n20036 = n3178 ^ n1352 ^ 1'b0 ;
  assign n20037 = ~n8666 & n20036 ;
  assign n20038 = ( ~n321 & n7093 ) | ( ~n321 & n8383 ) | ( n7093 & n8383 ) ;
  assign n20039 = n20038 ^ n4801 ^ 1'b0 ;
  assign n20040 = n20037 & n20039 ;
  assign n20041 = n20040 ^ n5875 ^ 1'b0 ;
  assign n20042 = ( n995 & n5314 ) | ( n995 & ~n8691 ) | ( n5314 & ~n8691 ) ;
  assign n20043 = n4905 & n20042 ;
  assign n20044 = n20043 ^ n4795 ^ 1'b0 ;
  assign n20045 = n20044 ^ n14376 ^ n1423 ;
  assign n20046 = ( ~n6397 & n20041 ) | ( ~n6397 & n20045 ) | ( n20041 & n20045 ) ;
  assign n20047 = n17329 ^ n12240 ^ n2427 ;
  assign n20048 = ~n1224 & n4552 ;
  assign n20049 = ~n466 & n20048 ;
  assign n20050 = ( n1275 & ~n4748 ) | ( n1275 & n20049 ) | ( ~n4748 & n20049 ) ;
  assign n20051 = n11988 & n20050 ;
  assign n20052 = n20051 ^ n13088 ^ n12260 ;
  assign n20053 = ( n4432 & ~n20047 ) | ( n4432 & n20052 ) | ( ~n20047 & n20052 ) ;
  assign n20054 = ( n9655 & n11933 ) | ( n9655 & n20053 ) | ( n11933 & n20053 ) ;
  assign n20055 = n16089 ^ n9499 ^ 1'b0 ;
  assign n20056 = n6506 & n8967 ;
  assign n20057 = n20055 & n20056 ;
  assign n20058 = n10660 & ~n12188 ;
  assign n20059 = n1692 & ~n18320 ;
  assign n20060 = ~n20058 & n20059 ;
  assign n20061 = n10014 | n12256 ;
  assign n20062 = n20061 ^ n2561 ^ 1'b0 ;
  assign n20063 = n20062 ^ n8786 ^ 1'b0 ;
  assign n20064 = ~n11802 & n20063 ;
  assign n20065 = ~n3272 & n7504 ;
  assign n20066 = n6336 & n20065 ;
  assign n20067 = ( n6723 & n16088 ) | ( n6723 & n20066 ) | ( n16088 & n20066 ) ;
  assign n20068 = n5199 ^ n536 ^ n317 ;
  assign n20069 = ~n720 & n20068 ;
  assign n20070 = ~n11455 & n20069 ;
  assign n20071 = ( n5241 & n20067 ) | ( n5241 & n20070 ) | ( n20067 & n20070 ) ;
  assign n20072 = n12158 ^ n9695 ^ 1'b0 ;
  assign n20073 = n295 & ~n20072 ;
  assign n20074 = ( n8842 & n15141 ) | ( n8842 & n20073 ) | ( n15141 & n20073 ) ;
  assign n20075 = n1605 & n11830 ;
  assign n20076 = ~n20074 & n20075 ;
  assign n20077 = n2298 | n10678 ;
  assign n20078 = ( n2093 & n2378 ) | ( n2093 & n20077 ) | ( n2378 & n20077 ) ;
  assign n20080 = ~n701 & n1775 ;
  assign n20081 = n20080 ^ n12338 ^ n6966 ;
  assign n20079 = n8904 & ~n11195 ;
  assign n20082 = n20081 ^ n20079 ^ 1'b0 ;
  assign n20083 = ~n20078 & n20082 ;
  assign n20085 = ( x152 & n4840 ) | ( x152 & n6463 ) | ( n4840 & n6463 ) ;
  assign n20084 = n14036 ^ n9546 ^ 1'b0 ;
  assign n20086 = n20085 ^ n20084 ^ n15832 ;
  assign n20087 = n20086 ^ n17315 ^ n15191 ;
  assign n20088 = n20087 ^ n18983 ^ n1085 ;
  assign n20090 = n9601 ^ n5552 ^ n3196 ;
  assign n20091 = n3954 | n20090 ;
  assign n20092 = n20091 ^ n7058 ^ 1'b0 ;
  assign n20089 = n14720 ^ n1535 ^ n823 ;
  assign n20093 = n20092 ^ n20089 ^ n4738 ;
  assign n20094 = ( n7656 & n8795 ) | ( n7656 & ~n10370 ) | ( n8795 & ~n10370 ) ;
  assign n20095 = n11920 & ~n12711 ;
  assign n20096 = n20095 ^ n7230 ^ 1'b0 ;
  assign n20097 = n20096 ^ n11026 ^ 1'b0 ;
  assign n20098 = ( ~n11461 & n20094 ) | ( ~n11461 & n20097 ) | ( n20094 & n20097 ) ;
  assign n20099 = n18666 ^ n6884 ^ 1'b0 ;
  assign n20100 = n8631 | n20099 ;
  assign n20101 = n15792 ^ n6247 ^ n2838 ;
  assign n20102 = ( n10177 & ~n20100 ) | ( n10177 & n20101 ) | ( ~n20100 & n20101 ) ;
  assign n20103 = n20102 ^ n8339 ^ 1'b0 ;
  assign n20104 = n10303 | n17066 ;
  assign n20105 = n20104 ^ n9183 ^ 1'b0 ;
  assign n20106 = n20105 ^ n8150 ^ 1'b0 ;
  assign n20107 = ~n12975 & n20106 ;
  assign n20108 = ( n11152 & n12619 ) | ( n11152 & n14608 ) | ( n12619 & n14608 ) ;
  assign n20109 = n8684 ^ n4108 ^ n1218 ;
  assign n20110 = ( ~n272 & n20108 ) | ( ~n272 & n20109 ) | ( n20108 & n20109 ) ;
  assign n20111 = n4037 ^ n720 ^ 1'b0 ;
  assign n20112 = n13865 | n20111 ;
  assign n20113 = ( n3708 & n15244 ) | ( n3708 & n20112 ) | ( n15244 & n20112 ) ;
  assign n20114 = n2082 | n7564 ;
  assign n20115 = n20113 & ~n20114 ;
  assign n20116 = n20115 ^ n12623 ^ n10987 ;
  assign n20117 = n888 & n3232 ;
  assign n20118 = n5959 ^ n2602 ^ n2467 ;
  assign n20119 = ( n8475 & n13702 ) | ( n8475 & n20118 ) | ( n13702 & n20118 ) ;
  assign n20123 = n10153 ^ n10123 ^ 1'b0 ;
  assign n20120 = n3417 & n5785 ;
  assign n20121 = n8408 & ~n20120 ;
  assign n20122 = n20121 ^ n1155 ^ 1'b0 ;
  assign n20124 = n20123 ^ n20122 ^ x209 ;
  assign n20125 = ( n1007 & n20119 ) | ( n1007 & ~n20124 ) | ( n20119 & ~n20124 ) ;
  assign n20126 = n6463 | n15805 ;
  assign n20127 = n1692 & ~n5565 ;
  assign n20128 = n20127 ^ n7019 ^ 1'b0 ;
  assign n20129 = n20128 ^ n17566 ^ n14360 ;
  assign n20130 = n11807 ^ n11142 ^ n9211 ;
  assign n20131 = n20130 ^ n19513 ^ n7153 ;
  assign n20132 = ( n9695 & n15286 ) | ( n9695 & ~n17823 ) | ( n15286 & ~n17823 ) ;
  assign n20133 = ( n4894 & n9419 ) | ( n4894 & n13783 ) | ( n9419 & n13783 ) ;
  assign n20134 = ~n10237 & n20133 ;
  assign n20135 = ~n20132 & n20134 ;
  assign n20136 = n2803 & ~n11706 ;
  assign n20137 = ~n4521 & n20136 ;
  assign n20138 = n4215 | n20137 ;
  assign n20139 = x28 | n13286 ;
  assign n20141 = ( ~n2412 & n6206 ) | ( ~n2412 & n6574 ) | ( n6206 & n6574 ) ;
  assign n20142 = n2350 ^ n681 ^ 1'b0 ;
  assign n20143 = n2717 & ~n20142 ;
  assign n20144 = ~n3691 & n20143 ;
  assign n20145 = ( n13903 & n20141 ) | ( n13903 & n20144 ) | ( n20141 & n20144 ) ;
  assign n20140 = n18559 ^ n10323 ^ n6996 ;
  assign n20146 = n20145 ^ n20140 ^ 1'b0 ;
  assign n20147 = n20139 & n20146 ;
  assign n20148 = n17492 | n18113 ;
  assign n20149 = n14557 | n20148 ;
  assign n20150 = n838 & ~n20149 ;
  assign n20151 = ( n15880 & n19288 ) | ( n15880 & ~n20150 ) | ( n19288 & ~n20150 ) ;
  assign n20152 = n3369 ^ n2823 ^ 1'b0 ;
  assign n20153 = n7850 | n11263 ;
  assign n20154 = n14894 ^ n6402 ^ n3486 ;
  assign n20155 = n3187 | n11541 ;
  assign n20156 = n20154 | n20155 ;
  assign n20157 = ( n20152 & ~n20153 ) | ( n20152 & n20156 ) | ( ~n20153 & n20156 ) ;
  assign n20158 = n7060 ^ n3324 ^ 1'b0 ;
  assign n20159 = ( n14176 & ~n16689 ) | ( n14176 & n20158 ) | ( ~n16689 & n20158 ) ;
  assign n20160 = ~n830 & n20159 ;
  assign n20161 = ~n2456 & n20160 ;
  assign n20165 = ( n2115 & n5133 ) | ( n2115 & ~n6156 ) | ( n5133 & ~n6156 ) ;
  assign n20162 = ~n5558 & n7932 ;
  assign n20163 = ~n12932 & n20162 ;
  assign n20164 = n20163 ^ n675 ^ 1'b0 ;
  assign n20166 = n20165 ^ n20164 ^ n10189 ;
  assign n20167 = n5774 & ~n9054 ;
  assign n20168 = n20167 ^ n3480 ^ 1'b0 ;
  assign n20169 = ( n1519 & ~n6913 ) | ( n1519 & n12754 ) | ( ~n6913 & n12754 ) ;
  assign n20170 = n20169 ^ n8834 ^ n6813 ;
  assign n20171 = ( n2659 & n9988 ) | ( n2659 & n20170 ) | ( n9988 & n20170 ) ;
  assign n20172 = ( ~n4482 & n20168 ) | ( ~n4482 & n20171 ) | ( n20168 & n20171 ) ;
  assign n20173 = n20166 & n20172 ;
  assign n20174 = ( ~n3085 & n20161 ) | ( ~n3085 & n20173 ) | ( n20161 & n20173 ) ;
  assign n20175 = ( n1116 & n5413 ) | ( n1116 & n20170 ) | ( n5413 & n20170 ) ;
  assign n20176 = n9435 ^ n4948 ^ 1'b0 ;
  assign n20177 = n20175 & n20176 ;
  assign n20178 = ( ~n778 & n8360 ) | ( ~n778 & n9794 ) | ( n8360 & n9794 ) ;
  assign n20181 = n7082 ^ n4997 ^ n2898 ;
  assign n20179 = ( ~n1481 & n4452 ) | ( ~n1481 & n14215 ) | ( n4452 & n14215 ) ;
  assign n20180 = ( n11004 & ~n15860 ) | ( n11004 & n20179 ) | ( ~n15860 & n20179 ) ;
  assign n20182 = n20181 ^ n20180 ^ n2971 ;
  assign n20183 = ( n6160 & n20178 ) | ( n6160 & ~n20182 ) | ( n20178 & ~n20182 ) ;
  assign n20185 = n19263 ^ n11777 ^ 1'b0 ;
  assign n20186 = n6250 & n20185 ;
  assign n20184 = n17778 ^ n12887 ^ n5697 ;
  assign n20187 = n20186 ^ n20184 ^ n9185 ;
  assign n20188 = ( n542 & n1393 ) | ( n542 & n17889 ) | ( n1393 & n17889 ) ;
  assign n20189 = n20188 ^ n15904 ^ n1839 ;
  assign n20190 = n20189 ^ n15433 ^ n4765 ;
  assign n20191 = ( ~n9749 & n12168 ) | ( ~n9749 & n20190 ) | ( n12168 & n20190 ) ;
  assign n20192 = n9296 ^ n5245 ^ 1'b0 ;
  assign n20193 = n16700 & ~n20192 ;
  assign n20194 = n4907 ^ n2514 ^ 1'b0 ;
  assign n20195 = n20194 ^ n18822 ^ n9725 ;
  assign n20196 = n16237 ^ n3110 ^ 1'b0 ;
  assign n20197 = n18410 & ~n20196 ;
  assign n20198 = x140 & n20197 ;
  assign n20199 = ~n2231 & n20198 ;
  assign n20200 = n5278 ^ n2608 ^ n1390 ;
  assign n20201 = ( n1218 & n9942 ) | ( n1218 & n20200 ) | ( n9942 & n20200 ) ;
  assign n20202 = ( n7609 & n19146 ) | ( n7609 & n20201 ) | ( n19146 & n20201 ) ;
  assign n20206 = n4399 ^ n1431 ^ n475 ;
  assign n20207 = n3620 & n6860 ;
  assign n20208 = ( n15016 & n20206 ) | ( n15016 & n20207 ) | ( n20206 & n20207 ) ;
  assign n20203 = n13127 ^ n5183 ^ 1'b0 ;
  assign n20204 = ( ~n960 & n18449 ) | ( ~n960 & n20203 ) | ( n18449 & n20203 ) ;
  assign n20205 = ( n9809 & n19717 ) | ( n9809 & n20204 ) | ( n19717 & n20204 ) ;
  assign n20209 = n20208 ^ n20205 ^ n14573 ;
  assign n20210 = n20209 ^ n19451 ^ n10786 ;
  assign n20211 = ( ~n14166 & n20202 ) | ( ~n14166 & n20210 ) | ( n20202 & n20210 ) ;
  assign n20212 = ( ~n16136 & n20199 ) | ( ~n16136 & n20211 ) | ( n20199 & n20211 ) ;
  assign n20213 = ( n407 & n1414 ) | ( n407 & n13819 ) | ( n1414 & n13819 ) ;
  assign n20214 = ~n4062 & n20213 ;
  assign n20215 = n20214 ^ n9011 ^ 1'b0 ;
  assign n20216 = ~n3660 & n18427 ;
  assign n20217 = n20216 ^ n10249 ^ 1'b0 ;
  assign n20218 = n14016 ^ n12665 ^ n1592 ;
  assign n20219 = n1390 & n20218 ;
  assign n20220 = ( n1288 & n12992 ) | ( n1288 & ~n15288 ) | ( n12992 & ~n15288 ) ;
  assign n20221 = n20220 ^ n10746 ^ n2517 ;
  assign n20222 = n4670 & ~n5613 ;
  assign n20223 = n20222 ^ x170 ^ 1'b0 ;
  assign n20224 = n9694 ^ n6470 ^ n5516 ;
  assign n20225 = ( n14824 & n20223 ) | ( n14824 & ~n20224 ) | ( n20223 & ~n20224 ) ;
  assign n20226 = n10618 ^ n4234 ^ n3624 ;
  assign n20227 = n17666 ^ n4408 ^ n2810 ;
  assign n20228 = ( n2286 & ~n20226 ) | ( n2286 & n20227 ) | ( ~n20226 & n20227 ) ;
  assign n20229 = n12479 ^ n1686 ^ n1677 ;
  assign n20230 = n20229 ^ n2183 ^ n872 ;
  assign n20233 = n12307 ^ n2859 ^ 1'b0 ;
  assign n20234 = n9255 & n20233 ;
  assign n20231 = ( n7099 & ~n11038 ) | ( n7099 & n11540 ) | ( ~n11038 & n11540 ) ;
  assign n20232 = ( n13022 & ~n16456 ) | ( n13022 & n20231 ) | ( ~n16456 & n20231 ) ;
  assign n20235 = n20234 ^ n20232 ^ n18378 ;
  assign n20240 = n6658 & ~n17059 ;
  assign n20236 = ( n3234 & ~n6077 ) | ( n3234 & n16341 ) | ( ~n6077 & n16341 ) ;
  assign n20237 = n20236 ^ n4755 ^ x97 ;
  assign n20238 = ( n4574 & n9193 ) | ( n4574 & n20237 ) | ( n9193 & n20237 ) ;
  assign n20239 = ( n3950 & n6554 ) | ( n3950 & ~n20238 ) | ( n6554 & ~n20238 ) ;
  assign n20241 = n20240 ^ n20239 ^ n3004 ;
  assign n20242 = ( n4537 & ~n4933 ) | ( n4537 & n20141 ) | ( ~n4933 & n20141 ) ;
  assign n20243 = n20242 ^ n7433 ^ n7300 ;
  assign n20246 = ( n4749 & n10837 ) | ( n4749 & ~n17093 ) | ( n10837 & ~n17093 ) ;
  assign n20244 = ( ~n6830 & n17421 ) | ( ~n6830 & n17424 ) | ( n17421 & n17424 ) ;
  assign n20245 = ( n15867 & ~n19714 ) | ( n15867 & n20244 ) | ( ~n19714 & n20244 ) ;
  assign n20247 = n20246 ^ n20245 ^ n8124 ;
  assign n20248 = ( ~n2293 & n9968 ) | ( ~n2293 & n20247 ) | ( n9968 & n20247 ) ;
  assign n20249 = ( ~n6517 & n20243 ) | ( ~n6517 & n20248 ) | ( n20243 & n20248 ) ;
  assign n20250 = n18029 ^ n2392 ^ n417 ;
  assign n20251 = ( n1446 & ~n2465 ) | ( n1446 & n20250 ) | ( ~n2465 & n20250 ) ;
  assign n20254 = n18119 ^ n11061 ^ 1'b0 ;
  assign n20252 = ~n5849 & n8858 ;
  assign n20253 = n20252 ^ n15099 ^ 1'b0 ;
  assign n20255 = n20254 ^ n20253 ^ n10007 ;
  assign n20256 = ( n2466 & ~n20251 ) | ( n2466 & n20255 ) | ( ~n20251 & n20255 ) ;
  assign n20257 = n1897 & ~n9938 ;
  assign n20258 = ( n653 & ~n9451 ) | ( n653 & n20257 ) | ( ~n9451 & n20257 ) ;
  assign n20259 = ~n5848 & n20258 ;
  assign n20260 = n20259 ^ n9258 ^ 1'b0 ;
  assign n20261 = n12179 ^ n10435 ^ 1'b0 ;
  assign n20262 = n20149 & n20261 ;
  assign n20263 = n1849 | n9635 ;
  assign n20264 = n2518 & ~n20263 ;
  assign n20265 = n20264 ^ n10505 ^ n889 ;
  assign n20266 = ( ~n5580 & n18223 ) | ( ~n5580 & n20265 ) | ( n18223 & n20265 ) ;
  assign n20267 = n9364 & ~n18958 ;
  assign n20268 = n17131 | n20267 ;
  assign n20269 = n20268 ^ n594 ^ 1'b0 ;
  assign n20270 = ( n276 & n6917 ) | ( n276 & ~n20269 ) | ( n6917 & ~n20269 ) ;
  assign n20271 = ( n7905 & n15963 ) | ( n7905 & n20270 ) | ( n15963 & n20270 ) ;
  assign n20272 = ( ~n5257 & n5728 ) | ( ~n5257 & n11939 ) | ( n5728 & n11939 ) ;
  assign n20273 = ( n5246 & ~n9091 ) | ( n5246 & n20272 ) | ( ~n9091 & n20272 ) ;
  assign n20279 = n6928 & ~n7991 ;
  assign n20280 = n20279 ^ n15003 ^ 1'b0 ;
  assign n20274 = ( x153 & ~n506 ) | ( x153 & n2351 ) | ( ~n506 & n2351 ) ;
  assign n20275 = ( n10965 & n17425 ) | ( n10965 & n20274 ) | ( n17425 & n20274 ) ;
  assign n20276 = ( n1372 & ~n9539 ) | ( n1372 & n20275 ) | ( ~n9539 & n20275 ) ;
  assign n20277 = n20265 ^ n5012 ^ n2070 ;
  assign n20278 = ( n3379 & ~n20276 ) | ( n3379 & n20277 ) | ( ~n20276 & n20277 ) ;
  assign n20281 = n20280 ^ n20278 ^ n14449 ;
  assign n20282 = n9897 & ~n18047 ;
  assign n20283 = n17934 ^ n5701 ^ 1'b0 ;
  assign n20284 = n3421 ^ n673 ^ 1'b0 ;
  assign n20285 = ( n475 & n6489 ) | ( n475 & ~n20284 ) | ( n6489 & ~n20284 ) ;
  assign n20286 = n7828 ^ n3084 ^ 1'b0 ;
  assign n20287 = ~n20285 & n20286 ;
  assign n20288 = n9628 ^ n5558 ^ n4781 ;
  assign n20289 = ( n3056 & n20287 ) | ( n3056 & ~n20288 ) | ( n20287 & ~n20288 ) ;
  assign n20291 = n3345 & ~n18143 ;
  assign n20292 = n20291 ^ n14121 ^ 1'b0 ;
  assign n20290 = n9402 | n13906 ;
  assign n20293 = n20292 ^ n20290 ^ n388 ;
  assign n20294 = n16879 ^ n12884 ^ 1'b0 ;
  assign n20295 = n2607 | n20294 ;
  assign n20296 = ( ~n367 & n1173 ) | ( ~n367 & n4867 ) | ( n1173 & n4867 ) ;
  assign n20297 = n20296 ^ n15775 ^ n1611 ;
  assign n20298 = ( n15265 & ~n20295 ) | ( n15265 & n20297 ) | ( ~n20295 & n20297 ) ;
  assign n20299 = n20298 ^ n16646 ^ 1'b0 ;
  assign n20300 = ( n4521 & n10868 ) | ( n4521 & ~n11490 ) | ( n10868 & ~n11490 ) ;
  assign n20301 = ( n2433 & ~n19735 ) | ( n2433 & n20300 ) | ( ~n19735 & n20300 ) ;
  assign n20302 = ~n4370 & n8762 ;
  assign n20303 = n20302 ^ n2052 ^ 1'b0 ;
  assign n20304 = n20303 ^ n18011 ^ n15524 ;
  assign n20305 = n20304 ^ n15065 ^ n8737 ;
  assign n20306 = ~n6616 & n12940 ;
  assign n20307 = ~n14977 & n20306 ;
  assign n20308 = n20166 ^ n16450 ^ n13017 ;
  assign n20309 = ( n8375 & ~n10139 ) | ( n8375 & n17795 ) | ( ~n10139 & n17795 ) ;
  assign n20310 = n20309 ^ n5055 ^ 1'b0 ;
  assign n20311 = ~n20308 & n20310 ;
  assign n20312 = ~n7454 & n10205 ;
  assign n20313 = n16130 ^ n2296 ^ 1'b0 ;
  assign n20314 = n20313 ^ n19500 ^ n19323 ;
  assign n20315 = n19057 ^ n10122 ^ n2459 ;
  assign n20316 = ( ~n6167 & n19267 ) | ( ~n6167 & n20315 ) | ( n19267 & n20315 ) ;
  assign n20317 = ( n10136 & ~n10725 ) | ( n10136 & n12766 ) | ( ~n10725 & n12766 ) ;
  assign n20318 = ( n10175 & n20316 ) | ( n10175 & n20317 ) | ( n20316 & n20317 ) ;
  assign n20319 = ( ~n3334 & n8821 ) | ( ~n3334 & n14511 ) | ( n8821 & n14511 ) ;
  assign n20320 = ( n13947 & ~n20318 ) | ( n13947 & n20319 ) | ( ~n20318 & n20319 ) ;
  assign n20321 = n10225 ^ n10057 ^ n3458 ;
  assign n20322 = ( x148 & ~n5296 ) | ( x148 & n20321 ) | ( ~n5296 & n20321 ) ;
  assign n20323 = ~n7169 & n20322 ;
  assign n20324 = ~n10725 & n20323 ;
  assign n20328 = n14422 ^ n1823 ^ 1'b0 ;
  assign n20325 = ~n1777 & n2385 ;
  assign n20326 = n12284 & n20325 ;
  assign n20327 = ( n14323 & ~n19515 ) | ( n14323 & n20326 ) | ( ~n19515 & n20326 ) ;
  assign n20329 = n20328 ^ n20327 ^ 1'b0 ;
  assign n20330 = n17944 ^ n6917 ^ n1722 ;
  assign n20331 = n12388 ^ n9339 ^ 1'b0 ;
  assign n20332 = n20002 | n20331 ;
  assign n20333 = ( n302 & n6151 ) | ( n302 & n20332 ) | ( n6151 & n20332 ) ;
  assign n20334 = ~n15079 & n20333 ;
  assign n20335 = ( x3 & n999 ) | ( x3 & ~n1306 ) | ( n999 & ~n1306 ) ;
  assign n20336 = n20335 ^ n17967 ^ n7612 ;
  assign n20337 = n10568 ^ n9295 ^ n796 ;
  assign n20338 = n11182 ^ n10777 ^ n1747 ;
  assign n20339 = ( ~n5126 & n9088 ) | ( ~n5126 & n20338 ) | ( n9088 & n20338 ) ;
  assign n20340 = ( n1369 & ~n20337 ) | ( n1369 & n20339 ) | ( ~n20337 & n20339 ) ;
  assign n20341 = n1749 ^ n894 ^ 1'b0 ;
  assign n20342 = ( n3275 & n5866 ) | ( n3275 & n20341 ) | ( n5866 & n20341 ) ;
  assign n20343 = n15680 ^ n7337 ^ n1965 ;
  assign n20344 = n20343 ^ n5103 ^ 1'b0 ;
  assign n20345 = n19711 | n20344 ;
  assign n20348 = n13632 ^ n6603 ^ x178 ;
  assign n20349 = ( n5836 & ~n6282 ) | ( n5836 & n20348 ) | ( ~n6282 & n20348 ) ;
  assign n20346 = n9382 | n14879 ;
  assign n20347 = n3743 & n20346 ;
  assign n20350 = n20349 ^ n20347 ^ 1'b0 ;
  assign n20351 = n3253 & ~n20350 ;
  assign n20352 = n20351 ^ n5805 ^ 1'b0 ;
  assign n20353 = n13545 & ~n18390 ;
  assign n20354 = ~n1305 & n20353 ;
  assign n20355 = n20354 ^ n18042 ^ n2167 ;
  assign n20356 = ( n8953 & n11491 ) | ( n8953 & n18840 ) | ( n11491 & n18840 ) ;
  assign n20357 = ~n4208 & n15013 ;
  assign n20358 = n20356 & n20357 ;
  assign n20361 = n10380 ^ n6792 ^ n4872 ;
  assign n20362 = n20361 ^ n12904 ^ 1'b0 ;
  assign n20359 = ( n2174 & n3605 ) | ( n2174 & n18784 ) | ( n3605 & n18784 ) ;
  assign n20360 = n12012 | n20359 ;
  assign n20363 = n20362 ^ n20360 ^ n17035 ;
  assign n20364 = n8221 ^ n6975 ^ 1'b0 ;
  assign n20365 = ( n1546 & n4200 ) | ( n1546 & n18498 ) | ( n4200 & n18498 ) ;
  assign n20366 = x87 & ~n9990 ;
  assign n20367 = n1326 & ~n5138 ;
  assign n20368 = n20367 ^ n15884 ^ 1'b0 ;
  assign n20369 = n5290 ^ n3909 ^ 1'b0 ;
  assign n20370 = ~n20368 & n20369 ;
  assign n20371 = ( ~n5429 & n20366 ) | ( ~n5429 & n20370 ) | ( n20366 & n20370 ) ;
  assign n20372 = ( ~n2661 & n4134 ) | ( ~n2661 & n5472 ) | ( n4134 & n5472 ) ;
  assign n20373 = ( n1834 & n6167 ) | ( n1834 & ~n10813 ) | ( n6167 & ~n10813 ) ;
  assign n20374 = n6027 ^ n3584 ^ 1'b0 ;
  assign n20375 = ( ~n20372 & n20373 ) | ( ~n20372 & n20374 ) | ( n20373 & n20374 ) ;
  assign n20376 = n20375 ^ n18306 ^ n16011 ;
  assign n20377 = x253 & n18965 ;
  assign n20378 = ( x136 & n1619 ) | ( x136 & ~n5247 ) | ( n1619 & ~n5247 ) ;
  assign n20379 = n20378 ^ n12865 ^ n10744 ;
  assign n20380 = n20379 ^ n6102 ^ 1'b0 ;
  assign n20381 = n6082 | n20380 ;
  assign n20385 = n15207 ^ n14232 ^ n6238 ;
  assign n20382 = n3354 & n8981 ;
  assign n20383 = ~n2408 & n20382 ;
  assign n20384 = n645 & ~n20383 ;
  assign n20386 = n20385 ^ n20384 ^ 1'b0 ;
  assign n20387 = n16712 ^ n6997 ^ 1'b0 ;
  assign n20388 = n20386 & ~n20387 ;
  assign n20389 = n914 & ~n12980 ;
  assign n20390 = n5521 & n20389 ;
  assign n20391 = n3661 & ~n20390 ;
  assign n20392 = ~n6339 & n20391 ;
  assign n20393 = n19659 ^ n430 ^ 1'b0 ;
  assign n20398 = n8721 ^ n8486 ^ n904 ;
  assign n20396 = ( n2115 & n10605 ) | ( n2115 & n11359 ) | ( n10605 & n11359 ) ;
  assign n20394 = n5551 ^ n1272 ^ 1'b0 ;
  assign n20395 = ~n7476 & n20394 ;
  assign n20397 = n20396 ^ n20395 ^ n5110 ;
  assign n20399 = n20398 ^ n20397 ^ n5469 ;
  assign n20400 = n20399 ^ n3437 ^ n1733 ;
  assign n20401 = ( x161 & n6525 ) | ( x161 & ~n7237 ) | ( n6525 & ~n7237 ) ;
  assign n20402 = n20401 ^ n6039 ^ n2576 ;
  assign n20403 = ( n833 & n1030 ) | ( n833 & ~n6870 ) | ( n1030 & ~n6870 ) ;
  assign n20404 = n20402 & ~n20403 ;
  assign n20405 = ( n2054 & ~n8216 ) | ( n2054 & n17803 ) | ( ~n8216 & n17803 ) ;
  assign n20406 = ~n8670 & n20405 ;
  assign n20407 = n20406 ^ n14775 ^ 1'b0 ;
  assign n20408 = ( n9265 & ~n15273 ) | ( n9265 & n16193 ) | ( ~n15273 & n16193 ) ;
  assign n20409 = n3294 & n5413 ;
  assign n20410 = n20409 ^ n2385 ^ 1'b0 ;
  assign n20411 = ( ~n3151 & n7309 ) | ( ~n3151 & n20410 ) | ( n7309 & n20410 ) ;
  assign n20422 = n9706 ^ n4627 ^ n2225 ;
  assign n20418 = ( n1549 & n3477 ) | ( n1549 & ~n17472 ) | ( n3477 & ~n17472 ) ;
  assign n20419 = n4161 & n14252 ;
  assign n20420 = ( n19089 & n20418 ) | ( n19089 & ~n20419 ) | ( n20418 & ~n20419 ) ;
  assign n20421 = n20420 ^ n18067 ^ 1'b0 ;
  assign n20415 = n9514 | n10682 ;
  assign n20416 = n5335 | n20415 ;
  assign n20413 = ( n7943 & n13339 ) | ( n7943 & ~n17749 ) | ( n13339 & ~n17749 ) ;
  assign n20414 = ( n5218 & n14546 ) | ( n5218 & n20413 ) | ( n14546 & n20413 ) ;
  assign n20412 = n18843 & n19262 ;
  assign n20417 = n20416 ^ n20414 ^ n20412 ;
  assign n20423 = n20422 ^ n20421 ^ n20417 ;
  assign n20424 = n8658 ^ n797 ^ 1'b0 ;
  assign n20425 = ~n10368 & n20424 ;
  assign n20426 = n19424 ^ n13462 ^ n12838 ;
  assign n20427 = ( n3517 & n5383 ) | ( n3517 & ~n20426 ) | ( n5383 & ~n20426 ) ;
  assign n20428 = ( n11387 & n16709 ) | ( n11387 & n20427 ) | ( n16709 & n20427 ) ;
  assign n20429 = n1754 & n8964 ;
  assign n20430 = n7570 ^ n4843 ^ 1'b0 ;
  assign n20431 = ( n3229 & n7418 ) | ( n3229 & ~n20430 ) | ( n7418 & ~n20430 ) ;
  assign n20432 = ( n7731 & n20429 ) | ( n7731 & ~n20431 ) | ( n20429 & ~n20431 ) ;
  assign n20438 = n16830 ^ n8884 ^ n8197 ;
  assign n20437 = ( n8804 & n15492 ) | ( n8804 & ~n17646 ) | ( n15492 & ~n17646 ) ;
  assign n20434 = ( ~n1208 & n2265 ) | ( ~n1208 & n11427 ) | ( n2265 & n11427 ) ;
  assign n20433 = ~n10728 & n12492 ;
  assign n20435 = n20434 ^ n20433 ^ 1'b0 ;
  assign n20436 = ( n1194 & n6337 ) | ( n1194 & n20435 ) | ( n6337 & n20435 ) ;
  assign n20439 = n20438 ^ n20437 ^ n20436 ;
  assign n20442 = n7984 & n19256 ;
  assign n20443 = n20442 ^ n4844 ^ 1'b0 ;
  assign n20440 = n1022 & n1410 ;
  assign n20441 = n20440 ^ n5613 ^ 1'b0 ;
  assign n20444 = n20443 ^ n20441 ^ 1'b0 ;
  assign n20445 = ( n3512 & n5838 ) | ( n3512 & ~n9803 ) | ( n5838 & ~n9803 ) ;
  assign n20446 = ( n14237 & n14589 ) | ( n14237 & ~n20445 ) | ( n14589 & ~n20445 ) ;
  assign n20450 = n14279 ^ n12745 ^ n10141 ;
  assign n20447 = n2784 & n5810 ;
  assign n20448 = n20447 ^ n4481 ^ x15 ;
  assign n20449 = n20448 ^ n14572 ^ n7688 ;
  assign n20451 = n20450 ^ n20449 ^ n2414 ;
  assign n20452 = ( ~n872 & n3728 ) | ( ~n872 & n8678 ) | ( n3728 & n8678 ) ;
  assign n20453 = ( n439 & n3715 ) | ( n439 & ~n15284 ) | ( n3715 & ~n15284 ) ;
  assign n20454 = n20453 ^ n9186 ^ n622 ;
  assign n20455 = n8440 ^ n8116 ^ 1'b0 ;
  assign n20456 = ( ~n8286 & n14503 ) | ( ~n8286 & n20455 ) | ( n14503 & n20455 ) ;
  assign n20460 = n1667 & n8876 ;
  assign n20457 = n7315 & ~n20141 ;
  assign n20458 = n9499 & n20457 ;
  assign n20459 = n20458 ^ n19165 ^ n950 ;
  assign n20461 = n20460 ^ n20459 ^ n9793 ;
  assign n20462 = n18475 ^ n17629 ^ n15734 ;
  assign n20463 = n5696 | n20462 ;
  assign n20464 = ( n14422 & ~n14578 ) | ( n14422 & n16280 ) | ( ~n14578 & n16280 ) ;
  assign n20465 = ( ~n15521 & n18817 ) | ( ~n15521 & n20464 ) | ( n18817 & n20464 ) ;
  assign n20466 = ( n3745 & n7175 ) | ( n3745 & n11041 ) | ( n7175 & n11041 ) ;
  assign n20468 = n9755 ^ n3495 ^ 1'b0 ;
  assign n20469 = n1290 & n20468 ;
  assign n20467 = n6238 | n8325 ;
  assign n20470 = n20469 ^ n20467 ^ n15918 ;
  assign n20471 = n6520 & n12916 ;
  assign n20472 = n13264 & n20471 ;
  assign n20476 = x50 & n5528 ;
  assign n20477 = n20476 ^ n14833 ^ 1'b0 ;
  assign n20478 = ~n2356 & n20477 ;
  assign n20479 = n1044 & n20478 ;
  assign n20473 = ( n1935 & n1953 ) | ( n1935 & ~n13994 ) | ( n1953 & ~n13994 ) ;
  assign n20474 = ( n891 & n7567 ) | ( n891 & ~n20473 ) | ( n7567 & ~n20473 ) ;
  assign n20475 = ( ~n4974 & n8588 ) | ( ~n4974 & n20474 ) | ( n8588 & n20474 ) ;
  assign n20480 = n20479 ^ n20475 ^ n11779 ;
  assign n20481 = n9244 ^ n9016 ^ n1324 ;
  assign n20482 = n10176 & ~n11302 ;
  assign n20483 = n20482 ^ n9183 ^ 1'b0 ;
  assign n20484 = n15195 ^ n4093 ^ n2699 ;
  assign n20485 = n10971 | n15031 ;
  assign n20486 = n20484 | n20485 ;
  assign n20487 = ~x39 & n5732 ;
  assign n20488 = ~n737 & n3795 ;
  assign n20489 = n20488 ^ n13627 ^ 1'b0 ;
  assign n20490 = n8352 ^ n4920 ^ 1'b0 ;
  assign n20491 = ~n14538 & n20490 ;
  assign n20492 = ( ~n2826 & n20489 ) | ( ~n2826 & n20491 ) | ( n20489 & n20491 ) ;
  assign n20493 = ( n10269 & ~n16215 ) | ( n10269 & n20492 ) | ( ~n16215 & n20492 ) ;
  assign n20494 = ( n11189 & n20487 ) | ( n11189 & ~n20493 ) | ( n20487 & ~n20493 ) ;
  assign n20495 = ( ~n5052 & n12489 ) | ( ~n5052 & n18328 ) | ( n12489 & n18328 ) ;
  assign n20496 = n2441 | n14351 ;
  assign n20497 = n259 | n20496 ;
  assign n20498 = ( ~n2963 & n5132 ) | ( ~n2963 & n5406 ) | ( n5132 & n5406 ) ;
  assign n20499 = n20498 ^ n17675 ^ n13940 ;
  assign n20500 = n5178 ^ x126 ^ 1'b0 ;
  assign n20501 = n2263 | n20500 ;
  assign n20502 = ( n18716 & n20499 ) | ( n18716 & ~n20501 ) | ( n20499 & ~n20501 ) ;
  assign n20503 = n17056 ^ n14352 ^ n6090 ;
  assign n20504 = ~n426 & n3395 ;
  assign n20507 = ( n5146 & ~n10386 ) | ( n5146 & n12390 ) | ( ~n10386 & n12390 ) ;
  assign n20508 = ( n3298 & ~n4401 ) | ( n3298 & n20507 ) | ( ~n4401 & n20507 ) ;
  assign n20506 = n1891 & n5948 ;
  assign n20505 = n16995 ^ n7683 ^ 1'b0 ;
  assign n20509 = n20508 ^ n20506 ^ n20505 ;
  assign n20510 = n14064 ^ n535 ^ 1'b0 ;
  assign n20511 = ( n3154 & n3990 ) | ( n3154 & ~n7089 ) | ( n3990 & ~n7089 ) ;
  assign n20512 = ~n11876 & n20511 ;
  assign n20513 = n20512 ^ n16957 ^ 1'b0 ;
  assign n20514 = ~n20510 & n20513 ;
  assign n20515 = n3157 ^ n2000 ^ n986 ;
  assign n20516 = n15592 ^ n13233 ^ n3906 ;
  assign n20517 = ( n10161 & n20515 ) | ( n10161 & n20516 ) | ( n20515 & n20516 ) ;
  assign n20518 = n20517 ^ n9025 ^ n7277 ;
  assign n20519 = n19532 ^ n1015 ^ 1'b0 ;
  assign n20520 = ( n9641 & n10072 ) | ( n9641 & n20519 ) | ( n10072 & n20519 ) ;
  assign n20521 = n20520 ^ n19449 ^ n12183 ;
  assign n20522 = n4292 ^ n885 ^ 1'b0 ;
  assign n20523 = n8933 | n20522 ;
  assign n20524 = n16533 & ~n20523 ;
  assign n20525 = ( n14790 & n18893 ) | ( n14790 & ~n20524 ) | ( n18893 & ~n20524 ) ;
  assign n20526 = ( ~n1549 & n2318 ) | ( ~n1549 & n5368 ) | ( n2318 & n5368 ) ;
  assign n20527 = n3702 & n20526 ;
  assign n20528 = n20527 ^ n8525 ^ n1075 ;
  assign n20529 = n11481 ^ n891 ^ 1'b0 ;
  assign n20530 = n15055 ^ n5975 ^ n1440 ;
  assign n20531 = n20529 | n20530 ;
  assign n20532 = n20528 & ~n20531 ;
  assign n20533 = ( ~n849 & n15741 ) | ( ~n849 & n19037 ) | ( n15741 & n19037 ) ;
  assign n20534 = n20533 ^ n15399 ^ n11386 ;
  assign n20535 = n20534 ^ n10015 ^ n5307 ;
  assign n20536 = n19863 ^ n5938 ^ 1'b0 ;
  assign n20537 = n6874 & n20536 ;
  assign n20538 = n15220 ^ n4407 ^ n2677 ;
  assign n20539 = n2589 ^ n851 ^ n334 ;
  assign n20540 = n20539 ^ n15256 ^ n7873 ;
  assign n20541 = ( n1848 & n20538 ) | ( n1848 & ~n20540 ) | ( n20538 & ~n20540 ) ;
  assign n20542 = n18292 ^ n3526 ^ 1'b0 ;
  assign n20543 = n7341 & ~n20542 ;
  assign n20549 = n9371 | n13649 ;
  assign n20550 = n20549 ^ n2000 ^ 1'b0 ;
  assign n20551 = n14113 & ~n20550 ;
  assign n20552 = n20551 ^ n14734 ^ 1'b0 ;
  assign n20548 = ( n10029 & ~n11409 ) | ( n10029 & n12807 ) | ( ~n11409 & n12807 ) ;
  assign n20544 = n10264 ^ n5761 ^ n3500 ;
  assign n20545 = ( n4712 & n11395 ) | ( n4712 & ~n20544 ) | ( n11395 & ~n20544 ) ;
  assign n20546 = n16091 ^ n11918 ^ 1'b0 ;
  assign n20547 = ( n5828 & n20545 ) | ( n5828 & n20546 ) | ( n20545 & n20546 ) ;
  assign n20553 = n20552 ^ n20548 ^ n20547 ;
  assign n20554 = n9672 & ~n16398 ;
  assign n20559 = n11429 ^ n11105 ^ n9318 ;
  assign n20556 = n5024 ^ n4719 ^ x247 ;
  assign n20557 = n20556 ^ n15409 ^ 1'b0 ;
  assign n20558 = ( n5618 & ~n9545 ) | ( n5618 & n20557 ) | ( ~n9545 & n20557 ) ;
  assign n20555 = ( n5683 & n15770 ) | ( n5683 & ~n18671 ) | ( n15770 & ~n18671 ) ;
  assign n20560 = n20559 ^ n20558 ^ n20555 ;
  assign n20561 = n17931 | n19461 ;
  assign n20562 = ( n1226 & n8789 ) | ( n1226 & n18609 ) | ( n8789 & n18609 ) ;
  assign n20563 = n12135 & n20562 ;
  assign n20564 = n20563 ^ n12831 ^ 1'b0 ;
  assign n20565 = ~n3796 & n9432 ;
  assign n20566 = ~n4295 & n20565 ;
  assign n20567 = n611 & ~n2022 ;
  assign n20568 = n20567 ^ n13198 ^ 1'b0 ;
  assign n20569 = n5898 ^ n1305 ^ n766 ;
  assign n20570 = n20569 ^ n8906 ^ 1'b0 ;
  assign n20571 = n4165 | n4898 ;
  assign n20576 = n7786 ^ n3731 ^ 1'b0 ;
  assign n20577 = n20576 ^ n18667 ^ 1'b0 ;
  assign n20572 = ( ~n1784 & n10301 ) | ( ~n1784 & n14506 ) | ( n10301 & n14506 ) ;
  assign n20573 = ( n714 & n2162 ) | ( n714 & ~n19392 ) | ( n2162 & ~n19392 ) ;
  assign n20574 = n20573 ^ n2510 ^ 1'b0 ;
  assign n20575 = n20572 & n20574 ;
  assign n20578 = n20577 ^ n20575 ^ 1'b0 ;
  assign n20579 = n1553 | n6579 ;
  assign n20583 = ( ~n383 & n1930 ) | ( ~n383 & n3578 ) | ( n1930 & n3578 ) ;
  assign n20580 = n6122 ^ n267 ^ 1'b0 ;
  assign n20581 = n14041 & n20580 ;
  assign n20582 = n20581 ^ n13812 ^ 1'b0 ;
  assign n20584 = n20583 ^ n20582 ^ n482 ;
  assign n20585 = n5734 ^ n3235 ^ x58 ;
  assign n20586 = ( n5139 & ~n10214 ) | ( n5139 & n20585 ) | ( ~n10214 & n20585 ) ;
  assign n20587 = n11044 & ~n20586 ;
  assign n20588 = n19259 ^ n9034 ^ n4512 ;
  assign n20591 = n3193 & n13136 ;
  assign n20592 = ( ~n5264 & n7750 ) | ( ~n5264 & n20591 ) | ( n7750 & n20591 ) ;
  assign n20593 = n9766 & ~n20592 ;
  assign n20589 = n13507 ^ n2456 ^ 1'b0 ;
  assign n20590 = n19243 & ~n20589 ;
  assign n20594 = n20593 ^ n20590 ^ n14331 ;
  assign n20595 = n20594 ^ n2952 ^ 1'b0 ;
  assign n20596 = n5844 & ~n20595 ;
  assign n20597 = n4072 ^ n3469 ^ n614 ;
  assign n20598 = n20597 ^ n14584 ^ 1'b0 ;
  assign n20599 = n14635 & n20598 ;
  assign n20600 = n20445 ^ n18731 ^ n16520 ;
  assign n20601 = n17260 ^ n7019 ^ 1'b0 ;
  assign n20602 = n8175 & n20601 ;
  assign n20603 = ( n3923 & n13358 ) | ( n3923 & n20602 ) | ( n13358 & n20602 ) ;
  assign n20604 = ( x61 & n9347 ) | ( x61 & ~n20603 ) | ( n9347 & ~n20603 ) ;
  assign n20605 = n5159 ^ n535 ^ n487 ;
  assign n20606 = n17432 & n19818 ;
  assign n20607 = n10926 & n20606 ;
  assign n20608 = ( n8491 & n10649 ) | ( n8491 & ~n14078 ) | ( n10649 & ~n14078 ) ;
  assign n20609 = n20608 ^ n11666 ^ n7107 ;
  assign n20610 = n20607 | n20609 ;
  assign n20611 = ( ~n3569 & n11189 ) | ( ~n3569 & n11392 ) | ( n11189 & n11392 ) ;
  assign n20612 = n20611 ^ n15403 ^ n2637 ;
  assign n20613 = ( n1092 & n8206 ) | ( n1092 & n16922 ) | ( n8206 & n16922 ) ;
  assign n20614 = ( n2152 & n20510 ) | ( n2152 & ~n20613 ) | ( n20510 & ~n20613 ) ;
  assign n20616 = ( n2302 & n4099 ) | ( n2302 & n7293 ) | ( n4099 & n7293 ) ;
  assign n20615 = n6240 ^ n5355 ^ n568 ;
  assign n20617 = n20616 ^ n20615 ^ n12426 ;
  assign n20618 = ( n426 & n10668 ) | ( n426 & ~n20617 ) | ( n10668 & ~n20617 ) ;
  assign n20619 = n6539 ^ n1829 ^ n334 ;
  assign n20620 = x166 & ~n20619 ;
  assign n20621 = n6192 ^ n4059 ^ n2395 ;
  assign n20623 = n19822 ^ n8238 ^ n6886 ;
  assign n20622 = n11888 ^ n10624 ^ n1870 ;
  assign n20624 = n20623 ^ n20622 ^ n12439 ;
  assign n20625 = n20621 & n20624 ;
  assign n20626 = n20620 & n20625 ;
  assign n20627 = n20626 ^ n20615 ^ n1518 ;
  assign n20631 = n1199 | n1344 ;
  assign n20632 = n20631 ^ n3892 ^ 1'b0 ;
  assign n20628 = n14671 ^ n4677 ^ n2978 ;
  assign n20629 = ( n1477 & ~n11888 ) | ( n1477 & n20628 ) | ( ~n11888 & n20628 ) ;
  assign n20630 = n20629 ^ n20190 ^ n18116 ;
  assign n20633 = n20632 ^ n20630 ^ 1'b0 ;
  assign n20634 = n16099 | n20633 ;
  assign n20635 = n13894 ^ n11679 ^ n6715 ;
  assign n20636 = x25 & n6240 ;
  assign n20637 = n14913 & n20636 ;
  assign n20638 = n20637 ^ n12752 ^ n7181 ;
  assign n20639 = ( ~n7560 & n10993 ) | ( ~n7560 & n20638 ) | ( n10993 & n20638 ) ;
  assign n20640 = ( n10606 & n19936 ) | ( n10606 & ~n20639 ) | ( n19936 & ~n20639 ) ;
  assign n20641 = ( ~n20246 & n20635 ) | ( ~n20246 & n20640 ) | ( n20635 & n20640 ) ;
  assign n20642 = n15141 ^ n11962 ^ n3524 ;
  assign n20643 = n20642 ^ n14412 ^ 1'b0 ;
  assign n20644 = n17392 & ~n20643 ;
  assign n20645 = n20644 ^ n4970 ^ 1'b0 ;
  assign n20646 = n20645 ^ n14385 ^ 1'b0 ;
  assign n20647 = n19180 ^ n2376 ^ n431 ;
  assign n20648 = n20647 ^ n15138 ^ n7984 ;
  assign n20649 = n14025 ^ n5394 ^ n1736 ;
  assign n20650 = n20649 ^ n7510 ^ n277 ;
  assign n20651 = n3998 | n20650 ;
  assign n20652 = ~n551 & n14665 ;
  assign n20653 = n9094 & n20652 ;
  assign n20654 = n14759 ^ n8075 ^ 1'b0 ;
  assign n20655 = ~n1074 & n20654 ;
  assign n20656 = n14503 & n20655 ;
  assign n20657 = n17485 ^ n16515 ^ n14576 ;
  assign n20658 = n15055 ^ n10936 ^ n4993 ;
  assign n20659 = ( n5101 & n19838 ) | ( n5101 & n20658 ) | ( n19838 & n20658 ) ;
  assign n20660 = ( n992 & n5793 ) | ( n992 & ~n7067 ) | ( n5793 & ~n7067 ) ;
  assign n20661 = ( ~n1216 & n4164 ) | ( ~n1216 & n10241 ) | ( n4164 & n10241 ) ;
  assign n20662 = ( n9481 & ~n20660 ) | ( n9481 & n20661 ) | ( ~n20660 & n20661 ) ;
  assign n20663 = n7133 ^ n4795 ^ 1'b0 ;
  assign n20664 = n12995 ^ n12286 ^ n7716 ;
  assign n20665 = n15941 & n20664 ;
  assign n20666 = n8881 ^ n4376 ^ x19 ;
  assign n20667 = ~n8269 & n20666 ;
  assign n20668 = n20667 ^ n4910 ^ 1'b0 ;
  assign n20669 = ( n3945 & ~n9937 ) | ( n3945 & n20668 ) | ( ~n9937 & n20668 ) ;
  assign n20670 = ( ~n7791 & n20665 ) | ( ~n7791 & n20669 ) | ( n20665 & n20669 ) ;
  assign n20671 = ( n8925 & ~n11564 ) | ( n8925 & n20670 ) | ( ~n11564 & n20670 ) ;
  assign n20672 = n16598 ^ n14111 ^ n10300 ;
  assign n20673 = n20672 ^ n20004 ^ n16381 ;
  assign n20675 = n10946 ^ n9604 ^ n6439 ;
  assign n20676 = ~n956 & n20675 ;
  assign n20677 = n20676 ^ n17301 ^ 1'b0 ;
  assign n20674 = n16658 ^ n748 ^ 1'b0 ;
  assign n20678 = n20677 ^ n20674 ^ 1'b0 ;
  assign n20679 = ( n3189 & n4085 ) | ( n3189 & n20678 ) | ( n4085 & n20678 ) ;
  assign n20680 = n18982 ^ n10747 ^ n798 ;
  assign n20681 = n17250 ^ n923 ^ 1'b0 ;
  assign n20682 = ~n5142 & n5734 ;
  assign n20683 = n20682 ^ n5034 ^ n2725 ;
  assign n20684 = n20683 ^ n16416 ^ n7309 ;
  assign n20685 = n7667 ^ n1939 ^ 1'b0 ;
  assign n20686 = ~n20684 & n20685 ;
  assign n20692 = ( n604 & n2201 ) | ( n604 & ~n10449 ) | ( n2201 & ~n10449 ) ;
  assign n20687 = ( ~n4543 & n6487 ) | ( ~n4543 & n16486 ) | ( n6487 & n16486 ) ;
  assign n20688 = n20687 ^ n11877 ^ n1937 ;
  assign n20689 = ( n544 & n7124 ) | ( n544 & n8088 ) | ( n7124 & n8088 ) ;
  assign n20690 = n20689 ^ n5547 ^ 1'b0 ;
  assign n20691 = ~n20688 & n20690 ;
  assign n20693 = n20692 ^ n20691 ^ n18086 ;
  assign n20694 = ( x13 & ~n345 ) | ( x13 & n970 ) | ( ~n345 & n970 ) ;
  assign n20695 = n6468 & ~n10664 ;
  assign n20696 = n20695 ^ n11197 ^ 1'b0 ;
  assign n20697 = x211 & n20696 ;
  assign n20698 = n13983 & n20697 ;
  assign n20699 = n8575 ^ n7285 ^ n7070 ;
  assign n20700 = ( ~n3568 & n4335 ) | ( ~n3568 & n20699 ) | ( n4335 & n20699 ) ;
  assign n20701 = n18761 ^ n13127 ^ n12544 ;
  assign n20706 = n14034 ^ n13757 ^ 1'b0 ;
  assign n20707 = n371 & ~n20706 ;
  assign n20703 = ~n1690 & n16355 ;
  assign n20704 = n20292 & n20703 ;
  assign n20702 = n8283 & ~n15766 ;
  assign n20705 = n20704 ^ n20702 ^ 1'b0 ;
  assign n20708 = n20707 ^ n20705 ^ n10226 ;
  assign n20709 = n20708 ^ n18113 ^ 1'b0 ;
  assign n20710 = n414 & ~n3574 ;
  assign n20711 = ( n822 & n16093 ) | ( n822 & ~n20710 ) | ( n16093 & ~n20710 ) ;
  assign n20712 = ~n7450 & n20711 ;
  assign n20713 = ~n9226 & n20712 ;
  assign n20714 = ( n3851 & n13548 ) | ( n3851 & n20713 ) | ( n13548 & n20713 ) ;
  assign n20715 = ( n1193 & n13702 ) | ( n1193 & ~n19002 ) | ( n13702 & ~n19002 ) ;
  assign n20716 = ( ~n439 & n19088 ) | ( ~n439 & n20715 ) | ( n19088 & n20715 ) ;
  assign n20717 = n3027 | n5108 ;
  assign n20718 = n20717 ^ x176 ^ 1'b0 ;
  assign n20719 = n20718 ^ n15545 ^ 1'b0 ;
  assign n20720 = n8557 & n20719 ;
  assign n20721 = n14041 & ~n18114 ;
  assign n20722 = ( n9758 & ~n12221 ) | ( n9758 & n20721 ) | ( ~n12221 & n20721 ) ;
  assign n20723 = n20722 ^ n4298 ^ 1'b0 ;
  assign n20724 = n19795 ^ n14958 ^ n5645 ;
  assign n20725 = ( ~n14510 & n20723 ) | ( ~n14510 & n20724 ) | ( n20723 & n20724 ) ;
  assign n20731 = n19710 ^ n16745 ^ n13847 ;
  assign n20726 = ( n851 & n10521 ) | ( n851 & n14221 ) | ( n10521 & n14221 ) ;
  assign n20727 = n1921 & ~n3309 ;
  assign n20728 = ( n9100 & ~n20726 ) | ( n9100 & n20727 ) | ( ~n20726 & n20727 ) ;
  assign n20729 = n590 & n20728 ;
  assign n20730 = n11935 & n20729 ;
  assign n20732 = n20731 ^ n20730 ^ n647 ;
  assign n20733 = n20732 ^ n15889 ^ n4427 ;
  assign n20734 = ( n12844 & ~n14546 ) | ( n12844 & n20733 ) | ( ~n14546 & n20733 ) ;
  assign n20739 = ( n3705 & n7111 ) | ( n3705 & n8709 ) | ( n7111 & n8709 ) ;
  assign n20735 = n12045 ^ n3857 ^ 1'b0 ;
  assign n20736 = n6862 & n12920 ;
  assign n20737 = n20735 & n20736 ;
  assign n20738 = n5568 | n20737 ;
  assign n20740 = n20739 ^ n20738 ^ 1'b0 ;
  assign n20743 = n7370 ^ n2755 ^ x178 ;
  assign n20741 = ( n1257 & ~n2884 ) | ( n1257 & n10583 ) | ( ~n2884 & n10583 ) ;
  assign n20742 = n14614 & n20741 ;
  assign n20744 = n20743 ^ n20742 ^ n4414 ;
  assign n20745 = n4169 | n20744 ;
  assign n20746 = ( ~n678 & n1837 ) | ( ~n678 & n2850 ) | ( n1837 & n2850 ) ;
  assign n20747 = ( ~n1703 & n9268 ) | ( ~n1703 & n12488 ) | ( n9268 & n12488 ) ;
  assign n20748 = n20747 ^ n4140 ^ 1'b0 ;
  assign n20749 = ( n16436 & n20746 ) | ( n16436 & ~n20748 ) | ( n20746 & ~n20748 ) ;
  assign n20750 = n11688 ^ n3990 ^ n1814 ;
  assign n20751 = n20750 ^ n7128 ^ n579 ;
  assign n20752 = ( n3712 & n5247 ) | ( n3712 & ~n6378 ) | ( n5247 & ~n6378 ) ;
  assign n20753 = ( n8748 & n11305 ) | ( n8748 & ~n16093 ) | ( n11305 & ~n16093 ) ;
  assign n20756 = n4991 & ~n15376 ;
  assign n20757 = n20756 ^ n2949 ^ 1'b0 ;
  assign n20758 = ~n19182 & n20757 ;
  assign n20754 = n389 & ~n1044 ;
  assign n20755 = ( n2596 & n7906 ) | ( n2596 & n20754 ) | ( n7906 & n20754 ) ;
  assign n20759 = n20758 ^ n20755 ^ n4652 ;
  assign n20760 = ( n20752 & ~n20753 ) | ( n20752 & n20759 ) | ( ~n20753 & n20759 ) ;
  assign n20764 = ( n5886 & ~n5910 ) | ( n5886 & n8837 ) | ( ~n5910 & n8837 ) ;
  assign n20761 = ( n551 & n2218 ) | ( n551 & n7196 ) | ( n2218 & n7196 ) ;
  assign n20762 = n7775 & n20761 ;
  assign n20763 = n20762 ^ n11152 ^ n6890 ;
  assign n20765 = n20764 ^ n20763 ^ 1'b0 ;
  assign n20766 = n6855 & ~n20765 ;
  assign n20767 = n10396 ^ n2751 ^ n1439 ;
  assign n20768 = n20767 ^ n8272 ^ n3061 ;
  assign n20769 = n10300 ^ n577 ^ 1'b0 ;
  assign n20770 = ~n20768 & n20769 ;
  assign n20771 = n10065 | n18156 ;
  assign n20772 = n20771 ^ n5693 ^ 1'b0 ;
  assign n20773 = n19670 ^ n10735 ^ n4110 ;
  assign n20774 = ( n3308 & ~n20772 ) | ( n3308 & n20773 ) | ( ~n20772 & n20773 ) ;
  assign n20775 = n9850 ^ n5127 ^ 1'b0 ;
  assign n20776 = ~n8899 & n20775 ;
  assign n20782 = ~n4883 & n6063 ;
  assign n20783 = n20782 ^ n20632 ^ 1'b0 ;
  assign n20784 = n20783 ^ n8384 ^ 1'b0 ;
  assign n20781 = n9885 ^ n3309 ^ 1'b0 ;
  assign n20777 = n3838 & ~n14960 ;
  assign n20778 = n20777 ^ n11128 ^ 1'b0 ;
  assign n20779 = n20778 ^ n7906 ^ n3237 ;
  assign n20780 = n20779 ^ n801 ^ 1'b0 ;
  assign n20785 = n20784 ^ n20781 ^ n20780 ;
  assign n20786 = ( ~n20352 & n20776 ) | ( ~n20352 & n20785 ) | ( n20776 & n20785 ) ;
  assign n20787 = n20341 ^ n2258 ^ x182 ;
  assign n20788 = n20787 ^ n5782 ^ n4056 ;
  assign n20789 = n20788 ^ n14455 ^ n869 ;
  assign n20790 = n15290 ^ n6102 ^ 1'b0 ;
  assign n20791 = n20789 & ~n20790 ;
  assign n20792 = n20791 ^ n6255 ^ n1576 ;
  assign n20795 = n5279 ^ n4188 ^ n2643 ;
  assign n20796 = n20795 ^ n13334 ^ n6432 ;
  assign n20793 = n10004 ^ n4690 ^ n2659 ;
  assign n20794 = ( n6374 & n12219 ) | ( n6374 & ~n20793 ) | ( n12219 & ~n20793 ) ;
  assign n20797 = n20796 ^ n20794 ^ n7809 ;
  assign n20798 = n20797 ^ n16168 ^ 1'b0 ;
  assign n20799 = n18664 ^ n6901 ^ 1'b0 ;
  assign n20800 = n528 & n20799 ;
  assign n20801 = n20800 ^ n17530 ^ 1'b0 ;
  assign n20802 = n20801 ^ n16030 ^ n8070 ;
  assign n20803 = ( n6333 & n12705 ) | ( n6333 & ~n17960 ) | ( n12705 & ~n17960 ) ;
  assign n20804 = n7444 & ~n11466 ;
  assign n20827 = n6689 ^ x46 ^ 1'b0 ;
  assign n20828 = n12219 | n20827 ;
  assign n20821 = n6819 ^ n4566 ^ 1'b0 ;
  assign n20820 = ~n15821 & n16058 ;
  assign n20822 = n20821 ^ n20820 ^ 1'b0 ;
  assign n20823 = n20822 ^ n4526 ^ 1'b0 ;
  assign n20824 = n13778 & n20823 ;
  assign n20825 = ~n17376 & n20824 ;
  assign n20826 = n20825 ^ n2667 ^ 1'b0 ;
  assign n20805 = n12619 ^ n4704 ^ n3155 ;
  assign n20806 = n9943 ^ n1090 ^ 1'b0 ;
  assign n20811 = ( ~n2671 & n8346 ) | ( ~n2671 & n10189 ) | ( n8346 & n10189 ) ;
  assign n20812 = ( n1072 & n4810 ) | ( n1072 & n8048 ) | ( n4810 & n8048 ) ;
  assign n20813 = ~n20811 & n20812 ;
  assign n20814 = ~n15399 & n20813 ;
  assign n20815 = x83 | n6631 ;
  assign n20816 = ( n4365 & ~n20814 ) | ( n4365 & n20815 ) | ( ~n20814 & n20815 ) ;
  assign n20817 = n20816 ^ n17513 ^ n690 ;
  assign n20808 = n18513 ^ n18211 ^ 1'b0 ;
  assign n20809 = n2084 & ~n20808 ;
  assign n20807 = ( n2479 & n8438 ) | ( n2479 & n15719 ) | ( n8438 & n15719 ) ;
  assign n20810 = n20809 ^ n20807 ^ n1606 ;
  assign n20818 = n20817 ^ n20810 ^ n8259 ;
  assign n20819 = ( n20805 & ~n20806 ) | ( n20805 & n20818 ) | ( ~n20806 & n20818 ) ;
  assign n20829 = n20828 ^ n20826 ^ n20819 ;
  assign n20830 = n5498 & ~n18897 ;
  assign n20831 = n20830 ^ n3605 ^ 1'b0 ;
  assign n20832 = ( n4907 & n7992 ) | ( n4907 & ~n20831 ) | ( n7992 & ~n20831 ) ;
  assign n20833 = n20832 ^ n18864 ^ n2072 ;
  assign n20834 = x104 & n20833 ;
  assign n20835 = n16451 ^ n724 ^ x63 ;
  assign n20836 = n2637 & n19472 ;
  assign n20837 = n20836 ^ n12844 ^ 1'b0 ;
  assign n20838 = n17498 ^ n10681 ^ 1'b0 ;
  assign n20839 = n6078 | n20838 ;
  assign n20841 = n2484 & n2550 ;
  assign n20840 = n18190 ^ n3050 ^ 1'b0 ;
  assign n20842 = n20841 ^ n20840 ^ n3737 ;
  assign n20843 = n13142 ^ n10508 ^ n4769 ;
  assign n20845 = n16338 ^ n8461 ^ 1'b0 ;
  assign n20844 = ~n2590 & n3698 ;
  assign n20846 = n20845 ^ n20844 ^ 1'b0 ;
  assign n20847 = n4399 & n5706 ;
  assign n20848 = ( x43 & n6681 ) | ( x43 & n11885 ) | ( n6681 & n11885 ) ;
  assign n20849 = n20848 ^ n16585 ^ n2058 ;
  assign n20851 = ( n5591 & n8097 ) | ( n5591 & ~n13099 ) | ( n8097 & ~n13099 ) ;
  assign n20850 = n17217 ^ n8422 ^ n2821 ;
  assign n20852 = n20851 ^ n20850 ^ n4037 ;
  assign n20853 = n14213 ^ n10523 ^ 1'b0 ;
  assign n20854 = ~n3286 & n16681 ;
  assign n20855 = n20853 & n20854 ;
  assign n20856 = ( n20849 & n20852 ) | ( n20849 & n20855 ) | ( n20852 & n20855 ) ;
  assign n20865 = ( ~n6018 & n9557 ) | ( ~n6018 & n14376 ) | ( n9557 & n14376 ) ;
  assign n20860 = ( n1067 & ~n3397 ) | ( n1067 & n7417 ) | ( ~n3397 & n7417 ) ;
  assign n20861 = n20860 ^ n7180 ^ n2251 ;
  assign n20862 = n20861 ^ n4305 ^ 1'b0 ;
  assign n20863 = ( n2209 & n5984 ) | ( n2209 & ~n20862 ) | ( n5984 & ~n20862 ) ;
  assign n20857 = n10502 ^ n4336 ^ 1'b0 ;
  assign n20858 = n20857 ^ n20418 ^ n14434 ;
  assign n20859 = n3573 & n20858 ;
  assign n20864 = n20863 ^ n20859 ^ 1'b0 ;
  assign n20866 = n20865 ^ n20864 ^ n6590 ;
  assign n20867 = n6860 & ~n11084 ;
  assign n20868 = n20867 ^ n6694 ^ 1'b0 ;
  assign n20869 = n20868 ^ n332 ^ 1'b0 ;
  assign n20871 = ~n1604 & n3628 ;
  assign n20872 = ( n1514 & ~n17243 ) | ( n1514 & n20871 ) | ( ~n17243 & n20871 ) ;
  assign n20870 = n13568 ^ n10141 ^ x166 ;
  assign n20873 = n20872 ^ n20870 ^ n7588 ;
  assign n20874 = n20083 ^ n16276 ^ 1'b0 ;
  assign n20875 = n14690 & n20874 ;
  assign n20876 = n10126 ^ n1067 ^ x8 ;
  assign n20877 = n971 | n20876 ;
  assign n20878 = n2127 & ~n18446 ;
  assign n20879 = n6939 & ~n20878 ;
  assign n20880 = ~n7119 & n20879 ;
  assign n20881 = n11443 ^ n8965 ^ n2246 ;
  assign n20882 = ( n1961 & n2668 ) | ( n1961 & n18442 ) | ( n2668 & n18442 ) ;
  assign n20884 = ( n283 & n5288 ) | ( n283 & n15060 ) | ( n5288 & n15060 ) ;
  assign n20883 = n16713 ^ n10652 ^ 1'b0 ;
  assign n20885 = n20884 ^ n20883 ^ 1'b0 ;
  assign n20886 = ~n15437 & n20885 ;
  assign n20887 = n13340 ^ n8301 ^ n5244 ;
  assign n20888 = n20887 ^ n12139 ^ n5408 ;
  assign n20890 = n4382 | n16948 ;
  assign n20889 = n10059 & n11176 ;
  assign n20891 = n20890 ^ n20889 ^ 1'b0 ;
  assign n20892 = n1414 ^ n479 ^ 1'b0 ;
  assign n20893 = n20892 ^ n14426 ^ n1897 ;
  assign n20894 = n20893 ^ n11804 ^ n1052 ;
  assign n20895 = ( n4579 & n6923 ) | ( n4579 & ~n20894 ) | ( n6923 & ~n20894 ) ;
  assign n20899 = n385 | n7576 ;
  assign n20900 = n20899 ^ n16600 ^ 1'b0 ;
  assign n20901 = ( n3117 & ~n19953 ) | ( n3117 & n20900 ) | ( ~n19953 & n20900 ) ;
  assign n20898 = n6177 & n7763 ;
  assign n20902 = n20901 ^ n20898 ^ n17890 ;
  assign n20896 = n11585 & n13748 ;
  assign n20897 = n20896 ^ n5084 ^ 1'b0 ;
  assign n20903 = n20902 ^ n20897 ^ 1'b0 ;
  assign n20906 = n11404 ^ n2786 ^ n2559 ;
  assign n20907 = ~n409 & n827 ;
  assign n20908 = ~n11845 & n20907 ;
  assign n20909 = ~n20906 & n20908 ;
  assign n20904 = ( n5709 & n6661 ) | ( n5709 & n7262 ) | ( n6661 & n7262 ) ;
  assign n20905 = n20904 ^ n8454 ^ n2213 ;
  assign n20910 = n20909 ^ n20905 ^ 1'b0 ;
  assign n20911 = n6926 ^ n1925 ^ n256 ;
  assign n20912 = n13210 ^ n875 ^ n316 ;
  assign n20913 = n20912 ^ n17408 ^ n1337 ;
  assign n20914 = ~n20911 & n20913 ;
  assign n20915 = n15420 ^ n5673 ^ 1'b0 ;
  assign n20916 = n20915 ^ n18336 ^ n7040 ;
  assign n20917 = ~n5429 & n10322 ;
  assign n20918 = ( n2857 & n20916 ) | ( n2857 & n20917 ) | ( n20916 & n20917 ) ;
  assign n20919 = ( n2900 & ~n9714 ) | ( n2900 & n10144 ) | ( ~n9714 & n10144 ) ;
  assign n20920 = n20919 ^ n5420 ^ x27 ;
  assign n20921 = n979 & n7706 ;
  assign n20922 = n8393 & n20921 ;
  assign n20923 = ( n5551 & n9133 ) | ( n5551 & ~n20922 ) | ( n9133 & ~n20922 ) ;
  assign n20924 = n20923 ^ n1343 ^ 1'b0 ;
  assign n20925 = n16549 & n20924 ;
  assign n20926 = n20920 & n20925 ;
  assign n20927 = ~n5976 & n20926 ;
  assign n20928 = ( ~n7570 & n11779 ) | ( ~n7570 & n13455 ) | ( n11779 & n13455 ) ;
  assign n20929 = n9760 ^ n9216 ^ 1'b0 ;
  assign n20930 = ( ~n14129 & n20928 ) | ( ~n14129 & n20929 ) | ( n20928 & n20929 ) ;
  assign n20931 = ( n2818 & n7656 ) | ( n2818 & n15642 ) | ( n7656 & n15642 ) ;
  assign n20932 = ( n6640 & ~n8111 ) | ( n6640 & n20176 ) | ( ~n8111 & n20176 ) ;
  assign n20933 = ( n12037 & n16542 ) | ( n12037 & ~n20932 ) | ( n16542 & ~n20932 ) ;
  assign n20934 = ( n15886 & n19327 ) | ( n15886 & n20933 ) | ( n19327 & n20933 ) ;
  assign n20935 = n11023 ^ n6166 ^ n4662 ;
  assign n20936 = ( n7658 & ~n10010 ) | ( n7658 & n20935 ) | ( ~n10010 & n20935 ) ;
  assign n20937 = n20936 ^ n9418 ^ 1'b0 ;
  assign n20938 = n20934 | n20937 ;
  assign n20939 = ( ~n6998 & n7202 ) | ( ~n6998 & n20862 ) | ( n7202 & n20862 ) ;
  assign n20949 = n16849 ^ n3459 ^ 1'b0 ;
  assign n20950 = n9237 & n20949 ;
  assign n20940 = ( n2931 & ~n5383 ) | ( n2931 & n19908 ) | ( ~n5383 & n19908 ) ;
  assign n20941 = ( n855 & n19800 ) | ( n855 & ~n20940 ) | ( n19800 & ~n20940 ) ;
  assign n20942 = n17242 ^ n8080 ^ n2018 ;
  assign n20943 = ( n4858 & n9972 ) | ( n4858 & ~n20942 ) | ( n9972 & ~n20942 ) ;
  assign n20944 = ( n3538 & n18557 ) | ( n3538 & n20943 ) | ( n18557 & n20943 ) ;
  assign n20945 = n20944 ^ n20697 ^ n14581 ;
  assign n20946 = ( n5418 & n20941 ) | ( n5418 & n20945 ) | ( n20941 & n20945 ) ;
  assign n20947 = n7605 & n20946 ;
  assign n20948 = n20947 ^ n8600 ^ 1'b0 ;
  assign n20951 = n20950 ^ n20948 ^ n4545 ;
  assign n20952 = n5944 ^ n4753 ^ n3956 ;
  assign n20953 = n20952 ^ n13314 ^ n9689 ;
  assign n20954 = n20953 ^ n11798 ^ n4710 ;
  assign n20959 = n14984 ^ n10345 ^ n1478 ;
  assign n20960 = n20959 ^ n6458 ^ n4918 ;
  assign n20955 = n1437 ^ n1137 ^ n1043 ;
  assign n20956 = ( ~n2478 & n12984 ) | ( ~n2478 & n20955 ) | ( n12984 & n20955 ) ;
  assign n20957 = ( n13167 & ~n16785 ) | ( n13167 & n20956 ) | ( ~n16785 & n20956 ) ;
  assign n20958 = n20957 ^ n3603 ^ n2231 ;
  assign n20961 = n20960 ^ n20958 ^ n17530 ;
  assign n20962 = n5770 | n20961 ;
  assign n20965 = ( n1555 & n2330 ) | ( n1555 & n3950 ) | ( n2330 & n3950 ) ;
  assign n20963 = n5442 ^ n2833 ^ x20 ;
  assign n20964 = ~n15355 & n20963 ;
  assign n20966 = n20965 ^ n20964 ^ 1'b0 ;
  assign n20972 = ~n3400 & n4057 ;
  assign n20971 = n15968 ^ n4407 ^ n423 ;
  assign n20973 = n20972 ^ n20971 ^ n10897 ;
  assign n20967 = n16129 ^ n9427 ^ n3418 ;
  assign n20968 = n20967 ^ n2152 ^ 1'b0 ;
  assign n20969 = n20968 ^ n2248 ^ 1'b0 ;
  assign n20970 = ~n4489 & n20969 ;
  assign n20974 = n20973 ^ n20970 ^ n20791 ;
  assign n20975 = ( ~n295 & n7139 ) | ( ~n295 & n14448 ) | ( n7139 & n14448 ) ;
  assign n20976 = n11531 ^ n2716 ^ 1'b0 ;
  assign n20977 = n6825 ^ n3212 ^ 1'b0 ;
  assign n20978 = n20976 | n20977 ;
  assign n20979 = ( n10197 & n12480 ) | ( n10197 & ~n20978 ) | ( n12480 & ~n20978 ) ;
  assign n20980 = n3229 | n16734 ;
  assign n20981 = n2313 | n20980 ;
  assign n20982 = n11459 & n20981 ;
  assign n20983 = ( n5614 & ~n7078 ) | ( n5614 & n18484 ) | ( ~n7078 & n18484 ) ;
  assign n20998 = n12992 ^ n9510 ^ n8225 ;
  assign n20991 = ( n1094 & ~n1804 ) | ( n1094 & n5175 ) | ( ~n1804 & n5175 ) ;
  assign n20993 = n1155 & ~n8822 ;
  assign n20994 = n20993 ^ n3293 ^ 1'b0 ;
  assign n20992 = n10477 ^ n2313 ^ 1'b0 ;
  assign n20995 = n20994 ^ n20992 ^ n5408 ;
  assign n20996 = ( ~n1224 & n20991 ) | ( ~n1224 & n20995 ) | ( n20991 & n20995 ) ;
  assign n20989 = ( n2442 & ~n7611 ) | ( n2442 & n20922 ) | ( ~n7611 & n20922 ) ;
  assign n20984 = n9455 & n17003 ;
  assign n20985 = ~n756 & n6134 ;
  assign n20986 = ( n2786 & ~n6036 ) | ( n2786 & n20985 ) | ( ~n6036 & n20985 ) ;
  assign n20987 = n20984 | n20986 ;
  assign n20988 = ( n3264 & ~n10698 ) | ( n3264 & n20987 ) | ( ~n10698 & n20987 ) ;
  assign n20990 = n20989 ^ n20988 ^ n16338 ;
  assign n20997 = n20996 ^ n20990 ^ n8720 ;
  assign n20999 = n20998 ^ n20997 ^ 1'b0 ;
  assign n21000 = ~n20983 & n20999 ;
  assign n21001 = n12662 ^ n7786 ^ 1'b0 ;
  assign n21002 = n11405 & n21001 ;
  assign n21003 = n21002 ^ n18541 ^ n13192 ;
  assign n21004 = n21003 ^ n7248 ^ 1'b0 ;
  assign n21005 = ( n3820 & n5016 ) | ( n3820 & n11338 ) | ( n5016 & n11338 ) ;
  assign n21006 = ( n1126 & n1216 ) | ( n1126 & n6870 ) | ( n1216 & n6870 ) ;
  assign n21007 = n21006 ^ n7224 ^ n4062 ;
  assign n21008 = n21007 ^ n6119 ^ n2759 ;
  assign n21009 = n9326 | n9808 ;
  assign n21010 = ( n21005 & n21008 ) | ( n21005 & ~n21009 ) | ( n21008 & ~n21009 ) ;
  assign n21011 = n21010 ^ n6301 ^ n3687 ;
  assign n21012 = ( n6209 & n8345 ) | ( n6209 & ~n11846 ) | ( n8345 & ~n11846 ) ;
  assign n21013 = n21012 ^ n18065 ^ n17813 ;
  assign n21014 = n16819 ^ n9184 ^ n5157 ;
  assign n21015 = n21014 ^ n11594 ^ n8886 ;
  assign n21016 = n4057 ^ n2448 ^ n1791 ;
  assign n21017 = ( n1644 & n5890 ) | ( n1644 & n21016 ) | ( n5890 & n21016 ) ;
  assign n21018 = n1699 & n6410 ;
  assign n21019 = n21018 ^ n12133 ^ 1'b0 ;
  assign n21020 = n21019 ^ n3526 ^ x222 ;
  assign n21021 = n20746 ^ n9283 ^ n4457 ;
  assign n21022 = n21021 ^ n12655 ^ 1'b0 ;
  assign n21023 = n21020 | n21022 ;
  assign n21024 = ( n2292 & ~n14182 ) | ( n2292 & n21023 ) | ( ~n14182 & n21023 ) ;
  assign n21028 = n13462 | n14258 ;
  assign n21027 = ~n7246 & n12873 ;
  assign n21025 = n5618 ^ n2394 ^ n1856 ;
  assign n21026 = n21025 ^ n6362 ^ 1'b0 ;
  assign n21029 = n21028 ^ n21027 ^ n21026 ;
  assign n21030 = n16867 ^ n12136 ^ n6319 ;
  assign n21031 = n11607 & n21030 ;
  assign n21032 = n21031 ^ n5922 ^ 1'b0 ;
  assign n21033 = n21032 ^ n19905 ^ 1'b0 ;
  assign n21034 = n2605 & n11539 ;
  assign n21035 = n21034 ^ n10029 ^ n8322 ;
  assign n21043 = n3650 & ~n4755 ;
  assign n21044 = ~n12587 & n21043 ;
  assign n21045 = n21044 ^ n13524 ^ n6500 ;
  assign n21039 = ( ~n9841 & n11413 ) | ( ~n9841 & n15758 ) | ( n11413 & n15758 ) ;
  assign n21036 = n19323 ^ n3093 ^ 1'b0 ;
  assign n21037 = n2759 | n21036 ;
  assign n21038 = n21037 ^ n18831 ^ n1756 ;
  assign n21040 = n21039 ^ n21038 ^ n440 ;
  assign n21041 = n21040 ^ n1609 ^ 1'b0 ;
  assign n21042 = ~n15038 & n21041 ;
  assign n21046 = n21045 ^ n21042 ^ n4780 ;
  assign n21047 = n2902 & ~n4457 ;
  assign n21048 = ( n2987 & n7708 ) | ( n2987 & n21047 ) | ( n7708 & n21047 ) ;
  assign n21049 = n20498 ^ n11109 ^ 1'b0 ;
  assign n21050 = n21049 ^ n2512 ^ n2126 ;
  assign n21051 = n2093 & n21050 ;
  assign n21052 = ( n3270 & ~n6432 ) | ( n3270 & n20576 ) | ( ~n6432 & n20576 ) ;
  assign n21053 = ( n9820 & ~n9904 ) | ( n9820 & n11046 ) | ( ~n9904 & n11046 ) ;
  assign n21054 = n2731 & n21053 ;
  assign n21055 = n21054 ^ n5177 ^ 1'b0 ;
  assign n21056 = n21052 & n21055 ;
  assign n21058 = n1741 ^ n567 ^ 1'b0 ;
  assign n21059 = n761 & n21058 ;
  assign n21057 = n4406 ^ n3618 ^ n555 ;
  assign n21060 = n21059 ^ n21057 ^ n11513 ;
  assign n21061 = n1961 | n12775 ;
  assign n21062 = n9684 ^ n8532 ^ n3714 ;
  assign n21063 = ( n15613 & n21061 ) | ( n15613 & ~n21062 ) | ( n21061 & ~n21062 ) ;
  assign n21064 = ( ~n5616 & n15865 ) | ( ~n5616 & n21063 ) | ( n15865 & n21063 ) ;
  assign n21065 = n14719 ^ n5457 ^ n703 ;
  assign n21066 = n21065 ^ n3056 ^ 1'b0 ;
  assign n21067 = ~n7979 & n21066 ;
  assign n21068 = n10455 ^ n6260 ^ n1278 ;
  assign n21069 = n21068 ^ n4911 ^ n2777 ;
  assign n21072 = n1122 & ~n5780 ;
  assign n21073 = n21072 ^ n7560 ^ n5887 ;
  assign n21071 = n17806 ^ n13142 ^ n711 ;
  assign n21070 = ( x235 & n11876 ) | ( x235 & ~n15371 ) | ( n11876 & ~n15371 ) ;
  assign n21074 = n21073 ^ n21071 ^ n21070 ;
  assign n21075 = n13845 ^ n7850 ^ n363 ;
  assign n21077 = ~n1173 & n4252 ;
  assign n21078 = n21077 ^ n17442 ^ 1'b0 ;
  assign n21076 = n5027 & ~n13211 ;
  assign n21079 = n21078 ^ n21076 ^ 1'b0 ;
  assign n21080 = n21079 ^ n14287 ^ n8305 ;
  assign n21082 = ~n2226 & n9655 ;
  assign n21083 = n14351 & n21082 ;
  assign n21084 = n21083 ^ n17891 ^ 1'b0 ;
  assign n21081 = n2651 ^ n1471 ^ x226 ;
  assign n21085 = n21084 ^ n21081 ^ n10522 ;
  assign n21087 = ( ~n3172 & n4459 ) | ( ~n3172 & n8521 ) | ( n4459 & n8521 ) ;
  assign n21086 = ( n1806 & n2815 ) | ( n1806 & n3493 ) | ( n2815 & n3493 ) ;
  assign n21088 = n21087 ^ n21086 ^ n4759 ;
  assign n21089 = n5166 & ~n7462 ;
  assign n21090 = n12835 ^ n4926 ^ 1'b0 ;
  assign n21091 = n8035 ^ n4272 ^ n2679 ;
  assign n21092 = ( n7192 & ~n21090 ) | ( n7192 & n21091 ) | ( ~n21090 & n21091 ) ;
  assign n21093 = ( n12620 & ~n13592 ) | ( n12620 & n21092 ) | ( ~n13592 & n21092 ) ;
  assign n21096 = ~n3512 & n6040 ;
  assign n21097 = n21096 ^ n9960 ^ 1'b0 ;
  assign n21094 = n11869 ^ n2617 ^ 1'b0 ;
  assign n21095 = ~n12673 & n21094 ;
  assign n21098 = n21097 ^ n21095 ^ n16132 ;
  assign n21099 = ~n8735 & n10037 ;
  assign n21100 = n21099 ^ n311 ^ 1'b0 ;
  assign n21101 = n13756 | n21100 ;
  assign n21102 = n7126 & ~n21101 ;
  assign n21103 = n21102 ^ n10803 ^ n6544 ;
  assign n21104 = n16650 ^ n11266 ^ n1870 ;
  assign n21105 = ( n10996 & n13007 ) | ( n10996 & n15095 ) | ( n13007 & n15095 ) ;
  assign n21106 = n16492 ^ n3759 ^ x124 ;
  assign n21107 = ( n10922 & n15891 ) | ( n10922 & n21106 ) | ( n15891 & n21106 ) ;
  assign n21108 = ( n7060 & n14657 ) | ( n7060 & ~n21107 ) | ( n14657 & ~n21107 ) ;
  assign n21109 = n17905 ^ n13420 ^ n6103 ;
  assign n21110 = n21109 ^ n9148 ^ n7883 ;
  assign n21113 = n6861 ^ n6175 ^ 1'b0 ;
  assign n21111 = ( n8260 & ~n18298 ) | ( n8260 & n18828 ) | ( ~n18298 & n18828 ) ;
  assign n21112 = ( n13236 & n18350 ) | ( n13236 & ~n21111 ) | ( n18350 & ~n21111 ) ;
  assign n21114 = n21113 ^ n21112 ^ n14148 ;
  assign n21115 = n5146 & n12157 ;
  assign n21116 = ~n2723 & n21115 ;
  assign n21117 = n583 | n1856 ;
  assign n21118 = n10444 ^ n9596 ^ n6232 ;
  assign n21126 = n10018 ^ n4375 ^ n2384 ;
  assign n21124 = n15929 ^ n5055 ^ n4198 ;
  assign n21119 = n3605 & n4625 ;
  assign n21120 = n6950 & n21119 ;
  assign n21121 = n7535 & ~n14586 ;
  assign n21122 = n15487 | n21121 ;
  assign n21123 = n21120 & ~n21122 ;
  assign n21125 = n21124 ^ n21123 ^ n1962 ;
  assign n21127 = n21126 ^ n21125 ^ n3667 ;
  assign n21131 = n8746 ^ n4413 ^ 1'b0 ;
  assign n21132 = ~n10809 & n21131 ;
  assign n21130 = n14185 ^ n11930 ^ n5831 ;
  assign n21128 = n3106 & n14295 ;
  assign n21129 = ( n3469 & n16044 ) | ( n3469 & n21128 ) | ( n16044 & n21128 ) ;
  assign n21133 = n21132 ^ n21130 ^ n21129 ;
  assign n21134 = ( n4616 & n9991 ) | ( n4616 & ~n10711 ) | ( n9991 & ~n10711 ) ;
  assign n21135 = n21134 ^ n1716 ^ x184 ;
  assign n21136 = n15420 ^ n12864 ^ n11420 ;
  assign n21137 = n21136 ^ n11221 ^ x182 ;
  assign n21138 = n10537 | n14978 ;
  assign n21139 = n21138 ^ n6424 ^ 1'b0 ;
  assign n21140 = ( n7425 & n15701 ) | ( n7425 & n21139 ) | ( n15701 & n21139 ) ;
  assign n21143 = ( n5985 & n9944 ) | ( n5985 & n11565 ) | ( n9944 & n11565 ) ;
  assign n21141 = n3345 & n15607 ;
  assign n21142 = n21141 ^ n20624 ^ n10177 ;
  assign n21144 = n21143 ^ n21142 ^ n826 ;
  assign n21145 = n6574 ^ n5663 ^ 1'b0 ;
  assign n21146 = n18513 ^ n17305 ^ n8937 ;
  assign n21147 = ( ~n7878 & n11524 ) | ( ~n7878 & n21146 ) | ( n11524 & n21146 ) ;
  assign n21148 = n21145 & ~n21147 ;
  assign n21149 = n21148 ^ n18770 ^ 1'b0 ;
  assign n21151 = ( n2688 & ~n3142 ) | ( n2688 & n5422 ) | ( ~n3142 & n5422 ) ;
  assign n21152 = ( n15960 & ~n19951 ) | ( n15960 & n21151 ) | ( ~n19951 & n21151 ) ;
  assign n21150 = n5918 ^ n5864 ^ n1419 ;
  assign n21153 = n21152 ^ n21150 ^ 1'b0 ;
  assign n21154 = n18250 ^ n14596 ^ n6964 ;
  assign n21155 = n21154 ^ n8661 ^ 1'b0 ;
  assign n21156 = n21155 ^ n20232 ^ n2025 ;
  assign n21157 = n1099 & n6599 ;
  assign n21158 = ~n13799 & n21157 ;
  assign n21159 = n21158 ^ n17458 ^ n10573 ;
  assign n21160 = x239 & ~n18044 ;
  assign n21161 = ~n1642 & n21160 ;
  assign n21162 = n21161 ^ n12543 ^ 1'b0 ;
  assign n21163 = n400 | n3305 ;
  assign n21164 = n21163 ^ n5653 ^ 1'b0 ;
  assign n21165 = n5146 ^ n1967 ^ n353 ;
  assign n21166 = ( n9172 & ~n9550 ) | ( n9172 & n21165 ) | ( ~n9550 & n21165 ) ;
  assign n21167 = n11349 ^ n10763 ^ n539 ;
  assign n21168 = n21167 ^ n16198 ^ 1'b0 ;
  assign n21169 = n21168 ^ n20421 ^ n13672 ;
  assign n21170 = n5811 & ~n16493 ;
  assign n21171 = n21170 ^ n5908 ^ 1'b0 ;
  assign n21172 = n15972 ^ n4595 ^ n4288 ;
  assign n21173 = ( n8685 & n20661 ) | ( n8685 & n21172 ) | ( n20661 & n21172 ) ;
  assign n21174 = n21173 ^ n768 ^ 1'b0 ;
  assign n21177 = n1625 & ~n8036 ;
  assign n21178 = n21177 ^ n19356 ^ n5479 ;
  assign n21175 = n7686 ^ n6327 ^ 1'b0 ;
  assign n21176 = n20849 & ~n21175 ;
  assign n21179 = n21178 ^ n21176 ^ n10833 ;
  assign n21180 = n16940 ^ n15536 ^ n10259 ;
  assign n21181 = n21180 ^ n16548 ^ 1'b0 ;
  assign n21182 = ( n5565 & n17545 ) | ( n5565 & ~n20124 ) | ( n17545 & ~n20124 ) ;
  assign n21183 = ( ~n8226 & n8263 ) | ( ~n8226 & n11836 ) | ( n8263 & n11836 ) ;
  assign n21184 = n21183 ^ n1117 ^ 1'b0 ;
  assign n21185 = ( n10170 & n19188 ) | ( n10170 & ~n20038 ) | ( n19188 & ~n20038 ) ;
  assign n21186 = n21185 ^ n14117 ^ n11417 ;
  assign n21187 = ( n910 & n3573 ) | ( n910 & n15689 ) | ( n3573 & n15689 ) ;
  assign n21190 = n4017 ^ n2167 ^ 1'b0 ;
  assign n21191 = ~n6383 & n21190 ;
  assign n21188 = n4379 ^ n3707 ^ n2048 ;
  assign n21189 = n19552 & n21188 ;
  assign n21192 = n21191 ^ n21189 ^ 1'b0 ;
  assign n21193 = ( n20130 & n21187 ) | ( n20130 & ~n21192 ) | ( n21187 & ~n21192 ) ;
  assign n21194 = n9532 & n17963 ;
  assign n21195 = ~n4265 & n21194 ;
  assign n21196 = ( n5926 & n21193 ) | ( n5926 & n21195 ) | ( n21193 & n21195 ) ;
  assign n21197 = n2495 | n14649 ;
  assign n21198 = n17946 ^ n16890 ^ n3767 ;
  assign n21199 = n1846 & n9013 ;
  assign n21200 = ~n5008 & n21199 ;
  assign n21201 = n1010 | n9623 ;
  assign n21202 = ( n8442 & n13196 ) | ( n8442 & n21201 ) | ( n13196 & n21201 ) ;
  assign n21203 = ( n14759 & n21200 ) | ( n14759 & n21202 ) | ( n21200 & n21202 ) ;
  assign n21204 = ( n892 & n12042 ) | ( n892 & ~n12384 ) | ( n12042 & ~n12384 ) ;
  assign n21205 = ( ~n9561 & n13896 ) | ( ~n9561 & n21204 ) | ( n13896 & n21204 ) ;
  assign n21206 = n4186 ^ n2004 ^ 1'b0 ;
  assign n21207 = n8561 & n21206 ;
  assign n21208 = ( n6990 & n21205 ) | ( n6990 & n21207 ) | ( n21205 & n21207 ) ;
  assign n21213 = n6766 ^ n495 ^ x143 ;
  assign n21211 = ( n408 & ~n4218 ) | ( n408 & n18924 ) | ( ~n4218 & n18924 ) ;
  assign n21209 = n6573 & n14007 ;
  assign n21210 = n21209 ^ n11046 ^ n3014 ;
  assign n21212 = n21211 ^ n21210 ^ 1'b0 ;
  assign n21214 = n21213 ^ n21212 ^ n6502 ;
  assign n21215 = n13415 ^ n5330 ^ 1'b0 ;
  assign n21216 = n21215 ^ n13159 ^ n9380 ;
  assign n21217 = n21216 ^ n19085 ^ n18593 ;
  assign n21218 = n21217 ^ n10052 ^ n7447 ;
  assign n21219 = ( n732 & n1414 ) | ( n732 & ~n7018 ) | ( n1414 & ~n7018 ) ;
  assign n21220 = n5035 & ~n21219 ;
  assign n21221 = n21220 ^ n16879 ^ 1'b0 ;
  assign n21222 = n21221 ^ n8075 ^ n1835 ;
  assign n21223 = ~n7121 & n21222 ;
  assign n21224 = n21218 & n21223 ;
  assign n21225 = n11005 ^ n4989 ^ n2383 ;
  assign n21226 = ( ~n8878 & n9450 ) | ( ~n8878 & n19800 ) | ( n9450 & n19800 ) ;
  assign n21227 = ( ~n11475 & n21225 ) | ( ~n11475 & n21226 ) | ( n21225 & n21226 ) ;
  assign n21228 = n12226 ^ n10075 ^ n3385 ;
  assign n21229 = n20664 ^ n16892 ^ n7462 ;
  assign n21230 = n21229 ^ n13573 ^ n5725 ;
  assign n21231 = n19945 ^ n2317 ^ 1'b0 ;
  assign n21236 = n521 & ~n8674 ;
  assign n21237 = ( ~n806 & n5091 ) | ( ~n806 & n21236 ) | ( n5091 & n21236 ) ;
  assign n21235 = ( n2773 & n5367 ) | ( n2773 & ~n6112 ) | ( n5367 & ~n6112 ) ;
  assign n21232 = n9237 ^ n6156 ^ n884 ;
  assign n21233 = ( ~n7393 & n16166 ) | ( ~n7393 & n21232 ) | ( n16166 & n21232 ) ;
  assign n21234 = n21233 ^ n15952 ^ n4045 ;
  assign n21238 = n21237 ^ n21235 ^ n21234 ;
  assign n21246 = n16101 ^ n11627 ^ n7547 ;
  assign n21239 = n20580 ^ n2747 ^ n2275 ;
  assign n21240 = ( n2430 & n2710 ) | ( n2430 & ~n21239 ) | ( n2710 & ~n21239 ) ;
  assign n21241 = n16498 ^ n4775 ^ n2708 ;
  assign n21242 = n12170 ^ n2952 ^ 1'b0 ;
  assign n21243 = n2895 | n21242 ;
  assign n21244 = n5558 & ~n21243 ;
  assign n21245 = ( n21240 & n21241 ) | ( n21240 & ~n21244 ) | ( n21241 & ~n21244 ) ;
  assign n21247 = n21246 ^ n21245 ^ n1558 ;
  assign n21248 = n21247 ^ n3869 ^ 1'b0 ;
  assign n21249 = n21238 & ~n21248 ;
  assign n21250 = n13209 ^ n2590 ^ 1'b0 ;
  assign n21256 = n1520 & n2364 ;
  assign n21251 = ~n12274 & n14635 ;
  assign n21252 = n21251 ^ n6716 ^ 1'b0 ;
  assign n21253 = ( n1550 & n5820 ) | ( n1550 & n21252 ) | ( n5820 & n21252 ) ;
  assign n21254 = n12786 ^ n9385 ^ n1547 ;
  assign n21255 = ( n15261 & n21253 ) | ( n15261 & n21254 ) | ( n21253 & n21254 ) ;
  assign n21257 = n21256 ^ n21255 ^ n752 ;
  assign n21258 = ( ~n3439 & n4035 ) | ( ~n3439 & n7887 ) | ( n4035 & n7887 ) ;
  assign n21259 = ( n12671 & n21257 ) | ( n12671 & n21258 ) | ( n21257 & n21258 ) ;
  assign n21260 = n20971 ^ n9025 ^ n7440 ;
  assign n21261 = n21260 ^ n8359 ^ n4633 ;
  assign n21262 = n21261 ^ n12179 ^ n8118 ;
  assign n21263 = x147 & n21262 ;
  assign n21264 = ( n21250 & n21259 ) | ( n21250 & ~n21263 ) | ( n21259 & ~n21263 ) ;
  assign n21265 = n19207 ^ n7426 ^ n4853 ;
  assign n21266 = n7759 ^ n5333 ^ n5253 ;
  assign n21267 = ( ~n1796 & n6820 ) | ( ~n1796 & n21266 ) | ( n6820 & n21266 ) ;
  assign n21268 = n21267 ^ n13841 ^ n1173 ;
  assign n21269 = ( n18033 & ~n21265 ) | ( n18033 & n21268 ) | ( ~n21265 & n21268 ) ;
  assign n21271 = ~n7211 & n8867 ;
  assign n21272 = n16753 ^ n3874 ^ n1357 ;
  assign n21273 = ~n2946 & n21272 ;
  assign n21274 = n13994 & n21273 ;
  assign n21275 = ( n9503 & ~n21271 ) | ( n9503 & n21274 ) | ( ~n21271 & n21274 ) ;
  assign n21270 = n345 & n8096 ;
  assign n21276 = n21275 ^ n21270 ^ 1'b0 ;
  assign n21277 = ( n1212 & n21269 ) | ( n1212 & n21276 ) | ( n21269 & n21276 ) ;
  assign n21278 = n6841 ^ n6657 ^ n2180 ;
  assign n21279 = n10859 ^ n3788 ^ n1692 ;
  assign n21280 = ( n7019 & n8905 ) | ( n7019 & ~n21279 ) | ( n8905 & ~n21279 ) ;
  assign n21281 = ~n21278 & n21280 ;
  assign n21282 = n15085 ^ n15007 ^ n9493 ;
  assign n21283 = ( n9307 & ~n20746 ) | ( n9307 & n21282 ) | ( ~n20746 & n21282 ) ;
  assign n21284 = ( n6765 & ~n7671 ) | ( n6765 & n20526 ) | ( ~n7671 & n20526 ) ;
  assign n21286 = n6068 ^ n4737 ^ n1186 ;
  assign n21287 = x4 & ~n21286 ;
  assign n21288 = n21287 ^ n18132 ^ 1'b0 ;
  assign n21289 = ( n2756 & n7440 ) | ( n2756 & n21288 ) | ( n7440 & n21288 ) ;
  assign n21285 = ( ~n3158 & n15318 ) | ( ~n3158 & n20447 ) | ( n15318 & n20447 ) ;
  assign n21290 = n21289 ^ n21285 ^ n15814 ;
  assign n21291 = n2764 & n10511 ;
  assign n21292 = n7220 ^ n5582 ^ n1875 ;
  assign n21293 = ~n3166 & n11717 ;
  assign n21294 = ~n17624 & n21293 ;
  assign n21295 = ( n19863 & ~n21292 ) | ( n19863 & n21294 ) | ( ~n21292 & n21294 ) ;
  assign n21296 = ( n6031 & n6252 ) | ( n6031 & ~n9451 ) | ( n6252 & ~n9451 ) ;
  assign n21297 = n1355 & ~n15692 ;
  assign n21298 = ~n7433 & n21297 ;
  assign n21299 = ( ~n11305 & n21296 ) | ( ~n11305 & n21298 ) | ( n21296 & n21298 ) ;
  assign n21300 = n16355 ^ n8662 ^ n5370 ;
  assign n21301 = n7373 & ~n21300 ;
  assign n21302 = n21301 ^ n1395 ^ 1'b0 ;
  assign n21303 = n21302 ^ n12391 ^ n4528 ;
  assign n21304 = ( ~n3824 & n21299 ) | ( ~n3824 & n21303 ) | ( n21299 & n21303 ) ;
  assign n21305 = n15570 ^ n11050 ^ 1'b0 ;
  assign n21306 = n12396 ^ n8703 ^ n2223 ;
  assign n21307 = ( n18785 & n21305 ) | ( n18785 & n21306 ) | ( n21305 & n21306 ) ;
  assign n21308 = n10582 ^ n2448 ^ n2421 ;
  assign n21309 = ( ~n10952 & n13632 ) | ( ~n10952 & n21308 ) | ( n13632 & n21308 ) ;
  assign n21310 = ( n2773 & n10144 ) | ( n2773 & n21309 ) | ( n10144 & n21309 ) ;
  assign n21311 = n2786 | n10017 ;
  assign n21312 = ( n6061 & n7165 ) | ( n6061 & n21311 ) | ( n7165 & n21311 ) ;
  assign n21313 = n9311 & n21312 ;
  assign n21322 = n9550 ^ n2799 ^ 1'b0 ;
  assign n21323 = n1138 & n21322 ;
  assign n21324 = ~n12635 & n21323 ;
  assign n21315 = ( n3655 & n7401 ) | ( n3655 & n8936 ) | ( n7401 & n8936 ) ;
  assign n21314 = n14676 ^ n6136 ^ n5731 ;
  assign n21316 = n21315 ^ n21314 ^ n703 ;
  assign n21317 = n21316 ^ n19798 ^ n16446 ;
  assign n21318 = n4681 ^ n3470 ^ n1649 ;
  assign n21319 = n21318 ^ n13329 ^ n11925 ;
  assign n21320 = n832 & n21319 ;
  assign n21321 = ~n21317 & n21320 ;
  assign n21325 = n21324 ^ n21321 ^ n10889 ;
  assign n21326 = ( n4075 & n6450 ) | ( n4075 & ~n8237 ) | ( n6450 & ~n8237 ) ;
  assign n21327 = n21326 ^ n3520 ^ n3366 ;
  assign n21328 = n13802 ^ n8833 ^ n412 ;
  assign n21329 = n21327 & n21328 ;
  assign n21330 = n8355 & n11585 ;
  assign n21331 = ~n5560 & n21330 ;
  assign n21332 = ~n7453 & n15206 ;
  assign n21333 = n21332 ^ n8926 ^ 1'b0 ;
  assign n21335 = ~n1447 & n11515 ;
  assign n21334 = n10297 & ~n14527 ;
  assign n21336 = n21335 ^ n21334 ^ n7352 ;
  assign n21337 = n18842 ^ n8705 ^ n6045 ;
  assign n21338 = ( n8402 & n18374 ) | ( n8402 & n21337 ) | ( n18374 & n21337 ) ;
  assign n21339 = ~n9531 & n12166 ;
  assign n21340 = ( n3753 & n8787 ) | ( n3753 & ~n15857 ) | ( n8787 & ~n15857 ) ;
  assign n21341 = n21340 ^ n17123 ^ n2976 ;
  assign n21342 = ( n18604 & ~n21339 ) | ( n18604 & n21341 ) | ( ~n21339 & n21341 ) ;
  assign n21343 = ( ~n2383 & n6636 ) | ( ~n2383 & n8286 ) | ( n6636 & n8286 ) ;
  assign n21344 = n19127 ^ n15759 ^ n10320 ;
  assign n21345 = n6824 | n13381 ;
  assign n21346 = n580 | n21345 ;
  assign n21347 = ( n21343 & n21344 ) | ( n21343 & n21346 ) | ( n21344 & n21346 ) ;
  assign n21349 = n10867 ^ n6335 ^ n1844 ;
  assign n21348 = ( ~x191 & n2859 ) | ( ~x191 & n9229 ) | ( n2859 & n9229 ) ;
  assign n21350 = n21349 ^ n21348 ^ n6036 ;
  assign n21351 = ( n3320 & n5927 ) | ( n3320 & ~n21350 ) | ( n5927 & ~n21350 ) ;
  assign n21352 = ( n4117 & n4783 ) | ( n4117 & n7955 ) | ( n4783 & n7955 ) ;
  assign n21353 = n21352 ^ n16342 ^ 1'b0 ;
  assign n21354 = n21353 ^ n19036 ^ n13190 ;
  assign n21355 = n9203 ^ n3784 ^ n3739 ;
  assign n21356 = n21355 ^ n12615 ^ 1'b0 ;
  assign n21358 = ( n3379 & n5267 ) | ( n3379 & n6565 ) | ( n5267 & n6565 ) ;
  assign n21357 = ( n4337 & n5748 ) | ( n4337 & n10600 ) | ( n5748 & n10600 ) ;
  assign n21359 = n21358 ^ n21357 ^ n21132 ;
  assign n21360 = ( n13159 & ~n14044 ) | ( n13159 & n21359 ) | ( ~n14044 & n21359 ) ;
  assign n21361 = n3921 & ~n17895 ;
  assign n21362 = ~x73 & n21361 ;
  assign n21363 = ~n2728 & n3286 ;
  assign n21364 = ( n4298 & ~n21362 ) | ( n4298 & n21363 ) | ( ~n21362 & n21363 ) ;
  assign n21365 = n7225 ^ n6909 ^ n5537 ;
  assign n21366 = ( n11291 & n21364 ) | ( n11291 & ~n21365 ) | ( n21364 & ~n21365 ) ;
  assign n21369 = n11742 ^ n10832 ^ 1'b0 ;
  assign n21370 = n14393 & n21369 ;
  assign n21367 = ( n3054 & n3660 ) | ( n3054 & ~n11550 ) | ( n3660 & ~n11550 ) ;
  assign n21368 = n21367 ^ n12532 ^ n5252 ;
  assign n21371 = n21370 ^ n21368 ^ n13226 ;
  assign n21386 = ( n5964 & n9821 ) | ( n5964 & n19033 ) | ( n9821 & n19033 ) ;
  assign n21385 = ( n3189 & ~n6733 ) | ( n3189 & n15096 ) | ( ~n6733 & n15096 ) ;
  assign n21387 = n21386 ^ n21385 ^ n15619 ;
  assign n21388 = n14322 ^ n4231 ^ 1'b0 ;
  assign n21389 = n21387 & n21388 ;
  assign n21381 = ( n2046 & ~n2361 ) | ( n2046 & n7324 ) | ( ~n2361 & n7324 ) ;
  assign n21382 = n21381 ^ n2173 ^ n498 ;
  assign n21379 = n6019 ^ n5287 ^ 1'b0 ;
  assign n21380 = n9092 & n21379 ;
  assign n21377 = n2712 & n8160 ;
  assign n21378 = n21377 ^ n6895 ^ x128 ;
  assign n21383 = n21382 ^ n21380 ^ n21378 ;
  assign n21384 = n21383 ^ n16732 ^ n15780 ;
  assign n21372 = n2791 ^ n2342 ^ 1'b0 ;
  assign n21373 = n3116 | n21372 ;
  assign n21374 = n2308 & ~n21373 ;
  assign n21375 = n21374 ^ n15139 ^ 1'b0 ;
  assign n21376 = n21375 ^ n19148 ^ 1'b0 ;
  assign n21390 = n21389 ^ n21384 ^ n21376 ;
  assign n21391 = n7182 & ~n18654 ;
  assign n21392 = ~n3470 & n21391 ;
  assign n21393 = n21392 ^ n6907 ^ 1'b0 ;
  assign n21394 = n11347 & n21393 ;
  assign n21395 = n21394 ^ n8011 ^ 1'b0 ;
  assign n21396 = ( n1588 & n17424 ) | ( n1588 & ~n17883 ) | ( n17424 & ~n17883 ) ;
  assign n21397 = ( n13273 & ~n15301 ) | ( n13273 & n21396 ) | ( ~n15301 & n21396 ) ;
  assign n21398 = ( n4004 & n19121 ) | ( n4004 & n19452 ) | ( n19121 & n19452 ) ;
  assign n21399 = n9529 ^ n7171 ^ 1'b0 ;
  assign n21400 = n13354 ^ n6928 ^ 1'b0 ;
  assign n21401 = ( ~n10590 & n21399 ) | ( ~n10590 & n21400 ) | ( n21399 & n21400 ) ;
  assign n21402 = ( n2271 & n6330 ) | ( n2271 & ~n9727 ) | ( n6330 & ~n9727 ) ;
  assign n21403 = n21402 ^ n11593 ^ 1'b0 ;
  assign n21404 = ( n2496 & n16616 ) | ( n2496 & ~n19971 ) | ( n16616 & ~n19971 ) ;
  assign n21405 = ( n7964 & n11115 ) | ( n7964 & ~n15844 ) | ( n11115 & ~n15844 ) ;
  assign n21407 = ( n1479 & n2090 ) | ( n1479 & n8800 ) | ( n2090 & n8800 ) ;
  assign n21408 = n21407 ^ n7701 ^ n6732 ;
  assign n21406 = n11547 ^ n5429 ^ n3096 ;
  assign n21409 = n21408 ^ n21406 ^ n11298 ;
  assign n21410 = ( n4412 & n6863 ) | ( n4412 & ~n21409 ) | ( n6863 & ~n21409 ) ;
  assign n21411 = ( n13102 & n21405 ) | ( n13102 & ~n21410 ) | ( n21405 & ~n21410 ) ;
  assign n21412 = n7641 ^ n7436 ^ n4910 ;
  assign n21413 = ( n2345 & n9910 ) | ( n2345 & n10383 ) | ( n9910 & n10383 ) ;
  assign n21414 = ( ~n525 & n21412 ) | ( ~n525 & n21413 ) | ( n21412 & n21413 ) ;
  assign n21415 = ( n716 & n4361 ) | ( n716 & ~n4424 ) | ( n4361 & ~n4424 ) ;
  assign n21416 = n7073 ^ n6424 ^ n4669 ;
  assign n21419 = n18497 ^ n9938 ^ n7893 ;
  assign n21418 = n10014 ^ n5670 ^ x233 ;
  assign n21420 = n21419 ^ n21418 ^ n2525 ;
  assign n21421 = ( ~n4224 & n14795 ) | ( ~n4224 & n21420 ) | ( n14795 & n21420 ) ;
  assign n21417 = n5462 & n6701 ;
  assign n21422 = n21421 ^ n21417 ^ 1'b0 ;
  assign n21423 = ( n19582 & n21416 ) | ( n19582 & n21422 ) | ( n21416 & n21422 ) ;
  assign n21424 = n18258 ^ n13603 ^ n8102 ;
  assign n21425 = ( n15448 & n20569 ) | ( n15448 & n21424 ) | ( n20569 & n21424 ) ;
  assign n21426 = ( n2131 & n3234 ) | ( n2131 & ~n7927 ) | ( n3234 & ~n7927 ) ;
  assign n21427 = ~n21425 & n21426 ;
  assign n21428 = ( n900 & n3627 ) | ( n900 & ~n12595 ) | ( n3627 & ~n12595 ) ;
  assign n21429 = n1135 & n4159 ;
  assign n21430 = n5039 & n21429 ;
  assign n21431 = ( ~n3083 & n10816 ) | ( ~n3083 & n21430 ) | ( n10816 & n21430 ) ;
  assign n21432 = ( n4938 & ~n21428 ) | ( n4938 & n21431 ) | ( ~n21428 & n21431 ) ;
  assign n21433 = ( n6417 & n11325 ) | ( n6417 & n20459 ) | ( n11325 & n20459 ) ;
  assign n21434 = n21433 ^ n12977 ^ 1'b0 ;
  assign n21435 = n8743 ^ n3087 ^ n2556 ;
  assign n21436 = n21435 ^ n17295 ^ n6442 ;
  assign n21437 = ( n9010 & n15770 ) | ( n9010 & ~n21436 ) | ( n15770 & ~n21436 ) ;
  assign n21441 = n15226 ^ n14017 ^ n8932 ;
  assign n21439 = n18394 ^ n17699 ^ n997 ;
  assign n21440 = n21439 ^ n5720 ^ x69 ;
  assign n21438 = n8951 ^ n7424 ^ n3192 ;
  assign n21442 = n21441 ^ n21440 ^ n21438 ;
  assign n21443 = ( ~n20373 & n21437 ) | ( ~n20373 & n21442 ) | ( n21437 & n21442 ) ;
  assign n21445 = ( ~n653 & n5370 ) | ( ~n653 & n9670 ) | ( n5370 & n9670 ) ;
  assign n21444 = n4398 ^ n3932 ^ n1326 ;
  assign n21446 = n21445 ^ n21444 ^ n5046 ;
  assign n21447 = n10988 ^ n4205 ^ n1493 ;
  assign n21448 = n21447 ^ n6898 ^ n1465 ;
  assign n21449 = ( n7654 & ~n16450 ) | ( n7654 & n21448 ) | ( ~n16450 & n21448 ) ;
  assign n21451 = n15852 ^ n13620 ^ n2204 ;
  assign n21450 = ( ~n5246 & n9508 ) | ( ~n5246 & n10454 ) | ( n9508 & n10454 ) ;
  assign n21452 = n21451 ^ n21450 ^ 1'b0 ;
  assign n21453 = n21449 & ~n21452 ;
  assign n21454 = ~n21446 & n21453 ;
  assign n21455 = n12470 ^ n8056 ^ n3547 ;
  assign n21456 = ( n11316 & n14981 ) | ( n11316 & ~n21455 ) | ( n14981 & ~n21455 ) ;
  assign n21460 = ( n959 & n1865 ) | ( n959 & n13556 ) | ( n1865 & n13556 ) ;
  assign n21457 = n8728 ^ n7583 ^ n7021 ;
  assign n21458 = n16811 ^ n5146 ^ 1'b0 ;
  assign n21459 = ( n19977 & ~n21457 ) | ( n19977 & n21458 ) | ( ~n21457 & n21458 ) ;
  assign n21461 = n21460 ^ n21459 ^ n13423 ;
  assign n21462 = ( n7341 & ~n21456 ) | ( n7341 & n21461 ) | ( ~n21456 & n21461 ) ;
  assign n21463 = ( n9299 & n10546 ) | ( n9299 & ~n14849 ) | ( n10546 & ~n14849 ) ;
  assign n21464 = n9752 | n21463 ;
  assign n21465 = ( ~n1153 & n9088 ) | ( ~n1153 & n21464 ) | ( n9088 & n21464 ) ;
  assign n21466 = n6543 ^ n522 ^ 1'b0 ;
  assign n21467 = ( n2954 & n16936 ) | ( n2954 & n21466 ) | ( n16936 & n21466 ) ;
  assign n21468 = n21467 ^ n13313 ^ n11894 ;
  assign n21471 = n17191 ^ n15724 ^ n1424 ;
  assign n21469 = ( n916 & ~n8193 ) | ( n916 & n17249 ) | ( ~n8193 & n17249 ) ;
  assign n21470 = n21469 ^ n16610 ^ n14915 ;
  assign n21472 = n21471 ^ n21470 ^ n13900 ;
  assign n21473 = ( ~n13512 & n13837 ) | ( ~n13512 & n17315 ) | ( n13837 & n17315 ) ;
  assign n21474 = n21473 ^ n8271 ^ n5497 ;
  assign n21475 = n8064 ^ n6321 ^ 1'b0 ;
  assign n21476 = n1796 | n21475 ;
  assign n21477 = ( n12019 & n13935 ) | ( n12019 & ~n18067 ) | ( n13935 & ~n18067 ) ;
  assign n21478 = n21477 ^ n20176 ^ n18219 ;
  assign n21488 = n9965 ^ n6813 ^ n6673 ;
  assign n21485 = n15993 ^ n1716 ^ 1'b0 ;
  assign n21486 = n21485 ^ n11355 ^ 1'b0 ;
  assign n21487 = n11134 & ~n21486 ;
  assign n21480 = n1228 & ~n4148 ;
  assign n21481 = n2688 & n21480 ;
  assign n21479 = n18471 ^ n3883 ^ n327 ;
  assign n21482 = n21481 ^ n21479 ^ n551 ;
  assign n21483 = n17042 ^ n16097 ^ n8075 ;
  assign n21484 = n21482 & ~n21483 ;
  assign n21489 = n21488 ^ n21487 ^ n21484 ;
  assign n21491 = n6214 ^ n486 ^ 1'b0 ;
  assign n21492 = ~n5276 & n21491 ;
  assign n21493 = n17336 ^ n4039 ^ n3581 ;
  assign n21494 = n12387 ^ n5271 ^ 1'b0 ;
  assign n21495 = n21493 & n21494 ;
  assign n21496 = n21495 ^ n5574 ^ n4673 ;
  assign n21497 = ( n10954 & n21492 ) | ( n10954 & ~n21496 ) | ( n21492 & ~n21496 ) ;
  assign n21490 = n17505 ^ n13333 ^ n3162 ;
  assign n21498 = n21497 ^ n21490 ^ n16476 ;
  assign n21499 = n19659 ^ n6984 ^ 1'b0 ;
  assign n21500 = ~n20983 & n21499 ;
  assign n21501 = n21500 ^ n17531 ^ n7700 ;
  assign n21502 = ( n1045 & ~n14170 ) | ( n1045 & n21501 ) | ( ~n14170 & n21501 ) ;
  assign n21503 = ( n1637 & ~n8633 ) | ( n1637 & n11085 ) | ( ~n8633 & n11085 ) ;
  assign n21504 = ( n9164 & n17002 ) | ( n9164 & n21503 ) | ( n17002 & n21503 ) ;
  assign n21508 = n5001 & ~n6765 ;
  assign n21506 = n15356 ^ n9930 ^ n5043 ;
  assign n21507 = n459 | n21506 ;
  assign n21505 = n17446 ^ n5716 ^ n3639 ;
  assign n21509 = n21508 ^ n21507 ^ n21505 ;
  assign n21510 = n21466 ^ n13812 ^ n661 ;
  assign n21511 = ~n14385 & n21510 ;
  assign n21512 = ( n12386 & n21268 ) | ( n12386 & n21511 ) | ( n21268 & n21511 ) ;
  assign n21513 = ( n929 & n8278 ) | ( n929 & n21512 ) | ( n8278 & n21512 ) ;
  assign n21514 = ( ~n5173 & n15112 ) | ( ~n5173 & n15371 ) | ( n15112 & n15371 ) ;
  assign n21515 = n21514 ^ n10151 ^ n6581 ;
  assign n21516 = n5637 & ~n21515 ;
  assign n21517 = n21516 ^ n12462 ^ 1'b0 ;
  assign n21519 = n19985 ^ n15711 ^ n1635 ;
  assign n21520 = ( n1197 & n3488 ) | ( n1197 & ~n21519 ) | ( n3488 & ~n21519 ) ;
  assign n21518 = n19339 & n20580 ;
  assign n21521 = n21520 ^ n21518 ^ 1'b0 ;
  assign n21522 = n18967 ^ n9305 ^ n895 ;
  assign n21523 = ( n5889 & ~n10876 ) | ( n5889 & n21522 ) | ( ~n10876 & n21522 ) ;
  assign n21524 = n3298 & ~n10835 ;
  assign n21525 = n21524 ^ n11646 ^ 1'b0 ;
  assign n21526 = ( n8087 & n10219 ) | ( n8087 & n21525 ) | ( n10219 & n21525 ) ;
  assign n21527 = ( n6410 & n14761 ) | ( n6410 & ~n21526 ) | ( n14761 & ~n21526 ) ;
  assign n21528 = ( n2595 & n4095 ) | ( n2595 & ~n8364 ) | ( n4095 & ~n8364 ) ;
  assign n21529 = n8112 | n21528 ;
  assign n21530 = ( n8854 & n14247 ) | ( n8854 & ~n21529 ) | ( n14247 & ~n21529 ) ;
  assign n21531 = n18906 ^ n10996 ^ 1'b0 ;
  assign n21532 = ( ~n9933 & n11341 ) | ( ~n9933 & n13675 ) | ( n11341 & n13675 ) ;
  assign n21533 = ( ~n6314 & n9842 ) | ( ~n6314 & n21532 ) | ( n9842 & n21532 ) ;
  assign n21534 = n6361 ^ n5083 ^ n5003 ;
  assign n21535 = ~n7550 & n21534 ;
  assign n21536 = n21533 & ~n21535 ;
  assign n21537 = n12218 ^ n961 ^ n363 ;
  assign n21538 = n21537 ^ n9336 ^ n6299 ;
  assign n21539 = n11055 ^ n6938 ^ 1'b0 ;
  assign n21540 = n21539 ^ n16533 ^ n7903 ;
  assign n21543 = ( ~n4544 & n7523 ) | ( ~n4544 & n8243 ) | ( n7523 & n8243 ) ;
  assign n21544 = n13213 & n21543 ;
  assign n21545 = n9660 & ~n21544 ;
  assign n21541 = ( n3813 & ~n10380 ) | ( n3813 & n17750 ) | ( ~n10380 & n17750 ) ;
  assign n21542 = n21541 ^ n18214 ^ n973 ;
  assign n21546 = n21545 ^ n21542 ^ n11929 ;
  assign n21547 = ( n5164 & ~n8487 ) | ( n5164 & n19453 ) | ( ~n8487 & n19453 ) ;
  assign n21548 = n9770 ^ n5929 ^ 1'b0 ;
  assign n21549 = n21548 ^ n20312 ^ 1'b0 ;
  assign n21550 = ~n6902 & n21549 ;
  assign n21557 = ( n2436 & n3293 ) | ( n2436 & n4505 ) | ( n3293 & n4505 ) ;
  assign n21551 = n5519 & n12300 ;
  assign n21552 = n4231 & n21551 ;
  assign n21553 = n21552 ^ n13755 ^ n7319 ;
  assign n21554 = n16317 ^ n374 ^ 1'b0 ;
  assign n21555 = n21553 | n21554 ;
  assign n21556 = ( ~n11512 & n16345 ) | ( ~n11512 & n21555 ) | ( n16345 & n21555 ) ;
  assign n21558 = n21557 ^ n21556 ^ n3313 ;
  assign n21559 = n5070 & ~n10940 ;
  assign n21560 = n21559 ^ n11306 ^ 1'b0 ;
  assign n21561 = n21560 ^ n12462 ^ n916 ;
  assign n21567 = n12666 ^ n2859 ^ n1684 ;
  assign n21568 = n21567 ^ n11160 ^ n5600 ;
  assign n21569 = n21568 ^ n11214 ^ 1'b0 ;
  assign n21570 = n10197 & ~n21569 ;
  assign n21562 = n3470 & ~n4385 ;
  assign n21563 = n12525 ^ n11532 ^ 1'b0 ;
  assign n21564 = ( n11285 & n13627 ) | ( n11285 & n21563 ) | ( n13627 & n21563 ) ;
  assign n21565 = ( ~n21456 & n21562 ) | ( ~n21456 & n21564 ) | ( n21562 & n21564 ) ;
  assign n21566 = n21565 ^ n12302 ^ n11579 ;
  assign n21571 = n21570 ^ n21566 ^ n14704 ;
  assign n21574 = ~n5717 & n11582 ;
  assign n21575 = n21574 ^ n3106 ^ 1'b0 ;
  assign n21572 = n11755 ^ n4837 ^ 1'b0 ;
  assign n21573 = n5290 & ~n21572 ;
  assign n21576 = n21575 ^ n21573 ^ n1554 ;
  assign n21577 = n18639 ^ n11322 ^ n793 ;
  assign n21578 = ( n7371 & n10478 ) | ( n7371 & n16699 ) | ( n10478 & n16699 ) ;
  assign n21579 = n14033 ^ n3893 ^ 1'b0 ;
  assign n21580 = n21578 | n21579 ;
  assign n21581 = ( n2681 & ~n11970 ) | ( n2681 & n21580 ) | ( ~n11970 & n21580 ) ;
  assign n21593 = n21298 ^ n12438 ^ n4199 ;
  assign n21594 = n10291 & ~n21130 ;
  assign n21595 = ~n21593 & n21594 ;
  assign n21587 = n6141 ^ n1757 ^ n915 ;
  assign n21588 = n21587 ^ n1204 ^ n1087 ;
  assign n21589 = n3693 | n21588 ;
  assign n21590 = ( n11953 & n20050 ) | ( n11953 & ~n21589 ) | ( n20050 & ~n21589 ) ;
  assign n21585 = n3548 ^ n617 ^ 1'b0 ;
  assign n21586 = ( n10075 & n18935 ) | ( n10075 & ~n21585 ) | ( n18935 & ~n21585 ) ;
  assign n21582 = n9691 ^ n6465 ^ n1152 ;
  assign n21583 = ( x107 & n9937 ) | ( x107 & n21582 ) | ( n9937 & n21582 ) ;
  assign n21584 = ( n3147 & n14922 ) | ( n3147 & n21583 ) | ( n14922 & n21583 ) ;
  assign n21591 = n21590 ^ n21586 ^ n21584 ;
  assign n21592 = ( n1555 & ~n5402 ) | ( n1555 & n21591 ) | ( ~n5402 & n21591 ) ;
  assign n21596 = n21595 ^ n21592 ^ n9874 ;
  assign n21597 = n3072 ^ n1590 ^ 1'b0 ;
  assign n21598 = n21597 ^ n8798 ^ 1'b0 ;
  assign n21599 = n1919 | n21598 ;
  assign n21600 = n368 & ~n21599 ;
  assign n21601 = n21600 ^ n8470 ^ 1'b0 ;
  assign n21602 = ( ~n5199 & n11359 ) | ( ~n5199 & n18184 ) | ( n11359 & n18184 ) ;
  assign n21603 = n21602 ^ n17504 ^ n13925 ;
  assign n21604 = ( ~n311 & n15805 ) | ( ~n311 & n21603 ) | ( n15805 & n21603 ) ;
  assign n21605 = ( n15778 & n21601 ) | ( n15778 & n21604 ) | ( n21601 & n21604 ) ;
  assign n21606 = n16956 ^ n14998 ^ n4049 ;
  assign n21609 = ( n1072 & n12670 ) | ( n1072 & ~n17662 ) | ( n12670 & ~n17662 ) ;
  assign n21610 = ( n1188 & n7252 ) | ( n1188 & ~n21609 ) | ( n7252 & ~n21609 ) ;
  assign n21611 = n21610 ^ n17820 ^ n14773 ;
  assign n21607 = ( n4133 & n6913 ) | ( n4133 & n18342 ) | ( n6913 & n18342 ) ;
  assign n21608 = ( n12984 & ~n15423 ) | ( n12984 & n21607 ) | ( ~n15423 & n21607 ) ;
  assign n21612 = n21611 ^ n21608 ^ n9396 ;
  assign n21613 = n21606 | n21612 ;
  assign n21614 = n19085 ^ n12624 ^ x45 ;
  assign n21615 = n18859 & ~n21614 ;
  assign n21616 = n9342 ^ n6685 ^ n409 ;
  assign n21617 = ( n3702 & n7316 ) | ( n3702 & n21616 ) | ( n7316 & n21616 ) ;
  assign n21618 = n21617 ^ n12900 ^ n10378 ;
  assign n21619 = n15557 ^ n7911 ^ n4036 ;
  assign n21620 = n14427 ^ n666 ^ 1'b0 ;
  assign n21621 = n17360 ^ n9177 ^ n3846 ;
  assign n21623 = n8252 & ~n11113 ;
  assign n21624 = n12686 & n21623 ;
  assign n21622 = ~n810 & n7648 ;
  assign n21625 = n21624 ^ n21622 ^ 1'b0 ;
  assign n21626 = n11504 ^ n7122 ^ n1767 ;
  assign n21627 = ( x236 & ~n5253 ) | ( x236 & n21626 ) | ( ~n5253 & n21626 ) ;
  assign n21628 = ( n1285 & ~n1654 ) | ( n1285 & n12723 ) | ( ~n1654 & n12723 ) ;
  assign n21629 = n21628 ^ n5774 ^ n1263 ;
  assign n21630 = ( n13055 & ~n20615 ) | ( n13055 & n21629 ) | ( ~n20615 & n21629 ) ;
  assign n21631 = n11724 ^ n11490 ^ n6853 ;
  assign n21632 = n16058 ^ n14546 ^ n4749 ;
  assign n21633 = ( n7882 & ~n21311 ) | ( n7882 & n21632 ) | ( ~n21311 & n21632 ) ;
  assign n21634 = n21633 ^ n5848 ^ n2894 ;
  assign n21635 = ( ~n1020 & n4452 ) | ( ~n1020 & n6365 ) | ( n4452 & n6365 ) ;
  assign n21636 = ( n6721 & n13301 ) | ( n6721 & n17388 ) | ( n13301 & n17388 ) ;
  assign n21637 = ( n13656 & n21635 ) | ( n13656 & n21636 ) | ( n21635 & n21636 ) ;
  assign n21638 = ( n6752 & ~n10070 ) | ( n6752 & n21637 ) | ( ~n10070 & n21637 ) ;
  assign n21640 = n2050 | n9361 ;
  assign n21641 = n13946 & ~n21640 ;
  assign n21642 = n21641 ^ n17853 ^ 1'b0 ;
  assign n21639 = n4039 & n11749 ;
  assign n21643 = n21642 ^ n21639 ^ 1'b0 ;
  assign n21644 = ~n766 & n1262 ;
  assign n21645 = ~x135 & n21644 ;
  assign n21646 = ( n8082 & ~n10876 ) | ( n8082 & n21645 ) | ( ~n10876 & n21645 ) ;
  assign n21647 = x153 & n8504 ;
  assign n21648 = n2027 & n21647 ;
  assign n21649 = ( n1120 & ~n1131 ) | ( n1120 & n3407 ) | ( ~n1131 & n3407 ) ;
  assign n21650 = n21649 ^ n13926 ^ n1915 ;
  assign n21651 = ( n441 & n21648 ) | ( n441 & n21650 ) | ( n21648 & n21650 ) ;
  assign n21652 = n20242 ^ n4081 ^ 1'b0 ;
  assign n21653 = n21652 ^ n21588 ^ n6993 ;
  assign n21654 = ( n3721 & ~n4677 ) | ( n3721 & n8453 ) | ( ~n4677 & n8453 ) ;
  assign n21655 = n21654 ^ n16081 ^ x107 ;
  assign n21656 = n15944 ^ n10557 ^ n2834 ;
  assign n21657 = n21656 ^ n4156 ^ n1264 ;
  assign n21658 = n21657 ^ n18060 ^ n16339 ;
  assign n21659 = n21340 & n21658 ;
  assign n21660 = ~n18172 & n21659 ;
  assign n21661 = ( ~n4197 & n7438 ) | ( ~n4197 & n8205 ) | ( n7438 & n8205 ) ;
  assign n21662 = n17366 ^ n8575 ^ 1'b0 ;
  assign n21663 = n21662 ^ n14061 ^ n6159 ;
  assign n21665 = n2610 ^ x55 ^ 1'b0 ;
  assign n21664 = n12692 ^ n7673 ^ x33 ;
  assign n21666 = n21665 ^ n21664 ^ n17699 ;
  assign n21667 = ( n21661 & n21663 ) | ( n21661 & ~n21666 ) | ( n21663 & ~n21666 ) ;
  assign n21668 = ( n2810 & n14640 ) | ( n2810 & n19045 ) | ( n14640 & n19045 ) ;
  assign n21669 = n21668 ^ n10313 ^ n9754 ;
  assign n21670 = n10189 ^ n7199 ^ n588 ;
  assign n21671 = n18038 ^ n3672 ^ n1664 ;
  assign n21672 = ( ~n14518 & n21670 ) | ( ~n14518 & n21671 ) | ( n21670 & n21671 ) ;
  assign n21673 = n21672 ^ n3316 ^ 1'b0 ;
  assign n21686 = n16499 | n18155 ;
  assign n21687 = n21686 ^ n3249 ^ 1'b0 ;
  assign n21684 = n3514 & ~n7390 ;
  assign n21681 = n13393 ^ n3541 ^ n1261 ;
  assign n21682 = n21681 ^ n4338 ^ n2410 ;
  assign n21683 = ( n1701 & n10777 ) | ( n1701 & ~n21682 ) | ( n10777 & ~n21682 ) ;
  assign n21685 = n21684 ^ n21683 ^ 1'b0 ;
  assign n21674 = n5358 ^ n4157 ^ n2222 ;
  assign n21675 = n21674 ^ n8900 ^ n5454 ;
  assign n21676 = ( n2914 & ~n4283 ) | ( n2914 & n21675 ) | ( ~n4283 & n21675 ) ;
  assign n21677 = ( n6262 & n14767 ) | ( n6262 & ~n21254 ) | ( n14767 & ~n21254 ) ;
  assign n21678 = ( n9563 & n18243 ) | ( n9563 & ~n21677 ) | ( n18243 & ~n21677 ) ;
  assign n21679 = n18758 ^ n11664 ^ n1989 ;
  assign n21680 = ( n21676 & n21678 ) | ( n21676 & ~n21679 ) | ( n21678 & ~n21679 ) ;
  assign n21688 = n21687 ^ n21685 ^ n21680 ;
  assign n21691 = ( n7998 & n11386 ) | ( n7998 & ~n14473 ) | ( n11386 & ~n14473 ) ;
  assign n21692 = ( ~n4066 & n9227 ) | ( ~n4066 & n21691 ) | ( n9227 & n21691 ) ;
  assign n21689 = n20915 ^ n16784 ^ n4428 ;
  assign n21690 = n21689 ^ n12019 ^ n7809 ;
  assign n21693 = n21692 ^ n21690 ^ n7999 ;
  assign n21694 = ( ~n14637 & n17530 ) | ( ~n14637 & n19851 ) | ( n17530 & n19851 ) ;
  assign n21695 = n15107 ^ n13113 ^ 1'b0 ;
  assign n21696 = n13973 | n21695 ;
  assign n21697 = n21340 ^ n12241 ^ n5581 ;
  assign n21698 = n5097 ^ n4354 ^ n2721 ;
  assign n21699 = ( n7058 & ~n18645 ) | ( n7058 & n21698 ) | ( ~n18645 & n21698 ) ;
  assign n21700 = n17261 ^ n16883 ^ n6891 ;
  assign n21701 = ( ~n5698 & n14947 ) | ( ~n5698 & n21700 ) | ( n14947 & n21700 ) ;
  assign n21702 = n21701 ^ n17965 ^ n11137 ;
  assign n21703 = n21702 ^ n4186 ^ n3002 ;
  assign n21704 = ( ~n1140 & n1446 ) | ( ~n1140 & n14907 ) | ( n1446 & n14907 ) ;
  assign n21719 = ( n2620 & ~n3509 ) | ( n2620 & n8065 ) | ( ~n3509 & n8065 ) ;
  assign n21717 = n7708 ^ n1226 ^ 1'b0 ;
  assign n21718 = n1752 & n21717 ;
  assign n21720 = n21719 ^ n21718 ^ n2651 ;
  assign n21705 = n3236 & ~n4793 ;
  assign n21706 = ( ~n5811 & n5956 ) | ( ~n5811 & n21705 ) | ( n5956 & n21705 ) ;
  assign n21707 = n21706 ^ n11314 ^ n1432 ;
  assign n21713 = ( n868 & n10247 ) | ( n868 & n10350 ) | ( n10247 & n10350 ) ;
  assign n21714 = ( ~n6313 & n10709 ) | ( ~n6313 & n21713 ) | ( n10709 & n21713 ) ;
  assign n21710 = n6862 ^ n6813 ^ n3767 ;
  assign n21711 = ( n13006 & ~n18328 ) | ( n13006 & n21710 ) | ( ~n18328 & n21710 ) ;
  assign n21708 = ( n397 & ~n10111 ) | ( n397 & n10893 ) | ( ~n10111 & n10893 ) ;
  assign n21709 = n21708 ^ n21120 ^ n8818 ;
  assign n21712 = n21711 ^ n21709 ^ n8643 ;
  assign n21715 = n21714 ^ n21712 ^ n1381 ;
  assign n21716 = ( ~n5993 & n21707 ) | ( ~n5993 & n21715 ) | ( n21707 & n21715 ) ;
  assign n21721 = n21720 ^ n21716 ^ n14586 ;
  assign n21722 = n1684 & n8168 ;
  assign n21723 = n2162 & ~n21722 ;
  assign n21728 = ( ~n804 & n15414 ) | ( ~n804 & n15592 ) | ( n15414 & n15592 ) ;
  assign n21724 = n6720 ^ n1889 ^ 1'b0 ;
  assign n21725 = n21724 ^ n7567 ^ 1'b0 ;
  assign n21726 = n8989 | n21725 ;
  assign n21727 = n21726 ^ n10885 ^ n1262 ;
  assign n21729 = n21728 ^ n21727 ^ n8744 ;
  assign n21730 = n7479 ^ n3771 ^ 1'b0 ;
  assign n21731 = n21730 ^ n10568 ^ n2555 ;
  assign n21732 = ( n2059 & n12202 ) | ( n2059 & ~n17512 ) | ( n12202 & ~n17512 ) ;
  assign n21733 = n21732 ^ n2609 ^ n2235 ;
  assign n21734 = n6577 | n8681 ;
  assign n21735 = n7120 | n21734 ;
  assign n21736 = ~n8810 & n21735 ;
  assign n21737 = n21733 & n21736 ;
  assign n21738 = ( n8113 & n20441 ) | ( n8113 & ~n21737 ) | ( n20441 & ~n21737 ) ;
  assign n21739 = n21738 ^ n20985 ^ n10705 ;
  assign n21740 = n6828 ^ n5993 ^ n1983 ;
  assign n21742 = ( ~n6235 & n10912 ) | ( ~n6235 & n14517 ) | ( n10912 & n14517 ) ;
  assign n21743 = n21742 ^ n12124 ^ n1588 ;
  assign n21741 = n10309 ^ n6841 ^ n2729 ;
  assign n21744 = n21743 ^ n21741 ^ n617 ;
  assign n21745 = n10884 ^ n7997 ^ n675 ;
  assign n21749 = ( n11408 & n14339 ) | ( n11408 & n20811 ) | ( n14339 & n20811 ) ;
  assign n21746 = n11963 ^ n10375 ^ n7674 ;
  assign n21747 = n21746 ^ n12588 ^ 1'b0 ;
  assign n21748 = n12702 & ~n21747 ;
  assign n21750 = n21749 ^ n21748 ^ 1'b0 ;
  assign n21751 = n12612 ^ n5668 ^ 1'b0 ;
  assign n21752 = ( n2715 & n3200 ) | ( n2715 & ~n16950 ) | ( n3200 & ~n16950 ) ;
  assign n21753 = n21752 ^ n21660 ^ n12403 ;
  assign n21755 = n6284 ^ n2954 ^ n1471 ;
  assign n21756 = ( n2581 & n3406 ) | ( n2581 & n21755 ) | ( n3406 & n21755 ) ;
  assign n21754 = n6192 & ~n14212 ;
  assign n21757 = n21756 ^ n21754 ^ 1'b0 ;
  assign n21758 = ( ~n4353 & n14392 ) | ( ~n4353 & n21757 ) | ( n14392 & n21757 ) ;
  assign n21759 = n12459 ^ n2498 ^ 1'b0 ;
  assign n21760 = n21759 ^ n19008 ^ n18455 ;
  assign n21761 = n2987 & n3035 ;
  assign n21762 = n21761 ^ n2759 ^ 1'b0 ;
  assign n21763 = ( ~n4816 & n11541 ) | ( ~n4816 & n21762 ) | ( n11541 & n21762 ) ;
  assign n21768 = ( n1355 & n1758 ) | ( n1355 & n13098 ) | ( n1758 & n13098 ) ;
  assign n21764 = n9545 ^ n3551 ^ n346 ;
  assign n21765 = n21764 ^ n9396 ^ n1432 ;
  assign n21766 = n6885 & ~n21765 ;
  assign n21767 = n9964 & n21766 ;
  assign n21769 = n21768 ^ n21767 ^ 1'b0 ;
  assign n21770 = n8766 & ~n21769 ;
  assign n21771 = ( n7163 & ~n21763 ) | ( n7163 & n21770 ) | ( ~n21763 & n21770 ) ;
  assign n21772 = ~n2860 & n10765 ;
  assign n21773 = n21772 ^ n17874 ^ n12962 ;
  assign n21774 = n21773 ^ n18495 ^ 1'b0 ;
  assign n21775 = n21774 ^ n17120 ^ n13813 ;
  assign n21776 = n12858 ^ n4034 ^ n2243 ;
  assign n21780 = n16644 ^ n14231 ^ n7194 ;
  assign n21777 = n5925 ^ x108 ^ 1'b0 ;
  assign n21778 = ( n6977 & n19477 ) | ( n6977 & n21777 ) | ( n19477 & n21777 ) ;
  assign n21779 = n21778 ^ n10122 ^ x141 ;
  assign n21781 = n21780 ^ n21779 ^ n2171 ;
  assign n21782 = n21781 ^ n19667 ^ n6734 ;
  assign n21783 = n12261 & n21676 ;
  assign n21785 = ( n9879 & n12682 ) | ( n9879 & n20152 ) | ( n12682 & n20152 ) ;
  assign n21786 = n21785 ^ n17075 ^ n2067 ;
  assign n21784 = ( n3745 & n7536 ) | ( n3745 & n10365 ) | ( n7536 & n10365 ) ;
  assign n21787 = n21786 ^ n21784 ^ n17489 ;
  assign n21788 = ( n1905 & n13032 ) | ( n1905 & n15667 ) | ( n13032 & n15667 ) ;
  assign n21789 = n17178 ^ n13834 ^ 1'b0 ;
  assign n21794 = n6231 & n15793 ;
  assign n21795 = n21794 ^ n4675 ^ 1'b0 ;
  assign n21792 = ~n1283 & n2265 ;
  assign n21793 = n21792 ^ n11566 ^ 1'b0 ;
  assign n21790 = n3742 | n19611 ;
  assign n21791 = n21790 ^ n1531 ^ 1'b0 ;
  assign n21796 = n21795 ^ n21793 ^ n21791 ;
  assign n21797 = ~n15948 & n16071 ;
  assign n21798 = n15145 ^ n6575 ^ 1'b0 ;
  assign n21799 = ( n4270 & ~n9478 ) | ( n4270 & n21798 ) | ( ~n9478 & n21798 ) ;
  assign n21800 = n21799 ^ n21793 ^ 1'b0 ;
  assign n21801 = n21797 & n21800 ;
  assign n21802 = n21801 ^ n7816 ^ 1'b0 ;
  assign n21806 = ( ~n555 & n9803 ) | ( ~n555 & n10558 ) | ( n9803 & n10558 ) ;
  assign n21803 = ~n3404 & n8338 ;
  assign n21804 = n6910 & n21803 ;
  assign n21805 = n10205 | n21804 ;
  assign n21807 = n21806 ^ n21805 ^ 1'b0 ;
  assign n21808 = n2507 ^ n2247 ^ n1451 ;
  assign n21809 = ~n4582 & n21808 ;
  assign n21810 = ~n8919 & n21809 ;
  assign n21811 = ( n4119 & n5762 ) | ( n4119 & ~n21810 ) | ( n5762 & ~n21810 ) ;
  assign n21812 = n21811 ^ n6506 ^ n2874 ;
  assign n21813 = n6743 & ~n8778 ;
  assign n21814 = ( ~n7016 & n10989 ) | ( ~n7016 & n21813 ) | ( n10989 & n21813 ) ;
  assign n21815 = ( ~n8747 & n10638 ) | ( ~n8747 & n21814 ) | ( n10638 & n21814 ) ;
  assign n21816 = n9756 | n15659 ;
  assign n21817 = n21815 | n21816 ;
  assign n21819 = n12667 ^ n8110 ^ n295 ;
  assign n21818 = ( n7476 & n8142 ) | ( n7476 & ~n18764 ) | ( n8142 & ~n18764 ) ;
  assign n21820 = n21819 ^ n21818 ^ n12213 ;
  assign n21821 = n9243 ^ n508 ^ 1'b0 ;
  assign n21822 = n21820 & n21821 ;
  assign n21823 = n11470 & ~n21381 ;
  assign n21824 = ( ~n9953 & n19995 ) | ( ~n9953 & n21823 ) | ( n19995 & n21823 ) ;
  assign n21825 = n6959 & ~n21824 ;
  assign n21826 = ~n17287 & n21825 ;
  assign n21836 = ( n6687 & n7810 ) | ( n6687 & n17196 ) | ( n7810 & n17196 ) ;
  assign n21827 = n5975 ^ n1357 ^ 1'b0 ;
  assign n21828 = n3425 & n21827 ;
  assign n21829 = ( n465 & n8813 ) | ( n465 & n10572 ) | ( n8813 & n10572 ) ;
  assign n21830 = ( n9435 & n21828 ) | ( n9435 & n21829 ) | ( n21828 & n21829 ) ;
  assign n21831 = n16587 ^ n9456 ^ n2164 ;
  assign n21832 = n10892 & ~n21831 ;
  assign n21833 = ~n21830 & n21832 ;
  assign n21834 = n21833 ^ n9202 ^ n7388 ;
  assign n21835 = n21834 ^ n15008 ^ n6904 ;
  assign n21837 = n21836 ^ n21835 ^ n3557 ;
  assign n21838 = n18614 ^ n15750 ^ n9499 ;
  assign n21843 = n6947 & n17566 ;
  assign n21839 = n4884 & ~n10718 ;
  assign n21840 = ~n20085 & n21839 ;
  assign n21841 = n21840 ^ n21482 ^ n3869 ;
  assign n21842 = ( n1970 & n7329 ) | ( n1970 & n21841 ) | ( n7329 & n21841 ) ;
  assign n21844 = n21843 ^ n21842 ^ n1685 ;
  assign n21846 = n14374 ^ n9827 ^ 1'b0 ;
  assign n21847 = n21846 ^ n12274 ^ 1'b0 ;
  assign n21845 = n17340 ^ n4128 ^ n3056 ;
  assign n21848 = n21847 ^ n21845 ^ n20170 ;
  assign n21849 = ( n13909 & n14485 ) | ( n13909 & ~n21240 ) | ( n14485 & ~n21240 ) ;
  assign n21850 = n14902 ^ n4575 ^ x201 ;
  assign n21851 = ~n3376 & n21850 ;
  assign n21852 = n21851 ^ n17889 ^ n11471 ;
  assign n21853 = ( n1118 & ~n6204 ) | ( n1118 & n12670 ) | ( ~n6204 & n12670 ) ;
  assign n21854 = n1904 & n7512 ;
  assign n21855 = n21854 ^ n1136 ^ 1'b0 ;
  assign n21856 = n21855 ^ n7692 ^ n4158 ;
  assign n21857 = n21856 ^ n1979 ^ 1'b0 ;
  assign n21858 = ( n2582 & ~n16768 ) | ( n2582 & n21857 ) | ( ~n16768 & n21857 ) ;
  assign n21859 = n19035 | n21858 ;
  assign n21860 = ( n5354 & ~n6746 ) | ( n5354 & n7589 ) | ( ~n6746 & n7589 ) ;
  assign n21861 = ( n702 & n1032 ) | ( n702 & n11189 ) | ( n1032 & n11189 ) ;
  assign n21862 = n21860 & n21861 ;
  assign n21863 = n21862 ^ n2591 ^ 1'b0 ;
  assign n21864 = n4156 | n14570 ;
  assign n21865 = ( n5755 & ~n21863 ) | ( n5755 & n21864 ) | ( ~n21863 & n21864 ) ;
  assign n21866 = n21865 ^ n18664 ^ n4084 ;
  assign n21867 = n17092 ^ n7540 ^ n2833 ;
  assign n21868 = ( n5237 & ~n10015 ) | ( n5237 & n21867 ) | ( ~n10015 & n21867 ) ;
  assign n21869 = n21868 ^ n16980 ^ n2479 ;
  assign n21870 = n10502 ^ n7379 ^ n5782 ;
  assign n21871 = n8920 ^ n6204 ^ x192 ;
  assign n21872 = ( n8766 & n21870 ) | ( n8766 & ~n21871 ) | ( n21870 & ~n21871 ) ;
  assign n21873 = ( n13452 & n21869 ) | ( n13452 & ~n21872 ) | ( n21869 & ~n21872 ) ;
  assign n21874 = n16147 ^ n9086 ^ n2566 ;
  assign n21875 = n18634 ^ n4924 ^ n2671 ;
  assign n21876 = ( n3355 & n7029 ) | ( n3355 & ~n11952 ) | ( n7029 & ~n11952 ) ;
  assign n21877 = ( n7684 & ~n12438 ) | ( n7684 & n21876 ) | ( ~n12438 & n21876 ) ;
  assign n21882 = n4948 & ~n7426 ;
  assign n21883 = n21882 ^ n4797 ^ 1'b0 ;
  assign n21884 = ( ~n13074 & n19477 ) | ( ~n13074 & n21883 ) | ( n19477 & n21883 ) ;
  assign n21880 = n19633 ^ n9585 ^ n3363 ;
  assign n21878 = n18195 ^ n12727 ^ 1'b0 ;
  assign n21879 = ( ~n8579 & n16036 ) | ( ~n8579 & n21878 ) | ( n16036 & n21878 ) ;
  assign n21881 = n21880 ^ n21879 ^ 1'b0 ;
  assign n21885 = n21884 ^ n21881 ^ n1131 ;
  assign n21890 = ( n821 & ~n12023 ) | ( n821 & n13282 ) | ( ~n12023 & n13282 ) ;
  assign n21887 = n12141 ^ n760 ^ x154 ;
  assign n21886 = n557 & ~n11281 ;
  assign n21888 = n21887 ^ n21886 ^ 1'b0 ;
  assign n21889 = ( n12918 & ~n16321 ) | ( n12918 & n21888 ) | ( ~n16321 & n21888 ) ;
  assign n21891 = n21890 ^ n21889 ^ n1095 ;
  assign n21895 = n16690 ^ n16109 ^ n4990 ;
  assign n21894 = n15269 ^ n11935 ^ n3718 ;
  assign n21892 = ~n835 & n14763 ;
  assign n21893 = n21892 ^ n5377 ^ n4251 ;
  assign n21896 = n21895 ^ n21894 ^ n21893 ;
  assign n21897 = n9743 & n12737 ;
  assign n21898 = n12942 ^ n11141 ^ n1531 ;
  assign n21899 = ~n2914 & n16336 ;
  assign n21900 = n21899 ^ n8409 ^ 1'b0 ;
  assign n21901 = n21898 & ~n21900 ;
  assign n21902 = n21901 ^ n13644 ^ 1'b0 ;
  assign n21903 = ~n16799 & n21902 ;
  assign n21904 = ( n1022 & n6911 ) | ( n1022 & n18503 ) | ( n6911 & n18503 ) ;
  assign n21905 = n21904 ^ n15515 ^ n430 ;
  assign n21906 = n21905 ^ n13175 ^ n1159 ;
  assign n21907 = ( n3699 & ~n3957 ) | ( n3699 & n17180 ) | ( ~n3957 & n17180 ) ;
  assign n21911 = ( ~n1152 & n1902 ) | ( ~n1152 & n4637 ) | ( n1902 & n4637 ) ;
  assign n21908 = ~n7002 & n8398 ;
  assign n21909 = n21908 ^ n14313 ^ 1'b0 ;
  assign n21910 = ~n11234 & n21909 ;
  assign n21912 = n21911 ^ n21910 ^ 1'b0 ;
  assign n21913 = n21912 ^ n14728 ^ n5583 ;
  assign n21914 = ( ~n18743 & n21907 ) | ( ~n18743 & n21913 ) | ( n21907 & n21913 ) ;
  assign n21916 = ( ~n1139 & n12801 ) | ( ~n1139 & n15618 ) | ( n12801 & n15618 ) ;
  assign n21915 = n7628 & n12635 ;
  assign n21917 = n21916 ^ n21915 ^ 1'b0 ;
  assign n21918 = n5570 ^ n767 ^ 1'b0 ;
  assign n21919 = ~n16827 & n21918 ;
  assign n21920 = n2654 & n9279 ;
  assign n21921 = n2074 & n21920 ;
  assign n21922 = n4717 | n21921 ;
  assign n21923 = n21919 | n21922 ;
  assign n21924 = n14258 ^ n7207 ^ n5097 ;
  assign n21925 = ( n5819 & n7354 ) | ( n5819 & n16376 ) | ( n7354 & n16376 ) ;
  assign n21926 = n1692 & ~n5415 ;
  assign n21927 = n21926 ^ n9983 ^ 1'b0 ;
  assign n21928 = ( n5581 & ~n20784 ) | ( n5581 & n21927 ) | ( ~n20784 & n21927 ) ;
  assign n21929 = n15582 & ~n21928 ;
  assign n21930 = n19388 & n21929 ;
  assign n21931 = ( n10845 & n21925 ) | ( n10845 & n21930 ) | ( n21925 & n21930 ) ;
  assign n21933 = n1075 ^ n768 ^ 1'b0 ;
  assign n21932 = ~n4994 & n9066 ;
  assign n21934 = n21933 ^ n21932 ^ n18959 ;
  assign n21935 = n14872 | n21934 ;
  assign n21936 = n13877 ^ n10393 ^ n1272 ;
  assign n21937 = ( n5669 & ~n8595 ) | ( n5669 & n9284 ) | ( ~n8595 & n9284 ) ;
  assign n21938 = ( n14854 & ~n21936 ) | ( n14854 & n21937 ) | ( ~n21936 & n21937 ) ;
  assign n21939 = n4502 ^ n2992 ^ n1316 ;
  assign n21940 = n21939 ^ n13457 ^ n7492 ;
  assign n21941 = ( n2404 & n3478 ) | ( n2404 & ~n3981 ) | ( n3478 & ~n3981 ) ;
  assign n21942 = ( n523 & n21940 ) | ( n523 & ~n21941 ) | ( n21940 & ~n21941 ) ;
  assign n21943 = n18783 & n21349 ;
  assign n21944 = ~n3190 & n21943 ;
  assign n21945 = ( n7791 & n15079 ) | ( n7791 & ~n21944 ) | ( n15079 & ~n21944 ) ;
  assign n21946 = ( ~n20019 & n21942 ) | ( ~n20019 & n21945 ) | ( n21942 & n21945 ) ;
  assign n21947 = n9668 ^ n3143 ^ x245 ;
  assign n21948 = n21947 ^ n15992 ^ n6720 ;
  assign n21949 = n21948 ^ n11729 ^ 1'b0 ;
  assign n21950 = ( n8293 & ~n14326 ) | ( n8293 & n18012 ) | ( ~n14326 & n18012 ) ;
  assign n21951 = n15617 ^ n9617 ^ n1722 ;
  assign n21952 = n5797 & ~n21951 ;
  assign n21953 = ~n21950 & n21952 ;
  assign n21954 = n12668 | n19829 ;
  assign n21955 = n21954 ^ n9482 ^ 1'b0 ;
  assign n21956 = n21955 ^ n11491 ^ n4868 ;
  assign n21957 = ( x152 & ~n2640 ) | ( x152 & n11739 ) | ( ~n2640 & n11739 ) ;
  assign n21958 = n21957 ^ n6800 ^ 1'b0 ;
  assign n21959 = ~n5296 & n21958 ;
  assign n21960 = ( n2827 & n5870 ) | ( n2827 & ~n7713 ) | ( n5870 & ~n7713 ) ;
  assign n21961 = ( ~n1714 & n6915 ) | ( ~n1714 & n8307 ) | ( n6915 & n8307 ) ;
  assign n21962 = n21960 & ~n21961 ;
  assign n21970 = ( x67 & n5055 ) | ( x67 & n7240 ) | ( n5055 & n7240 ) ;
  assign n21963 = ( n620 & n4993 ) | ( n620 & ~n7178 ) | ( n4993 & ~n7178 ) ;
  assign n21966 = n7874 ^ n3239 ^ n2987 ;
  assign n21964 = n4508 ^ n3695 ^ 1'b0 ;
  assign n21965 = n6739 & n21964 ;
  assign n21967 = n21966 ^ n21965 ^ n13692 ;
  assign n21968 = n21963 & ~n21967 ;
  assign n21969 = ~n1756 & n21968 ;
  assign n21971 = n21970 ^ n21969 ^ n8102 ;
  assign n21972 = ( n6330 & n6390 ) | ( n6330 & n6856 ) | ( n6390 & n6856 ) ;
  assign n21973 = ( ~n3982 & n10356 ) | ( ~n3982 & n21972 ) | ( n10356 & n21972 ) ;
  assign n21974 = ( n18212 & n21971 ) | ( n18212 & n21973 ) | ( n21971 & n21973 ) ;
  assign n21975 = n21974 ^ n20460 ^ n9278 ;
  assign n21976 = n8555 ^ n4895 ^ 1'b0 ;
  assign n21979 = ( n1704 & n4628 ) | ( n1704 & n13884 ) | ( n4628 & n13884 ) ;
  assign n21978 = ( n1624 & ~n2217 ) | ( n1624 & n8279 ) | ( ~n2217 & n8279 ) ;
  assign n21977 = ( n13176 & ~n16644 ) | ( n13176 & n20822 ) | ( ~n16644 & n20822 ) ;
  assign n21980 = n21979 ^ n21978 ^ n21977 ;
  assign n21982 = n6970 ^ n1453 ^ 1'b0 ;
  assign n21983 = n21982 ^ n6389 ^ x141 ;
  assign n21981 = ~n399 & n8957 ;
  assign n21984 = n21983 ^ n21981 ^ 1'b0 ;
  assign n21985 = n21984 ^ n3309 ^ 1'b0 ;
  assign n21986 = n1370 & n21985 ;
  assign n21987 = n21986 ^ n9583 ^ n1293 ;
  assign n21988 = ( ~n21976 & n21980 ) | ( ~n21976 & n21987 ) | ( n21980 & n21987 ) ;
  assign n21989 = ( ~n2453 & n4219 ) | ( ~n2453 & n6981 ) | ( n4219 & n6981 ) ;
  assign n21990 = ( n16250 & n20770 ) | ( n16250 & n21989 ) | ( n20770 & n21989 ) ;
  assign n21991 = n21983 ^ n12585 ^ n2772 ;
  assign n21992 = n5546 | n15828 ;
  assign n21993 = n10057 & ~n10167 ;
  assign n21994 = ~n12665 & n21288 ;
  assign n21995 = n21994 ^ n982 ^ 1'b0 ;
  assign n21996 = n21995 ^ n17487 ^ n2835 ;
  assign n21997 = n18203 ^ n8946 ^ n3720 ;
  assign n21998 = ( n3793 & n3951 ) | ( n3793 & ~n7546 ) | ( n3951 & ~n7546 ) ;
  assign n21999 = n21997 | n21998 ;
  assign n22000 = n21996 & ~n21999 ;
  assign n22001 = n15741 ^ n14287 ^ n4489 ;
  assign n22005 = n8905 & n14123 ;
  assign n22002 = n2113 & ~n12102 ;
  assign n22003 = n22002 ^ n14593 ^ n9505 ;
  assign n22004 = n22003 ^ n2649 ^ 1'b0 ;
  assign n22006 = n22005 ^ n22004 ^ n16469 ;
  assign n22010 = n17087 ^ n3836 ^ 1'b0 ;
  assign n22008 = ( n12107 & ~n13860 ) | ( n12107 & n17070 ) | ( ~n13860 & n17070 ) ;
  assign n22009 = n17781 | n22008 ;
  assign n22007 = ( ~n2081 & n15362 ) | ( ~n2081 & n15484 ) | ( n15362 & n15484 ) ;
  assign n22011 = n22010 ^ n22009 ^ n22007 ;
  assign n22012 = ( n5462 & n5710 ) | ( n5462 & n19002 ) | ( n5710 & n19002 ) ;
  assign n22013 = n15822 ^ n5574 ^ 1'b0 ;
  assign n22014 = ~n11841 & n22013 ;
  assign n22015 = ~n22012 & n22014 ;
  assign n22016 = n22015 ^ n18452 ^ n11302 ;
  assign n22017 = ( n6185 & n17509 ) | ( n6185 & ~n22016 ) | ( n17509 & ~n22016 ) ;
  assign n22018 = ( n7638 & n9155 ) | ( n7638 & ~n14382 ) | ( n9155 & ~n14382 ) ;
  assign n22019 = n22018 ^ n19014 ^ n13728 ;
  assign n22020 = ~n13251 & n22019 ;
  assign n22026 = n11203 ^ x144 ^ 1'b0 ;
  assign n22023 = n3725 ^ x157 ^ 1'b0 ;
  assign n22022 = n20498 ^ n2939 ^ 1'b0 ;
  assign n22021 = n19110 ^ n9902 ^ 1'b0 ;
  assign n22024 = n22023 ^ n22022 ^ n22021 ;
  assign n22025 = ( n2258 & n15661 ) | ( n2258 & ~n22024 ) | ( n15661 & ~n22024 ) ;
  assign n22027 = n22026 ^ n22025 ^ x27 ;
  assign n22028 = n11924 ^ n766 ^ 1'b0 ;
  assign n22029 = ~n19530 & n22028 ;
  assign n22030 = ~n623 & n15648 ;
  assign n22031 = n22030 ^ n3189 ^ 1'b0 ;
  assign n22032 = n22031 ^ n7990 ^ 1'b0 ;
  assign n22033 = n22032 ^ n19226 ^ n17229 ;
  assign n22034 = n22029 | n22033 ;
  assign n22035 = ( n8427 & n16268 ) | ( n8427 & n20755 ) | ( n16268 & n20755 ) ;
  assign n22036 = n22035 ^ n5769 ^ n4004 ;
  assign n22037 = n9141 & n10444 ;
  assign n22038 = ~n7984 & n22037 ;
  assign n22039 = n14759 ^ n269 ^ 1'b0 ;
  assign n22040 = ~n22038 & n22039 ;
  assign n22041 = n22040 ^ n15371 ^ 1'b0 ;
  assign n22042 = ( ~n19081 & n22036 ) | ( ~n19081 & n22041 ) | ( n22036 & n22041 ) ;
  assign n22043 = n858 | n17728 ;
  assign n22044 = n17166 & ~n22043 ;
  assign n22045 = n1731 & n12159 ;
  assign n22046 = n22045 ^ n11135 ^ 1'b0 ;
  assign n22047 = ( n7361 & ~n7366 ) | ( n7361 & n9053 ) | ( ~n7366 & n9053 ) ;
  assign n22048 = n1398 & ~n18185 ;
  assign n22049 = n22048 ^ n8629 ^ 1'b0 ;
  assign n22050 = n22049 ^ n13110 ^ n8464 ;
  assign n22051 = ~n12545 & n16920 ;
  assign n22052 = n16700 ^ n12025 ^ n1896 ;
  assign n22053 = n959 & ~n3287 ;
  assign n22054 = n22052 & n22053 ;
  assign n22055 = n951 | n4530 ;
  assign n22056 = ( ~n6303 & n15657 ) | ( ~n6303 & n22055 ) | ( n15657 & n22055 ) ;
  assign n22057 = n22056 ^ n13658 ^ n3048 ;
  assign n22058 = n22057 ^ n3052 ^ n663 ;
  assign n22059 = ~n6026 & n22058 ;
  assign n22060 = n22059 ^ n7786 ^ 1'b0 ;
  assign n22061 = ( n371 & n17742 ) | ( n371 & n22060 ) | ( n17742 & n22060 ) ;
  assign n22062 = n4941 ^ n1512 ^ 1'b0 ;
  assign n22063 = n2459 & n22062 ;
  assign n22064 = ( ~n1724 & n5270 ) | ( ~n1724 & n22063 ) | ( n5270 & n22063 ) ;
  assign n22065 = n22064 ^ n9782 ^ n962 ;
  assign n22066 = ( n7947 & n16672 ) | ( n7947 & ~n22065 ) | ( n16672 & ~n22065 ) ;
  assign n22067 = n22066 ^ n9865 ^ n4859 ;
  assign n22068 = ( n11622 & n20254 ) | ( n11622 & n22067 ) | ( n20254 & n22067 ) ;
  assign n22069 = ( n702 & n6401 ) | ( n702 & n12089 ) | ( n6401 & n12089 ) ;
  assign n22070 = n22069 ^ n716 ^ 1'b0 ;
  assign n22071 = n22068 & n22070 ;
  assign n22072 = ( n22061 & ~n22067 ) | ( n22061 & n22071 ) | ( ~n22067 & n22071 ) ;
  assign n22075 = n10711 ^ n5710 ^ 1'b0 ;
  assign n22073 = n8449 & ~n11809 ;
  assign n22074 = n22073 ^ n16195 ^ 1'b0 ;
  assign n22076 = n22075 ^ n22074 ^ n4347 ;
  assign n22077 = ( n7085 & ~n14107 ) | ( n7085 & n14356 ) | ( ~n14107 & n14356 ) ;
  assign n22078 = n22077 ^ n2258 ^ 1'b0 ;
  assign n22079 = n19310 & n22078 ;
  assign n22080 = ( ~n4209 & n4863 ) | ( ~n4209 & n5930 ) | ( n4863 & n5930 ) ;
  assign n22081 = n22080 ^ n18548 ^ 1'b0 ;
  assign n22082 = n11401 & ~n22081 ;
  assign n22087 = n17201 ^ n12737 ^ 1'b0 ;
  assign n22088 = n16689 | n22087 ;
  assign n22089 = n2931 & ~n22088 ;
  assign n22083 = n19956 ^ n12044 ^ 1'b0 ;
  assign n22084 = ( ~n1811 & n3366 ) | ( ~n1811 & n8872 ) | ( n3366 & n8872 ) ;
  assign n22085 = n22083 & ~n22084 ;
  assign n22086 = n844 & n22085 ;
  assign n22090 = n22089 ^ n22086 ^ n1082 ;
  assign n22091 = n11928 & ~n16136 ;
  assign n22092 = n18639 ^ n15422 ^ 1'b0 ;
  assign n22093 = n3359 & n6169 ;
  assign n22094 = ~n2659 & n22093 ;
  assign n22095 = n22094 ^ n3932 ^ 1'b0 ;
  assign n22096 = ( n9586 & ~n12173 ) | ( n9586 & n22095 ) | ( ~n12173 & n22095 ) ;
  assign n22097 = n1527 ^ x4 ^ 1'b0 ;
  assign n22098 = ( x55 & ~n6569 ) | ( x55 & n22097 ) | ( ~n6569 & n22097 ) ;
  assign n22099 = ~n4131 & n14113 ;
  assign n22100 = n22098 & n22099 ;
  assign n22101 = n8923 ^ n1291 ^ 1'b0 ;
  assign n22102 = n6848 & n22101 ;
  assign n22103 = n22100 & n22102 ;
  assign n22104 = n17683 ^ n10045 ^ 1'b0 ;
  assign n22105 = n12972 ^ n587 ^ 1'b0 ;
  assign n22106 = ( n2801 & ~n7235 ) | ( n2801 & n20715 ) | ( ~n7235 & n20715 ) ;
  assign n22112 = ( n892 & ~n959 ) | ( n892 & n9097 ) | ( ~n959 & n9097 ) ;
  assign n22107 = n1257 & n3975 ;
  assign n22108 = ( n7224 & n9655 ) | ( n7224 & ~n16185 ) | ( n9655 & ~n16185 ) ;
  assign n22109 = ~n14421 & n22108 ;
  assign n22110 = n22109 ^ n3538 ^ 1'b0 ;
  assign n22111 = n22107 | n22110 ;
  assign n22113 = n22112 ^ n22111 ^ 1'b0 ;
  assign n22114 = ( n9225 & n16269 ) | ( n9225 & ~n22113 ) | ( n16269 & ~n22113 ) ;
  assign n22115 = n2514 | n22114 ;
  assign n22116 = n20730 & ~n22115 ;
  assign n22117 = n2646 | n8681 ;
  assign n22118 = n2465 & ~n10463 ;
  assign n22119 = n22118 ^ n12026 ^ 1'b0 ;
  assign n22120 = n9698 ^ n5162 ^ n1450 ;
  assign n22121 = ( n2364 & n11465 ) | ( n2364 & n22120 ) | ( n11465 & n22120 ) ;
  assign n22122 = ( ~n1055 & n3268 ) | ( ~n1055 & n11867 ) | ( n3268 & n11867 ) ;
  assign n22123 = ( n22119 & n22121 ) | ( n22119 & ~n22122 ) | ( n22121 & ~n22122 ) ;
  assign n22125 = ( n1807 & ~n3231 ) | ( n1807 & n5065 ) | ( ~n3231 & n5065 ) ;
  assign n22126 = n15982 | n22125 ;
  assign n22124 = n2985 & ~n15703 ;
  assign n22127 = n22126 ^ n22124 ^ n1606 ;
  assign n22136 = n2628 ^ n2037 ^ 1'b0 ;
  assign n22137 = n2188 & ~n22136 ;
  assign n22133 = n1787 & ~n6059 ;
  assign n22134 = n775 & n22133 ;
  assign n22135 = n1895 & ~n22134 ;
  assign n22138 = n22137 ^ n22135 ^ 1'b0 ;
  assign n22139 = n2448 & ~n22138 ;
  assign n22132 = n12384 ^ n11385 ^ n3249 ;
  assign n22129 = n9009 & ~n10785 ;
  assign n22130 = n7539 & n22129 ;
  assign n22128 = ~n415 & n1455 ;
  assign n22131 = n22130 ^ n22128 ^ n9225 ;
  assign n22140 = n22139 ^ n22132 ^ n22131 ;
  assign n22141 = n22140 ^ n21678 ^ n5056 ;
  assign n22142 = ( ~n12204 & n21421 ) | ( ~n12204 & n21604 ) | ( n21421 & n21604 ) ;
  assign n22143 = n6273 | n22142 ;
  assign n22144 = n22143 ^ n9146 ^ 1'b0 ;
  assign n22146 = n14462 & ~n14945 ;
  assign n22147 = ~n4329 & n22146 ;
  assign n22145 = ( n1107 & n2109 ) | ( n1107 & n9474 ) | ( n2109 & n9474 ) ;
  assign n22148 = n22147 ^ n22145 ^ n282 ;
  assign n22149 = ( n7836 & ~n10796 ) | ( n7836 & n13112 ) | ( ~n10796 & n13112 ) ;
  assign n22150 = n19431 ^ n13569 ^ 1'b0 ;
  assign n22151 = n15780 & n22150 ;
  assign n22152 = ~n4298 & n15195 ;
  assign n22153 = n22152 ^ n1827 ^ 1'b0 ;
  assign n22154 = n7153 ^ n1443 ^ 1'b0 ;
  assign n22155 = ~n22153 & n22154 ;
  assign n22156 = n17901 ^ n16956 ^ n5772 ;
  assign n22159 = n18236 ^ n1828 ^ 1'b0 ;
  assign n22160 = ( n5966 & ~n8082 ) | ( n5966 & n22159 ) | ( ~n8082 & n22159 ) ;
  assign n22157 = n15923 ^ n2258 ^ n820 ;
  assign n22158 = n22157 ^ n9328 ^ x124 ;
  assign n22161 = n22160 ^ n22158 ^ n16533 ;
  assign n22162 = n4080 & n19640 ;
  assign n22163 = n22162 ^ n14473 ^ 1'b0 ;
  assign n22164 = n9972 | n22163 ;
  assign n22165 = n18335 | n22164 ;
  assign n22166 = n1873 & ~n7140 ;
  assign n22167 = n22166 ^ n1414 ^ 1'b0 ;
  assign n22168 = ( n1597 & ~n15266 ) | ( n1597 & n19907 ) | ( ~n15266 & n19907 ) ;
  assign n22169 = n17682 ^ n6852 ^ 1'b0 ;
  assign n22170 = ( ~n3350 & n5153 ) | ( ~n3350 & n5284 ) | ( n5153 & n5284 ) ;
  assign n22171 = n22170 ^ n19365 ^ n1365 ;
  assign n22172 = ( ~n1370 & n22169 ) | ( ~n1370 & n22171 ) | ( n22169 & n22171 ) ;
  assign n22173 = n22172 ^ n13735 ^ n2954 ;
  assign n22174 = n3495 ^ n1858 ^ n364 ;
  assign n22175 = n7047 ^ n3479 ^ 1'b0 ;
  assign n22176 = n22175 ^ n7348 ^ n694 ;
  assign n22177 = ( n441 & ~n22174 ) | ( n441 & n22176 ) | ( ~n22174 & n22176 ) ;
  assign n22178 = n10757 | n13592 ;
  assign n22179 = n22178 ^ n5774 ^ 1'b0 ;
  assign n22180 = n22179 ^ n11399 ^ n2161 ;
  assign n22181 = n16750 ^ n6714 ^ n5004 ;
  assign n22182 = ( ~n18592 & n22180 ) | ( ~n18592 & n22181 ) | ( n22180 & n22181 ) ;
  assign n22184 = n15199 ^ n14659 ^ n5834 ;
  assign n22185 = ( n4730 & n13745 ) | ( n4730 & n22184 ) | ( n13745 & n22184 ) ;
  assign n22183 = n9350 & ~n16004 ;
  assign n22186 = n22185 ^ n22183 ^ 1'b0 ;
  assign n22187 = n3453 ^ n2998 ^ n997 ;
  assign n22188 = ( n1840 & n9323 ) | ( n1840 & n22187 ) | ( n9323 & n22187 ) ;
  assign n22189 = ( n5741 & n9902 ) | ( n5741 & n11114 ) | ( n9902 & n11114 ) ;
  assign n22190 = n22189 ^ n17127 ^ n549 ;
  assign n22191 = n17446 ^ n2278 ^ n1272 ;
  assign n22192 = n7639 & ~n18276 ;
  assign n22193 = ( ~n20727 & n22191 ) | ( ~n20727 & n22192 ) | ( n22191 & n22192 ) ;
  assign n22194 = ~n9157 & n17776 ;
  assign n22195 = n2066 & n22194 ;
  assign n22196 = ( ~n8410 & n15483 ) | ( ~n8410 & n21235 ) | ( n15483 & n21235 ) ;
  assign n22197 = n22196 ^ n10645 ^ 1'b0 ;
  assign n22198 = ~n4186 & n22197 ;
  assign n22201 = n19226 ^ n9149 ^ n6351 ;
  assign n22199 = ( n3169 & n5505 ) | ( n3169 & n7468 ) | ( n5505 & n7468 ) ;
  assign n22200 = ( n2026 & n2064 ) | ( n2026 & n22199 ) | ( n2064 & n22199 ) ;
  assign n22202 = n22201 ^ n22200 ^ n9156 ;
  assign n22203 = n22202 ^ n7418 ^ n5089 ;
  assign n22204 = n5238 ^ n697 ^ 1'b0 ;
  assign n22205 = ~n18363 & n22204 ;
  assign n22206 = n12506 ^ n9718 ^ n2092 ;
  assign n22207 = ( ~n413 & n1288 ) | ( ~n413 & n22206 ) | ( n1288 & n22206 ) ;
  assign n22208 = n17180 ^ n6076 ^ n3451 ;
  assign n22209 = n9842 ^ n2638 ^ 1'b0 ;
  assign n22210 = n2196 | n22209 ;
  assign n22211 = n16890 ^ n11103 ^ n9268 ;
  assign n22212 = ( ~n22208 & n22210 ) | ( ~n22208 & n22211 ) | ( n22210 & n22211 ) ;
  assign n22213 = n15935 ^ n2413 ^ 1'b0 ;
  assign n22216 = n3246 ^ n2920 ^ x43 ;
  assign n22217 = n2275 | n11871 ;
  assign n22218 = n22217 ^ n21808 ^ 1'b0 ;
  assign n22219 = n22218 ^ n16986 ^ n5872 ;
  assign n22220 = ( ~n10487 & n22216 ) | ( ~n10487 & n22219 ) | ( n22216 & n22219 ) ;
  assign n22214 = n20018 ^ n3660 ^ 1'b0 ;
  assign n22215 = n18917 & n22214 ;
  assign n22221 = n22220 ^ n22215 ^ n4029 ;
  assign n22222 = ( ~n2554 & n14287 ) | ( ~n2554 & n22221 ) | ( n14287 & n22221 ) ;
  assign n22229 = ( n5090 & n7603 ) | ( n5090 & n17663 ) | ( n7603 & n17663 ) ;
  assign n22223 = n7181 ^ n4491 ^ 1'b0 ;
  assign n22224 = n4417 | n22223 ;
  assign n22225 = n20871 ^ n3115 ^ 1'b0 ;
  assign n22226 = ~n383 & n22225 ;
  assign n22227 = n22226 ^ n11980 ^ n2066 ;
  assign n22228 = ( n7723 & ~n22224 ) | ( n7723 & n22227 ) | ( ~n22224 & n22227 ) ;
  assign n22230 = n22229 ^ n22228 ^ n17450 ;
  assign n22232 = n8170 | n14034 ;
  assign n22231 = ( n2491 & n3625 ) | ( n2491 & ~n16565 ) | ( n3625 & ~n16565 ) ;
  assign n22233 = n22232 ^ n22231 ^ n3314 ;
  assign n22234 = n3300 & ~n22233 ;
  assign n22235 = ~n11869 & n19753 ;
  assign n22236 = n12904 & n22235 ;
  assign n22237 = ~n2966 & n9630 ;
  assign n22238 = ( n3562 & n5742 ) | ( n3562 & ~n8647 ) | ( n5742 & ~n8647 ) ;
  assign n22239 = n8567 & ~n22238 ;
  assign n22240 = n22237 & n22239 ;
  assign n22241 = n9832 ^ n7962 ^ n7542 ;
  assign n22242 = n6344 ^ n1722 ^ n905 ;
  assign n22243 = ( ~n7674 & n14751 ) | ( ~n7674 & n22242 ) | ( n14751 & n22242 ) ;
  assign n22244 = n14070 ^ n8666 ^ 1'b0 ;
  assign n22245 = ~n536 & n22244 ;
  assign n22246 = ( n903 & ~n12665 ) | ( n903 & n22245 ) | ( ~n12665 & n22245 ) ;
  assign n22247 = ~n11605 & n19690 ;
  assign n22248 = ( n22243 & ~n22246 ) | ( n22243 & n22247 ) | ( ~n22246 & n22247 ) ;
  assign n22256 = n20295 ^ n6264 ^ n4793 ;
  assign n22257 = ( x206 & n15213 ) | ( x206 & ~n22256 ) | ( n15213 & ~n22256 ) ;
  assign n22249 = n7383 ^ n7042 ^ n5402 ;
  assign n22250 = ~n14965 & n21132 ;
  assign n22251 = n22249 & n22250 ;
  assign n22252 = ( n1107 & n8193 ) | ( n1107 & ~n22251 ) | ( n8193 & ~n22251 ) ;
  assign n22253 = n22252 ^ n11736 ^ n691 ;
  assign n22254 = n16096 ^ n4637 ^ 1'b0 ;
  assign n22255 = n22253 & n22254 ;
  assign n22258 = n22257 ^ n22255 ^ n17816 ;
  assign n22259 = ( n2575 & n15419 ) | ( n2575 & ~n21814 ) | ( n15419 & ~n21814 ) ;
  assign n22260 = n16118 ^ n12472 ^ n12411 ;
  assign n22261 = n11894 ^ n7198 ^ n5997 ;
  assign n22262 = n4464 & ~n22261 ;
  assign n22263 = ( n3876 & n6297 ) | ( n3876 & n7367 ) | ( n6297 & n7367 ) ;
  assign n22264 = ( n8971 & n11105 ) | ( n8971 & n22263 ) | ( n11105 & n22263 ) ;
  assign n22265 = ( n6477 & n11606 ) | ( n6477 & ~n22264 ) | ( n11606 & ~n22264 ) ;
  assign n22279 = n5402 ^ n1914 ^ 1'b0 ;
  assign n22276 = n9605 ^ n3637 ^ n1313 ;
  assign n22277 = ( n3287 & n13407 ) | ( n3287 & n22276 ) | ( n13407 & n22276 ) ;
  assign n22278 = n22277 ^ n15906 ^ n7454 ;
  assign n22266 = ~n6617 & n21982 ;
  assign n22267 = n22266 ^ n16884 ^ n14921 ;
  assign n22268 = ~n5526 & n22267 ;
  assign n22269 = n22268 ^ n4788 ^ 1'b0 ;
  assign n22270 = ( n681 & ~n10457 ) | ( n681 & n12667 ) | ( ~n10457 & n12667 ) ;
  assign n22271 = ( ~x97 & n8286 ) | ( ~x97 & n18109 ) | ( n8286 & n18109 ) ;
  assign n22272 = n5656 & n10524 ;
  assign n22273 = n22271 & n22272 ;
  assign n22274 = ( n10524 & n22270 ) | ( n10524 & n22273 ) | ( n22270 & n22273 ) ;
  assign n22275 = ( n2120 & n22269 ) | ( n2120 & ~n22274 ) | ( n22269 & ~n22274 ) ;
  assign n22280 = n22279 ^ n22278 ^ n22275 ;
  assign n22281 = ( ~n2680 & n3548 ) | ( ~n2680 & n4415 ) | ( n3548 & n4415 ) ;
  assign n22282 = ( ~n2066 & n3973 ) | ( ~n2066 & n5546 ) | ( n3973 & n5546 ) ;
  assign n22283 = n10289 | n11030 ;
  assign n22284 = n2814 & ~n22283 ;
  assign n22285 = ( n849 & n22282 ) | ( n849 & n22284 ) | ( n22282 & n22284 ) ;
  assign n22286 = ( n15648 & ~n22281 ) | ( n15648 & n22285 ) | ( ~n22281 & n22285 ) ;
  assign n22294 = n9844 ^ n6473 ^ 1'b0 ;
  assign n22293 = ( n10946 & n14154 ) | ( n10946 & ~n15034 ) | ( n14154 & ~n15034 ) ;
  assign n22290 = n1143 & n12652 ;
  assign n22291 = n22290 ^ n17543 ^ 1'b0 ;
  assign n22287 = ( n688 & n2804 ) | ( n688 & n5194 ) | ( n2804 & n5194 ) ;
  assign n22288 = n22287 ^ n15716 ^ 1'b0 ;
  assign n22289 = n22288 ^ n6160 ^ n476 ;
  assign n22292 = n22291 ^ n22289 ^ n17363 ;
  assign n22295 = n22294 ^ n22293 ^ n22292 ;
  assign n22296 = n5917 & n7406 ;
  assign n22297 = n22296 ^ n8534 ^ 1'b0 ;
  assign n22298 = n19691 | n22297 ;
  assign n22299 = n4359 | n22298 ;
  assign n22303 = n2709 & ~n19997 ;
  assign n22300 = n18083 ^ n15314 ^ n4100 ;
  assign n22301 = n17563 ^ n749 ^ n296 ;
  assign n22302 = n22300 & ~n22301 ;
  assign n22304 = n22303 ^ n22302 ^ 1'b0 ;
  assign n22305 = n21044 ^ n13003 ^ n757 ;
  assign n22306 = n5672 ^ n3506 ^ n847 ;
  assign n22307 = n9467 & n19929 ;
  assign n22308 = n22307 ^ n5512 ^ n5498 ;
  assign n22309 = ( n2124 & n18489 ) | ( n2124 & ~n22308 ) | ( n18489 & ~n22308 ) ;
  assign n22310 = ( n2424 & n7469 ) | ( n2424 & n22309 ) | ( n7469 & n22309 ) ;
  assign n22311 = ( ~n3958 & n14839 ) | ( ~n3958 & n22310 ) | ( n14839 & n22310 ) ;
  assign n22312 = n6137 ^ n5172 ^ 1'b0 ;
  assign n22313 = n699 & ~n22312 ;
  assign n22314 = n12718 ^ n4195 ^ n793 ;
  assign n22315 = ( ~n3298 & n21500 ) | ( ~n3298 & n22314 ) | ( n21500 & n22314 ) ;
  assign n22316 = ~n9217 & n13680 ;
  assign n22317 = n16178 ^ n14833 ^ n1208 ;
  assign n22321 = n11370 ^ n10513 ^ n939 ;
  assign n22318 = ~n3077 & n9401 ;
  assign n22319 = n22318 ^ n8059 ^ 1'b0 ;
  assign n22320 = n22319 ^ n17336 ^ n2842 ;
  assign n22322 = n22321 ^ n22320 ^ n5001 ;
  assign n22323 = n21083 ^ n3736 ^ n1990 ;
  assign n22324 = ( n19620 & ~n22322 ) | ( n19620 & n22323 ) | ( ~n22322 & n22323 ) ;
  assign n22325 = ( n11645 & ~n22317 ) | ( n11645 & n22324 ) | ( ~n22317 & n22324 ) ;
  assign n22326 = n16096 & n21326 ;
  assign n22327 = ~n12200 & n22326 ;
  assign n22328 = ( n9384 & ~n10269 ) | ( n9384 & n22327 ) | ( ~n10269 & n22327 ) ;
  assign n22329 = ( n1675 & n16267 ) | ( n1675 & ~n22328 ) | ( n16267 & ~n22328 ) ;
  assign n22330 = n20169 ^ n14518 ^ n3169 ;
  assign n22331 = ( n406 & n8081 ) | ( n406 & ~n22330 ) | ( n8081 & ~n22330 ) ;
  assign n22332 = n19704 | n22331 ;
  assign n22333 = n22329 | n22332 ;
  assign n22334 = n17973 ^ n3391 ^ 1'b0 ;
  assign n22335 = n2173 & ~n22334 ;
  assign n22336 = n22335 ^ n16267 ^ n8237 ;
  assign n22337 = n22336 ^ n2199 ^ 1'b0 ;
  assign n22338 = n15342 ^ n10531 ^ 1'b0 ;
  assign n22339 = n22337 & n22338 ;
  assign n22341 = n1463 ^ n1384 ^ x56 ;
  assign n22340 = ( n2682 & ~n8341 ) | ( n2682 & n11109 ) | ( ~n8341 & n11109 ) ;
  assign n22342 = n22341 ^ n22340 ^ n14762 ;
  assign n22348 = n4734 ^ n1939 ^ 1'b0 ;
  assign n22343 = n8611 | n13984 ;
  assign n22344 = n11936 | n22343 ;
  assign n22345 = n22344 ^ n22210 ^ 1'b0 ;
  assign n22346 = n10011 | n22345 ;
  assign n22347 = n22346 ^ n8678 ^ 1'b0 ;
  assign n22349 = n22348 ^ n22347 ^ n2897 ;
  assign n22351 = ( x48 & n2751 ) | ( x48 & n4464 ) | ( n2751 & n4464 ) ;
  assign n22350 = ( n3725 & n15943 ) | ( n3725 & ~n20991 ) | ( n15943 & ~n20991 ) ;
  assign n22352 = n22351 ^ n22350 ^ n15374 ;
  assign n22353 = n3028 & ~n8456 ;
  assign n22354 = n14913 ^ n14176 ^ 1'b0 ;
  assign n22355 = n11488 & ~n22354 ;
  assign n22356 = ( ~n14563 & n22353 ) | ( ~n14563 & n22355 ) | ( n22353 & n22355 ) ;
  assign n22357 = n6854 ^ n2162 ^ 1'b0 ;
  assign n22358 = n22357 ^ n8742 ^ 1'b0 ;
  assign n22359 = n9550 | n22358 ;
  assign n22360 = n2338 & ~n3302 ;
  assign n22361 = n1737 & n22360 ;
  assign n22362 = n22361 ^ n11507 ^ n4774 ;
  assign n22363 = n22362 ^ n17592 ^ n3094 ;
  assign n22364 = ~n4131 & n22363 ;
  assign n22365 = ~n8315 & n22364 ;
  assign n22366 = ( n3679 & n17418 ) | ( n3679 & n20601 ) | ( n17418 & n20601 ) ;
  assign n22367 = n13556 & ~n14421 ;
  assign n22368 = n22367 ^ n19407 ^ n8186 ;
  assign n22369 = ( n2471 & n8909 ) | ( n2471 & n16801 ) | ( n8909 & n16801 ) ;
  assign n22370 = ( n13869 & n16617 ) | ( n13869 & ~n22369 ) | ( n16617 & ~n22369 ) ;
  assign n22371 = n15078 ^ n4349 ^ n2900 ;
  assign n22372 = ( n5332 & n17891 ) | ( n5332 & n22371 ) | ( n17891 & n22371 ) ;
  assign n22373 = n16117 ^ n11118 ^ 1'b0 ;
  assign n22374 = ~n14145 & n22373 ;
  assign n22375 = ( n3526 & n6210 ) | ( n3526 & n22374 ) | ( n6210 & n22374 ) ;
  assign n22376 = ( n2494 & n11159 ) | ( n2494 & n12087 ) | ( n11159 & n12087 ) ;
  assign n22377 = n22376 ^ n19124 ^ n2578 ;
  assign n22378 = n22377 ^ n9182 ^ n4053 ;
  assign n22379 = ~n10514 & n20945 ;
  assign n22380 = n22379 ^ n4157 ^ 1'b0 ;
  assign n22381 = n3859 ^ n3284 ^ n874 ;
  assign n22382 = ( n3924 & n6286 ) | ( n3924 & n22381 ) | ( n6286 & n22381 ) ;
  assign n22383 = n22380 & n22382 ;
  assign n22384 = ( n2374 & n13117 ) | ( n2374 & ~n21829 ) | ( n13117 & ~n21829 ) ;
  assign n22385 = n22384 ^ n6479 ^ 1'b0 ;
  assign n22386 = n11372 ^ n11195 ^ n1724 ;
  assign n22387 = n20150 & ~n22386 ;
  assign n22395 = n20735 ^ n12718 ^ n5658 ;
  assign n22389 = ( n443 & ~n1253 ) | ( n443 & n10554 ) | ( ~n1253 & n10554 ) ;
  assign n22390 = ( n879 & n3629 ) | ( n879 & ~n22389 ) | ( n3629 & ~n22389 ) ;
  assign n22391 = n11780 | n22390 ;
  assign n22392 = ( ~n1639 & n7171 ) | ( ~n1639 & n22391 ) | ( n7171 & n22391 ) ;
  assign n22393 = n22392 ^ n12515 ^ n5100 ;
  assign n22394 = ( n7032 & ~n16755 ) | ( n7032 & n22393 ) | ( ~n16755 & n22393 ) ;
  assign n22388 = n21756 ^ n4120 ^ n2254 ;
  assign n22396 = n22395 ^ n22394 ^ n22388 ;
  assign n22397 = ( n4300 & n10850 ) | ( n4300 & ~n13191 ) | ( n10850 & ~n13191 ) ;
  assign n22398 = n22397 ^ n16492 ^ n3416 ;
  assign n22399 = n19246 ^ n3705 ^ 1'b0 ;
  assign n22404 = n15919 ^ n8867 ^ n8320 ;
  assign n22405 = n22404 ^ n1897 ^ n1691 ;
  assign n22402 = n15040 ^ n2996 ^ 1'b0 ;
  assign n22403 = n4016 & n22402 ;
  assign n22400 = n10093 ^ n5435 ^ 1'b0 ;
  assign n22401 = ~n21545 & n22400 ;
  assign n22406 = n22405 ^ n22403 ^ n22401 ;
  assign n22407 = n10077 ^ n6183 ^ n839 ;
  assign n22408 = n9761 & n21470 ;
  assign n22409 = n22407 & n22408 ;
  assign n22414 = n2609 | n7525 ;
  assign n22415 = n22414 ^ n18451 ^ 1'b0 ;
  assign n22410 = n10642 ^ n8269 ^ n3754 ;
  assign n22411 = n22410 ^ n17691 ^ n9818 ;
  assign n22412 = n4900 | n22411 ;
  assign n22413 = n22412 ^ n7749 ^ 1'b0 ;
  assign n22416 = n22415 ^ n22413 ^ n15488 ;
  assign n22417 = ( n3785 & n13799 ) | ( n3785 & ~n22276 ) | ( n13799 & ~n22276 ) ;
  assign n22418 = ( n706 & ~n12157 ) | ( n706 & n15419 ) | ( ~n12157 & n15419 ) ;
  assign n22419 = n22418 ^ n19289 ^ 1'b0 ;
  assign n22420 = ( n7479 & ~n22417 ) | ( n7479 & n22419 ) | ( ~n22417 & n22419 ) ;
  assign n22421 = n3194 & n4864 ;
  assign n22422 = n22421 ^ n4163 ^ 1'b0 ;
  assign n22423 = n1262 & n16400 ;
  assign n22424 = ~n7468 & n22423 ;
  assign n22425 = ( n16006 & n22422 ) | ( n16006 & ~n22424 ) | ( n22422 & ~n22424 ) ;
  assign n22426 = ( n3008 & n4190 ) | ( n3008 & ~n7918 ) | ( n4190 & ~n7918 ) ;
  assign n22427 = ( n1298 & n11270 ) | ( n1298 & n22426 ) | ( n11270 & n22426 ) ;
  assign n22428 = n12580 ^ n5771 ^ n2141 ;
  assign n22429 = n11014 & ~n22428 ;
  assign n22430 = n17604 ^ n6726 ^ n2286 ;
  assign n22431 = n22430 ^ n15624 ^ n5603 ;
  assign n22432 = ( n20688 & n22429 ) | ( n20688 & ~n22431 ) | ( n22429 & ~n22431 ) ;
  assign n22433 = n12335 ^ n11410 ^ 1'b0 ;
  assign n22434 = n5552 & ~n12097 ;
  assign n22435 = n22434 ^ n16610 ^ 1'b0 ;
  assign n22436 = n20316 ^ n13424 ^ 1'b0 ;
  assign n22437 = n14112 & ~n22436 ;
  assign n22438 = ~n19933 & n22437 ;
  assign n22439 = ( n3631 & n9780 ) | ( n3631 & n22438 ) | ( n9780 & n22438 ) ;
  assign n22440 = n5819 ^ n5702 ^ n3753 ;
  assign n22441 = n21733 ^ n13120 ^ n3258 ;
  assign n22442 = n18776 & ~n19584 ;
  assign n22443 = ~n10115 & n22442 ;
  assign n22444 = n22443 ^ n16984 ^ 1'b0 ;
  assign n22445 = n22441 & ~n22444 ;
  assign n22446 = n22445 ^ n11331 ^ 1'b0 ;
  assign n22447 = ( ~n2914 & n7259 ) | ( ~n2914 & n7300 ) | ( n7259 & n7300 ) ;
  assign n22448 = n19688 & n22447 ;
  assign n22449 = n22448 ^ n14510 ^ 1'b0 ;
  assign n22450 = n22449 ^ n2898 ^ 1'b0 ;
  assign n22451 = ~n1620 & n19555 ;
  assign n22452 = ~n22450 & n22451 ;
  assign n22453 = n13931 ^ n4298 ^ n3808 ;
  assign n22454 = ( ~n16227 & n17639 ) | ( ~n16227 & n22453 ) | ( n17639 & n22453 ) ;
  assign n22457 = n19791 ^ n12617 ^ n3675 ;
  assign n22455 = ( n3451 & ~n8636 ) | ( n3451 & n12953 ) | ( ~n8636 & n12953 ) ;
  assign n22456 = ( n1598 & ~n6745 ) | ( n1598 & n22455 ) | ( ~n6745 & n22455 ) ;
  assign n22458 = n22457 ^ n22456 ^ 1'b0 ;
  assign n22459 = n21493 ^ n10392 ^ n9755 ;
  assign n22460 = ( n5056 & n19413 ) | ( n5056 & n22459 ) | ( n19413 & n22459 ) ;
  assign n22461 = ( n1034 & ~n13140 ) | ( n1034 & n19405 ) | ( ~n13140 & n19405 ) ;
  assign n22462 = n12274 ^ n7573 ^ n927 ;
  assign n22463 = ( n2981 & n17507 ) | ( n2981 & n22462 ) | ( n17507 & n22462 ) ;
  assign n22464 = ( ~n3634 & n19484 ) | ( ~n3634 & n22463 ) | ( n19484 & n22463 ) ;
  assign n22465 = ( n3398 & ~n12701 ) | ( n3398 & n22464 ) | ( ~n12701 & n22464 ) ;
  assign n22466 = n6477 ^ n536 ^ 1'b0 ;
  assign n22467 = n20163 ^ n18395 ^ n3108 ;
  assign n22468 = n22467 ^ n11638 ^ n7045 ;
  assign n22469 = n17272 ^ n4314 ^ 1'b0 ;
  assign n22470 = ( ~n22466 & n22468 ) | ( ~n22466 & n22469 ) | ( n22468 & n22469 ) ;
  assign n22471 = ( n1476 & n5664 ) | ( n1476 & n12063 ) | ( n5664 & n12063 ) ;
  assign n22472 = n22471 ^ n4994 ^ n4919 ;
  assign n22473 = n2067 & n22472 ;
  assign n22474 = n19721 & n22473 ;
  assign n22475 = n17702 ^ n13219 ^ 1'b0 ;
  assign n22476 = n22390 & ~n22475 ;
  assign n22477 = n6971 ^ n6874 ^ n2945 ;
  assign n22478 = ( ~n2770 & n5755 ) | ( ~n2770 & n22477 ) | ( n5755 & n22477 ) ;
  assign n22479 = ( n2376 & n9153 ) | ( n2376 & n22478 ) | ( n9153 & n22478 ) ;
  assign n22480 = n16382 ^ n7837 ^ n5712 ;
  assign n22481 = n8915 ^ n8391 ^ n6522 ;
  assign n22482 = ( n1445 & ~n8017 ) | ( n1445 & n22481 ) | ( ~n8017 & n22481 ) ;
  assign n22483 = ( ~n526 & n5457 ) | ( ~n526 & n22482 ) | ( n5457 & n22482 ) ;
  assign n22484 = ( ~n6501 & n10176 ) | ( ~n6501 & n13785 ) | ( n10176 & n13785 ) ;
  assign n22485 = n22484 ^ n17139 ^ 1'b0 ;
  assign n22486 = ( n2539 & n4827 ) | ( n2539 & n22485 ) | ( n4827 & n22485 ) ;
  assign n22487 = n6285 ^ n5756 ^ 1'b0 ;
  assign n22488 = ~n11912 & n22487 ;
  assign n22489 = n22488 ^ n11865 ^ 1'b0 ;
  assign n22490 = n22486 | n22489 ;
  assign n22491 = n16477 ^ n10014 ^ n3016 ;
  assign n22492 = ( n4774 & ~n22490 ) | ( n4774 & n22491 ) | ( ~n22490 & n22491 ) ;
  assign n22493 = n18225 ^ n12947 ^ 1'b0 ;
  assign n22495 = n16357 ^ n13319 ^ n7222 ;
  assign n22494 = ~n4246 & n8091 ;
  assign n22496 = n22495 ^ n22494 ^ 1'b0 ;
  assign n22497 = ( n1060 & n11758 ) | ( n1060 & n22496 ) | ( n11758 & n22496 ) ;
  assign n22501 = ~n2200 & n21552 ;
  assign n22500 = n10961 ^ n6435 ^ n2092 ;
  assign n22502 = n22501 ^ n22500 ^ n19181 ;
  assign n22498 = n10815 ^ n7329 ^ 1'b0 ;
  assign n22499 = n16605 | n22498 ;
  assign n22503 = n22502 ^ n22499 ^ n7198 ;
  assign n22504 = ( n5363 & n8642 ) | ( n5363 & ~n11674 ) | ( n8642 & ~n11674 ) ;
  assign n22505 = n22504 ^ n10792 ^ n10439 ;
  assign n22506 = ( ~n6838 & n12693 ) | ( ~n6838 & n22505 ) | ( n12693 & n22505 ) ;
  assign n22507 = ( n9415 & ~n21084 ) | ( n9415 & n22506 ) | ( ~n21084 & n22506 ) ;
  assign n22508 = n10521 & ~n22507 ;
  assign n22509 = ( n590 & n21172 ) | ( n590 & n22508 ) | ( n21172 & n22508 ) ;
  assign n22514 = n17537 ^ n12911 ^ 1'b0 ;
  assign n22515 = n22495 & ~n22514 ;
  assign n22516 = ( n1078 & n4463 ) | ( n1078 & ~n15443 ) | ( n4463 & ~n15443 ) ;
  assign n22517 = ( n10140 & n22515 ) | ( n10140 & n22516 ) | ( n22515 & n22516 ) ;
  assign n22510 = ( ~n1500 & n4274 ) | ( ~n1500 & n5470 ) | ( n4274 & n5470 ) ;
  assign n22511 = n7729 ^ n3925 ^ n2816 ;
  assign n22512 = n22511 ^ n10437 ^ 1'b0 ;
  assign n22513 = n22510 & n22512 ;
  assign n22518 = n22517 ^ n22513 ^ n16145 ;
  assign n22519 = n15499 ^ n12970 ^ n719 ;
  assign n22520 = n22519 ^ n5489 ^ 1'b0 ;
  assign n22521 = n22518 & n22520 ;
  assign n22522 = n20029 ^ n12259 ^ n9378 ;
  assign n22523 = n22522 ^ n11683 ^ n8836 ;
  assign n22525 = n5937 ^ n3261 ^ n1875 ;
  assign n22524 = n14984 ^ n10420 ^ n3620 ;
  assign n22526 = n22525 ^ n22524 ^ n18669 ;
  assign n22534 = ( n15550 & ~n18780 ) | ( n15550 & n21593 ) | ( ~n18780 & n21593 ) ;
  assign n22527 = ( n708 & n1278 ) | ( n708 & n5429 ) | ( n1278 & n5429 ) ;
  assign n22528 = ( n9172 & ~n10594 ) | ( n9172 & n22527 ) | ( ~n10594 & n22527 ) ;
  assign n22529 = n4397 & n13006 ;
  assign n22530 = ~n5390 & n22529 ;
  assign n22531 = n22530 ^ n6145 ^ n4536 ;
  assign n22532 = ( n320 & n22528 ) | ( n320 & n22531 ) | ( n22528 & n22531 ) ;
  assign n22533 = ~n13812 & n22532 ;
  assign n22535 = n22534 ^ n22533 ^ 1'b0 ;
  assign n22536 = n21532 ^ n7698 ^ 1'b0 ;
  assign n22537 = n1675 ^ n1646 ^ n690 ;
  assign n22538 = n22537 ^ n8585 ^ n7042 ;
  assign n22539 = n7829 ^ n4404 ^ 1'b0 ;
  assign n22540 = ~n16062 & n22539 ;
  assign n22541 = ( n5309 & n22538 ) | ( n5309 & n22540 ) | ( n22538 & n22540 ) ;
  assign n22542 = ( ~n2474 & n16600 ) | ( ~n2474 & n22541 ) | ( n16600 & n22541 ) ;
  assign n22543 = n22542 ^ n20208 ^ n18771 ;
  assign n22544 = ( n6391 & n11561 ) | ( n6391 & ~n22543 ) | ( n11561 & ~n22543 ) ;
  assign n22545 = n20539 ^ n12778 ^ n4362 ;
  assign n22546 = n687 & n14165 ;
  assign n22547 = n2658 & n22546 ;
  assign n22548 = ( n4685 & n17574 ) | ( n4685 & ~n22547 ) | ( n17574 & ~n22547 ) ;
  assign n22549 = n22548 ^ n13634 ^ x121 ;
  assign n22550 = n22549 ^ n13472 ^ n986 ;
  assign n22551 = n22550 ^ n8912 ^ n1118 ;
  assign n22552 = ~n1012 & n7387 ;
  assign n22553 = n22552 ^ n981 ^ 1'b0 ;
  assign n22554 = n2415 & ~n22553 ;
  assign n22555 = n16826 ^ n9404 ^ 1'b0 ;
  assign n22556 = ~n20123 & n22555 ;
  assign n22557 = n12835 & n22556 ;
  assign n22558 = ( n11798 & n22554 ) | ( n11798 & n22557 ) | ( n22554 & n22557 ) ;
  assign n22561 = ( n4564 & n5943 ) | ( n4564 & n10835 ) | ( n5943 & n10835 ) ;
  assign n22559 = n12076 ^ n4884 ^ x215 ;
  assign n22560 = ~n5572 & n22559 ;
  assign n22562 = n22561 ^ n22560 ^ n11299 ;
  assign n22563 = n16603 ^ n8901 ^ 1'b0 ;
  assign n22564 = ( ~n8660 & n12205 ) | ( ~n8660 & n22563 ) | ( n12205 & n22563 ) ;
  assign n22567 = n8742 | n16524 ;
  assign n22568 = n22567 ^ n5785 ^ 1'b0 ;
  assign n22569 = n8678 | n22568 ;
  assign n22565 = n14497 ^ n7722 ^ n1092 ;
  assign n22566 = ( n6167 & n9507 ) | ( n6167 & n22565 ) | ( n9507 & n22565 ) ;
  assign n22570 = n22569 ^ n22566 ^ n15460 ;
  assign n22571 = n22564 & ~n22570 ;
  assign n22572 = n22571 ^ n8567 ^ 1'b0 ;
  assign n22573 = ( n11341 & n15951 ) | ( n11341 & ~n22572 ) | ( n15951 & ~n22572 ) ;
  assign n22574 = n12754 ^ n6164 ^ n3355 ;
  assign n22575 = x210 | n2881 ;
  assign n22576 = n22575 ^ n4066 ^ n1813 ;
  assign n22577 = ( ~n2589 & n12059 ) | ( ~n2589 & n22576 ) | ( n12059 & n22576 ) ;
  assign n22578 = n22577 ^ n17894 ^ 1'b0 ;
  assign n22579 = n22574 | n22578 ;
  assign n22580 = n5406 ^ n4260 ^ 1'b0 ;
  assign n22581 = n11098 & ~n22580 ;
  assign n22582 = n943 | n20884 ;
  assign n22583 = n22582 ^ n7272 ^ 1'b0 ;
  assign n22584 = ( n12564 & ~n17308 ) | ( n12564 & n22583 ) | ( ~n17308 & n22583 ) ;
  assign n22586 = n14331 ^ n5361 ^ n2651 ;
  assign n22585 = ~n12723 & n16998 ;
  assign n22587 = n22586 ^ n22585 ^ 1'b0 ;
  assign n22588 = ~n22584 & n22587 ;
  assign n22589 = n18239 ^ n18064 ^ n12821 ;
  assign n22590 = ( n8816 & n11634 ) | ( n8816 & ~n22589 ) | ( n11634 & ~n22589 ) ;
  assign n22591 = n2210 | n22590 ;
  assign n22592 = n22588 & ~n22591 ;
  assign n22597 = n18147 ^ n10262 ^ n5450 ;
  assign n22593 = n20989 ^ n18841 ^ n13053 ;
  assign n22594 = ( n7144 & n15139 ) | ( n7144 & ~n22593 ) | ( n15139 & ~n22593 ) ;
  assign n22595 = ( n2305 & n11331 ) | ( n2305 & n22594 ) | ( n11331 & n22594 ) ;
  assign n22596 = ~n20794 & n22595 ;
  assign n22598 = n22597 ^ n22596 ^ 1'b0 ;
  assign n22599 = n12143 ^ n10124 ^ 1'b0 ;
  assign n22600 = n2862 | n22599 ;
  assign n22601 = ( n367 & n8129 ) | ( n367 & n22600 ) | ( n8129 & n22600 ) ;
  assign n22602 = ( n408 & n10386 ) | ( n408 & n12030 ) | ( n10386 & n12030 ) ;
  assign n22603 = ~n9662 & n19438 ;
  assign n22604 = n22603 ^ n13316 ^ n5565 ;
  assign n22605 = n22604 ^ n20963 ^ n9090 ;
  assign n22606 = ( n3190 & n22602 ) | ( n3190 & ~n22605 ) | ( n22602 & ~n22605 ) ;
  assign n22607 = n16928 ^ n6749 ^ n462 ;
  assign n22608 = n22607 ^ n13011 ^ x249 ;
  assign n22609 = n22608 ^ n10417 ^ 1'b0 ;
  assign n22610 = n22609 ^ n9333 ^ n3651 ;
  assign n22611 = ( n6309 & n10576 ) | ( n6309 & n19470 ) | ( n10576 & n19470 ) ;
  assign n22612 = ( n9185 & ~n16429 ) | ( n9185 & n22611 ) | ( ~n16429 & n22611 ) ;
  assign n22613 = n3759 & ~n10548 ;
  assign n22614 = n14622 & n22613 ;
  assign n22615 = n13946 ^ n3054 ^ n2050 ;
  assign n22616 = ( n10494 & ~n15934 ) | ( n10494 & n22615 ) | ( ~n15934 & n22615 ) ;
  assign n22617 = n1291 ^ n548 ^ 1'b0 ;
  assign n22618 = ~n22616 & n22617 ;
  assign n22619 = ~n9589 & n10459 ;
  assign n22620 = ~n5956 & n22619 ;
  assign n22621 = n22620 ^ n17471 ^ 1'b0 ;
  assign n22622 = ~n8034 & n22621 ;
  assign n22623 = ( n2548 & ~n11219 ) | ( n2548 & n22622 ) | ( ~n11219 & n22622 ) ;
  assign n22624 = n22623 ^ n10136 ^ n764 ;
  assign n22625 = ( n448 & n6199 ) | ( n448 & ~n10209 ) | ( n6199 & ~n10209 ) ;
  assign n22626 = n5429 & ~n10600 ;
  assign n22627 = n690 & ~n14185 ;
  assign n22628 = n14164 & n22627 ;
  assign n22629 = n22628 ^ n1443 ^ n846 ;
  assign n22630 = ( n9353 & n17052 ) | ( n9353 & n19813 ) | ( n17052 & n19813 ) ;
  assign n22631 = n19071 | n22630 ;
  assign n22632 = ( n2933 & n5331 ) | ( n2933 & ~n9892 ) | ( n5331 & ~n9892 ) ;
  assign n22633 = ( n3735 & ~n17794 ) | ( n3735 & n22632 ) | ( ~n17794 & n22632 ) ;
  assign n22634 = n22633 ^ n17398 ^ n1150 ;
  assign n22635 = ( n2740 & n5413 ) | ( n2740 & n8807 ) | ( n5413 & n8807 ) ;
  assign n22636 = ( ~n5661 & n7169 ) | ( ~n5661 & n12344 ) | ( n7169 & n12344 ) ;
  assign n22637 = ( n4378 & ~n22635 ) | ( n4378 & n22636 ) | ( ~n22635 & n22636 ) ;
  assign n22638 = n22637 ^ n9351 ^ n1497 ;
  assign n22639 = n10347 ^ n948 ^ 1'b0 ;
  assign n22640 = n22638 & ~n22639 ;
  assign n22643 = n5143 ^ n2379 ^ 1'b0 ;
  assign n22642 = n22323 ^ n13301 ^ n5908 ;
  assign n22641 = n13605 & n16867 ;
  assign n22644 = n22643 ^ n22642 ^ n22641 ;
  assign n22645 = n5832 ^ n4278 ^ 1'b0 ;
  assign n22646 = n12142 ^ n6281 ^ n3278 ;
  assign n22647 = ( n5981 & n13318 ) | ( n5981 & ~n22646 ) | ( n13318 & ~n22646 ) ;
  assign n22648 = n4217 | n22647 ;
  assign n22649 = n22648 ^ n11925 ^ 1'b0 ;
  assign n22650 = n20176 ^ n11527 ^ 1'b0 ;
  assign n22651 = ( n6130 & n20326 ) | ( n6130 & ~n22650 ) | ( n20326 & ~n22650 ) ;
  assign n22652 = n10558 | n14616 ;
  assign n22653 = n22651 & ~n22652 ;
  assign n22658 = n21843 ^ n15719 ^ n7704 ;
  assign n22654 = n18024 ^ n1475 ^ n660 ;
  assign n22655 = n22654 ^ n16251 ^ n8787 ;
  assign n22656 = n22655 ^ n3223 ^ n1297 ;
  assign n22657 = ~n21418 & n22656 ;
  assign n22659 = n22658 ^ n22657 ^ 1'b0 ;
  assign n22660 = n10301 & n17258 ;
  assign n22661 = ( n2368 & n7152 ) | ( n2368 & n22660 ) | ( n7152 & n22660 ) ;
  assign n22666 = ( n9725 & n13561 ) | ( n9725 & n14167 ) | ( n13561 & n14167 ) ;
  assign n22664 = ( ~n6609 & n7504 ) | ( ~n6609 & n10809 ) | ( n7504 & n10809 ) ;
  assign n22665 = n22664 ^ n4939 ^ n2405 ;
  assign n22667 = n22666 ^ n22665 ^ n11164 ;
  assign n22662 = n9929 & ~n20265 ;
  assign n22663 = n21584 & n22662 ;
  assign n22668 = n22667 ^ n22663 ^ n18529 ;
  assign n22669 = n11220 ^ n7742 ^ n6845 ;
  assign n22670 = n3727 ^ n1629 ^ 1'b0 ;
  assign n22671 = n15824 ^ n9958 ^ n1464 ;
  assign n22672 = n19816 ^ n9479 ^ n2280 ;
  assign n22673 = ( n22670 & ~n22671 ) | ( n22670 & n22672 ) | ( ~n22671 & n22672 ) ;
  assign n22674 = n9092 ^ n4179 ^ n982 ;
  assign n22675 = n18402 ^ n1013 ^ 1'b0 ;
  assign n22676 = ( n6281 & n17508 ) | ( n6281 & ~n22675 ) | ( n17508 & ~n22675 ) ;
  assign n22677 = ( ~n6654 & n11279 ) | ( ~n6654 & n22676 ) | ( n11279 & n22676 ) ;
  assign n22680 = n694 | n2194 ;
  assign n22681 = n3433 & ~n22680 ;
  assign n22678 = n6780 ^ n1148 ^ 1'b0 ;
  assign n22679 = n287 & ~n22678 ;
  assign n22682 = n22681 ^ n22679 ^ n18277 ;
  assign n22685 = n4807 ^ n2791 ^ n1118 ;
  assign n22686 = n5810 & n22685 ;
  assign n22687 = n8324 & n12834 ;
  assign n22688 = ( ~n21296 & n22686 ) | ( ~n21296 & n22687 ) | ( n22686 & n22687 ) ;
  assign n22683 = n1600 & n6461 ;
  assign n22684 = n22683 ^ n16353 ^ 1'b0 ;
  assign n22689 = n22688 ^ n22684 ^ n10275 ;
  assign n22692 = n17066 & ~n18225 ;
  assign n22690 = ~n1697 & n10532 ;
  assign n22691 = n22690 ^ n3729 ^ 1'b0 ;
  assign n22693 = n22692 ^ n22691 ^ n12193 ;
  assign n22694 = n6295 & n14808 ;
  assign n22696 = n9306 & n13412 ;
  assign n22697 = n1162 & n22696 ;
  assign n22698 = ( n1343 & ~n8410 ) | ( n1343 & n22697 ) | ( ~n8410 & n22697 ) ;
  assign n22695 = n2188 & n2670 ;
  assign n22699 = n22698 ^ n22695 ^ 1'b0 ;
  assign n22708 = n8593 & n12959 ;
  assign n22709 = ( n2484 & n11944 ) | ( n2484 & ~n22708 ) | ( n11944 & ~n22708 ) ;
  assign n22706 = n6892 ^ n710 ^ 1'b0 ;
  assign n22707 = n271 & n22706 ;
  assign n22703 = n20240 ^ n9132 ^ 1'b0 ;
  assign n22704 = ~n19390 & n22703 ;
  assign n22700 = n1015 | n6054 ;
  assign n22701 = n11965 | n22700 ;
  assign n22702 = ( n4980 & n13329 ) | ( n4980 & n22701 ) | ( n13329 & n22701 ) ;
  assign n22705 = n22704 ^ n22702 ^ n1078 ;
  assign n22710 = n22709 ^ n22707 ^ n22705 ;
  assign n22713 = n2846 & ~n22052 ;
  assign n22711 = n18974 ^ n4281 ^ 1'b0 ;
  assign n22712 = n3698 | n22711 ;
  assign n22714 = n22713 ^ n22712 ^ n1950 ;
  assign n22715 = n6928 & n9533 ;
  assign n22716 = n22715 ^ n22061 ^ 1'b0 ;
  assign n22717 = n884 & ~n12728 ;
  assign n22718 = n2951 & n18950 ;
  assign n22719 = ~n22717 & n22718 ;
  assign n22720 = n19119 ^ n16205 ^ n10616 ;
  assign n22721 = ( ~n2874 & n5283 ) | ( ~n2874 & n13230 ) | ( n5283 & n13230 ) ;
  assign n22722 = n5881 | n10963 ;
  assign n22723 = ~n2608 & n8051 ;
  assign n22724 = n22723 ^ n9403 ^ 1'b0 ;
  assign n22725 = n22724 ^ n19000 ^ n15563 ;
  assign n22726 = ( ~n6939 & n15762 ) | ( ~n6939 & n17591 ) | ( n15762 & n17591 ) ;
  assign n22727 = n22726 ^ n9758 ^ n4754 ;
  assign n22728 = n22727 ^ n5089 ^ 1'b0 ;
  assign n22729 = ~n2167 & n22728 ;
  assign n22730 = n22729 ^ n6564 ^ 1'b0 ;
  assign n22731 = ( n15331 & ~n22725 ) | ( n15331 & n22730 ) | ( ~n22725 & n22730 ) ;
  assign n22736 = n2521 ^ n689 ^ x200 ;
  assign n22732 = ( n1927 & ~n4474 ) | ( n1927 & n13142 ) | ( ~n4474 & n13142 ) ;
  assign n22733 = n7313 & n7657 ;
  assign n22734 = n22733 ^ n14104 ^ 1'b0 ;
  assign n22735 = ( n1997 & n22732 ) | ( n1997 & n22734 ) | ( n22732 & n22734 ) ;
  assign n22737 = n22736 ^ n22735 ^ n22287 ;
  assign n22738 = n1671 & n8162 ;
  assign n22742 = ~n14712 & n22391 ;
  assign n22739 = n9877 | n14012 ;
  assign n22740 = n2087 | n22739 ;
  assign n22741 = n22740 ^ n6633 ^ 1'b0 ;
  assign n22743 = n22742 ^ n22741 ^ n14772 ;
  assign n22744 = ( ~n1581 & n11004 ) | ( ~n1581 & n13053 ) | ( n11004 & n13053 ) ;
  assign n22745 = ~n16438 & n22744 ;
  assign n22746 = n13660 & n22745 ;
  assign n22747 = ( n8112 & n14238 ) | ( n8112 & ~n15657 ) | ( n14238 & ~n15657 ) ;
  assign n22748 = n2480 & n3119 ;
  assign n22749 = n22748 ^ n3455 ^ 1'b0 ;
  assign n22750 = n22747 & ~n22749 ;
  assign n22751 = n18276 & n22750 ;
  assign n22752 = ( n9566 & n16791 ) | ( n9566 & ~n17117 ) | ( n16791 & ~n17117 ) ;
  assign n22753 = ( n792 & n9791 ) | ( n792 & ~n22752 ) | ( n9791 & ~n22752 ) ;
  assign n22754 = n17432 ^ n2192 ^ 1'b0 ;
  assign n22755 = n22754 ^ n11816 ^ n4797 ;
  assign n22760 = n12963 ^ n11885 ^ 1'b0 ;
  assign n22761 = n20580 & ~n22760 ;
  assign n22757 = n7070 & n8839 ;
  assign n22758 = n22757 ^ n5095 ^ 1'b0 ;
  assign n22759 = ( n6102 & n6706 ) | ( n6102 & n22758 ) | ( n6706 & n22758 ) ;
  assign n22756 = n20661 ^ n11541 ^ n7808 ;
  assign n22762 = n22761 ^ n22759 ^ n22756 ;
  assign n22763 = n20526 ^ n794 ^ 1'b0 ;
  assign n22764 = n7630 ^ n1782 ^ x102 ;
  assign n22765 = n21349 ^ n4606 ^ n1657 ;
  assign n22766 = ( n1761 & n22764 ) | ( n1761 & ~n22765 ) | ( n22764 & ~n22765 ) ;
  assign n22767 = n22766 ^ n21459 ^ n17080 ;
  assign n22768 = n3443 & ~n22274 ;
  assign n22769 = n22768 ^ n16495 ^ 1'b0 ;
  assign n22770 = ( n5143 & ~n10461 ) | ( n5143 & n18079 ) | ( ~n10461 & n18079 ) ;
  assign n22771 = ( n1081 & n17682 ) | ( n1081 & ~n22770 ) | ( n17682 & ~n22770 ) ;
  assign n22772 = n22771 ^ n12357 ^ n12002 ;
  assign n22773 = n16529 ^ n12869 ^ n5890 ;
  assign n22774 = n478 & n22773 ;
  assign n22775 = n22774 ^ n15666 ^ 1'b0 ;
  assign n22776 = n4425 & ~n5849 ;
  assign n22777 = n701 & n22776 ;
  assign n22778 = ( ~n4040 & n6223 ) | ( ~n4040 & n10867 ) | ( n6223 & n10867 ) ;
  assign n22779 = n9970 ^ n2035 ^ 1'b0 ;
  assign n22780 = n1308 & n22779 ;
  assign n22781 = ( n3166 & n7973 ) | ( n3166 & n22780 ) | ( n7973 & n22780 ) ;
  assign n22782 = n22781 ^ n17388 ^ n506 ;
  assign n22783 = ( n4136 & n22778 ) | ( n4136 & ~n22782 ) | ( n22778 & ~n22782 ) ;
  assign n22784 = ( n7206 & n7731 ) | ( n7206 & n22783 ) | ( n7731 & n22783 ) ;
  assign n22785 = n22777 & ~n22784 ;
  assign n22786 = n4668 & n11739 ;
  assign n22790 = n6801 & ~n8980 ;
  assign n22791 = n22790 ^ n1233 ^ 1'b0 ;
  assign n22787 = ~n1091 & n7162 ;
  assign n22788 = ~n1835 & n22787 ;
  assign n22789 = n20205 & ~n22788 ;
  assign n22792 = n22791 ^ n22789 ^ 1'b0 ;
  assign n22796 = n22226 ^ n9640 ^ n5574 ;
  assign n22797 = ( n1936 & ~n21151 ) | ( n1936 & n22796 ) | ( ~n21151 & n22796 ) ;
  assign n22798 = n22797 ^ n22358 ^ n18713 ;
  assign n22793 = n8224 ^ n1411 ^ x236 ;
  assign n22794 = n22793 ^ n8963 ^ 1'b0 ;
  assign n22795 = n11199 & ~n22794 ;
  assign n22799 = n22798 ^ n22795 ^ n9000 ;
  assign n22803 = n13234 ^ n13167 ^ n3948 ;
  assign n22802 = n4235 | n11601 ;
  assign n22804 = n22803 ^ n22802 ^ 1'b0 ;
  assign n22800 = n5507 ^ n3045 ^ 1'b0 ;
  assign n22801 = ~n6347 & n22800 ;
  assign n22805 = n22804 ^ n22801 ^ n10877 ;
  assign n22806 = n22805 ^ n16366 ^ n15149 ;
  assign n22808 = ( n8963 & n11025 ) | ( n8963 & n15706 ) | ( n11025 & n15706 ) ;
  assign n22809 = n22808 ^ n11440 ^ n561 ;
  assign n22807 = n4655 & ~n19821 ;
  assign n22810 = n22809 ^ n22807 ^ n15087 ;
  assign n22811 = ( n2596 & ~n3364 ) | ( n2596 & n5983 ) | ( ~n3364 & n5983 ) ;
  assign n22812 = n22811 ^ n18672 ^ n9246 ;
  assign n22813 = n15116 ^ n13186 ^ n9259 ;
  assign n22814 = n8161 & ~n11399 ;
  assign n22815 = n22813 & n22814 ;
  assign n22816 = n22815 ^ n18744 ^ n15138 ;
  assign n22817 = n6790 & n20327 ;
  assign n22818 = n22817 ^ n19496 ^ 1'b0 ;
  assign n22819 = ( n5368 & n9874 ) | ( n5368 & n11161 ) | ( n9874 & n11161 ) ;
  assign n22825 = ( n350 & n1460 ) | ( n350 & ~n15354 ) | ( n1460 & ~n15354 ) ;
  assign n22823 = n12679 ^ n1954 ^ n1207 ;
  assign n22820 = ( n6062 & n8810 ) | ( n6062 & ~n9318 ) | ( n8810 & ~n9318 ) ;
  assign n22821 = ( ~n8274 & n21050 ) | ( ~n8274 & n22820 ) | ( n21050 & n22820 ) ;
  assign n22822 = n8755 & ~n22821 ;
  assign n22824 = n22823 ^ n22822 ^ 1'b0 ;
  assign n22826 = n22825 ^ n22824 ^ 1'b0 ;
  assign n22827 = ~n5154 & n22826 ;
  assign n22828 = ( n14694 & ~n14734 ) | ( n14694 & n16354 ) | ( ~n14734 & n16354 ) ;
  assign n22829 = ( ~n10558 & n22827 ) | ( ~n10558 & n22828 ) | ( n22827 & n22828 ) ;
  assign n22830 = ( n5433 & n9829 ) | ( n5433 & n15056 ) | ( n9829 & n15056 ) ;
  assign n22831 = n22830 ^ n19871 ^ n9612 ;
  assign n22832 = n16709 & n22831 ;
  assign n22833 = ( ~n4756 & n7284 ) | ( ~n4756 & n9192 ) | ( n7284 & n9192 ) ;
  assign n22834 = ( n8902 & ~n17243 ) | ( n8902 & n22833 ) | ( ~n17243 & n22833 ) ;
  assign n22835 = ( n2931 & n22795 ) | ( n2931 & n22834 ) | ( n22795 & n22834 ) ;
  assign n22836 = n18717 ^ n17909 ^ n4197 ;
  assign n22837 = ~n8463 & n22836 ;
  assign n22838 = ( n8260 & ~n10017 ) | ( n8260 & n11656 ) | ( ~n10017 & n11656 ) ;
  assign n22839 = n17545 ^ n6835 ^ 1'b0 ;
  assign n22840 = n22839 ^ n2531 ^ 1'b0 ;
  assign n22841 = ( x31 & n14432 ) | ( x31 & n20184 ) | ( n14432 & n20184 ) ;
  assign n22842 = n22841 ^ n22778 ^ n1888 ;
  assign n22843 = ( n1983 & n16942 ) | ( n1983 & n18805 ) | ( n16942 & n18805 ) ;
  assign n22844 = n18370 ^ n3990 ^ n3404 ;
  assign n22845 = n22844 ^ n10384 ^ n7413 ;
  assign n22846 = n22845 ^ n9743 ^ n4094 ;
  assign n22847 = ( x104 & n12009 ) | ( x104 & ~n22846 ) | ( n12009 & ~n22846 ) ;
  assign n22851 = n6732 ^ n1027 ^ 1'b0 ;
  assign n22852 = n14834 | n22851 ;
  assign n22848 = n6458 & n20021 ;
  assign n22849 = n22848 ^ n4306 ^ 1'b0 ;
  assign n22850 = ( n7555 & n9657 ) | ( n7555 & ~n22849 ) | ( n9657 & ~n22849 ) ;
  assign n22853 = n22852 ^ n22850 ^ n14271 ;
  assign n22854 = ( n22843 & ~n22847 ) | ( n22843 & n22853 ) | ( ~n22847 & n22853 ) ;
  assign n22855 = n6691 ^ n5250 ^ n4422 ;
  assign n22856 = ( n770 & ~n12951 ) | ( n770 & n22855 ) | ( ~n12951 & n22855 ) ;
  assign n22857 = n16161 | n22856 ;
  assign n22858 = n20909 & ~n22857 ;
  assign n22859 = n19186 ^ n12709 ^ 1'b0 ;
  assign n22860 = ( n17613 & n22858 ) | ( n17613 & n22859 ) | ( n22858 & n22859 ) ;
  assign n22861 = n9081 & ~n20168 ;
  assign n22862 = n22861 ^ n6581 ^ 1'b0 ;
  assign n22863 = n22862 ^ n22122 ^ n19660 ;
  assign n22864 = n22193 ^ n7535 ^ n3520 ;
  assign n22866 = n10896 ^ n5788 ^ n4170 ;
  assign n22867 = ~n17652 & n22866 ;
  assign n22868 = n22867 ^ n12575 ^ 1'b0 ;
  assign n22865 = n22620 ^ n19818 ^ n19169 ;
  assign n22869 = n22868 ^ n22865 ^ n4987 ;
  assign n22872 = n3746 ^ n2143 ^ n1588 ;
  assign n22873 = ( n6587 & ~n9635 ) | ( n6587 & n22872 ) | ( ~n9635 & n22872 ) ;
  assign n22870 = ( ~x142 & n2401 ) | ( ~x142 & n5772 ) | ( n2401 & n5772 ) ;
  assign n22871 = ( ~n14007 & n21806 ) | ( ~n14007 & n22870 ) | ( n21806 & n22870 ) ;
  assign n22874 = n22873 ^ n22871 ^ n7490 ;
  assign n22875 = n20092 ^ n4472 ^ 1'b0 ;
  assign n22876 = n22875 ^ n7693 ^ n3214 ;
  assign n22877 = ( ~n15907 & n22874 ) | ( ~n15907 & n22876 ) | ( n22874 & n22876 ) ;
  assign n22881 = ( n1326 & n8980 ) | ( n1326 & n10082 ) | ( n8980 & n10082 ) ;
  assign n22880 = n16865 ^ n12544 ^ n6623 ;
  assign n22878 = n21225 ^ n3685 ^ n1053 ;
  assign n22879 = n22878 ^ n13845 ^ n897 ;
  assign n22882 = n22881 ^ n22880 ^ n22879 ;
  assign n22884 = ( n2894 & ~n9471 ) | ( n2894 & n18260 ) | ( ~n9471 & n18260 ) ;
  assign n22883 = ( n1293 & ~n1938 ) | ( n1293 & n2224 ) | ( ~n1938 & n2224 ) ;
  assign n22885 = n22884 ^ n22883 ^ 1'b0 ;
  assign n22886 = n706 & ~n22885 ;
  assign n22887 = ( n4934 & n8803 ) | ( n4934 & ~n10402 ) | ( n8803 & ~n10402 ) ;
  assign n22888 = ~n8750 & n22887 ;
  assign n22889 = ~n2113 & n16230 ;
  assign n22890 = n22889 ^ n16443 ^ n13242 ;
  assign n22891 = n6632 ^ n4539 ^ n2776 ;
  assign n22892 = n22891 ^ n13753 ^ n3807 ;
  assign n22893 = n6509 | n22892 ;
  assign n22894 = n14014 & ~n22893 ;
  assign n22895 = ( n7299 & n12126 ) | ( n7299 & n12252 ) | ( n12126 & n12252 ) ;
  assign n22896 = n15847 & n20019 ;
  assign n22897 = n22895 & n22896 ;
  assign n22898 = n22897 ^ n18598 ^ n1564 ;
  assign n22899 = n22894 | n22898 ;
  assign n22900 = n517 | n22899 ;
  assign n22901 = n11425 & n12178 ;
  assign n22902 = ( n11665 & n18510 ) | ( n11665 & n21272 ) | ( n18510 & n21272 ) ;
  assign n22903 = n5201 ^ n4604 ^ n4286 ;
  assign n22904 = ( n4667 & n7262 ) | ( n4667 & n22903 ) | ( n7262 & n22903 ) ;
  assign n22905 = ( n17734 & n22902 ) | ( n17734 & n22904 ) | ( n22902 & n22904 ) ;
  assign n22911 = n16649 ^ n11174 ^ 1'b0 ;
  assign n22912 = ( n7076 & n13030 ) | ( n7076 & n22911 ) | ( n13030 & n22911 ) ;
  assign n22910 = n2861 & ~n2957 ;
  assign n22913 = n22912 ^ n22910 ^ 1'b0 ;
  assign n22914 = n22913 ^ n14482 ^ n8002 ;
  assign n22906 = n6124 ^ n4836 ^ 1'b0 ;
  assign n22907 = n6803 & n22906 ;
  assign n22908 = n16078 ^ n15811 ^ x44 ;
  assign n22909 = ( n9257 & n22907 ) | ( n9257 & n22908 ) | ( n22907 & n22908 ) ;
  assign n22915 = n22914 ^ n22909 ^ n8662 ;
  assign n22916 = ( n16499 & ~n16903 ) | ( n16499 & n20517 ) | ( ~n16903 & n20517 ) ;
  assign n22917 = n4215 ^ n2744 ^ x232 ;
  assign n22918 = n12370 ^ n2004 ^ 1'b0 ;
  assign n22919 = ~n7940 & n22918 ;
  assign n22920 = ~n22917 & n22919 ;
  assign n22921 = ~n11337 & n22920 ;
  assign n22922 = ( n1784 & n8315 ) | ( n1784 & ~n8690 ) | ( n8315 & ~n8690 ) ;
  assign n22923 = n22922 ^ n17736 ^ n15423 ;
  assign n22924 = n21471 ^ n20066 ^ n14894 ;
  assign n22925 = n16302 | n22758 ;
  assign n22926 = n8181 & ~n22925 ;
  assign n22927 = n22926 ^ n5572 ^ 1'b0 ;
  assign n22928 = n4746 & n22927 ;
  assign n22929 = n22928 ^ n17236 ^ n4149 ;
  assign n22930 = ( n6285 & ~n8025 ) | ( n6285 & n10236 ) | ( ~n8025 & n10236 ) ;
  assign n22931 = n21663 ^ n9936 ^ n6690 ;
  assign n22932 = n19448 ^ n16492 ^ n4108 ;
  assign n22933 = n22932 ^ n20805 ^ n8260 ;
  assign n22934 = ( n20903 & n22931 ) | ( n20903 & ~n22933 ) | ( n22931 & ~n22933 ) ;
  assign n22936 = ( n5485 & n14789 ) | ( n5485 & ~n18389 ) | ( n14789 & ~n18389 ) ;
  assign n22935 = ~n4464 & n12261 ;
  assign n22937 = n22936 ^ n22935 ^ n13689 ;
  assign n22939 = ( n10142 & n16968 ) | ( n10142 & n19795 ) | ( n16968 & n19795 ) ;
  assign n22938 = n13364 ^ n8181 ^ 1'b0 ;
  assign n22940 = n22939 ^ n22938 ^ n10509 ;
  assign n22941 = n5778 ^ n2200 ^ n1402 ;
  assign n22942 = ~n14237 & n15593 ;
  assign n22943 = n22942 ^ n4133 ^ 1'b0 ;
  assign n22944 = n12205 ^ n3511 ^ 1'b0 ;
  assign n22945 = n17022 & ~n22944 ;
  assign n22946 = ( n752 & n5201 ) | ( n752 & n8034 ) | ( n5201 & n8034 ) ;
  assign n22947 = n4299 | n5415 ;
  assign n22948 = n22946 & ~n22947 ;
  assign n22949 = n9082 | n16768 ;
  assign n22950 = n22949 ^ n3462 ^ 1'b0 ;
  assign n22951 = ( ~n18706 & n22948 ) | ( ~n18706 & n22950 ) | ( n22948 & n22950 ) ;
  assign n22952 = ( ~n22943 & n22945 ) | ( ~n22943 & n22951 ) | ( n22945 & n22951 ) ;
  assign n22953 = n22941 & ~n22952 ;
  assign n22954 = ~n6095 & n7804 ;
  assign n22955 = n22954 ^ n6282 ^ 1'b0 ;
  assign n22956 = ( n5637 & n8203 ) | ( n5637 & ~n22955 ) | ( n8203 & ~n22955 ) ;
  assign n22957 = ( n6762 & n11193 ) | ( n6762 & ~n17578 ) | ( n11193 & ~n17578 ) ;
  assign n22958 = n22957 ^ n19460 ^ n11274 ;
  assign n22959 = ( ~n8451 & n15164 ) | ( ~n8451 & n17803 ) | ( n15164 & n17803 ) ;
  assign n22960 = ( n13369 & n16272 ) | ( n13369 & ~n22959 ) | ( n16272 & ~n22959 ) ;
  assign n22961 = n22960 ^ n12150 ^ 1'b0 ;
  assign n22962 = n22958 | n22961 ;
  assign n22965 = n14843 ^ n8772 ^ n1030 ;
  assign n22964 = n9051 ^ n5602 ^ n4894 ;
  assign n22963 = ( n4821 & n13025 ) | ( n4821 & ~n20871 ) | ( n13025 & ~n20871 ) ;
  assign n22966 = n22965 ^ n22964 ^ n22963 ;
  assign n22967 = ( n6021 & n7591 ) | ( n6021 & ~n21483 ) | ( n7591 & ~n21483 ) ;
  assign n22968 = n13645 ^ n10381 ^ n320 ;
  assign n22969 = ( n2244 & n4343 ) | ( n2244 & ~n22289 ) | ( n4343 & ~n22289 ) ;
  assign n22970 = ( n6170 & n22968 ) | ( n6170 & n22969 ) | ( n22968 & n22969 ) ;
  assign n22971 = n4092 | n7343 ;
  assign n22972 = n22971 ^ n4082 ^ 1'b0 ;
  assign n22973 = ( n460 & ~n12172 ) | ( n460 & n22972 ) | ( ~n12172 & n22972 ) ;
  assign n22974 = n12077 ^ n6026 ^ n3056 ;
  assign n22975 = ( n13088 & ~n18619 ) | ( n13088 & n22974 ) | ( ~n18619 & n22974 ) ;
  assign n22976 = n22975 ^ n10918 ^ n8462 ;
  assign n22977 = n13278 ^ n3539 ^ 1'b0 ;
  assign n22978 = ( n5041 & n13430 ) | ( n5041 & ~n22977 ) | ( n13430 & ~n22977 ) ;
  assign n22979 = n22978 ^ n12488 ^ n3808 ;
  assign n22980 = n15208 ^ n9966 ^ 1'b0 ;
  assign n22981 = n13228 & ~n22980 ;
  assign n22982 = ( ~n9593 & n18637 ) | ( ~n9593 & n22981 ) | ( n18637 & n22981 ) ;
  assign n22983 = ( n1685 & n2294 ) | ( n1685 & n8934 ) | ( n2294 & n8934 ) ;
  assign n22984 = ( ~n10544 & n18813 ) | ( ~n10544 & n22983 ) | ( n18813 & n22983 ) ;
  assign n22985 = n8980 & n22984 ;
  assign n22986 = n22985 ^ n3367 ^ 1'b0 ;
  assign n22987 = n22986 ^ n17909 ^ n10735 ;
  assign n22988 = n22987 ^ n12634 ^ n4503 ;
  assign n22989 = n12823 ^ n9456 ^ 1'b0 ;
  assign n22990 = n5861 & n22989 ;
  assign n22991 = n1567 & ~n1834 ;
  assign n22992 = ~n18532 & n22991 ;
  assign n22993 = ~n10272 & n20762 ;
  assign n22994 = ( ~n2283 & n11660 ) | ( ~n2283 & n19549 ) | ( n11660 & n19549 ) ;
  assign n22995 = ( n6087 & ~n17183 ) | ( n6087 & n17331 ) | ( ~n17183 & n17331 ) ;
  assign n22996 = n22995 ^ n4130 ^ 1'b0 ;
  assign n22997 = n22996 ^ n17393 ^ 1'b0 ;
  assign n22998 = n2564 & n19365 ;
  assign n22999 = ( n4991 & ~n8864 ) | ( n4991 & n22998 ) | ( ~n8864 & n22998 ) ;
  assign n23000 = ~n1529 & n4626 ;
  assign n23001 = n23000 ^ n9409 ^ 1'b0 ;
  assign n23002 = ( ~n1838 & n10372 ) | ( ~n1838 & n23001 ) | ( n10372 & n23001 ) ;
  assign n23003 = n8444 & n23002 ;
  assign n23004 = n23003 ^ n8251 ^ 1'b0 ;
  assign n23005 = n23004 ^ n19729 ^ n7673 ;
  assign n23006 = ( n10289 & n15536 ) | ( n10289 & n22660 ) | ( n15536 & n22660 ) ;
  assign n23007 = ( n2051 & n3969 ) | ( n2051 & n13221 ) | ( n3969 & n13221 ) ;
  assign n23008 = n2591 ^ n924 ^ 1'b0 ;
  assign n23009 = n23007 | n23008 ;
  assign n23010 = n14649 ^ n10613 ^ 1'b0 ;
  assign n23011 = ~n15362 & n23010 ;
  assign n23014 = n8051 ^ n5445 ^ x42 ;
  assign n23015 = ( ~n3476 & n7849 ) | ( ~n3476 & n23014 ) | ( n7849 & n23014 ) ;
  assign n23016 = n23015 ^ n6993 ^ 1'b0 ;
  assign n23017 = ( n8244 & n9797 ) | ( n8244 & ~n23016 ) | ( n9797 & ~n23016 ) ;
  assign n23018 = n6575 & n17650 ;
  assign n23019 = ( n5498 & n23017 ) | ( n5498 & n23018 ) | ( n23017 & n23018 ) ;
  assign n23012 = n8053 & n12170 ;
  assign n23013 = ( n4391 & n22655 ) | ( n4391 & n23012 ) | ( n22655 & n23012 ) ;
  assign n23020 = n23019 ^ n23013 ^ n18154 ;
  assign n23021 = n16806 & ~n19266 ;
  assign n23022 = n826 & n23021 ;
  assign n23024 = n19111 ^ n7896 ^ n4771 ;
  assign n23025 = n5762 ^ n5713 ^ 1'b0 ;
  assign n23026 = n1787 & n23025 ;
  assign n23027 = n23026 ^ n11227 ^ n3180 ;
  assign n23028 = ( ~n867 & n5708 ) | ( ~n867 & n7037 ) | ( n5708 & n7037 ) ;
  assign n23029 = n23028 ^ n9303 ^ n6247 ;
  assign n23030 = n23029 ^ n17361 ^ n11080 ;
  assign n23031 = n23027 | n23030 ;
  assign n23032 = n23024 & ~n23031 ;
  assign n23033 = n18412 ^ n9184 ^ 1'b0 ;
  assign n23034 = ( n8537 & ~n23032 ) | ( n8537 & n23033 ) | ( ~n23032 & n23033 ) ;
  assign n23023 = n19879 & n21627 ;
  assign n23035 = n23034 ^ n23023 ^ 1'b0 ;
  assign n23036 = n3450 ^ n2454 ^ x37 ;
  assign n23037 = n18024 ^ n6270 ^ n3075 ;
  assign n23038 = ~n3197 & n23037 ;
  assign n23039 = ( n8563 & ~n23036 ) | ( n8563 & n23038 ) | ( ~n23036 & n23038 ) ;
  assign n23040 = n21014 ^ n5893 ^ 1'b0 ;
  assign n23041 = ~n1987 & n23040 ;
  assign n23042 = n23041 ^ n20438 ^ 1'b0 ;
  assign n23044 = n19180 ^ n15780 ^ 1'b0 ;
  assign n23043 = ~n3898 & n8107 ;
  assign n23045 = n23044 ^ n23043 ^ n20833 ;
  assign n23046 = ( n4991 & n14978 ) | ( n4991 & n19446 ) | ( n14978 & n19446 ) ;
  assign n23047 = n2711 ^ n1840 ^ n1699 ;
  assign n23048 = n23047 ^ n19904 ^ n16823 ;
  assign n23051 = n18631 ^ n10082 ^ n4327 ;
  assign n23049 = ( n9456 & ~n10389 ) | ( n9456 & n16800 ) | ( ~n10389 & n16800 ) ;
  assign n23050 = n23049 ^ n11661 ^ n506 ;
  assign n23052 = n23051 ^ n23050 ^ 1'b0 ;
  assign n23053 = ~n1912 & n4109 ;
  assign n23054 = ~n2148 & n23053 ;
  assign n23055 = ( ~n3369 & n21142 ) | ( ~n3369 & n23054 ) | ( n21142 & n23054 ) ;
  assign n23056 = n6290 ^ n5889 ^ n4763 ;
  assign n23057 = ( ~n3680 & n13054 ) | ( ~n3680 & n19462 ) | ( n13054 & n19462 ) ;
  assign n23058 = n7253 ^ n2440 ^ 1'b0 ;
  assign n23059 = n12350 & n23058 ;
  assign n23060 = n795 & n23059 ;
  assign n23061 = n23057 & n23060 ;
  assign n23062 = ( ~x6 & n21510 ) | ( ~x6 & n23061 ) | ( n21510 & n23061 ) ;
  assign n23063 = n23062 ^ n13610 ^ 1'b0 ;
  assign n23064 = ( ~n4251 & n7638 ) | ( ~n4251 & n23063 ) | ( n7638 & n23063 ) ;
  assign n23065 = n23064 ^ n16018 ^ n11922 ;
  assign n23066 = n12542 ^ n10453 ^ n839 ;
  assign n23067 = n8631 & ~n23066 ;
  assign n23068 = ( n10176 & n23065 ) | ( n10176 & n23067 ) | ( n23065 & n23067 ) ;
  assign n23069 = n9001 ^ n2876 ^ 1'b0 ;
  assign n23070 = x136 & n23069 ;
  assign n23080 = ( n7105 & n9267 ) | ( n7105 & n17563 ) | ( n9267 & n17563 ) ;
  assign n23071 = ( ~n5811 & n10596 ) | ( ~n5811 & n19301 ) | ( n10596 & n19301 ) ;
  assign n23072 = n23071 ^ n18081 ^ n5194 ;
  assign n23073 = ( n2147 & n6134 ) | ( n2147 & ~n23072 ) | ( n6134 & ~n23072 ) ;
  assign n23074 = n6536 | n14926 ;
  assign n23075 = n23074 ^ n6641 ^ 1'b0 ;
  assign n23076 = n20620 | n23075 ;
  assign n23077 = ( ~n21063 & n23073 ) | ( ~n21063 & n23076 ) | ( n23073 & n23076 ) ;
  assign n23078 = n23077 ^ n9625 ^ 1'b0 ;
  assign n23079 = ~n5723 & n23078 ;
  assign n23081 = n23080 ^ n23079 ^ n15195 ;
  assign n23082 = n5000 ^ n4497 ^ 1'b0 ;
  assign n23083 = n1495 & ~n23082 ;
  assign n23084 = n23083 ^ n10145 ^ n8728 ;
  assign n23085 = ( n5771 & n9672 ) | ( n5771 & ~n11378 ) | ( n9672 & ~n11378 ) ;
  assign n23086 = ( n9166 & n23084 ) | ( n9166 & ~n23085 ) | ( n23084 & ~n23085 ) ;
  assign n23090 = n3318 | n16321 ;
  assign n23091 = n6305 | n23090 ;
  assign n23087 = n19359 ^ n15689 ^ n6788 ;
  assign n23088 = ( n5285 & n9589 ) | ( n5285 & ~n23087 ) | ( n9589 & ~n23087 ) ;
  assign n23089 = n23088 ^ n19869 ^ n5452 ;
  assign n23092 = n23091 ^ n23089 ^ n3610 ;
  assign n23093 = n23092 ^ n20810 ^ n2358 ;
  assign n23094 = ( n17280 & n23086 ) | ( n17280 & n23093 ) | ( n23086 & n23093 ) ;
  assign n23095 = n6222 | n10308 ;
  assign n23096 = n23095 ^ n6965 ^ n2641 ;
  assign n23097 = n16730 | n23096 ;
  assign n23098 = n23097 ^ n5983 ^ 1'b0 ;
  assign n23099 = ( n4396 & n10698 ) | ( n4396 & n10788 ) | ( n10698 & n10788 ) ;
  assign n23100 = n1758 & n8129 ;
  assign n23101 = n23100 ^ n3183 ^ 1'b0 ;
  assign n23102 = ( n3937 & n7875 ) | ( n3937 & ~n16289 ) | ( n7875 & ~n16289 ) ;
  assign n23103 = n23101 & ~n23102 ;
  assign n23104 = n23103 ^ n5664 ^ n4247 ;
  assign n23105 = ( n10402 & ~n11791 ) | ( n10402 & n23104 ) | ( ~n11791 & n23104 ) ;
  assign n23106 = ( n8660 & ~n23099 ) | ( n8660 & n23105 ) | ( ~n23099 & n23105 ) ;
  assign n23107 = n16008 ^ n3828 ^ 1'b0 ;
  assign n23108 = ~n18476 & n23107 ;
  assign n23109 = n2063 ^ n2024 ^ 1'b0 ;
  assign n23110 = n1172 & n23109 ;
  assign n23111 = n13231 & ~n23110 ;
  assign n23112 = ( n6293 & ~n8238 ) | ( n6293 & n14672 ) | ( ~n8238 & n14672 ) ;
  assign n23113 = n23112 ^ n2416 ^ 1'b0 ;
  assign n23114 = n9067 ^ n5064 ^ n4199 ;
  assign n23115 = n10950 ^ n6472 ^ n851 ;
  assign n23116 = n23115 ^ n20087 ^ 1'b0 ;
  assign n23119 = n13444 ^ n10341 ^ n2718 ;
  assign n23117 = ( ~n2855 & n5926 ) | ( ~n2855 & n12338 ) | ( n5926 & n12338 ) ;
  assign n23118 = ~n20285 & n23117 ;
  assign n23120 = n23119 ^ n23118 ^ 1'b0 ;
  assign n23121 = n14261 ^ n1905 ^ 1'b0 ;
  assign n23122 = ~n9497 & n23121 ;
  assign n23123 = n23122 ^ n17476 ^ n7376 ;
  assign n23124 = ( n20037 & n23120 ) | ( n20037 & ~n23123 ) | ( n23120 & ~n23123 ) ;
  assign n23125 = ( n7497 & n10845 ) | ( n7497 & n18957 ) | ( n10845 & n18957 ) ;
  assign n23138 = n12115 ^ n6278 ^ 1'b0 ;
  assign n23139 = n23138 ^ n13505 ^ n7696 ;
  assign n23136 = ( n5258 & n7495 ) | ( n5258 & ~n16268 ) | ( n7495 & ~n16268 ) ;
  assign n23126 = n1625 & n15832 ;
  assign n23127 = n19876 & ~n23126 ;
  assign n23128 = ~n10815 & n23127 ;
  assign n23129 = ( n5389 & n8309 ) | ( n5389 & n14198 ) | ( n8309 & n14198 ) ;
  assign n23130 = ( ~n3333 & n3833 ) | ( ~n3333 & n13109 ) | ( n3833 & n13109 ) ;
  assign n23131 = ( n5612 & n7467 ) | ( n5612 & n23130 ) | ( n7467 & n23130 ) ;
  assign n23132 = ( ~n11921 & n19915 ) | ( ~n11921 & n23131 ) | ( n19915 & n23131 ) ;
  assign n23133 = n23132 ^ n22707 ^ 1'b0 ;
  assign n23134 = ( n9083 & ~n23129 ) | ( n9083 & n23133 ) | ( ~n23129 & n23133 ) ;
  assign n23135 = ( n1627 & n23128 ) | ( n1627 & n23134 ) | ( n23128 & n23134 ) ;
  assign n23137 = n23136 ^ n23135 ^ 1'b0 ;
  assign n23140 = n23139 ^ n23137 ^ 1'b0 ;
  assign n23141 = ( ~n2446 & n3290 ) | ( ~n2446 & n10576 ) | ( n3290 & n10576 ) ;
  assign n23142 = ~n3384 & n6737 ;
  assign n23143 = n23142 ^ n6687 ^ n1600 ;
  assign n23144 = n11857 ^ n7745 ^ n2285 ;
  assign n23145 = ( n16374 & n19156 ) | ( n16374 & ~n23144 ) | ( n19156 & ~n23144 ) ;
  assign n23146 = n23145 ^ n13059 ^ n5772 ;
  assign n23147 = n23143 & n23146 ;
  assign n23148 = n23147 ^ n22773 ^ n18005 ;
  assign n23149 = n18648 ^ n4985 ^ n4603 ;
  assign n23150 = n10269 ^ n6654 ^ n318 ;
  assign n23151 = ( ~n2049 & n14130 ) | ( ~n2049 & n18173 ) | ( n14130 & n18173 ) ;
  assign n23152 = ( n23149 & ~n23150 ) | ( n23149 & n23151 ) | ( ~n23150 & n23151 ) ;
  assign n23153 = n14000 ^ n8095 ^ 1'b0 ;
  assign n23154 = n19360 & n23153 ;
  assign n23155 = ( n14734 & ~n23152 ) | ( n14734 & n23154 ) | ( ~n23152 & n23154 ) ;
  assign n23156 = ( n3976 & n3999 ) | ( n3976 & n18788 ) | ( n3999 & n18788 ) ;
  assign n23161 = n22570 ^ n1012 ^ 1'b0 ;
  assign n23162 = ~n16575 & n23161 ;
  assign n23157 = n10683 ^ n7411 ^ n4370 ;
  assign n23158 = n11866 ^ n3095 ^ n729 ;
  assign n23159 = ( n13439 & n23157 ) | ( n13439 & ~n23158 ) | ( n23157 & ~n23158 ) ;
  assign n23160 = n17355 | n23159 ;
  assign n23163 = n23162 ^ n23160 ^ 1'b0 ;
  assign n23164 = n21656 ^ n16622 ^ n11183 ;
  assign n23166 = n17607 ^ n11033 ^ n6023 ;
  assign n23165 = n12306 ^ n11864 ^ n2404 ;
  assign n23167 = n23166 ^ n23165 ^ n15436 ;
  assign n23168 = n17624 ^ n5685 ^ n2701 ;
  assign n23169 = ( n1896 & n2666 ) | ( n1896 & n23168 ) | ( n2666 & n23168 ) ;
  assign n23170 = ( x215 & ~n3277 ) | ( x215 & n12425 ) | ( ~n3277 & n12425 ) ;
  assign n23171 = n23170 ^ n16585 ^ n3822 ;
  assign n23172 = n23171 ^ n11421 ^ n5619 ;
  assign n23173 = n16763 ^ n5271 ^ 1'b0 ;
  assign n23174 = n23173 ^ n19008 ^ n1060 ;
  assign n23175 = n12319 ^ n1370 ^ 1'b0 ;
  assign n23176 = ( ~n15056 & n23174 ) | ( ~n15056 & n23175 ) | ( n23174 & n23175 ) ;
  assign n23177 = n23176 ^ n19533 ^ n2009 ;
  assign n23178 = n4995 | n21646 ;
  assign n23179 = n1970 & ~n23178 ;
  assign n23180 = n1427 & n10541 ;
  assign n23181 = n4081 ^ n894 ^ 1'b0 ;
  assign n23182 = ( ~n14464 & n23180 ) | ( ~n14464 & n23181 ) | ( n23180 & n23181 ) ;
  assign n23183 = n13311 ^ n13017 ^ n11233 ;
  assign n23185 = ( ~x231 & n763 ) | ( ~x231 & n3929 ) | ( n763 & n3929 ) ;
  assign n23184 = ~n9179 & n18724 ;
  assign n23186 = n23185 ^ n23184 ^ 1'b0 ;
  assign n23187 = n8442 & n12970 ;
  assign n23188 = n23187 ^ n15809 ^ n13370 ;
  assign n23194 = n10068 ^ n985 ^ 1'b0 ;
  assign n23189 = n7229 ^ n1738 ^ n1503 ;
  assign n23190 = n23189 ^ n14387 ^ n7271 ;
  assign n23191 = n14075 ^ n5737 ^ n4943 ;
  assign n23192 = x28 & n23191 ;
  assign n23193 = ( n16708 & n23190 ) | ( n16708 & ~n23192 ) | ( n23190 & ~n23192 ) ;
  assign n23195 = n23194 ^ n23193 ^ n11786 ;
  assign n23200 = ~n5373 & n19762 ;
  assign n23201 = ( n412 & n990 ) | ( n412 & ~n23200 ) | ( n990 & ~n23200 ) ;
  assign n23196 = ( n1407 & n4006 ) | ( n1407 & n7701 ) | ( n4006 & n7701 ) ;
  assign n23197 = ( ~n8497 & n8650 ) | ( ~n8497 & n22482 ) | ( n8650 & n22482 ) ;
  assign n23198 = n23196 & n23197 ;
  assign n23199 = ~n7683 & n23198 ;
  assign n23202 = n23201 ^ n23199 ^ n18212 ;
  assign n23203 = n13484 ^ n10873 ^ n10521 ;
  assign n23204 = ( ~n1215 & n13457 ) | ( ~n1215 & n23203 ) | ( n13457 & n23203 ) ;
  assign n23205 = n10091 & n23204 ;
  assign n23206 = n23205 ^ n8610 ^ n5112 ;
  assign n23207 = n14118 ^ n12669 ^ n6001 ;
  assign n23208 = ( n1288 & n12951 ) | ( n1288 & ~n23207 ) | ( n12951 & ~n23207 ) ;
  assign n23209 = ( ~n6276 & n22240 ) | ( ~n6276 & n23208 ) | ( n22240 & n23208 ) ;
  assign n23210 = ( n4140 & n6240 ) | ( n4140 & n18777 ) | ( n6240 & n18777 ) ;
  assign n23211 = n23210 ^ n18704 ^ n10811 ;
  assign n23212 = n20010 ^ n6414 ^ n692 ;
  assign n23213 = n5686 ^ n4440 ^ 1'b0 ;
  assign n23214 = n7403 ^ n5725 ^ n5220 ;
  assign n23215 = n23214 ^ n21983 ^ n3492 ;
  assign n23216 = n23215 ^ n17315 ^ n14223 ;
  assign n23217 = ( n2119 & ~n2665 ) | ( n2119 & n16069 ) | ( ~n2665 & n16069 ) ;
  assign n23218 = ( ~n6534 & n21899 ) | ( ~n6534 & n22707 ) | ( n21899 & n22707 ) ;
  assign n23219 = ~n15480 & n23218 ;
  assign n23220 = ( n13098 & ~n18237 ) | ( n13098 & n20287 ) | ( ~n18237 & n20287 ) ;
  assign n23221 = ( n5630 & n7383 ) | ( n5630 & ~n23220 ) | ( n7383 & ~n23220 ) ;
  assign n23222 = n23221 ^ n3205 ^ 1'b0 ;
  assign n23223 = n16202 ^ n8946 ^ n1789 ;
  assign n23226 = n9074 ^ n5906 ^ n3780 ;
  assign n23227 = n4388 & ~n23226 ;
  assign n23224 = n15115 & n20448 ;
  assign n23225 = n23224 ^ n11330 ^ 1'b0 ;
  assign n23228 = n23227 ^ n23225 ^ 1'b0 ;
  assign n23229 = n22688 ^ n9983 ^ 1'b0 ;
  assign n23230 = n18483 | n23229 ;
  assign n23231 = n11772 ^ n10144 ^ n3606 ;
  assign n23232 = n23231 ^ n7073 ^ 1'b0 ;
  assign n23233 = ~n23230 & n23232 ;
  assign n23234 = n13006 ^ n1891 ^ n487 ;
  assign n23235 = ( n3447 & ~n6711 ) | ( n3447 & n23234 ) | ( ~n6711 & n23234 ) ;
  assign n23236 = ( ~n14183 & n15141 ) | ( ~n14183 & n23235 ) | ( n15141 & n23235 ) ;
  assign n23237 = ( n7221 & n13582 ) | ( n7221 & ~n23236 ) | ( n13582 & ~n23236 ) ;
  assign n23238 = n8172 ^ n7149 ^ n2307 ;
  assign n23239 = n23238 ^ n13960 ^ n7943 ;
  assign n23240 = n23239 ^ n21966 ^ n19767 ;
  assign n23241 = ( n21441 & n22615 ) | ( n21441 & n23240 ) | ( n22615 & n23240 ) ;
  assign n23242 = n23241 ^ n19432 ^ n17095 ;
  assign n23243 = n8616 ^ n4356 ^ 1'b0 ;
  assign n23244 = ~n14622 & n23243 ;
  assign n23245 = ~n9915 & n23244 ;
  assign n23246 = ~n12953 & n23245 ;
  assign n23247 = ( n2440 & ~n4901 ) | ( n2440 & n23246 ) | ( ~n4901 & n23246 ) ;
  assign n23250 = n7433 ^ n6953 ^ n4850 ;
  assign n23251 = ( x204 & n698 ) | ( x204 & ~n23250 ) | ( n698 & ~n23250 ) ;
  assign n23249 = n3172 | n13775 ;
  assign n23248 = n22931 ^ n3561 ^ 1'b0 ;
  assign n23252 = n23251 ^ n23249 ^ n23248 ;
  assign n23253 = ( n10502 & n16432 ) | ( n10502 & n17334 ) | ( n16432 & n17334 ) ;
  assign n23254 = ( n3115 & ~n8050 ) | ( n3115 & n23253 ) | ( ~n8050 & n23253 ) ;
  assign n23255 = ~x151 & n21259 ;
  assign n23256 = n6394 ^ n630 ^ 1'b0 ;
  assign n23257 = ~n12349 & n23256 ;
  assign n23258 = ~n2597 & n11343 ;
  assign n23259 = n9087 & n23258 ;
  assign n23260 = n2605 & n14329 ;
  assign n23261 = ~n23259 & n23260 ;
  assign n23262 = n23257 & ~n23261 ;
  assign n23263 = n23262 ^ n21034 ^ 1'b0 ;
  assign n23264 = ( n3304 & n3724 ) | ( n3304 & ~n11539 ) | ( n3724 & ~n11539 ) ;
  assign n23265 = n20898 ^ n9061 ^ n5438 ;
  assign n23266 = n23265 ^ n22701 ^ n15405 ;
  assign n23267 = ( n4230 & n17400 ) | ( n4230 & n23266 ) | ( n17400 & n23266 ) ;
  assign n23268 = n10538 ^ n5938 ^ n354 ;
  assign n23269 = n23268 ^ n6308 ^ n4356 ;
  assign n23270 = ~n13616 & n21534 ;
  assign n23271 = n16952 ^ n4850 ^ n3414 ;
  assign n23272 = n17171 ^ n17142 ^ n13060 ;
  assign n23273 = n23272 ^ n21539 ^ 1'b0 ;
  assign n23274 = n15590 ^ n9155 ^ 1'b0 ;
  assign n23275 = n5861 ^ n4044 ^ 1'b0 ;
  assign n23276 = n22554 ^ n10212 ^ n4437 ;
  assign n23277 = n23276 ^ n3992 ^ n644 ;
  assign n23278 = n23277 ^ n19286 ^ n11137 ;
  assign n23279 = ( n9430 & n23275 ) | ( n9430 & ~n23278 ) | ( n23275 & ~n23278 ) ;
  assign n23280 = n23279 ^ n20811 ^ 1'b0 ;
  assign n23281 = ~n21310 & n23280 ;
  assign n23282 = n23281 ^ n16084 ^ 1'b0 ;
  assign n23283 = ( n1671 & ~n15559 ) | ( n1671 & n20156 ) | ( ~n15559 & n20156 ) ;
  assign n23284 = n12959 ^ n5882 ^ n3774 ;
  assign n23285 = n23284 ^ n7715 ^ 1'b0 ;
  assign n23286 = n14626 & ~n23285 ;
  assign n23287 = n8827 & n10522 ;
  assign n23288 = n20234 ^ n2102 ^ 1'b0 ;
  assign n23289 = ~n23287 & n23288 ;
  assign n23290 = n23289 ^ n21911 ^ n21420 ;
  assign n23291 = ( n2226 & n7217 ) | ( n2226 & n23290 ) | ( n7217 & n23290 ) ;
  assign n23292 = ( ~n3025 & n6875 ) | ( ~n3025 & n10358 ) | ( n6875 & n10358 ) ;
  assign n23294 = n15860 ^ n7822 ^ 1'b0 ;
  assign n23295 = n9178 | n23294 ;
  assign n23296 = n23295 ^ n5299 ^ n1288 ;
  assign n23293 = n3715 ^ n809 ^ 1'b0 ;
  assign n23297 = n23296 ^ n23293 ^ 1'b0 ;
  assign n23299 = n3761 ^ n2066 ^ n276 ;
  assign n23298 = n17931 ^ n9517 ^ n8173 ;
  assign n23300 = n23299 ^ n23298 ^ n16176 ;
  assign n23301 = ( n9514 & ~n13439 ) | ( n9514 & n21759 ) | ( ~n13439 & n21759 ) ;
  assign n23302 = ( n1312 & n8835 ) | ( n1312 & n10106 ) | ( n8835 & n10106 ) ;
  assign n23303 = n15994 | n23302 ;
  assign n23304 = n20873 | n23303 ;
  assign n23305 = ( ~n2516 & n9290 ) | ( ~n2516 & n13942 ) | ( n9290 & n13942 ) ;
  assign n23306 = ( n14290 & ~n16498 ) | ( n14290 & n23305 ) | ( ~n16498 & n23305 ) ;
  assign n23307 = n20573 ^ n19170 ^ 1'b0 ;
  assign n23308 = ~n8982 & n23307 ;
  assign n23309 = ( n13543 & n23306 ) | ( n13543 & ~n23308 ) | ( n23306 & ~n23308 ) ;
  assign n23310 = ( n653 & ~n1304 ) | ( n653 & n7618 ) | ( ~n1304 & n7618 ) ;
  assign n23311 = n7727 & ~n12183 ;
  assign n23312 = ~n12341 & n15028 ;
  assign n23313 = n23312 ^ n14767 ^ 1'b0 ;
  assign n23314 = ( n5183 & n23311 ) | ( n5183 & ~n23313 ) | ( n23311 & ~n23313 ) ;
  assign n23315 = ( n13363 & n23310 ) | ( n13363 & n23314 ) | ( n23310 & n23314 ) ;
  assign n23316 = n19453 ^ n3828 ^ n2521 ;
  assign n23320 = n17630 ^ n12716 ^ x92 ;
  assign n23317 = n15600 ^ n7381 ^ 1'b0 ;
  assign n23318 = n19057 ^ n14160 ^ 1'b0 ;
  assign n23319 = ( n15895 & n23317 ) | ( n15895 & n23318 ) | ( n23317 & n23318 ) ;
  assign n23321 = n23320 ^ n23319 ^ 1'b0 ;
  assign n23322 = ~n23316 & n23321 ;
  assign n23323 = ( ~n5010 & n15685 ) | ( ~n5010 & n17620 ) | ( n15685 & n17620 ) ;
  assign n23324 = n23323 ^ n626 ^ 1'b0 ;
  assign n23325 = ~n2850 & n15079 ;
  assign n23326 = ( n13463 & n15144 ) | ( n13463 & n23325 ) | ( n15144 & n23325 ) ;
  assign n23327 = ( n19190 & n23324 ) | ( n19190 & n23326 ) | ( n23324 & n23326 ) ;
  assign n23328 = n5583 ^ n2506 ^ n1378 ;
  assign n23329 = n1053 & n5674 ;
  assign n23330 = ( n11465 & n23328 ) | ( n11465 & ~n23329 ) | ( n23328 & ~n23329 ) ;
  assign n23336 = n21399 ^ n9537 ^ n5730 ;
  assign n23334 = n5400 & n10811 ;
  assign n23335 = ~n18766 & n23334 ;
  assign n23331 = ~n2134 & n10864 ;
  assign n23332 = n23331 ^ n9608 ^ n4907 ;
  assign n23333 = n23332 ^ n16396 ^ n3136 ;
  assign n23337 = n23336 ^ n23335 ^ n23333 ;
  assign n23338 = n11609 | n12108 ;
  assign n23339 = ( n4195 & n10356 ) | ( n4195 & n19344 ) | ( n10356 & n19344 ) ;
  assign n23340 = ( n3138 & ~n14976 ) | ( n3138 & n18102 ) | ( ~n14976 & n18102 ) ;
  assign n23341 = ( n341 & ~n8048 ) | ( n341 & n23340 ) | ( ~n8048 & n23340 ) ;
  assign n23342 = n15815 ^ n4166 ^ n2751 ;
  assign n23344 = n8202 ^ n4778 ^ n3087 ;
  assign n23343 = n7596 & ~n18067 ;
  assign n23345 = n23344 ^ n23343 ^ 1'b0 ;
  assign n23346 = ( n3313 & ~n9144 ) | ( n3313 & n13000 ) | ( ~n9144 & n13000 ) ;
  assign n23347 = n8805 & ~n23346 ;
  assign n23348 = n8906 ^ n4148 ^ n1958 ;
  assign n23349 = ( n10729 & n12932 ) | ( n10729 & ~n23348 ) | ( n12932 & ~n23348 ) ;
  assign n23350 = n20332 ^ n13148 ^ 1'b0 ;
  assign n23354 = ~n613 & n6432 ;
  assign n23355 = ( n1991 & ~n3223 ) | ( n1991 & n23354 ) | ( ~n3223 & n23354 ) ;
  assign n23356 = ( n2978 & n21009 ) | ( n2978 & ~n23355 ) | ( n21009 & ~n23355 ) ;
  assign n23352 = n14342 ^ n13340 ^ 1'b0 ;
  assign n23351 = n10809 ^ n6173 ^ 1'b0 ;
  assign n23353 = n23352 ^ n23351 ^ n5720 ;
  assign n23357 = n23356 ^ n23353 ^ n16546 ;
  assign n23360 = n8899 ^ n2700 ^ n1406 ;
  assign n23361 = n23360 ^ n6999 ^ n714 ;
  assign n23358 = ~n5006 & n7516 ;
  assign n23359 = n23358 ^ n15886 ^ 1'b0 ;
  assign n23362 = n23361 ^ n23359 ^ n23162 ;
  assign n23365 = ( x231 & n5127 ) | ( x231 & ~n13085 ) | ( n5127 & ~n13085 ) ;
  assign n23366 = n23365 ^ n18324 ^ n11246 ;
  assign n23363 = n14050 ^ n13344 ^ n10598 ;
  assign n23364 = n23363 ^ n8622 ^ n8591 ;
  assign n23367 = n23366 ^ n23364 ^ n16115 ;
  assign n23373 = n6514 | n10070 ;
  assign n23374 = n2443 & ~n23373 ;
  assign n23375 = ( ~n7240 & n14631 ) | ( ~n7240 & n23374 ) | ( n14631 & n23374 ) ;
  assign n23370 = ( n5384 & n6929 ) | ( n5384 & n9734 ) | ( n6929 & n9734 ) ;
  assign n23368 = n18997 ^ n1909 ^ 1'b0 ;
  assign n23369 = ~n12902 & n23368 ;
  assign n23371 = n23370 ^ n23369 ^ n3428 ;
  assign n23372 = ( n14586 & ~n22670 ) | ( n14586 & n23371 ) | ( ~n22670 & n23371 ) ;
  assign n23376 = n23375 ^ n23372 ^ n17024 ;
  assign n23379 = ~n2515 & n8057 ;
  assign n23380 = ( ~n10171 & n10356 ) | ( ~n10171 & n23379 ) | ( n10356 & n23379 ) ;
  assign n23377 = ( n2195 & ~n2567 ) | ( n2195 & n6754 ) | ( ~n2567 & n6754 ) ;
  assign n23378 = ( n2440 & n22685 ) | ( n2440 & n23377 ) | ( n22685 & n23377 ) ;
  assign n23381 = n23380 ^ n23378 ^ n17438 ;
  assign n23382 = ( n3427 & ~n4622 ) | ( n3427 & n7189 ) | ( ~n4622 & n7189 ) ;
  assign n23383 = n23382 ^ n12578 ^ n7191 ;
  assign n23384 = n7645 ^ n5819 ^ n1146 ;
  assign n23385 = n23384 ^ n7265 ^ n5156 ;
  assign n23386 = ~n15752 & n23385 ;
  assign n23387 = ~n23383 & n23386 ;
  assign n23388 = n1719 ^ n1638 ^ n774 ;
  assign n23389 = n12638 & n20904 ;
  assign n23390 = ( n11766 & n16769 ) | ( n11766 & n23389 ) | ( n16769 & n23389 ) ;
  assign n23391 = ~n23388 & n23390 ;
  assign n23392 = ~n12207 & n23391 ;
  assign n23393 = n763 | n1715 ;
  assign n23394 = n5836 & n12039 ;
  assign n23395 = n23393 & n23394 ;
  assign n23396 = n23395 ^ n13577 ^ n5228 ;
  assign n23397 = ( ~n5940 & n6452 ) | ( ~n5940 & n20628 ) | ( n6452 & n20628 ) ;
  assign n23398 = n16264 & n23397 ;
  assign n23399 = n21651 & n23398 ;
  assign n23400 = ( ~n3163 & n10259 ) | ( ~n3163 & n15592 ) | ( n10259 & n15592 ) ;
  assign n23401 = ( n3104 & n3946 ) | ( n3104 & n10681 ) | ( n3946 & n10681 ) ;
  assign n23402 = ~n3883 & n4806 ;
  assign n23403 = n7317 | n23402 ;
  assign n23404 = ~n2454 & n23403 ;
  assign n23405 = n23401 & n23404 ;
  assign n23406 = n14534 | n18940 ;
  assign n23407 = x33 | n23406 ;
  assign n23408 = n22833 ^ n7492 ^ n2622 ;
  assign n23409 = ~n10408 & n23408 ;
  assign n23417 = n2383 & n5143 ;
  assign n23414 = n8930 ^ n5502 ^ n799 ;
  assign n23415 = ( n8400 & ~n16138 ) | ( n8400 & n23414 ) | ( ~n16138 & n23414 ) ;
  assign n23412 = n12775 ^ n6737 ^ n5085 ;
  assign n23410 = n3913 & ~n6696 ;
  assign n23411 = n15025 & n23410 ;
  assign n23413 = n23412 ^ n23411 ^ n12162 ;
  assign n23416 = n23415 ^ n23413 ^ n8035 ;
  assign n23418 = n23417 ^ n23416 ^ n2885 ;
  assign n23419 = n23418 ^ n15953 ^ n7085 ;
  assign n23420 = ( n2870 & n10297 ) | ( n2870 & n14712 ) | ( n10297 & n14712 ) ;
  assign n23421 = n23420 ^ n9725 ^ 1'b0 ;
  assign n23422 = n21340 ^ n4729 ^ n961 ;
  assign n23423 = n21377 & n23422 ;
  assign n23424 = n23423 ^ n3771 ^ 1'b0 ;
  assign n23425 = n23424 ^ n911 ^ x79 ;
  assign n23432 = n13358 ^ n9972 ^ n1877 ;
  assign n23428 = n1846 & ~n4217 ;
  assign n23429 = n2729 & n23428 ;
  assign n23430 = n23429 ^ n22064 ^ 1'b0 ;
  assign n23431 = n23430 ^ n12496 ^ n11737 ;
  assign n23426 = ( ~n2608 & n11214 ) | ( ~n2608 & n19141 ) | ( n11214 & n19141 ) ;
  assign n23427 = n12634 & n23426 ;
  assign n23433 = n23432 ^ n23431 ^ n23427 ;
  assign n23434 = n11183 ^ n2177 ^ 1'b0 ;
  assign n23435 = n5566 & ~n23434 ;
  assign n23437 = ( n9011 & ~n12718 ) | ( n9011 & n18760 ) | ( ~n12718 & n18760 ) ;
  assign n23438 = ( x27 & n8353 ) | ( x27 & n23437 ) | ( n8353 & n23437 ) ;
  assign n23436 = ( n5974 & n12534 ) | ( n5974 & ~n14017 ) | ( n12534 & ~n14017 ) ;
  assign n23439 = n23438 ^ n23436 ^ n16841 ;
  assign n23440 = ( n20219 & n23435 ) | ( n20219 & ~n23439 ) | ( n23435 & ~n23439 ) ;
  assign n23441 = ( n5725 & ~n11324 ) | ( n5725 & n18857 ) | ( ~n11324 & n18857 ) ;
  assign n23442 = n22057 ^ n12693 ^ n10988 ;
  assign n23443 = n23442 ^ n22584 ^ n2526 ;
  assign n23444 = n23443 ^ n11126 ^ n2137 ;
  assign n23445 = n23444 ^ n16828 ^ n5427 ;
  assign n23446 = ( n2299 & ~n11486 ) | ( n2299 & n12508 ) | ( ~n11486 & n12508 ) ;
  assign n23447 = ( ~n4733 & n14310 ) | ( ~n4733 & n23446 ) | ( n14310 & n23446 ) ;
  assign n23448 = n23447 ^ n19839 ^ n15275 ;
  assign n23449 = ( n4178 & n12054 ) | ( n4178 & ~n23448 ) | ( n12054 & ~n23448 ) ;
  assign n23450 = ( n899 & ~n1758 ) | ( n899 & n12587 ) | ( ~n1758 & n12587 ) ;
  assign n23451 = n11989 ^ n8042 ^ n1455 ;
  assign n23452 = n23451 ^ n21130 ^ 1'b0 ;
  assign n23453 = n23450 & n23452 ;
  assign n23454 = n9964 & ~n22764 ;
  assign n23455 = n23454 ^ n21061 ^ n10912 ;
  assign n23456 = n9758 & n21925 ;
  assign n23457 = n321 & n23456 ;
  assign n23458 = n3625 & ~n23457 ;
  assign n23459 = ~n6963 & n23458 ;
  assign n23460 = n5149 & n23459 ;
  assign n23465 = ( n530 & ~n12159 ) | ( n530 & n15691 ) | ( ~n12159 & n15691 ) ;
  assign n23466 = n14673 & ~n23465 ;
  assign n23461 = n19531 ^ n8155 ^ 1'b0 ;
  assign n23462 = n8315 & ~n23461 ;
  assign n23463 = n23462 ^ n18837 ^ n16043 ;
  assign n23464 = n23463 ^ n2937 ^ n2660 ;
  assign n23467 = n23466 ^ n23464 ^ n2343 ;
  assign n23468 = n17878 ^ n2655 ^ 1'b0 ;
  assign n23469 = n3262 & n23468 ;
  assign n23470 = n1020 | n10578 ;
  assign n23471 = n7412 & ~n23470 ;
  assign n23472 = ( ~n8543 & n10455 ) | ( ~n8543 & n23471 ) | ( n10455 & n23471 ) ;
  assign n23474 = n4539 & ~n5698 ;
  assign n23473 = n17820 ^ n13635 ^ n1049 ;
  assign n23475 = n23474 ^ n23473 ^ 1'b0 ;
  assign n23477 = n1648 ^ n1598 ^ n1134 ;
  assign n23476 = ( n5655 & ~n11270 ) | ( n5655 & n19195 ) | ( ~n11270 & n19195 ) ;
  assign n23478 = n23477 ^ n23476 ^ n22636 ;
  assign n23479 = ( x200 & ~n5849 ) | ( x200 & n23478 ) | ( ~n5849 & n23478 ) ;
  assign n23480 = ( n4015 & n10557 ) | ( n4015 & ~n23479 ) | ( n10557 & ~n23479 ) ;
  assign n23481 = n17883 ^ n6632 ^ 1'b0 ;
  assign n23482 = n23481 ^ n13596 ^ n8438 ;
  assign n23483 = n23482 ^ n18308 ^ n12334 ;
  assign n23484 = ( ~n2119 & n9114 ) | ( ~n2119 & n13933 ) | ( n9114 & n13933 ) ;
  assign n23485 = n20058 ^ n16801 ^ n9654 ;
  assign n23486 = n23485 ^ n7808 ^ 1'b0 ;
  assign n23487 = ~n23484 & n23486 ;
  assign n23488 = n12026 ^ n2035 ^ 1'b0 ;
  assign n23489 = ( ~n4890 & n7002 ) | ( ~n4890 & n10259 ) | ( n7002 & n10259 ) ;
  assign n23490 = n23489 ^ n6572 ^ 1'b0 ;
  assign n23491 = n3063 ^ n2140 ^ 1'b0 ;
  assign n23494 = n2568 ^ n2389 ^ n2094 ;
  assign n23492 = ( x28 & ~n1896 ) | ( x28 & n8611 ) | ( ~n1896 & n8611 ) ;
  assign n23493 = ( ~n3767 & n17825 ) | ( ~n3767 & n23492 ) | ( n17825 & n23492 ) ;
  assign n23495 = n23494 ^ n23493 ^ n13105 ;
  assign n23496 = ( n21846 & n23491 ) | ( n21846 & n23495 ) | ( n23491 & n23495 ) ;
  assign n23497 = ( n10067 & ~n17454 ) | ( n10067 & n23496 ) | ( ~n17454 & n23496 ) ;
  assign n23498 = n19299 ^ n8681 ^ 1'b0 ;
  assign n23499 = n23498 ^ n22654 ^ n3661 ;
  assign n23502 = n3471 & n10608 ;
  assign n23503 = n23502 ^ n2081 ^ 1'b0 ;
  assign n23500 = n15399 ^ n12076 ^ n6597 ;
  assign n23501 = n20081 & n23500 ;
  assign n23504 = n23503 ^ n23501 ^ 1'b0 ;
  assign n23505 = n23504 ^ n19340 ^ n9578 ;
  assign n23506 = n23505 ^ n22066 ^ n3616 ;
  assign n23507 = ( ~n1923 & n4885 ) | ( ~n1923 & n23506 ) | ( n4885 & n23506 ) ;
  assign n23509 = n9535 ^ n5436 ^ n5237 ;
  assign n23510 = n2739 & ~n2741 ;
  assign n23511 = n23509 & n23510 ;
  assign n23508 = n22630 ^ n4554 ^ 1'b0 ;
  assign n23512 = n23511 ^ n23508 ^ n6527 ;
  assign n23513 = n16203 ^ n14613 ^ 1'b0 ;
  assign n23514 = n23513 ^ n5088 ^ n4624 ;
  assign n23515 = n23512 & n23514 ;
  assign n23516 = ~n9881 & n23515 ;
  assign n23519 = n13775 ^ n8569 ^ n5318 ;
  assign n23520 = n23519 ^ n18788 ^ 1'b0 ;
  assign n23517 = ( x222 & n1778 ) | ( x222 & ~n9905 ) | ( n1778 & ~n9905 ) ;
  assign n23518 = n23517 ^ n18243 ^ 1'b0 ;
  assign n23521 = n23520 ^ n23518 ^ n16153 ;
  assign n23522 = n1043 & ~n23521 ;
  assign n23523 = ~n4545 & n21377 ;
  assign n23524 = n23523 ^ n4210 ^ 1'b0 ;
  assign n23525 = n23524 ^ n6080 ^ n4899 ;
  assign n23526 = n23525 ^ n16466 ^ n1379 ;
  assign n23527 = n16729 ^ n9685 ^ n1057 ;
  assign n23528 = n19289 ^ n19165 ^ n13160 ;
  assign n23529 = n23119 ^ n21561 ^ n8332 ;
  assign n23530 = n13126 & ~n15865 ;
  assign n23531 = ( ~n11059 & n13115 ) | ( ~n11059 & n15570 ) | ( n13115 & n15570 ) ;
  assign n23532 = n2811 | n23531 ;
  assign n23533 = n23530 | n23532 ;
  assign n23534 = n17660 ^ n5591 ^ n3566 ;
  assign n23535 = ( n7784 & ~n8828 ) | ( n7784 & n9630 ) | ( ~n8828 & n9630 ) ;
  assign n23536 = n19671 ^ n15512 ^ x92 ;
  assign n23537 = ( ~n904 & n8856 ) | ( ~n904 & n9499 ) | ( n8856 & n9499 ) ;
  assign n23538 = n23537 ^ n8131 ^ n5720 ;
  assign n23539 = n23538 ^ n19962 ^ n18507 ;
  assign n23540 = n13594 ^ n8876 ^ 1'b0 ;
  assign n23541 = ( x189 & n13812 ) | ( x189 & n15353 ) | ( n13812 & n15353 ) ;
  assign n23542 = ( n13690 & n19706 ) | ( n13690 & n23541 ) | ( n19706 & n23541 ) ;
  assign n23543 = n10287 ^ n7744 ^ n3071 ;
  assign n23544 = n23543 ^ n20841 ^ n7962 ;
  assign n23550 = ( n3410 & n6516 ) | ( n3410 & n6909 ) | ( n6516 & n6909 ) ;
  assign n23545 = ( ~n876 & n13297 ) | ( ~n876 & n21719 ) | ( n13297 & n21719 ) ;
  assign n23546 = n22291 ^ n3987 ^ 1'b0 ;
  assign n23547 = n5895 & n23546 ;
  assign n23548 = n23547 ^ n10064 ^ n9625 ;
  assign n23549 = ( n9323 & n23545 ) | ( n9323 & ~n23548 ) | ( n23545 & ~n23548 ) ;
  assign n23551 = n23550 ^ n23549 ^ n12169 ;
  assign n23552 = ( n23036 & n23544 ) | ( n23036 & n23551 ) | ( n23544 & n23551 ) ;
  assign n23553 = n10319 ^ n4673 ^ n2174 ;
  assign n23554 = n23553 ^ n2344 ^ 1'b0 ;
  assign n23555 = n6655 & ~n23554 ;
  assign n23556 = n23555 ^ n10498 ^ 1'b0 ;
  assign n23557 = ( n5849 & n7990 ) | ( n5849 & ~n23556 ) | ( n7990 & ~n23556 ) ;
  assign n23558 = n23557 ^ n2275 ^ n2185 ;
  assign n23559 = n18611 ^ n16262 ^ n12228 ;
  assign n23560 = n21060 ^ n3916 ^ n3851 ;
  assign n23561 = ~n491 & n14336 ;
  assign n23562 = ~n20038 & n23561 ;
  assign n23563 = ( ~n4763 & n5898 ) | ( ~n4763 & n8582 ) | ( n5898 & n8582 ) ;
  assign n23564 = n19360 | n23563 ;
  assign n23565 = ( ~n3284 & n17555 ) | ( ~n3284 & n19226 ) | ( n17555 & n19226 ) ;
  assign n23566 = n23565 ^ n19039 ^ n6221 ;
  assign n23567 = ( n2245 & n8030 ) | ( n2245 & ~n12260 ) | ( n8030 & ~n12260 ) ;
  assign n23568 = n23567 ^ n6689 ^ n5887 ;
  assign n23569 = n23566 & ~n23568 ;
  assign n23570 = n1776 & ~n23569 ;
  assign n23571 = n23570 ^ n8346 ^ 1'b0 ;
  assign n23572 = ~n2686 & n23098 ;
  assign n23573 = ( n4894 & ~n6442 ) | ( n4894 & n11504 ) | ( ~n6442 & n11504 ) ;
  assign n23574 = n21791 ^ n1489 ^ 1'b0 ;
  assign n23575 = ~n23573 & n23574 ;
  assign n23576 = ~n21015 & n23575 ;
  assign n23577 = n23576 ^ n9884 ^ 1'b0 ;
  assign n23579 = ( n4590 & n6836 ) | ( n4590 & n19297 ) | ( n6836 & n19297 ) ;
  assign n23580 = n23579 ^ n22498 ^ n9220 ;
  assign n23578 = ~n1233 & n13145 ;
  assign n23581 = n23580 ^ n23578 ^ n19095 ;
  assign n23587 = ( ~n5861 & n8714 ) | ( ~n5861 & n12451 ) | ( n8714 & n12451 ) ;
  assign n23588 = n8910 ^ n8451 ^ n3561 ;
  assign n23589 = n23587 & ~n23588 ;
  assign n23590 = n23589 ^ n1529 ^ 1'b0 ;
  assign n23591 = n23590 ^ n15734 ^ n7058 ;
  assign n23582 = ~n637 & n21939 ;
  assign n23583 = ( n7493 & n21047 ) | ( n7493 & n23582 ) | ( n21047 & n23582 ) ;
  assign n23584 = n3410 & ~n5719 ;
  assign n23585 = n23583 | n23584 ;
  assign n23586 = n23585 ^ n13977 ^ 1'b0 ;
  assign n23592 = n23591 ^ n23586 ^ n9653 ;
  assign n23593 = n16855 ^ n3404 ^ n342 ;
  assign n23594 = n23593 ^ n1414 ^ 1'b0 ;
  assign n23595 = ( ~n8906 & n13984 ) | ( ~n8906 & n15479 ) | ( n13984 & n15479 ) ;
  assign n23598 = n11413 ^ n9396 ^ n401 ;
  assign n23599 = n4604 | n6624 ;
  assign n23600 = n2261 | n23599 ;
  assign n23601 = n23600 ^ n3595 ^ 1'b0 ;
  assign n23602 = n23598 & n23601 ;
  assign n23596 = n8573 ^ n548 ^ n436 ;
  assign n23597 = n6209 & ~n23596 ;
  assign n23603 = n23602 ^ n23597 ^ 1'b0 ;
  assign n23604 = n23603 ^ n18871 ^ n15960 ;
  assign n23605 = ( n18466 & n23595 ) | ( n18466 & n23604 ) | ( n23595 & n23604 ) ;
  assign n23607 = x34 & ~n2800 ;
  assign n23608 = n23607 ^ n8456 ^ 1'b0 ;
  assign n23606 = ( n4120 & n4227 ) | ( n4120 & ~n14240 ) | ( n4227 & ~n14240 ) ;
  assign n23609 = n23608 ^ n23606 ^ n9619 ;
  assign n23610 = n10274 ^ n3342 ^ 1'b0 ;
  assign n23611 = n1353 & n23610 ;
  assign n23612 = n15829 ^ n7152 ^ n1918 ;
  assign n23613 = n7727 ^ n3747 ^ n371 ;
  assign n23614 = n23613 ^ n15547 ^ n8533 ;
  assign n23615 = n22974 ^ n12957 ^ 1'b0 ;
  assign n23616 = n2400 | n23615 ;
  assign n23617 = n2056 & ~n5317 ;
  assign n23618 = ~n5462 & n23617 ;
  assign n23619 = n16149 ^ n394 ^ 1'b0 ;
  assign n23620 = n10292 | n23619 ;
  assign n23621 = ( n12597 & n23618 ) | ( n12597 & n23620 ) | ( n23618 & n23620 ) ;
  assign n23622 = n23621 ^ n13708 ^ n4389 ;
  assign n23623 = n23622 ^ n6935 ^ x107 ;
  assign n23637 = n6632 ^ n6050 ^ n3051 ;
  assign n23638 = ( ~n946 & n6841 ) | ( ~n946 & n19078 ) | ( n6841 & n19078 ) ;
  assign n23639 = n6977 | n23638 ;
  assign n23640 = n23637 & ~n23639 ;
  assign n23633 = ( n702 & ~n3841 ) | ( n702 & n8968 ) | ( ~n3841 & n8968 ) ;
  assign n23634 = ( ~n8048 & n14501 ) | ( ~n8048 & n23633 ) | ( n14501 & n23633 ) ;
  assign n23635 = n17128 ^ n11865 ^ n9345 ;
  assign n23636 = n23634 & ~n23635 ;
  assign n23624 = n19809 ^ n5504 ^ n1004 ;
  assign n23625 = n10320 ^ n1143 ^ 1'b0 ;
  assign n23626 = n23624 | n23625 ;
  assign n23627 = ( n5247 & ~n14116 ) | ( n5247 & n23626 ) | ( ~n14116 & n23626 ) ;
  assign n23628 = n23627 ^ n11207 ^ 1'b0 ;
  assign n23629 = n1135 & n1268 ;
  assign n23630 = ~n4388 & n23629 ;
  assign n23631 = n3378 & ~n23630 ;
  assign n23632 = n23628 & n23631 ;
  assign n23641 = n23640 ^ n23636 ^ n23632 ;
  assign n23642 = n9512 ^ n4308 ^ 1'b0 ;
  assign n23643 = ( ~n11126 & n12017 ) | ( ~n11126 & n20661 ) | ( n12017 & n20661 ) ;
  assign n23644 = n16926 & n23643 ;
  assign n23645 = n11624 ^ n10509 ^ n1561 ;
  assign n23646 = n23366 & ~n23645 ;
  assign n23647 = ~n14583 & n23646 ;
  assign n23648 = ( n7624 & n23222 ) | ( n7624 & ~n23647 ) | ( n23222 & ~n23647 ) ;
  assign n23649 = n5086 | n11018 ;
  assign n23650 = n23649 ^ n3810 ^ 1'b0 ;
  assign n23651 = n23650 ^ n3764 ^ n1696 ;
  assign n23652 = n23651 ^ n21109 ^ n2544 ;
  assign n23653 = n22266 ^ n9385 ^ n6256 ;
  assign n23654 = ( n2850 & n13406 ) | ( n2850 & ~n14111 ) | ( n13406 & ~n14111 ) ;
  assign n23657 = n7510 | n9220 ;
  assign n23658 = n23657 ^ n2328 ^ 1'b0 ;
  assign n23656 = n2024 & ~n7698 ;
  assign n23655 = n6347 ^ n2808 ^ 1'b0 ;
  assign n23659 = n23658 ^ n23656 ^ n23655 ;
  assign n23662 = ( n1634 & n2026 ) | ( n1634 & ~n12951 ) | ( n2026 & ~n12951 ) ;
  assign n23663 = ( n2335 & n12382 ) | ( n2335 & ~n23662 ) | ( n12382 & ~n23662 ) ;
  assign n23661 = ( n999 & n1943 ) | ( n999 & n8803 ) | ( n1943 & n8803 ) ;
  assign n23660 = ( n6123 & n11353 ) | ( n6123 & ~n18725 ) | ( n11353 & ~n18725 ) ;
  assign n23664 = n23663 ^ n23661 ^ n23660 ;
  assign n23665 = n9389 ^ n1873 ^ 1'b0 ;
  assign n23671 = n4359 ^ n1562 ^ 1'b0 ;
  assign n23669 = ( n7319 & ~n12090 ) | ( n7319 & n15541 ) | ( ~n12090 & n15541 ) ;
  assign n23670 = n23669 ^ n5073 ^ 1'b0 ;
  assign n23666 = n12063 ^ n2155 ^ 1'b0 ;
  assign n23667 = n1079 & n23666 ;
  assign n23668 = ( n11832 & n15214 ) | ( n11832 & ~n23667 ) | ( n15214 & ~n23667 ) ;
  assign n23672 = n23671 ^ n23670 ^ n23668 ;
  assign n23673 = ~n3790 & n7098 ;
  assign n23674 = n13854 | n23673 ;
  assign n23675 = n8290 & ~n23674 ;
  assign n23679 = n10045 ^ n4224 ^ 1'b0 ;
  assign n23680 = ( ~n3847 & n7011 ) | ( ~n3847 & n23679 ) | ( n7011 & n23679 ) ;
  assign n23676 = ( n1698 & n6267 ) | ( n1698 & ~n10117 ) | ( n6267 & ~n10117 ) ;
  assign n23677 = n23676 ^ n9718 ^ n1611 ;
  assign n23678 = ( n21905 & ~n22995 ) | ( n21905 & n23677 ) | ( ~n22995 & n23677 ) ;
  assign n23681 = n23680 ^ n23678 ^ n5509 ;
  assign n23682 = n17557 ^ n6482 ^ n476 ;
  assign n23683 = ( n4993 & ~n19399 ) | ( n4993 & n23682 ) | ( ~n19399 & n23682 ) ;
  assign n23692 = ( ~n6822 & n7837 ) | ( ~n6822 & n8178 ) | ( n7837 & n8178 ) ;
  assign n23684 = n3054 & ~n5869 ;
  assign n23685 = n23684 ^ x86 ^ 1'b0 ;
  assign n23686 = ( n6570 & n17691 ) | ( n6570 & ~n23685 ) | ( n17691 & ~n23685 ) ;
  assign n23687 = n9121 | n23686 ;
  assign n23688 = n23687 ^ n9270 ^ 1'b0 ;
  assign n23689 = ~n2223 & n23688 ;
  assign n23690 = ( n9421 & ~n12746 ) | ( n9421 & n23689 ) | ( ~n12746 & n23689 ) ;
  assign n23691 = ~n15011 & n23690 ;
  assign n23693 = n23692 ^ n23691 ^ 1'b0 ;
  assign n23695 = ( x121 & n271 ) | ( x121 & n412 ) | ( n271 & n412 ) ;
  assign n23694 = n14992 | n18980 ;
  assign n23696 = n23695 ^ n23694 ^ 1'b0 ;
  assign n23697 = n20172 ^ n500 ^ 1'b0 ;
  assign n23698 = ( n3673 & n5167 ) | ( n3673 & n13292 ) | ( n5167 & n13292 ) ;
  assign n23699 = ( n1226 & n7799 ) | ( n1226 & ~n8874 ) | ( n7799 & ~n8874 ) ;
  assign n23700 = n23699 ^ n9874 ^ n6087 ;
  assign n23705 = n14894 ^ n13325 ^ n9087 ;
  assign n23701 = n14922 ^ n856 ^ x15 ;
  assign n23702 = n22565 ^ n3550 ^ n362 ;
  assign n23703 = n23702 ^ n11668 ^ 1'b0 ;
  assign n23704 = ( n19198 & ~n23701 ) | ( n19198 & n23703 ) | ( ~n23701 & n23703 ) ;
  assign n23706 = n23705 ^ n23704 ^ n11038 ;
  assign n23707 = ~n9197 & n14645 ;
  assign n23708 = n7839 | n23707 ;
  assign n23709 = n23708 ^ n8352 ^ n4564 ;
  assign n23710 = n21860 ^ n19592 ^ n4939 ;
  assign n23711 = n23710 ^ n9166 ^ 1'b0 ;
  assign n23712 = n23709 & n23711 ;
  assign n23719 = n5034 | n16460 ;
  assign n23720 = n23719 ^ n18363 ^ 1'b0 ;
  assign n23718 = n6119 & ~n17383 ;
  assign n23721 = n23720 ^ n23718 ^ 1'b0 ;
  assign n23713 = ~n3620 & n10658 ;
  assign n23714 = n23713 ^ n9422 ^ 1'b0 ;
  assign n23715 = ( n6167 & n9844 ) | ( n6167 & n11561 ) | ( n9844 & n11561 ) ;
  assign n23716 = n19280 & n23715 ;
  assign n23717 = ~n23714 & n23716 ;
  assign n23722 = n23721 ^ n23717 ^ n23231 ;
  assign n23726 = ( n15706 & ~n16349 ) | ( n15706 & n22777 ) | ( ~n16349 & n22777 ) ;
  assign n23723 = ~n2633 & n2708 ;
  assign n23724 = n23723 ^ n5929 ^ 1'b0 ;
  assign n23725 = n23724 ^ n4015 ^ 1'b0 ;
  assign n23727 = n23726 ^ n23725 ^ n7784 ;
  assign n23728 = ( ~n320 & n1905 ) | ( ~n320 & n16094 ) | ( n1905 & n16094 ) ;
  assign n23729 = ( ~n8765 & n22208 ) | ( ~n8765 & n23728 ) | ( n22208 & n23728 ) ;
  assign n23730 = ( n1757 & n7061 ) | ( n1757 & n15947 ) | ( n7061 & n15947 ) ;
  assign n23731 = ( ~n5039 & n23729 ) | ( ~n5039 & n23730 ) | ( n23729 & n23730 ) ;
  assign n23732 = n11387 ^ n7684 ^ n3523 ;
  assign n23733 = n8489 & n17196 ;
  assign n23734 = n23733 ^ n18409 ^ 1'b0 ;
  assign n23735 = n13812 ^ n2773 ^ 1'b0 ;
  assign n23736 = n23734 & n23735 ;
  assign n23737 = ( n12099 & n23732 ) | ( n12099 & n23736 ) | ( n23732 & n23736 ) ;
  assign n23738 = n23737 ^ n10249 ^ n8091 ;
  assign n23739 = n1780 & n23738 ;
  assign n23740 = n12479 ^ n5115 ^ 1'b0 ;
  assign n23741 = ( n1891 & ~n4108 ) | ( n1891 & n5700 ) | ( ~n4108 & n5700 ) ;
  assign n23742 = n9714 | n23741 ;
  assign n23743 = n23740 | n23742 ;
  assign n23744 = n23743 ^ n20617 ^ n10050 ;
  assign n23745 = n9975 ^ n7975 ^ 1'b0 ;
  assign n23746 = ( ~n17123 & n22655 ) | ( ~n17123 & n23745 ) | ( n22655 & n23745 ) ;
  assign n23747 = ( ~n1046 & n10153 ) | ( ~n1046 & n23746 ) | ( n10153 & n23746 ) ;
  assign n23751 = n15541 ^ n12790 ^ n3448 ;
  assign n23748 = n2375 ^ n839 ^ 1'b0 ;
  assign n23749 = n3414 & n23748 ;
  assign n23750 = ( n572 & n18593 ) | ( n572 & ~n23749 ) | ( n18593 & ~n23749 ) ;
  assign n23752 = n23751 ^ n23750 ^ n7032 ;
  assign n23753 = n23752 ^ n9246 ^ n3923 ;
  assign n23754 = n18575 ^ n15821 ^ 1'b0 ;
  assign n23755 = n20750 & ~n23754 ;
  assign n23756 = n23755 ^ n15031 ^ 1'b0 ;
  assign n23757 = ( n8101 & n19023 ) | ( n8101 & ~n20184 ) | ( n19023 & ~n20184 ) ;
  assign n23758 = ( ~n9205 & n14573 ) | ( ~n9205 & n20448 ) | ( n14573 & n20448 ) ;
  assign n23759 = n23758 ^ n18457 ^ n12224 ;
  assign n23760 = ( ~n6030 & n8378 ) | ( ~n6030 & n22681 ) | ( n8378 & n22681 ) ;
  assign n23761 = ( n7066 & ~n7384 ) | ( n7066 & n21126 ) | ( ~n7384 & n21126 ) ;
  assign n23762 = ( n6556 & n6669 ) | ( n6556 & ~n23761 ) | ( n6669 & ~n23761 ) ;
  assign n23763 = ( ~n9692 & n11597 ) | ( ~n9692 & n23762 ) | ( n11597 & n23762 ) ;
  assign n23764 = n23760 | n23763 ;
  assign n23765 = ( n4388 & ~n20668 ) | ( n4388 & n23131 ) | ( ~n20668 & n23131 ) ;
  assign n23766 = ( n711 & n5529 ) | ( n711 & ~n20058 ) | ( n5529 & ~n20058 ) ;
  assign n23767 = ( ~n10269 & n14586 ) | ( ~n10269 & n23766 ) | ( n14586 & n23766 ) ;
  assign n23768 = ( ~n12281 & n23765 ) | ( ~n12281 & n23767 ) | ( n23765 & n23767 ) ;
  assign n23769 = ~n23764 & n23768 ;
  assign n23770 = n6493 ^ n4397 ^ 1'b0 ;
  assign n23771 = n23770 ^ n3459 ^ n2762 ;
  assign n23772 = ( n805 & n2313 ) | ( n805 & ~n3525 ) | ( n2313 & ~n3525 ) ;
  assign n23773 = ( ~n2700 & n23771 ) | ( ~n2700 & n23772 ) | ( n23771 & n23772 ) ;
  assign n23774 = ( n437 & n1278 ) | ( n437 & ~n6885 ) | ( n1278 & ~n6885 ) ;
  assign n23776 = n12138 ^ n6111 ^ n2260 ;
  assign n23777 = n20383 | n23776 ;
  assign n23778 = n23777 ^ n9734 ^ 1'b0 ;
  assign n23779 = ( n2988 & ~n3315 ) | ( n2988 & n3731 ) | ( ~n3315 & n3731 ) ;
  assign n23780 = ( ~n3115 & n23778 ) | ( ~n3115 & n23779 ) | ( n23778 & n23779 ) ;
  assign n23775 = ( n682 & n845 ) | ( n682 & ~n6932 ) | ( n845 & ~n6932 ) ;
  assign n23781 = n23780 ^ n23775 ^ n2325 ;
  assign n23782 = n21470 ^ n9067 ^ 1'b0 ;
  assign n23783 = n23781 | n23782 ;
  assign n23784 = ( n23773 & ~n23774 ) | ( n23773 & n23783 ) | ( ~n23774 & n23783 ) ;
  assign n23785 = ~n2724 & n12309 ;
  assign n23786 = ( ~n4837 & n5504 ) | ( ~n4837 & n23785 ) | ( n5504 & n23785 ) ;
  assign n23787 = n23786 ^ n15092 ^ n10498 ;
  assign n23788 = ( ~n8484 & n23784 ) | ( ~n8484 & n23787 ) | ( n23784 & n23787 ) ;
  assign n23789 = ( n5480 & n8253 ) | ( n5480 & n23714 ) | ( n8253 & n23714 ) ;
  assign n23790 = n3705 & n8282 ;
  assign n23791 = n23789 & n23790 ;
  assign n23792 = n17231 ^ n6798 ^ 1'b0 ;
  assign n23793 = ~n17890 & n23792 ;
  assign n23794 = ( ~n11026 & n12691 ) | ( ~n11026 & n14061 ) | ( n12691 & n14061 ) ;
  assign n23795 = ( n20102 & n23793 ) | ( n20102 & ~n23794 ) | ( n23793 & ~n23794 ) ;
  assign n23796 = n2197 ^ n798 ^ x48 ;
  assign n23797 = ( n6560 & n11311 ) | ( n6560 & n23796 ) | ( n11311 & n23796 ) ;
  assign n23798 = ( n2645 & n3509 ) | ( n2645 & ~n15489 ) | ( n3509 & ~n15489 ) ;
  assign n23800 = n8201 ^ n8002 ^ n1507 ;
  assign n23799 = ( n920 & ~n2600 ) | ( n920 & n3104 ) | ( ~n2600 & n3104 ) ;
  assign n23801 = n23800 ^ n23799 ^ n10304 ;
  assign n23802 = ( n9048 & ~n23798 ) | ( n9048 & n23801 ) | ( ~n23798 & n23801 ) ;
  assign n23803 = n23802 ^ n23189 ^ n21969 ;
  assign n23804 = n3054 & n4794 ;
  assign n23808 = ( ~n634 & n4252 ) | ( ~n634 & n7316 ) | ( n4252 & n7316 ) ;
  assign n23809 = ( n7044 & n19511 ) | ( n7044 & ~n23808 ) | ( n19511 & ~n23808 ) ;
  assign n23805 = n3186 & ~n20876 ;
  assign n23806 = n8899 & n23805 ;
  assign n23807 = n23806 ^ n3051 ^ n2368 ;
  assign n23810 = n23809 ^ n23807 ^ n18453 ;
  assign n23811 = ( n11840 & n12273 ) | ( n11840 & ~n14763 ) | ( n12273 & ~n14763 ) ;
  assign n23812 = ( n7469 & n9589 ) | ( n7469 & n11392 ) | ( n9589 & n11392 ) ;
  assign n23813 = ( ~n833 & n22040 ) | ( ~n833 & n23812 ) | ( n22040 & n23812 ) ;
  assign n23814 = n327 & ~n23813 ;
  assign n23815 = ~n7135 & n23814 ;
  assign n23816 = n23815 ^ n22094 ^ 1'b0 ;
  assign n23817 = ~n2222 & n23816 ;
  assign n23818 = n366 & ~n10435 ;
  assign n23819 = n23818 ^ n400 ^ 1'b0 ;
  assign n23820 = n23819 ^ n14488 ^ 1'b0 ;
  assign n23821 = n13612 ^ n1561 ^ n985 ;
  assign n23822 = n23821 ^ n7518 ^ 1'b0 ;
  assign n23823 = n19604 & ~n23822 ;
  assign n23824 = ( ~n1554 & n5872 ) | ( ~n1554 & n10944 ) | ( n5872 & n10944 ) ;
  assign n23825 = n20572 ^ n8285 ^ n2097 ;
  assign n23826 = n1502 | n15934 ;
  assign n23827 = n13996 & ~n23826 ;
  assign n23828 = ~n7240 & n17975 ;
  assign n23829 = n9424 & n23828 ;
  assign n23830 = ( ~n3621 & n10416 ) | ( ~n3621 & n23829 ) | ( n10416 & n23829 ) ;
  assign n23831 = ( ~n11203 & n23827 ) | ( ~n11203 & n23830 ) | ( n23827 & n23830 ) ;
  assign n23832 = ( n426 & n8808 ) | ( n426 & ~n19375 ) | ( n8808 & ~n19375 ) ;
  assign n23833 = n23832 ^ n20978 ^ n7561 ;
  assign n23834 = n17555 ^ n3145 ^ 1'b0 ;
  assign n23835 = ~n23833 & n23834 ;
  assign n23838 = n7697 ^ n400 ^ 1'b0 ;
  assign n23839 = n23838 ^ n17505 ^ n2368 ;
  assign n23840 = ( ~n7215 & n8685 ) | ( ~n7215 & n9734 ) | ( n8685 & n9734 ) ;
  assign n23841 = ( n14705 & n23839 ) | ( n14705 & n23840 ) | ( n23839 & n23840 ) ;
  assign n23842 = ( ~n2243 & n21778 ) | ( ~n2243 & n23841 ) | ( n21778 & n23841 ) ;
  assign n23836 = n14685 ^ n12634 ^ n5369 ;
  assign n23837 = n23836 ^ n3981 ^ n2012 ;
  assign n23843 = n23842 ^ n23837 ^ n2918 ;
  assign n23844 = ( n2442 & n18918 ) | ( n2442 & ~n23843 ) | ( n18918 & ~n23843 ) ;
  assign n23845 = ~n2686 & n15780 ;
  assign n23846 = ( n1822 & n6747 ) | ( n1822 & n15574 ) | ( n6747 & n15574 ) ;
  assign n23847 = n9629 & n20154 ;
  assign n23848 = n23847 ^ n21732 ^ 1'b0 ;
  assign n23849 = ( n2127 & ~n22977 ) | ( n2127 & n23848 ) | ( ~n22977 & n23848 ) ;
  assign n23850 = n11557 | n15277 ;
  assign n23851 = n23850 ^ n2054 ^ 1'b0 ;
  assign n23852 = ( n6612 & n13796 ) | ( n6612 & ~n17646 ) | ( n13796 & ~n17646 ) ;
  assign n23853 = n8579 ^ n7615 ^ 1'b0 ;
  assign n23854 = n7044 & n23853 ;
  assign n23855 = n22788 | n23854 ;
  assign n23856 = ( ~n2223 & n2479 ) | ( ~n2223 & n4361 ) | ( n2479 & n4361 ) ;
  assign n23857 = ( n4264 & n6729 ) | ( n4264 & ~n15766 ) | ( n6729 & ~n15766 ) ;
  assign n23858 = ( n9067 & n23856 ) | ( n9067 & n23857 ) | ( n23856 & n23857 ) ;
  assign n23860 = n11911 ^ n9813 ^ n9611 ;
  assign n23859 = ( n2864 & ~n6467 ) | ( n2864 & n6911 ) | ( ~n6467 & n6911 ) ;
  assign n23861 = n23860 ^ n23859 ^ n361 ;
  assign n23865 = ( n854 & n2895 ) | ( n854 & ~n5820 ) | ( n2895 & ~n5820 ) ;
  assign n23862 = ( n5722 & n7380 ) | ( n5722 & ~n20868 ) | ( n7380 & ~n20868 ) ;
  assign n23863 = n23862 ^ n20491 ^ n8218 ;
  assign n23864 = ( n14161 & n21020 ) | ( n14161 & ~n23863 ) | ( n21020 & ~n23863 ) ;
  assign n23866 = n23865 ^ n23864 ^ n19918 ;
  assign n23867 = ( n2976 & n4238 ) | ( n2976 & ~n7308 ) | ( n4238 & ~n7308 ) ;
  assign n23868 = n19077 & ~n23867 ;
  assign n23870 = n8839 ^ n4345 ^ n2235 ;
  assign n23871 = n23870 ^ n6404 ^ n387 ;
  assign n23872 = ( ~n1475 & n11554 ) | ( ~n1475 & n23871 ) | ( n11554 & n23871 ) ;
  assign n23869 = n9424 ^ n8689 ^ 1'b0 ;
  assign n23873 = n23872 ^ n23869 ^ n4097 ;
  assign n23874 = ( ~n8226 & n23868 ) | ( ~n8226 & n23873 ) | ( n23868 & n23873 ) ;
  assign n23875 = ( n5845 & ~n16466 ) | ( n5845 & n23149 ) | ( ~n16466 & n23149 ) ;
  assign n23876 = n23875 ^ n22903 ^ n16529 ;
  assign n23877 = ( n1376 & n7525 ) | ( n1376 & n23876 ) | ( n7525 & n23876 ) ;
  assign n23878 = n23877 ^ n10250 ^ n3025 ;
  assign n23884 = n8519 ^ n8014 ^ n1737 ;
  assign n23882 = n12333 ^ n8946 ^ n5138 ;
  assign n23883 = ~n8348 & n23882 ;
  assign n23885 = n23884 ^ n23883 ^ 1'b0 ;
  assign n23879 = x64 & ~n6463 ;
  assign n23880 = ~n2764 & n23879 ;
  assign n23881 = n23880 ^ n7872 ^ n4278 ;
  assign n23886 = n23885 ^ n23881 ^ n14807 ;
  assign n23887 = ( n2845 & ~n6554 ) | ( n2845 & n23886 ) | ( ~n6554 & n23886 ) ;
  assign n23889 = n5718 ^ n5117 ^ 1'b0 ;
  assign n23890 = x176 & n23889 ;
  assign n23891 = ( ~n3303 & n12788 ) | ( ~n3303 & n23890 ) | ( n12788 & n23890 ) ;
  assign n23888 = n4034 | n21037 ;
  assign n23892 = n23891 ^ n23888 ^ 1'b0 ;
  assign n23894 = ~n4503 & n17727 ;
  assign n23895 = n23894 ^ n9924 ^ 1'b0 ;
  assign n23893 = n13635 ^ n9248 ^ n1226 ;
  assign n23896 = n23895 ^ n23893 ^ n3726 ;
  assign n23897 = n15780 ^ n12941 ^ n6171 ;
  assign n23898 = n9422 ^ n8798 ^ 1'b0 ;
  assign n23899 = ~n20559 & n23898 ;
  assign n23900 = ( n1212 & ~n5558 ) | ( n1212 & n18001 ) | ( ~n5558 & n18001 ) ;
  assign n23908 = n6483 ^ n3444 ^ 1'b0 ;
  assign n23909 = n23908 ^ n6767 ^ 1'b0 ;
  assign n23910 = n17162 | n23909 ;
  assign n23911 = n23910 ^ n12438 ^ n3259 ;
  assign n23906 = ( n1483 & ~n2966 ) | ( n1483 & n10417 ) | ( ~n2966 & n10417 ) ;
  assign n23907 = ( n8282 & n11059 ) | ( n8282 & n23906 ) | ( n11059 & n23906 ) ;
  assign n23901 = ~n10954 & n13233 ;
  assign n23902 = n2229 & n4238 ;
  assign n23903 = n23902 ^ n2571 ^ 1'b0 ;
  assign n23904 = n23903 ^ x225 ^ 1'b0 ;
  assign n23905 = n23901 | n23904 ;
  assign n23912 = n23911 ^ n23907 ^ n23905 ;
  assign n23913 = n17821 ^ n11388 ^ n1598 ;
  assign n23914 = n21280 ^ n20998 ^ n13301 ;
  assign n23915 = n493 & n14793 ;
  assign n23916 = n22415 ^ n16755 ^ n6953 ;
  assign n23917 = n16573 ^ n7505 ^ n2446 ;
  assign n23923 = n9564 & ~n11487 ;
  assign n23924 = ( ~n1909 & n5264 ) | ( ~n1909 & n23923 ) | ( n5264 & n23923 ) ;
  assign n23921 = ( ~n1715 & n2271 ) | ( ~n1715 & n3754 ) | ( n2271 & n3754 ) ;
  assign n23919 = ( ~n318 & n11142 ) | ( ~n318 & n20002 ) | ( n11142 & n20002 ) ;
  assign n23918 = n12861 ^ n9737 ^ x123 ;
  assign n23920 = n23919 ^ n23918 ^ n2262 ;
  assign n23922 = n23921 ^ n23920 ^ x0 ;
  assign n23925 = n23924 ^ n23922 ^ n18291 ;
  assign n23927 = ( n4463 & ~n4992 ) | ( n4463 & n10696 ) | ( ~n4992 & n10696 ) ;
  assign n23928 = n7654 | n23927 ;
  assign n23929 = ( n1497 & ~n1664 ) | ( n1497 & n23928 ) | ( ~n1664 & n23928 ) ;
  assign n23926 = n12419 ^ n4248 ^ 1'b0 ;
  assign n23930 = n23929 ^ n23926 ^ n19020 ;
  assign n23931 = n3293 ^ n2165 ^ n812 ;
  assign n23932 = n21583 | n23931 ;
  assign n23934 = n13629 ^ n12015 ^ n5033 ;
  assign n23935 = ( n11304 & n17814 ) | ( n11304 & n23934 ) | ( n17814 & n23934 ) ;
  assign n23933 = ( n4742 & n14595 ) | ( n4742 & ~n23478 ) | ( n14595 & ~n23478 ) ;
  assign n23936 = n23935 ^ n23933 ^ n20081 ;
  assign n23937 = ( n12249 & ~n20491 ) | ( n12249 & n23936 ) | ( ~n20491 & n23936 ) ;
  assign n23938 = n9097 ^ x74 ^ 1'b0 ;
  assign n23939 = n18910 & n23938 ;
  assign n23940 = ( n3786 & n5795 ) | ( n3786 & ~n7478 ) | ( n5795 & ~n7478 ) ;
  assign n23941 = ( n2365 & n23939 ) | ( n2365 & n23940 ) | ( n23939 & n23940 ) ;
  assign n23942 = n22278 ^ n16753 ^ 1'b0 ;
  assign n23943 = n20207 | n23942 ;
  assign n23944 = n23943 ^ n22160 ^ n3227 ;
  assign n23946 = n7353 ^ n3350 ^ n2721 ;
  assign n23945 = n2564 & n17751 ;
  assign n23947 = n23946 ^ n23945 ^ n22974 ;
  assign n23950 = n17943 ^ n1528 ^ n742 ;
  assign n23951 = ( ~n4556 & n14455 ) | ( ~n4556 & n23950 ) | ( n14455 & n23950 ) ;
  assign n23948 = n16800 ^ n12588 ^ 1'b0 ;
  assign n23949 = ( n10271 & ~n11135 ) | ( n10271 & n23948 ) | ( ~n11135 & n23948 ) ;
  assign n23952 = n23951 ^ n23949 ^ n9866 ;
  assign n23953 = n15286 ^ n12635 ^ 1'b0 ;
  assign n23954 = n11516 ^ n11370 ^ 1'b0 ;
  assign n23955 = n6885 & ~n23954 ;
  assign n23956 = ( n11002 & n12845 ) | ( n11002 & n23955 ) | ( n12845 & n23955 ) ;
  assign n23957 = n10333 & n23956 ;
  assign n23958 = ~n23953 & n23957 ;
  assign n23959 = ( n16302 & n23714 ) | ( n16302 & n23958 ) | ( n23714 & n23958 ) ;
  assign n23960 = n11040 ^ n10735 ^ n4063 ;
  assign n23964 = n10657 ^ n6609 ^ n4724 ;
  assign n23961 = n19412 ^ n12678 ^ 1'b0 ;
  assign n23962 = n5287 | n23961 ;
  assign n23963 = n14419 & ~n23962 ;
  assign n23965 = n23964 ^ n23963 ^ 1'b0 ;
  assign n23966 = n13670 ^ n9315 ^ n1282 ;
  assign n23967 = n11414 ^ n8839 ^ n2776 ;
  assign n23968 = n15023 ^ n3210 ^ 1'b0 ;
  assign n23969 = n23967 & n23968 ;
  assign n23970 = n23969 ^ n14497 ^ n9935 ;
  assign n23971 = n2814 | n7112 ;
  assign n23972 = ( ~n2113 & n2959 ) | ( ~n2113 & n13603 ) | ( n2959 & n13603 ) ;
  assign n23973 = n23972 ^ n14464 ^ n3266 ;
  assign n23974 = n23973 ^ n9627 ^ n1221 ;
  assign n23975 = n23974 ^ n17855 ^ 1'b0 ;
  assign n23976 = n14621 | n23975 ;
  assign n23980 = n5032 & n12620 ;
  assign n23981 = n23980 ^ n1864 ^ 1'b0 ;
  assign n23982 = n23981 ^ n11246 ^ 1'b0 ;
  assign n23977 = ~n316 & n8336 ;
  assign n23978 = n4546 & n23977 ;
  assign n23979 = n23978 ^ n12511 ^ n9866 ;
  assign n23983 = n23982 ^ n23979 ^ n1412 ;
  assign n23984 = n5231 ^ x205 ^ 1'b0 ;
  assign n23985 = ( x31 & n6549 ) | ( x31 & ~n18928 ) | ( n6549 & ~n18928 ) ;
  assign n23988 = ( n12785 & ~n16707 ) | ( n12785 & n21225 ) | ( ~n16707 & n21225 ) ;
  assign n23987 = n5737 ^ n2012 ^ n720 ;
  assign n23986 = ~n9273 & n16866 ;
  assign n23989 = n23988 ^ n23987 ^ n23986 ;
  assign n23997 = ( n9906 & n12604 ) | ( n9906 & n18374 ) | ( n12604 & n18374 ) ;
  assign n23998 = ( n2129 & n2302 ) | ( n2129 & n3770 ) | ( n2302 & n3770 ) ;
  assign n23999 = n17077 ^ n14918 ^ 1'b0 ;
  assign n24000 = n23998 | n23999 ;
  assign n24001 = ( n842 & n13660 ) | ( n842 & ~n24000 ) | ( n13660 & ~n24000 ) ;
  assign n24002 = ( n9472 & n23997 ) | ( n9472 & ~n24001 ) | ( n23997 & ~n24001 ) ;
  assign n23994 = n7260 ^ n6059 ^ n1616 ;
  assign n23995 = ( n6122 & n12139 ) | ( n6122 & n23994 ) | ( n12139 & n23994 ) ;
  assign n23993 = n21471 ^ n8762 ^ n3625 ;
  assign n23996 = n23995 ^ n23993 ^ n6245 ;
  assign n23990 = n4295 & n7903 ;
  assign n23991 = ~n2744 & n23990 ;
  assign n23992 = ( ~n2459 & n18109 ) | ( ~n2459 & n23991 ) | ( n18109 & n23991 ) ;
  assign n24003 = n24002 ^ n23996 ^ n23992 ;
  assign n24004 = n23503 ^ n21120 ^ n5650 ;
  assign n24005 = ( n8356 & n13191 ) | ( n8356 & n24004 ) | ( n13191 & n24004 ) ;
  assign n24006 = ( n4821 & ~n6437 ) | ( n4821 & n7658 ) | ( ~n6437 & n7658 ) ;
  assign n24007 = n1520 & n24006 ;
  assign n24012 = n4771 | n4992 ;
  assign n24013 = n24012 ^ n20405 ^ 1'b0 ;
  assign n24011 = ( ~n9312 & n9929 ) | ( ~n9312 & n23275 ) | ( n9929 & n23275 ) ;
  assign n24014 = n24013 ^ n24011 ^ n1935 ;
  assign n24008 = ( n2339 & n14524 ) | ( n2339 & ~n17236 ) | ( n14524 & ~n17236 ) ;
  assign n24009 = n24008 ^ n9257 ^ 1'b0 ;
  assign n24010 = n8864 & ~n24009 ;
  assign n24015 = n24014 ^ n24010 ^ 1'b0 ;
  assign n24019 = n12472 ^ x141 ^ 1'b0 ;
  assign n24020 = n12295 | n24019 ;
  assign n24021 = ( n5743 & n23203 ) | ( n5743 & n24020 ) | ( n23203 & n24020 ) ;
  assign n24016 = n10905 ^ n4238 ^ n3875 ;
  assign n24017 = n10645 & n24016 ;
  assign n24018 = ~n14545 & n24017 ;
  assign n24022 = n24021 ^ n24018 ^ n4841 ;
  assign n24023 = n12077 ^ n8255 ^ n5497 ;
  assign n24024 = ( n2395 & n2970 ) | ( n2395 & n5161 ) | ( n2970 & n5161 ) ;
  assign n24025 = ( n23370 & n24023 ) | ( n23370 & ~n24024 ) | ( n24023 & ~n24024 ) ;
  assign n24027 = ( n436 & n1256 ) | ( n436 & ~n3446 ) | ( n1256 & ~n3446 ) ;
  assign n24028 = ( n5237 & n6671 ) | ( n5237 & n24027 ) | ( n6671 & n24027 ) ;
  assign n24029 = n19325 ^ n8750 ^ n8485 ;
  assign n24030 = ( n3131 & n3359 ) | ( n3131 & n4188 ) | ( n3359 & n4188 ) ;
  assign n24031 = n24030 ^ n14530 ^ n4513 ;
  assign n24032 = ( n14081 & ~n24029 ) | ( n14081 & n24031 ) | ( ~n24029 & n24031 ) ;
  assign n24033 = n24032 ^ n21698 ^ n5641 ;
  assign n24034 = n24028 & n24033 ;
  assign n24026 = n17260 ^ n4901 ^ n3443 ;
  assign n24035 = n24034 ^ n24026 ^ n1218 ;
  assign n24036 = ( n2185 & n5769 ) | ( n2185 & ~n10607 ) | ( n5769 & ~n10607 ) ;
  assign n24037 = n24036 ^ n16264 ^ n8463 ;
  assign n24038 = ( n11352 & ~n12149 ) | ( n11352 & n24037 ) | ( ~n12149 & n24037 ) ;
  assign n24039 = x219 | n13699 ;
  assign n24040 = ( n4368 & n24038 ) | ( n4368 & n24039 ) | ( n24038 & n24039 ) ;
  assign n24041 = ( n3726 & n10517 ) | ( n3726 & n24040 ) | ( n10517 & n24040 ) ;
  assign n24042 = ( n15422 & n20530 ) | ( n15422 & ~n21995 ) | ( n20530 & ~n21995 ) ;
  assign n24043 = n6979 & n22120 ;
  assign n24044 = n24043 ^ n22866 ^ n12839 ;
  assign n24045 = n19409 ^ n18931 ^ n1092 ;
  assign n24047 = n8677 & ~n11579 ;
  assign n24048 = n24047 ^ n1978 ^ 1'b0 ;
  assign n24049 = n24048 ^ n22879 ^ n18905 ;
  assign n24046 = n2255 | n5479 ;
  assign n24050 = n24049 ^ n24046 ^ n20726 ;
  assign n24051 = n22977 ^ n20197 ^ n18110 ;
  assign n24052 = n14818 ^ n2509 ^ 1'b0 ;
  assign n24053 = n17543 & n24052 ;
  assign n24059 = n303 & ~n6875 ;
  assign n24060 = n24059 ^ n16109 ^ 1'b0 ;
  assign n24054 = n7408 ^ n6997 ^ n4824 ;
  assign n24055 = n14066 ^ n10504 ^ n6904 ;
  assign n24056 = n13772 & ~n24055 ;
  assign n24057 = ( n23841 & n24054 ) | ( n23841 & n24056 ) | ( n24054 & n24056 ) ;
  assign n24058 = n24057 ^ n8769 ^ 1'b0 ;
  assign n24061 = n24060 ^ n24058 ^ n11053 ;
  assign n24062 = n24053 | n24061 ;
  assign n24064 = n7695 & ~n22273 ;
  assign n24065 = n24064 ^ n19046 ^ 1'b0 ;
  assign n24063 = n4506 & ~n20132 ;
  assign n24066 = n24065 ^ n24063 ^ n15269 ;
  assign n24067 = ( n9359 & n24062 ) | ( n9359 & n24066 ) | ( n24062 & n24066 ) ;
  assign n24068 = n23157 ^ n8867 ^ 1'b0 ;
  assign n24069 = n24068 ^ n19155 ^ n16285 ;
  assign n24070 = n24069 ^ n20871 ^ n10041 ;
  assign n24071 = n21406 ^ n12834 ^ 1'b0 ;
  assign n24072 = n2848 | n24071 ;
  assign n24073 = ( n1669 & n5952 ) | ( n1669 & ~n15964 ) | ( n5952 & ~n15964 ) ;
  assign n24080 = n11164 ^ n2574 ^ n464 ;
  assign n24076 = ( ~n3203 & n9813 ) | ( ~n3203 & n14383 ) | ( n9813 & n14383 ) ;
  assign n24077 = n7629 ^ n6984 ^ n5008 ;
  assign n24078 = ( ~n7483 & n24076 ) | ( ~n7483 & n24077 ) | ( n24076 & n24077 ) ;
  assign n24074 = n14393 ^ n5319 ^ n2404 ;
  assign n24075 = ( ~n3568 & n10554 ) | ( ~n3568 & n24074 ) | ( n10554 & n24074 ) ;
  assign n24079 = n24078 ^ n24075 ^ n8627 ;
  assign n24081 = n24080 ^ n24079 ^ n4612 ;
  assign n24082 = ( n6260 & n9203 ) | ( n6260 & ~n10207 ) | ( n9203 & ~n10207 ) ;
  assign n24083 = n8497 ^ n6616 ^ 1'b0 ;
  assign n24084 = n24082 & n24083 ;
  assign n24085 = ( n1373 & n6749 ) | ( n1373 & ~n9185 ) | ( n6749 & ~n9185 ) ;
  assign n24086 = n7870 & ~n10842 ;
  assign n24087 = n24086 ^ n6372 ^ 1'b0 ;
  assign n24088 = n24087 ^ n4907 ^ n3462 ;
  assign n24089 = n24088 ^ n16623 ^ n8757 ;
  assign n24090 = n24089 ^ n1582 ^ 1'b0 ;
  assign n24091 = n24085 & n24090 ;
  assign n24092 = ( ~n7438 & n24084 ) | ( ~n7438 & n24091 ) | ( n24084 & n24091 ) ;
  assign n24093 = n11084 ^ n5511 ^ n2020 ;
  assign n24096 = n8193 ^ n7490 ^ n7444 ;
  assign n24094 = ( ~n472 & n4093 ) | ( ~n472 & n4684 ) | ( n4093 & n4684 ) ;
  assign n24095 = ( n12757 & ~n17426 ) | ( n12757 & n24094 ) | ( ~n17426 & n24094 ) ;
  assign n24097 = n24096 ^ n24095 ^ n18044 ;
  assign n24098 = ( n2431 & n2916 ) | ( n2431 & ~n17594 ) | ( n2916 & ~n17594 ) ;
  assign n24099 = n24098 ^ n9991 ^ n7331 ;
  assign n24103 = n17213 ^ n4752 ^ n1851 ;
  assign n24100 = ( ~n5638 & n8976 ) | ( ~n5638 & n16044 ) | ( n8976 & n16044 ) ;
  assign n24101 = ( n1002 & n11914 ) | ( n1002 & ~n20431 ) | ( n11914 & ~n20431 ) ;
  assign n24102 = n24100 & n24101 ;
  assign n24104 = n24103 ^ n24102 ^ n3840 ;
  assign n24105 = n21921 ^ n21904 ^ n7304 ;
  assign n24106 = n24105 ^ n13647 ^ n1749 ;
  assign n24112 = ( ~n8064 & n11221 ) | ( ~n8064 & n23227 ) | ( n11221 & n23227 ) ;
  assign n24113 = n302 & ~n5742 ;
  assign n24114 = ~n10268 & n24113 ;
  assign n24115 = n24114 ^ n15168 ^ n13692 ;
  assign n24116 = n7632 & ~n24115 ;
  assign n24117 = ( n8687 & ~n24112 ) | ( n8687 & n24116 ) | ( ~n24112 & n24116 ) ;
  assign n24108 = n9609 ^ n6744 ^ n6563 ;
  assign n24109 = ( ~n9193 & n11144 ) | ( ~n9193 & n24108 ) | ( n11144 & n24108 ) ;
  assign n24107 = n5786 & ~n6888 ;
  assign n24110 = n24109 ^ n24107 ^ 1'b0 ;
  assign n24111 = n24110 ^ n12836 ^ n2592 ;
  assign n24118 = n24117 ^ n24111 ^ n1126 ;
  assign n24119 = ( ~n571 & n23214 ) | ( ~n571 & n24118 ) | ( n23214 & n24118 ) ;
  assign n24120 = ( ~n7478 & n15347 ) | ( ~n7478 & n19993 ) | ( n15347 & n19993 ) ;
  assign n24121 = n24120 ^ n2054 ^ n1495 ;
  assign n24122 = ( n1840 & ~n2454 ) | ( n1840 & n3561 ) | ( ~n2454 & n3561 ) ;
  assign n24123 = n24122 ^ n2880 ^ n2177 ;
  assign n24124 = n11231 ^ n3932 ^ n3083 ;
  assign n24125 = n18023 ^ n4650 ^ n2412 ;
  assign n24126 = n2397 & ~n24125 ;
  assign n24127 = n24126 ^ n8206 ^ 1'b0 ;
  assign n24128 = n24127 ^ n5888 ^ n3672 ;
  assign n24129 = ( n4458 & n23491 ) | ( n4458 & ~n24128 ) | ( n23491 & ~n24128 ) ;
  assign n24130 = ( n18853 & n24124 ) | ( n18853 & ~n24129 ) | ( n24124 & ~n24129 ) ;
  assign n24131 = n4430 & ~n16556 ;
  assign n24132 = ~n24130 & n24131 ;
  assign n24133 = n10633 & n13992 ;
  assign n24134 = n2302 | n11867 ;
  assign n24135 = ( n14590 & n19566 ) | ( n14590 & ~n23222 ) | ( n19566 & ~n23222 ) ;
  assign n24140 = n12785 ^ n11100 ^ n1504 ;
  assign n24141 = ( ~n4047 & n14814 ) | ( ~n4047 & n24140 ) | ( n14814 & n24140 ) ;
  assign n24142 = n24141 ^ n12081 ^ n11796 ;
  assign n24143 = n15552 & n24142 ;
  assign n24144 = n7355 & n24143 ;
  assign n24136 = n16145 ^ n8725 ^ 1'b0 ;
  assign n24137 = n20580 ^ n16189 ^ n10465 ;
  assign n24138 = n24137 ^ n14272 ^ 1'b0 ;
  assign n24139 = n24136 | n24138 ;
  assign n24145 = n24144 ^ n24139 ^ n21142 ;
  assign n24150 = ~n5899 & n7983 ;
  assign n24146 = n16615 ^ x241 ^ 1'b0 ;
  assign n24147 = n7837 ^ n5247 ^ n3989 ;
  assign n24148 = ( ~n1381 & n24146 ) | ( ~n1381 & n24147 ) | ( n24146 & n24147 ) ;
  assign n24149 = n8101 & ~n24148 ;
  assign n24151 = n24150 ^ n24149 ^ 1'b0 ;
  assign n24152 = n10328 ^ n7226 ^ n4223 ;
  assign n24153 = ( n5319 & ~n22009 ) | ( n5319 & n24152 ) | ( ~n22009 & n24152 ) ;
  assign n24154 = n7671 & ~n9262 ;
  assign n24155 = n15312 ^ n2220 ^ 1'b0 ;
  assign n24156 = ~n23553 & n24155 ;
  assign n24157 = n12929 ^ n8985 ^ n1189 ;
  assign n24158 = n24157 ^ n21327 ^ n6224 ;
  assign n24159 = ( n1674 & n3724 ) | ( n1674 & ~n18392 ) | ( n3724 & ~n18392 ) ;
  assign n24160 = ~n1384 & n24159 ;
  assign n24161 = n16297 & n24160 ;
  assign n24162 = ( ~n3257 & n3913 ) | ( ~n3257 & n19541 ) | ( n3913 & n19541 ) ;
  assign n24163 = ( n850 & n2232 ) | ( n850 & ~n4762 ) | ( n2232 & ~n4762 ) ;
  assign n24164 = n24163 ^ n12670 ^ n8660 ;
  assign n24165 = n24164 ^ n13524 ^ n11760 ;
  assign n24166 = ( n22630 & ~n24162 ) | ( n22630 & n24165 ) | ( ~n24162 & n24165 ) ;
  assign n24174 = n16007 ^ n12520 ^ 1'b0 ;
  assign n24175 = n16280 | n24174 ;
  assign n24170 = n11219 ^ n9048 ^ 1'b0 ;
  assign n24171 = n6676 | n24170 ;
  assign n24172 = ( ~n772 & n8293 ) | ( ~n772 & n18580 ) | ( n8293 & n18580 ) ;
  assign n24173 = ( n17059 & ~n24171 ) | ( n17059 & n24172 ) | ( ~n24171 & n24172 ) ;
  assign n24167 = ( x97 & n8537 ) | ( x97 & n8728 ) | ( n8537 & n8728 ) ;
  assign n24168 = n24167 ^ n9173 ^ 1'b0 ;
  assign n24169 = ~n16646 & n24168 ;
  assign n24176 = n24175 ^ n24173 ^ n24169 ;
  assign n24184 = n2585 & n9268 ;
  assign n24185 = n24184 ^ n2454 ^ 1'b0 ;
  assign n24186 = n24185 ^ n10439 ^ n6703 ;
  assign n24187 = n24186 ^ n16890 ^ n9838 ;
  assign n24179 = ~n1048 & n7075 ;
  assign n24178 = ~n2407 & n22083 ;
  assign n24180 = n24179 ^ n24178 ^ 1'b0 ;
  assign n24177 = n21713 ^ n2369 ^ n1352 ;
  assign n24181 = n24180 ^ n24177 ^ n4476 ;
  assign n24182 = n14008 ^ n4045 ^ 1'b0 ;
  assign n24183 = n24181 & ~n24182 ;
  assign n24188 = n24187 ^ n24183 ^ n22654 ;
  assign n24189 = ( n4571 & n9129 ) | ( n4571 & n9270 ) | ( n9129 & n9270 ) ;
  assign n24190 = n24189 ^ n5935 ^ n1749 ;
  assign n24195 = n16513 ^ n10094 ^ 1'b0 ;
  assign n24191 = n1478 | n17738 ;
  assign n24192 = n24191 ^ n5784 ^ 1'b0 ;
  assign n24193 = n21606 | n24192 ;
  assign n24194 = n24193 ^ n3487 ^ 1'b0 ;
  assign n24196 = n24195 ^ n24194 ^ n8227 ;
  assign n24197 = n18752 ^ n16717 ^ n15775 ;
  assign n24198 = ( n5852 & n9425 ) | ( n5852 & n24197 ) | ( n9425 & n24197 ) ;
  assign n24199 = n15243 | n24198 ;
  assign n24200 = ~n19429 & n24199 ;
  assign n24205 = n18208 ^ n464 ^ 1'b0 ;
  assign n24206 = n24205 ^ n8087 ^ n4516 ;
  assign n24201 = n7253 ^ n2143 ^ 1'b0 ;
  assign n24202 = ( n8346 & n12752 ) | ( n8346 & ~n15434 ) | ( n12752 & ~n15434 ) ;
  assign n24203 = n24201 & ~n24202 ;
  assign n24204 = n19413 | n24203 ;
  assign n24207 = n24206 ^ n24204 ^ 1'b0 ;
  assign n24208 = n8030 & ~n9613 ;
  assign n24209 = n24208 ^ n10341 ^ 1'b0 ;
  assign n24210 = n6940 & ~n24209 ;
  assign n24211 = n10188 & n24210 ;
  assign n24212 = n24211 ^ n11794 ^ n10187 ;
  assign n24213 = ( n6175 & ~n24207 ) | ( n6175 & n24212 ) | ( ~n24207 & n24212 ) ;
  assign n24215 = n7976 & ~n14945 ;
  assign n24214 = n18942 ^ n3221 ^ x176 ;
  assign n24216 = n24215 ^ n24214 ^ n22166 ;
  assign n24217 = ( n6128 & n7941 ) | ( n6128 & ~n14145 ) | ( n7941 & ~n14145 ) ;
  assign n24218 = n15706 | n24217 ;
  assign n24219 = n24218 ^ n1562 ^ 1'b0 ;
  assign n24220 = n24219 ^ n16789 ^ x83 ;
  assign n24221 = n24220 ^ n416 ^ 1'b0 ;
  assign n24222 = ~n7568 & n24221 ;
  assign n24223 = n24125 ^ n12274 ^ n3638 ;
  assign n24224 = ( n2442 & n4208 ) | ( n2442 & n5891 ) | ( n4208 & n5891 ) ;
  assign n24225 = ~n24223 & n24224 ;
  assign n24226 = n14185 & n24225 ;
  assign n24230 = n15989 ^ n14057 ^ n897 ;
  assign n24227 = n13314 ^ n10174 ^ n9915 ;
  assign n24228 = n24227 ^ n14278 ^ n8766 ;
  assign n24229 = n24228 ^ n6542 ^ n5000 ;
  assign n24231 = n24230 ^ n24229 ^ n21806 ;
  assign n24232 = n24231 ^ n23505 ^ n9727 ;
  assign n24233 = n19477 ^ n4035 ^ 1'b0 ;
  assign n24234 = n24233 ^ n8519 ^ 1'b0 ;
  assign n24235 = n24234 ^ n18835 ^ n5359 ;
  assign n24243 = n13493 ^ n8301 ^ n7942 ;
  assign n24242 = n9662 ^ n2416 ^ 1'b0 ;
  assign n24240 = ( n12511 & n14064 ) | ( n12511 & ~n14680 ) | ( n14064 & ~n14680 ) ;
  assign n24236 = ~n617 & n14530 ;
  assign n24237 = n1932 & n24236 ;
  assign n24238 = n6923 & ~n24237 ;
  assign n24239 = n24238 ^ n6087 ^ 1'b0 ;
  assign n24241 = n24240 ^ n24239 ^ n19207 ;
  assign n24244 = n24243 ^ n24242 ^ n24241 ;
  assign n24245 = n24244 ^ n23778 ^ n8647 ;
  assign n24246 = n12908 | n21853 ;
  assign n24247 = n5053 | n24246 ;
  assign n24248 = n20907 ^ n16594 ^ n12824 ;
  assign n24249 = n3759 & ~n22124 ;
  assign n24250 = ~n24248 & n24249 ;
  assign n24251 = n23279 ^ n14298 ^ n6001 ;
  assign n24252 = n5396 | n19628 ;
  assign n24253 = ( n12604 & ~n20918 ) | ( n12604 & n24252 ) | ( ~n20918 & n24252 ) ;
  assign n24254 = n8729 ^ n3281 ^ 1'b0 ;
  assign n24255 = n4920 & n24254 ;
  assign n24256 = ( n2242 & n9422 ) | ( n2242 & n24255 ) | ( n9422 & n24255 ) ;
  assign n24257 = n3123 & ~n24256 ;
  assign n24258 = ( n1781 & n1806 ) | ( n1781 & n4089 ) | ( n1806 & n4089 ) ;
  assign n24259 = ( ~n17851 & n23190 ) | ( ~n17851 & n24258 ) | ( n23190 & n24258 ) ;
  assign n24260 = ( x166 & n23650 ) | ( x166 & n24259 ) | ( n23650 & n24259 ) ;
  assign n24261 = ( ~n8506 & n13147 ) | ( ~n8506 & n15206 ) | ( n13147 & n15206 ) ;
  assign n24262 = n21496 ^ n5233 ^ 1'b0 ;
  assign n24263 = n24261 & ~n24262 ;
  assign n24267 = ~n1535 & n11396 ;
  assign n24268 = n4121 & n24267 ;
  assign n24265 = ~n2747 & n15198 ;
  assign n24266 = n24265 ^ n12078 ^ 1'b0 ;
  assign n24269 = n24268 ^ n24266 ^ n23115 ;
  assign n24264 = ~n6514 & n18625 ;
  assign n24270 = n24269 ^ n24264 ^ 1'b0 ;
  assign n24271 = n24270 ^ n7216 ^ 1'b0 ;
  assign n24272 = n24271 ^ n14220 ^ 1'b0 ;
  assign n24273 = n21795 & ~n24272 ;
  assign n24274 = n22471 ^ n15085 ^ n5261 ;
  assign n24275 = ( x227 & n16367 ) | ( x227 & n24274 ) | ( n16367 & n24274 ) ;
  assign n24276 = ( n2027 & n5277 ) | ( n2027 & n18738 ) | ( n5277 & n18738 ) ;
  assign n24277 = ( n2763 & ~n21420 ) | ( n2763 & n24276 ) | ( ~n21420 & n24276 ) ;
  assign n24278 = ( n601 & n4401 ) | ( n601 & n5766 ) | ( n4401 & n5766 ) ;
  assign n24279 = ~n22191 & n24278 ;
  assign n24280 = n24279 ^ n9634 ^ 1'b0 ;
  assign n24281 = x112 & n24280 ;
  assign n24282 = ( n1549 & ~n2014 ) | ( n1549 & n16565 ) | ( ~n2014 & n16565 ) ;
  assign n24283 = n24282 ^ n23870 ^ n13861 ;
  assign n24284 = n16774 ^ n8753 ^ n7806 ;
  assign n24285 = n12492 ^ n10383 ^ 1'b0 ;
  assign n24286 = ( n6621 & n24284 ) | ( n6621 & ~n24285 ) | ( n24284 & ~n24285 ) ;
  assign n24287 = ( ~n1825 & n7953 ) | ( ~n1825 & n9606 ) | ( n7953 & n9606 ) ;
  assign n24288 = ( n6514 & n7448 ) | ( n6514 & ~n8958 ) | ( n7448 & ~n8958 ) ;
  assign n24289 = n24288 ^ n4398 ^ n1510 ;
  assign n24290 = ( n5510 & n24287 ) | ( n5510 & n24289 ) | ( n24287 & n24289 ) ;
  assign n24291 = ( n5512 & n10443 ) | ( n5512 & ~n10639 ) | ( n10443 & ~n10639 ) ;
  assign n24292 = ( n3471 & n17666 ) | ( n3471 & n24291 ) | ( n17666 & n24291 ) ;
  assign n24293 = n2750 & ~n7582 ;
  assign n24294 = ~n14967 & n24293 ;
  assign n24295 = n12467 | n24294 ;
  assign n24296 = n24295 ^ n9874 ^ 1'b0 ;
  assign n24297 = ( ~n12470 & n12861 ) | ( ~n12470 & n24296 ) | ( n12861 & n24296 ) ;
  assign n24298 = ( n4899 & ~n13960 ) | ( n4899 & n19431 ) | ( ~n13960 & n19431 ) ;
  assign n24299 = ( n7810 & n10085 ) | ( n7810 & ~n12612 ) | ( n10085 & ~n12612 ) ;
  assign n24300 = n24299 ^ n16373 ^ n6930 ;
  assign n24301 = n24300 ^ n21996 ^ 1'b0 ;
  assign n24302 = ( ~n3454 & n11166 ) | ( ~n3454 & n16347 ) | ( n11166 & n16347 ) ;
  assign n24303 = n8676 ^ n7815 ^ n5100 ;
  assign n24304 = ~n5138 & n24303 ;
  assign n24305 = ~n24302 & n24304 ;
  assign n24306 = ( n11940 & ~n12892 ) | ( n11940 & n19840 ) | ( ~n12892 & n19840 ) ;
  assign n24307 = n23110 ^ n3880 ^ 1'b0 ;
  assign n24308 = n14330 & n15520 ;
  assign n24309 = ~n4103 & n24308 ;
  assign n24310 = n20037 ^ n18119 ^ 1'b0 ;
  assign n24311 = ( n17166 & n19201 ) | ( n17166 & n24310 ) | ( n19201 & n24310 ) ;
  assign n24312 = n20318 ^ n12432 ^ 1'b0 ;
  assign n24313 = ( n595 & n4671 ) | ( n595 & ~n9584 ) | ( n4671 & ~n9584 ) ;
  assign n24314 = n6627 | n24313 ;
  assign n24315 = n19584 ^ n13639 ^ n11711 ;
  assign n24317 = ( n2704 & ~n13348 ) | ( n2704 & n18930 ) | ( ~n13348 & n18930 ) ;
  assign n24316 = n21106 ^ n18693 ^ n11674 ;
  assign n24318 = n24317 ^ n24316 ^ 1'b0 ;
  assign n24319 = ~n24192 & n24318 ;
  assign n24320 = ( ~n16774 & n24315 ) | ( ~n16774 & n24319 ) | ( n24315 & n24319 ) ;
  assign n24321 = ( x3 & n1662 ) | ( x3 & ~n9147 ) | ( n1662 & ~n9147 ) ;
  assign n24322 = ( ~n6562 & n9025 ) | ( ~n6562 & n24321 ) | ( n9025 & n24321 ) ;
  assign n24323 = n24322 ^ n10492 ^ n6272 ;
  assign n24325 = ( x16 & n15145 ) | ( x16 & n17901 ) | ( n15145 & n17901 ) ;
  assign n24324 = ( n5776 & n11358 ) | ( n5776 & n17753 ) | ( n11358 & n17753 ) ;
  assign n24326 = n24325 ^ n24324 ^ x46 ;
  assign n24327 = ( n7334 & n11551 ) | ( n7334 & ~n24326 ) | ( n11551 & ~n24326 ) ;
  assign n24328 = ~n4609 & n6585 ;
  assign n24329 = n24328 ^ n2829 ^ 1'b0 ;
  assign n24330 = n8171 ^ n6177 ^ n327 ;
  assign n24331 = ( ~n23549 & n24329 ) | ( ~n23549 & n24330 ) | ( n24329 & n24330 ) ;
  assign n24332 = n11218 ^ n8342 ^ n4760 ;
  assign n24333 = ~n5867 & n14130 ;
  assign n24334 = n24332 & n24333 ;
  assign n24335 = ~n8423 & n10234 ;
  assign n24336 = n24335 ^ n13042 ^ n1830 ;
  assign n24340 = n7876 & ~n21951 ;
  assign n24337 = n7742 & ~n10806 ;
  assign n24338 = n20919 ^ n6287 ^ n4829 ;
  assign n24339 = ( n6645 & n24337 ) | ( n6645 & ~n24338 ) | ( n24337 & ~n24338 ) ;
  assign n24341 = n24340 ^ n24339 ^ x25 ;
  assign n24342 = ( ~n3123 & n11612 ) | ( ~n3123 & n13269 ) | ( n11612 & n13269 ) ;
  assign n24343 = n7189 ^ n4048 ^ 1'b0 ;
  assign n24344 = n24343 ^ n18104 ^ 1'b0 ;
  assign n24345 = n24344 ^ n14621 ^ n5907 ;
  assign n24346 = ( ~n453 & n24342 ) | ( ~n453 & n24345 ) | ( n24342 & n24345 ) ;
  assign n24347 = n18812 & n24346 ;
  assign n24348 = n4622 & n15915 ;
  assign n24349 = ~n464 & n24348 ;
  assign n24351 = ( n1188 & n1802 ) | ( n1188 & ~n6631 ) | ( n1802 & ~n6631 ) ;
  assign n24352 = n24351 ^ n12232 ^ n4705 ;
  assign n24350 = n9697 ^ n6197 ^ n5889 ;
  assign n24353 = n24352 ^ n24350 ^ n2091 ;
  assign n24354 = n24349 | n24353 ;
  assign n24355 = ( ~n4485 & n7503 ) | ( ~n4485 & n8938 ) | ( n7503 & n8938 ) ;
  assign n24356 = n23378 & n24355 ;
  assign n24357 = ~n8070 & n17819 ;
  assign n24358 = n24357 ^ n5145 ^ 1'b0 ;
  assign n24359 = n2836 ^ n2568 ^ n1296 ;
  assign n24360 = n5634 | n24359 ;
  assign n24361 = ( ~n5251 & n24358 ) | ( ~n5251 & n24360 ) | ( n24358 & n24360 ) ;
  assign n24362 = n8018 & ~n24361 ;
  assign n24363 = n24362 ^ n3752 ^ 1'b0 ;
  assign n24364 = n24363 ^ n10274 ^ n4662 ;
  assign n24365 = ( n8139 & n13039 ) | ( n8139 & ~n24364 ) | ( n13039 & ~n24364 ) ;
  assign n24366 = n24365 ^ n9691 ^ n8904 ;
  assign n24367 = n21585 ^ n12286 ^ n6628 ;
  assign n24368 = n24367 ^ n21334 ^ n6972 ;
  assign n24369 = n3580 ^ n742 ^ 1'b0 ;
  assign n24370 = n14785 & ~n24369 ;
  assign n24371 = n2362 & ~n5676 ;
  assign n24372 = n24371 ^ n6816 ^ n4362 ;
  assign n24373 = ( n7011 & n15822 ) | ( n7011 & n24372 ) | ( n15822 & n24372 ) ;
  assign n24374 = n19460 ^ n4759 ^ 1'b0 ;
  assign n24375 = n18194 ^ n3373 ^ 1'b0 ;
  assign n24376 = n24374 | n24375 ;
  assign n24377 = ( ~n5268 & n24373 ) | ( ~n5268 & n24376 ) | ( n24373 & n24376 ) ;
  assign n24378 = ( ~n14624 & n24370 ) | ( ~n14624 & n24377 ) | ( n24370 & n24377 ) ;
  assign n24379 = ( n3841 & ~n16367 ) | ( n3841 & n21765 ) | ( ~n16367 & n21765 ) ;
  assign n24380 = n4199 | n6952 ;
  assign n24381 = n465 | n24380 ;
  assign n24382 = ( n962 & ~n5862 ) | ( n962 & n17498 ) | ( ~n5862 & n17498 ) ;
  assign n24383 = ( ~n5754 & n14977 ) | ( ~n5754 & n19255 ) | ( n14977 & n19255 ) ;
  assign n24384 = n1217 & ~n24383 ;
  assign n24385 = ( n3445 & n12988 ) | ( n3445 & n19714 ) | ( n12988 & n19714 ) ;
  assign n24386 = n9509 ^ n7052 ^ n2087 ;
  assign n24387 = n4077 | n24386 ;
  assign n24388 = n24387 ^ n3928 ^ 1'b0 ;
  assign n24389 = n24388 ^ n9882 ^ n8585 ;
  assign n24390 = ( n464 & n2374 ) | ( n464 & n10962 ) | ( n2374 & n10962 ) ;
  assign n24391 = ( n1834 & ~n8599 ) | ( n1834 & n16734 ) | ( ~n8599 & n16734 ) ;
  assign n24395 = n2971 | n19008 ;
  assign n24396 = n24395 ^ n7556 ^ 1'b0 ;
  assign n24397 = ( ~n9170 & n9829 ) | ( ~n9170 & n24396 ) | ( n9829 & n24396 ) ;
  assign n24394 = n15312 ^ n9648 ^ 1'b0 ;
  assign n24392 = n688 | n18451 ;
  assign n24393 = n24392 ^ n19225 ^ 1'b0 ;
  assign n24398 = n24397 ^ n24394 ^ n24393 ;
  assign n24399 = ( n11016 & n24391 ) | ( n11016 & ~n24398 ) | ( n24391 & ~n24398 ) ;
  assign n24403 = n890 | n10494 ;
  assign n24401 = ( n2886 & ~n12596 ) | ( n2886 & n23714 ) | ( ~n12596 & n23714 ) ;
  assign n24402 = ( n6995 & n21487 ) | ( n6995 & ~n24401 ) | ( n21487 & ~n24401 ) ;
  assign n24400 = n12896 ^ n2173 ^ 1'b0 ;
  assign n24404 = n24403 ^ n24402 ^ n24400 ;
  assign n24405 = n22206 ^ n12042 ^ n4401 ;
  assign n24406 = ~n15079 & n23967 ;
  assign n24407 = ~n14150 & n24406 ;
  assign n24408 = n3659 | n24407 ;
  assign n24409 = n3293 & ~n24408 ;
  assign n24410 = n12767 & ~n19215 ;
  assign n24411 = n5842 & n24410 ;
  assign n24412 = n24411 ^ n20726 ^ n19469 ;
  assign n24413 = n23092 ^ n14439 ^ n10137 ;
  assign n24414 = n22782 ^ n10242 ^ n1009 ;
  assign n24415 = ( n17860 & n21339 ) | ( n17860 & ~n24414 ) | ( n21339 & ~n24414 ) ;
  assign n24416 = x174 & ~n22541 ;
  assign n24417 = ~n12630 & n24416 ;
  assign n24418 = n22506 ^ n5787 ^ 1'b0 ;
  assign n24419 = ~n6096 & n24418 ;
  assign n24420 = n12485 ^ n12395 ^ n6164 ;
  assign n24421 = ( n18285 & ~n24419 ) | ( n18285 & n24420 ) | ( ~n24419 & n24420 ) ;
  assign n24422 = n24421 ^ n10293 ^ n459 ;
  assign n24423 = n16040 ^ n3209 ^ 1'b0 ;
  assign n24424 = n451 | n24423 ;
  assign n24425 = n10543 & ~n11338 ;
  assign n24426 = n12071 & n24425 ;
  assign n24427 = ~n20656 & n21141 ;
  assign n24428 = n24426 & n24427 ;
  assign n24429 = ( n10545 & n12705 ) | ( n10545 & ~n13807 ) | ( n12705 & ~n13807 ) ;
  assign n24433 = n13887 ^ n11084 ^ n7755 ;
  assign n24434 = n24433 ^ n2308 ^ 1'b0 ;
  assign n24435 = n14273 & n24434 ;
  assign n24430 = ( n631 & ~n1657 ) | ( n631 & n8648 ) | ( ~n1657 & n8648 ) ;
  assign n24431 = n4095 ^ n2156 ^ 1'b0 ;
  assign n24432 = n24430 & n24431 ;
  assign n24436 = n24435 ^ n24432 ^ n13420 ;
  assign n24437 = ( n3328 & n24429 ) | ( n3328 & n24436 ) | ( n24429 & n24436 ) ;
  assign n24438 = n5815 ^ n5056 ^ n4658 ;
  assign n24439 = n13343 ^ n3232 ^ n1469 ;
  assign n24440 = n4366 ^ n1909 ^ n345 ;
  assign n24441 = n8850 & n24440 ;
  assign n24442 = n24441 ^ n19095 ^ 1'b0 ;
  assign n24443 = n24442 ^ n4323 ^ 1'b0 ;
  assign n24444 = n21515 | n24443 ;
  assign n24445 = n24439 | n24444 ;
  assign n24446 = ~n7781 & n24445 ;
  assign n24447 = n24446 ^ n17460 ^ 1'b0 ;
  assign n24448 = ( ~n1246 & n1361 ) | ( ~n1246 & n3778 ) | ( n1361 & n3778 ) ;
  assign n24449 = ( n778 & n1027 ) | ( n778 & n1274 ) | ( n1027 & n1274 ) ;
  assign n24450 = n24449 ^ n20903 ^ 1'b0 ;
  assign n24451 = n17754 ^ n13249 ^ 1'b0 ;
  assign n24452 = n22823 ^ n20539 ^ n1636 ;
  assign n24453 = n6613 & n24452 ;
  assign n24454 = n24453 ^ n15409 ^ 1'b0 ;
  assign n24455 = n23393 & ~n24454 ;
  assign n24456 = n4725 ^ n1328 ^ 1'b0 ;
  assign n24457 = ( n11252 & ~n14965 ) | ( n11252 & n20556 ) | ( ~n14965 & n20556 ) ;
  assign n24458 = ( n14584 & ~n21816 ) | ( n14584 & n22887 ) | ( ~n21816 & n22887 ) ;
  assign n24459 = ( n9924 & n13668 ) | ( n9924 & ~n13935 ) | ( n13668 & ~n13935 ) ;
  assign n24460 = n24459 ^ n3421 ^ n790 ;
  assign n24461 = x110 & ~n21930 ;
  assign n24462 = n24460 & n24461 ;
  assign n24463 = n23004 ^ n592 ^ 1'b0 ;
  assign n24466 = n8241 & n23220 ;
  assign n24465 = ( ~n3599 & n6001 ) | ( ~n3599 & n12511 ) | ( n6001 & n12511 ) ;
  assign n24464 = n20741 ^ n13747 ^ n9111 ;
  assign n24467 = n24466 ^ n24465 ^ n24464 ;
  assign n24468 = n15230 & n15843 ;
  assign n24469 = n24468 ^ n9539 ^ n6200 ;
  assign n24470 = ( n2020 & ~n8464 ) | ( n2020 & n21112 ) | ( ~n8464 & n21112 ) ;
  assign n24471 = n23226 ^ n20299 ^ n13896 ;
  assign n24472 = n6019 ^ n1181 ^ 1'b0 ;
  assign n24473 = ( n6134 & ~n6862 ) | ( n6134 & n24472 ) | ( ~n6862 & n24472 ) ;
  assign n24474 = n19637 | n24473 ;
  assign n24475 = n24474 ^ n2598 ^ 1'b0 ;
  assign n24476 = ( n3851 & n8162 ) | ( n3851 & ~n21966 ) | ( n8162 & ~n21966 ) ;
  assign n24477 = ( ~n1328 & n10449 ) | ( ~n1328 & n24476 ) | ( n10449 & n24476 ) ;
  assign n24478 = n23838 ^ n6262 ^ n4172 ;
  assign n24479 = n12045 ^ n7275 ^ 1'b0 ;
  assign n24480 = ( ~n20257 & n20473 ) | ( ~n20257 & n24479 ) | ( n20473 & n24479 ) ;
  assign n24481 = ( n12555 & ~n17808 ) | ( n12555 & n24480 ) | ( ~n17808 & n24480 ) ;
  assign n24482 = ( n1920 & ~n2826 ) | ( n1920 & n3805 ) | ( ~n2826 & n3805 ) ;
  assign n24483 = n15457 & ~n24482 ;
  assign n24484 = n15431 ^ x72 ^ 1'b0 ;
  assign n24485 = n24484 ^ n9835 ^ n6522 ;
  assign n24486 = n12228 ^ n1663 ^ 1'b0 ;
  assign n24487 = n16238 & ~n24486 ;
  assign n24488 = n24485 & n24487 ;
  assign n24489 = ( n3727 & ~n6308 ) | ( n3727 & n18848 ) | ( ~n6308 & n18848 ) ;
  assign n24490 = ~n17507 & n24489 ;
  assign n24491 = n24488 & n24490 ;
  assign n24500 = ( n5411 & n12848 ) | ( n5411 & n15364 ) | ( n12848 & n15364 ) ;
  assign n24496 = n9647 & n15813 ;
  assign n24497 = ( ~n5034 & n15058 ) | ( ~n5034 & n24496 ) | ( n15058 & n24496 ) ;
  assign n24498 = ( n10366 & n16388 ) | ( n10366 & n20326 ) | ( n16388 & n20326 ) ;
  assign n24499 = ( n708 & n24497 ) | ( n708 & n24498 ) | ( n24497 & n24498 ) ;
  assign n24492 = ( ~n5309 & n7738 ) | ( ~n5309 & n11656 ) | ( n7738 & n11656 ) ;
  assign n24493 = n24492 ^ n24063 ^ n11946 ;
  assign n24494 = n2474 & n24493 ;
  assign n24495 = ( n12370 & n13599 ) | ( n12370 & ~n24494 ) | ( n13599 & ~n24494 ) ;
  assign n24501 = n24500 ^ n24499 ^ n24495 ;
  assign n24502 = n21755 ^ n9791 ^ n1562 ;
  assign n24503 = n24502 ^ n18664 ^ n7850 ;
  assign n24504 = n24503 ^ n4120 ^ n4018 ;
  assign n24508 = n7648 | n11281 ;
  assign n24509 = ~n3544 & n24508 ;
  assign n24510 = n13465 & n24509 ;
  assign n24506 = ~n8022 & n19249 ;
  assign n24507 = n24506 ^ n21084 ^ 1'b0 ;
  assign n24505 = n13532 ^ n13221 ^ n9840 ;
  assign n24511 = n24510 ^ n24507 ^ n24505 ;
  assign n24512 = ~n20267 & n24511 ;
  assign n24513 = ~n13283 & n24512 ;
  assign n24514 = n14659 | n24513 ;
  assign n24515 = n6770 & ~n24514 ;
  assign n24516 = n24515 ^ n23329 ^ 1'b0 ;
  assign n24517 = n938 & ~n20629 ;
  assign n24518 = n24517 ^ n14899 ^ 1'b0 ;
  assign n24519 = n19839 & n24518 ;
  assign n24526 = ( n2474 & n6417 ) | ( n2474 & ~n10345 ) | ( n6417 & ~n10345 ) ;
  assign n24525 = n21191 ^ n1566 ^ 1'b0 ;
  assign n24521 = n17614 ^ n10335 ^ n4872 ;
  assign n24522 = n12995 ^ n4415 ^ 1'b0 ;
  assign n24523 = ~n24521 & n24522 ;
  assign n24520 = n12785 ^ n11883 ^ n4937 ;
  assign n24524 = n24523 ^ n24520 ^ n12682 ;
  assign n24527 = n24526 ^ n24525 ^ n24524 ;
  assign n24528 = ( n11090 & n18405 ) | ( n11090 & ~n22243 ) | ( n18405 & ~n22243 ) ;
  assign n24529 = n11404 ^ n9489 ^ n4810 ;
  assign n24530 = n24529 ^ n14704 ^ n4163 ;
  assign n24531 = ~n2036 & n5469 ;
  assign n24532 = ~n13325 & n24531 ;
  assign n24533 = n24532 ^ n8871 ^ n5259 ;
  assign n24534 = ( n3566 & ~n4035 ) | ( n3566 & n13135 ) | ( ~n4035 & n13135 ) ;
  assign n24535 = n24534 ^ n301 ^ 1'b0 ;
  assign n24536 = n24533 | n24535 ;
  assign n24537 = n23538 ^ n12399 ^ n6390 ;
  assign n24538 = ( ~n3682 & n18559 ) | ( ~n3682 & n24537 ) | ( n18559 & n24537 ) ;
  assign n24544 = n13946 ^ n6255 ^ n1219 ;
  assign n24539 = ~n1464 & n18705 ;
  assign n24540 = n24539 ^ n6035 ^ n1502 ;
  assign n24541 = n24540 ^ n15923 ^ 1'b0 ;
  assign n24542 = ~n3172 & n24541 ;
  assign n24543 = ( n826 & ~n13860 ) | ( n826 & n24542 ) | ( ~n13860 & n24542 ) ;
  assign n24545 = n24544 ^ n24543 ^ n531 ;
  assign n24546 = n17251 ^ n15817 ^ n8837 ;
  assign n24547 = n24546 ^ n7320 ^ n7135 ;
  assign n24548 = ( n2030 & n21815 ) | ( n2030 & n24547 ) | ( n21815 & n24547 ) ;
  assign n24549 = ( n5994 & n12200 ) | ( n5994 & ~n24548 ) | ( n12200 & ~n24548 ) ;
  assign n24550 = n6966 | n10509 ;
  assign n24551 = n24550 ^ n5394 ^ 1'b0 ;
  assign n24552 = n3354 ^ n2834 ^ n1529 ;
  assign n24553 = ( n24206 & n24551 ) | ( n24206 & ~n24552 ) | ( n24551 & ~n24552 ) ;
  assign n24554 = ( n2020 & n8561 ) | ( n2020 & n15343 ) | ( n8561 & n15343 ) ;
  assign n24555 = n13464 ^ n8163 ^ n6718 ;
  assign n24556 = n24555 ^ n24330 ^ 1'b0 ;
  assign n24557 = n2728 | n13173 ;
  assign n24558 = n24557 ^ n895 ^ 1'b0 ;
  assign n24559 = n24558 ^ n12826 ^ n10606 ;
  assign n24560 = n24559 ^ n22560 ^ n22447 ;
  assign n24561 = ( ~n12343 & n20158 ) | ( ~n12343 & n20711 ) | ( n20158 & n20711 ) ;
  assign n24562 = n24561 ^ n10749 ^ 1'b0 ;
  assign n24563 = n24562 ^ n9576 ^ n2800 ;
  assign n24565 = n17985 ^ n10580 ^ 1'b0 ;
  assign n24566 = n24565 ^ n6287 ^ 1'b0 ;
  assign n24564 = n6854 & ~n22604 ;
  assign n24567 = n24566 ^ n24564 ^ n10368 ;
  assign n24568 = n9041 ^ n7798 ^ n3375 ;
  assign n24569 = n18961 & n24568 ;
  assign n24570 = ( n1226 & n1899 ) | ( n1226 & n4251 ) | ( n1899 & n4251 ) ;
  assign n24571 = n6329 ^ n3066 ^ 1'b0 ;
  assign n24572 = n24570 | n24571 ;
  assign n24573 = n8381 ^ n6999 ^ n5778 ;
  assign n24574 = ( n4101 & n9845 ) | ( n4101 & n24573 ) | ( n9845 & n24573 ) ;
  assign n24575 = n23668 ^ n5940 ^ 1'b0 ;
  assign n24576 = ~n24574 & n24575 ;
  assign n24577 = n20204 ^ n20144 ^ n2729 ;
  assign n24578 = n13627 ^ n9734 ^ n715 ;
  assign n24579 = n24578 ^ n18143 ^ n18129 ;
  assign n24580 = n4071 | n12776 ;
  assign n24581 = n24579 & ~n24580 ;
  assign n24582 = n24581 ^ n14683 ^ n7398 ;
  assign n24583 = ( n10058 & ~n19937 ) | ( n10058 & n24582 ) | ( ~n19937 & n24582 ) ;
  assign n24585 = n14951 ^ n6583 ^ n4540 ;
  assign n24586 = n24585 ^ n16007 ^ n1794 ;
  assign n24584 = n16275 ^ n11567 ^ 1'b0 ;
  assign n24587 = n24586 ^ n24584 ^ n18931 ;
  assign n24588 = n21380 ^ n19135 ^ 1'b0 ;
  assign n24589 = n20793 ^ n7801 ^ n1215 ;
  assign n24590 = n7923 & ~n24589 ;
  assign n24591 = ~n3609 & n7039 ;
  assign n24592 = n24591 ^ n4921 ^ 1'b0 ;
  assign n24593 = ( n5718 & n17863 ) | ( n5718 & ~n24592 ) | ( n17863 & ~n24592 ) ;
  assign n24594 = n10639 & n24593 ;
  assign n24595 = ( n15255 & ~n24590 ) | ( n15255 & n24594 ) | ( ~n24590 & n24594 ) ;
  assign n24596 = n15817 ^ n13735 ^ 1'b0 ;
  assign n24597 = ( n8356 & n9203 ) | ( n8356 & n21495 ) | ( n9203 & n21495 ) ;
  assign n24598 = n24597 ^ n14879 ^ n8005 ;
  assign n24599 = n11591 | n24598 ;
  assign n24600 = n24599 ^ n14263 ^ 1'b0 ;
  assign n24601 = n23024 ^ n11048 ^ n8124 ;
  assign n24602 = n20354 ^ n14235 ^ n9600 ;
  assign n24603 = ~n9202 & n20175 ;
  assign n24604 = n24603 ^ n13163 ^ n5994 ;
  assign n24605 = n24604 ^ n7764 ^ n1717 ;
  assign n24606 = n17926 ^ n17731 ^ 1'b0 ;
  assign n24607 = ( n5110 & n8110 ) | ( n5110 & ~n18284 ) | ( n8110 & ~n18284 ) ;
  assign n24608 = ( n1094 & n14038 ) | ( n1094 & ~n24607 ) | ( n14038 & ~n24607 ) ;
  assign n24609 = ( ~n5864 & n5918 ) | ( ~n5864 & n16649 ) | ( n5918 & n16649 ) ;
  assign n24612 = ( n2555 & ~n12365 ) | ( n2555 & n13718 ) | ( ~n12365 & n13718 ) ;
  assign n24610 = n17229 ^ n10893 ^ n10764 ;
  assign n24611 = n17001 & ~n24610 ;
  assign n24613 = n24612 ^ n24611 ^ 1'b0 ;
  assign n24615 = ~n826 & n23383 ;
  assign n24616 = ( n8701 & n12627 ) | ( n8701 & n24615 ) | ( n12627 & n24615 ) ;
  assign n24614 = ~n5107 & n6911 ;
  assign n24617 = n24616 ^ n24614 ^ 1'b0 ;
  assign n24618 = n24617 ^ n22636 ^ n19904 ;
  assign n24619 = n10567 ^ n1897 ^ n956 ;
  assign n24620 = ( n1747 & ~n8417 ) | ( n1747 & n24619 ) | ( ~n8417 & n24619 ) ;
  assign n24621 = n24620 ^ n8669 ^ n3190 ;
  assign n24622 = n15763 ^ n10444 ^ 1'b0 ;
  assign n24623 = ( n8537 & n24621 ) | ( n8537 & ~n24622 ) | ( n24621 & ~n24622 ) ;
  assign n24624 = ( n5725 & n17987 ) | ( n5725 & ~n24623 ) | ( n17987 & ~n24623 ) ;
  assign n24625 = n23680 ^ n17579 ^ x222 ;
  assign n24630 = ( n9655 & n13231 ) | ( n9655 & n14776 ) | ( n13231 & n14776 ) ;
  assign n24627 = ~n11400 & n13314 ;
  assign n24628 = n5318 & n24627 ;
  assign n24626 = n4780 ^ n3504 ^ n883 ;
  assign n24629 = n24628 ^ n24626 ^ 1'b0 ;
  assign n24631 = n24630 ^ n24629 ^ n4017 ;
  assign n24632 = n23594 ^ n13697 ^ n4321 ;
  assign n24633 = n7793 | n17144 ;
  assign n24634 = n24633 ^ n1186 ^ 1'b0 ;
  assign n24635 = ~n12261 & n24634 ;
  assign n24636 = n6405 ^ n632 ^ 1'b0 ;
  assign n24637 = n11603 ^ n9284 ^ 1'b0 ;
  assign n24638 = n8757 & n24637 ;
  assign n24639 = n24638 ^ n18496 ^ n392 ;
  assign n24640 = n17814 ^ n15768 ^ n2407 ;
  assign n24641 = n15542 | n24640 ;
  assign n24642 = ( n12277 & ~n19779 ) | ( n12277 & n24641 ) | ( ~n19779 & n24641 ) ;
  assign n24643 = n24642 ^ n12141 ^ n9261 ;
  assign n24644 = n24643 ^ n20853 ^ n17556 ;
  assign n24652 = n7034 ^ n2693 ^ x48 ;
  assign n24651 = n3112 & ~n12649 ;
  assign n24653 = n24652 ^ n24651 ^ 1'b0 ;
  assign n24654 = ( ~n6776 & n12125 ) | ( ~n6776 & n24653 ) | ( n12125 & n24653 ) ;
  assign n24649 = n9060 ^ n4419 ^ n1571 ;
  assign n24645 = n12449 ^ n7765 ^ 1'b0 ;
  assign n24646 = ( ~n3545 & n7872 ) | ( ~n3545 & n24645 ) | ( n7872 & n24645 ) ;
  assign n24647 = ( ~n5699 & n12956 ) | ( ~n5699 & n24646 ) | ( n12956 & n24646 ) ;
  assign n24648 = ( n17184 & n21458 ) | ( n17184 & ~n24647 ) | ( n21458 & ~n24647 ) ;
  assign n24650 = n24649 ^ n24648 ^ n10819 ;
  assign n24655 = n24654 ^ n24650 ^ n8096 ;
  assign n24656 = ( n1828 & ~n8271 ) | ( n1828 & n10801 ) | ( ~n8271 & n10801 ) ;
  assign n24657 = ( n330 & ~n12238 ) | ( n330 & n16405 ) | ( ~n12238 & n16405 ) ;
  assign n24658 = ( n3877 & n24656 ) | ( n3877 & ~n24657 ) | ( n24656 & ~n24657 ) ;
  assign n24659 = ~n8983 & n24658 ;
  assign n24660 = n6767 ^ n3367 ^ n523 ;
  assign n24661 = n24374 ^ n6728 ^ n436 ;
  assign n24662 = ( n7169 & n24660 ) | ( n7169 & n24661 ) | ( n24660 & n24661 ) ;
  assign n24663 = ( n553 & n5970 ) | ( n553 & ~n6835 ) | ( n5970 & ~n6835 ) ;
  assign n24664 = n5632 & n24663 ;
  assign n24665 = n24664 ^ n375 ^ x133 ;
  assign n24666 = n24665 ^ n22926 ^ 1'b0 ;
  assign n24667 = n12984 ^ n10017 ^ n529 ;
  assign n24668 = n24667 ^ n17891 ^ n11429 ;
  assign n24669 = ( n5442 & n20453 ) | ( n5442 & ~n24668 ) | ( n20453 & ~n24668 ) ;
  assign n24670 = n24085 ^ n19244 ^ n17434 ;
  assign n24671 = n8910 & n24670 ;
  assign n24672 = n24499 ^ n18332 ^ n7986 ;
  assign n24673 = n24672 ^ n17257 ^ n12987 ;
  assign n24675 = n11375 ^ n7709 ^ n1170 ;
  assign n24674 = n17708 ^ n12983 ^ n6531 ;
  assign n24676 = n24675 ^ n24674 ^ n544 ;
  assign n24678 = n10036 & n14190 ;
  assign n24679 = n13407 & n24678 ;
  assign n24680 = ( n3733 & n12801 ) | ( n3733 & ~n24679 ) | ( n12801 & ~n24679 ) ;
  assign n24681 = n24680 ^ n21188 ^ 1'b0 ;
  assign n24682 = ~n502 & n24681 ;
  assign n24677 = ( n10038 & n17295 ) | ( n10038 & n23640 ) | ( n17295 & n23640 ) ;
  assign n24683 = n24682 ^ n24677 ^ n11185 ;
  assign n24687 = n9510 | n9549 ;
  assign n24684 = n12241 ^ n1896 ^ n1320 ;
  assign n24685 = ( n1630 & ~n23838 ) | ( n1630 & n24684 ) | ( ~n23838 & n24684 ) ;
  assign n24686 = ~n19741 & n24685 ;
  assign n24688 = n24687 ^ n24686 ^ 1'b0 ;
  assign n24689 = n20789 ^ n6574 ^ n1573 ;
  assign n24690 = ( n1235 & n12856 ) | ( n1235 & n24689 ) | ( n12856 & n24689 ) ;
  assign n24691 = n15014 ^ n14198 ^ 1'b0 ;
  assign n24692 = n24690 & ~n24691 ;
  assign n24693 = ( n3997 & ~n16762 ) | ( n3997 & n18749 ) | ( ~n16762 & n18749 ) ;
  assign n24694 = n19315 ^ n9290 ^ 1'b0 ;
  assign n24695 = n24694 ^ n9546 ^ 1'b0 ;
  assign n24696 = n5304 | n24695 ;
  assign n24697 = n24696 ^ n16854 ^ n8541 ;
  assign n24703 = ( n2717 & ~n2735 ) | ( n2717 & n5450 ) | ( ~n2735 & n5450 ) ;
  assign n24704 = n1901 & ~n24703 ;
  assign n24701 = ( n4027 & n13767 ) | ( n4027 & n14111 ) | ( n13767 & n14111 ) ;
  assign n24699 = n23848 ^ n16427 ^ n7774 ;
  assign n24700 = n5429 & n24699 ;
  assign n24702 = n24701 ^ n24700 ^ 1'b0 ;
  assign n24698 = n17113 ^ n11654 ^ n2786 ;
  assign n24705 = n24704 ^ n24702 ^ n24698 ;
  assign n24706 = n2882 & ~n24705 ;
  assign n24707 = n4428 | n18347 ;
  assign n24708 = n24707 ^ n17985 ^ n269 ;
  assign n24711 = n13798 & ~n17366 ;
  assign n24709 = ( n554 & ~n1997 ) | ( n554 & n2015 ) | ( ~n1997 & n2015 ) ;
  assign n24710 = ( n7658 & ~n15200 ) | ( n7658 & n24709 ) | ( ~n15200 & n24709 ) ;
  assign n24712 = n24711 ^ n24710 ^ n934 ;
  assign n24713 = ( n8263 & ~n13261 ) | ( n8263 & n24712 ) | ( ~n13261 & n24712 ) ;
  assign n24714 = ( n812 & ~n24708 ) | ( n812 & n24713 ) | ( ~n24708 & n24713 ) ;
  assign n24717 = ( ~n1868 & n3098 ) | ( ~n1868 & n5251 ) | ( n3098 & n5251 ) ;
  assign n24715 = ( n2296 & n8628 ) | ( n2296 & n21328 ) | ( n8628 & n21328 ) ;
  assign n24716 = n24715 ^ n6381 ^ n2167 ;
  assign n24718 = n24717 ^ n24716 ^ n15392 ;
  assign n24719 = n13123 ^ n6106 ^ 1'b0 ;
  assign n24720 = ( n1895 & ~n4288 ) | ( n1895 & n24719 ) | ( ~n4288 & n24719 ) ;
  assign n24723 = n698 | n11081 ;
  assign n24721 = n17100 ^ n2221 ^ 1'b0 ;
  assign n24722 = n5389 & n24721 ;
  assign n24724 = n24723 ^ n24722 ^ n9211 ;
  assign n24725 = n23210 ^ n7930 ^ n7499 ;
  assign n24726 = ( x148 & ~n3836 ) | ( x148 & n10330 ) | ( ~n3836 & n10330 ) ;
  assign n24727 = ( ~n6285 & n17295 ) | ( ~n6285 & n24726 ) | ( n17295 & n24726 ) ;
  assign n24728 = n24727 ^ n19856 ^ 1'b0 ;
  assign n24729 = ( ~n5275 & n17810 ) | ( ~n5275 & n24728 ) | ( n17810 & n24728 ) ;
  assign n24730 = ( ~n23331 & n24244 ) | ( ~n23331 & n24729 ) | ( n24244 & n24729 ) ;
  assign n24731 = n15052 & n17093 ;
  assign n24732 = ( n640 & n14357 ) | ( n640 & n24731 ) | ( n14357 & n24731 ) ;
  assign n24733 = n16053 ^ n13783 ^ n9819 ;
  assign n24734 = n20814 | n22574 ;
  assign n24735 = n24733 | n24734 ;
  assign n24736 = n14722 | n24735 ;
  assign n24737 = ( ~n7189 & n12125 ) | ( ~n7189 & n16052 ) | ( n12125 & n16052 ) ;
  assign n24738 = n24737 ^ n18308 ^ n13767 ;
  assign n24739 = n14235 ^ n5564 ^ n992 ;
  assign n24740 = ( n12382 & ~n14798 ) | ( n12382 & n20434 ) | ( ~n14798 & n20434 ) ;
  assign n24741 = n24739 | n24740 ;
  assign n24742 = n24741 ^ n13820 ^ n3053 ;
  assign n24743 = ~n2865 & n24742 ;
  assign n24745 = ( n1126 & n4277 ) | ( n1126 & ~n4336 ) | ( n4277 & ~n4336 ) ;
  assign n24746 = n24745 ^ n21898 ^ n6706 ;
  assign n24747 = ( n6597 & ~n10077 ) | ( n6597 & n11858 ) | ( ~n10077 & n11858 ) ;
  assign n24748 = n9658 | n24747 ;
  assign n24749 = n7654 & ~n24748 ;
  assign n24750 = n24749 ^ n10778 ^ 1'b0 ;
  assign n24751 = n24746 | n24750 ;
  assign n24744 = n6287 & ~n18868 ;
  assign n24752 = n24751 ^ n24744 ^ 1'b0 ;
  assign n24753 = n9501 ^ n442 ^ 1'b0 ;
  assign n24754 = ( n9257 & ~n24752 ) | ( n9257 & n24753 ) | ( ~n24752 & n24753 ) ;
  assign n24755 = n5807 & ~n9963 ;
  assign n24756 = ( n533 & n639 ) | ( n533 & ~n16811 ) | ( n639 & ~n16811 ) ;
  assign n24757 = n8183 & ~n24756 ;
  assign n24758 = n24755 & n24757 ;
  assign n24759 = n3681 | n17408 ;
  assign n24760 = n24759 ^ n19448 ^ 1'b0 ;
  assign n24761 = n5333 ^ n3650 ^ n2869 ;
  assign n24762 = ( n12768 & n21348 ) | ( n12768 & ~n24761 ) | ( n21348 & ~n24761 ) ;
  assign n24763 = ( n2717 & n18857 ) | ( n2717 & n24762 ) | ( n18857 & n24762 ) ;
  assign n24764 = n15720 ^ n7914 ^ n7770 ;
  assign n24765 = n2599 ^ n2238 ^ 1'b0 ;
  assign n24766 = n24311 ^ n21019 ^ n15427 ;
  assign n24767 = n6602 ^ n2625 ^ n848 ;
  assign n24768 = n24767 ^ n19594 ^ n14988 ;
  assign n24769 = n17368 ^ n14942 ^ n1951 ;
  assign n24770 = ( n1725 & ~n5156 ) | ( n1725 & n9123 ) | ( ~n5156 & n9123 ) ;
  assign n24771 = n24770 ^ n4015 ^ n792 ;
  assign n24772 = ( ~n19142 & n19294 ) | ( ~n19142 & n24771 ) | ( n19294 & n24771 ) ;
  assign n24773 = n24769 | n24772 ;
  assign n24774 = n24768 | n24773 ;
  assign n24777 = n11697 ^ n10375 ^ n6804 ;
  assign n24778 = n24777 ^ n21545 ^ n11361 ;
  assign n24775 = ~n16341 & n18622 ;
  assign n24776 = n24775 ^ n5472 ^ 1'b0 ;
  assign n24779 = n24778 ^ n24776 ^ n1876 ;
  assign n24785 = n3249 | n6574 ;
  assign n24786 = n24785 ^ n15733 ^ 1'b0 ;
  assign n24782 = ( ~n5274 & n10747 ) | ( ~n5274 & n12274 ) | ( n10747 & n12274 ) ;
  assign n24783 = ( n4599 & ~n11948 ) | ( n4599 & n24782 ) | ( ~n11948 & n24782 ) ;
  assign n24784 = n6297 & n24783 ;
  assign n24780 = ( n3086 & n14524 ) | ( n3086 & ~n24414 ) | ( n14524 & ~n24414 ) ;
  assign n24781 = n24780 ^ n16136 ^ n270 ;
  assign n24787 = n24786 ^ n24784 ^ n24781 ;
  assign n24788 = n2036 | n3088 ;
  assign n24789 = n24788 ^ n2982 ^ n2770 ;
  assign n24790 = n1031 | n6559 ;
  assign n24791 = n790 & ~n24790 ;
  assign n24792 = n24791 ^ n11772 ^ 1'b0 ;
  assign n24793 = n19183 & ~n24792 ;
  assign n24794 = ( ~n4186 & n5999 ) | ( ~n4186 & n12634 ) | ( n5999 & n12634 ) ;
  assign n24795 = n24794 ^ n19164 ^ 1'b0 ;
  assign n24796 = ( n12656 & ~n24793 ) | ( n12656 & n24795 ) | ( ~n24793 & n24795 ) ;
  assign n24797 = n24796 ^ n6019 ^ 1'b0 ;
  assign n24798 = ~n7194 & n24797 ;
  assign n24799 = n24798 ^ n6214 ^ n4662 ;
  assign n24800 = n1487 & ~n12446 ;
  assign n24801 = ( n3158 & n12927 ) | ( n3158 & n24800 ) | ( n12927 & n24800 ) ;
  assign n24802 = ~n5581 & n11917 ;
  assign n24803 = ~n24801 & n24802 ;
  assign n24807 = ( n521 & ~n1711 ) | ( n521 & n2727 ) | ( ~n1711 & n2727 ) ;
  assign n24805 = n2231 ^ n1256 ^ n851 ;
  assign n24804 = n5249 | n6142 ;
  assign n24806 = n24805 ^ n24804 ^ 1'b0 ;
  assign n24808 = n24807 ^ n24806 ^ n14661 ;
  assign n24809 = n4907 | n11186 ;
  assign n24810 = n24808 | n24809 ;
  assign n24811 = n6396 ^ n4992 ^ x142 ;
  assign n24812 = ( n19757 & ~n23469 ) | ( n19757 & n24811 ) | ( ~n23469 & n24811 ) ;
  assign n24813 = ( ~n15388 & n24810 ) | ( ~n15388 & n24812 ) | ( n24810 & n24812 ) ;
  assign n24814 = ( n4038 & ~n4101 ) | ( n4038 & n5630 ) | ( ~n4101 & n5630 ) ;
  assign n24815 = n24814 ^ n8986 ^ 1'b0 ;
  assign n24816 = n14519 & ~n24815 ;
  assign n24819 = ~n8827 & n19271 ;
  assign n24820 = n14061 & ~n24819 ;
  assign n24817 = n24227 ^ n9831 ^ n9672 ;
  assign n24818 = n24817 ^ n6069 ^ 1'b0 ;
  assign n24821 = n24820 ^ n24818 ^ n17792 ;
  assign n24822 = ( n4686 & ~n10129 ) | ( n4686 & n15199 ) | ( ~n10129 & n15199 ) ;
  assign n24823 = ( n14414 & ~n15443 ) | ( n14414 & n24822 ) | ( ~n15443 & n24822 ) ;
  assign n24824 = n7521 & n16429 ;
  assign n24825 = n1143 & n24824 ;
  assign n24826 = n13673 ^ n8475 ^ n4812 ;
  assign n24827 = ( ~n12291 & n15175 ) | ( ~n12291 & n21617 ) | ( n15175 & n21617 ) ;
  assign n24828 = ( ~n13775 & n24826 ) | ( ~n13775 & n24827 ) | ( n24826 & n24827 ) ;
  assign n24829 = ( n11989 & ~n20767 ) | ( n11989 & n21868 ) | ( ~n20767 & n21868 ) ;
  assign n24830 = n24829 ^ n20140 ^ 1'b0 ;
  assign n24831 = ~n11541 & n24830 ;
  assign n24832 = ( n4561 & n5623 ) | ( n4561 & ~n24831 ) | ( n5623 & ~n24831 ) ;
  assign n24833 = ( n24825 & n24828 ) | ( n24825 & ~n24832 ) | ( n24828 & ~n24832 ) ;
  assign n24834 = ( n4064 & n5140 ) | ( n4064 & n9281 ) | ( n5140 & n9281 ) ;
  assign n24835 = n3469 ^ n2932 ^ 1'b0 ;
  assign n24836 = ~n777 & n24835 ;
  assign n24837 = ( n8647 & ~n24834 ) | ( n8647 & n24836 ) | ( ~n24834 & n24836 ) ;
  assign n24839 = ( ~n3752 & n9254 ) | ( ~n3752 & n20372 ) | ( n9254 & n20372 ) ;
  assign n24838 = ( n2808 & ~n8707 ) | ( n2808 & n18683 ) | ( ~n8707 & n18683 ) ;
  assign n24840 = n24839 ^ n24838 ^ n18452 ;
  assign n24841 = n13065 ^ n2291 ^ 1'b0 ;
  assign n24842 = n14956 | n24841 ;
  assign n24846 = ( n271 & n4242 ) | ( n271 & n11511 ) | ( n4242 & n11511 ) ;
  assign n24847 = ( n982 & ~n8761 ) | ( n982 & n24846 ) | ( ~n8761 & n24846 ) ;
  assign n24845 = n11164 ^ n1660 ^ 1'b0 ;
  assign n24843 = n14744 ^ n6711 ^ 1'b0 ;
  assign n24844 = n24843 ^ n19340 ^ n7958 ;
  assign n24848 = n24847 ^ n24845 ^ n24844 ;
  assign n24849 = n10713 ^ n9872 ^ n7088 ;
  assign n24850 = n24849 ^ n18897 ^ n18328 ;
  assign n24851 = ( ~n12274 & n15185 ) | ( ~n12274 & n24850 ) | ( n15185 & n24850 ) ;
  assign n24852 = n12508 ^ n9564 ^ 1'b0 ;
  assign n24853 = n2345 ^ n1754 ^ 1'b0 ;
  assign n24854 = ~n10262 & n24853 ;
  assign n24855 = n24854 ^ n13658 ^ 1'b0 ;
  assign n24856 = ( ~n24851 & n24852 ) | ( ~n24851 & n24855 ) | ( n24852 & n24855 ) ;
  assign n24858 = n7733 ^ n7348 ^ n2784 ;
  assign n24857 = n22139 ^ n16004 ^ n10948 ;
  assign n24859 = n24858 ^ n24857 ^ n24288 ;
  assign n24860 = ( n3268 & n9828 ) | ( n3268 & n17007 ) | ( n9828 & n17007 ) ;
  assign n24861 = ( n12657 & n15644 ) | ( n12657 & n16854 ) | ( n15644 & n16854 ) ;
  assign n24862 = n24861 ^ n14937 ^ 1'b0 ;
  assign n24863 = n24860 & ~n24862 ;
  assign n24864 = n7435 ^ n5276 ^ 1'b0 ;
  assign n24866 = n8571 ^ n3286 ^ x242 ;
  assign n24865 = n22294 ^ n6769 ^ n1923 ;
  assign n24867 = n24866 ^ n24865 ^ n4105 ;
  assign n24868 = ( n13657 & ~n20878 ) | ( n13657 & n24867 ) | ( ~n20878 & n24867 ) ;
  assign n24869 = ( ~n4403 & n6056 ) | ( ~n4403 & n8390 ) | ( n6056 & n8390 ) ;
  assign n24870 = ~n20123 & n24869 ;
  assign n24871 = n17132 & n24870 ;
  assign n24872 = n12475 & ~n24871 ;
  assign n24873 = ~n1336 & n23036 ;
  assign n24874 = n24873 ^ n3060 ^ 1'b0 ;
  assign n24875 = n24874 ^ n276 ^ 1'b0 ;
  assign n24876 = ~n18770 & n24875 ;
  assign n24877 = ( n2322 & ~n10240 ) | ( n2322 & n11131 ) | ( ~n10240 & n11131 ) ;
  assign n24878 = ( n9551 & ~n23537 ) | ( n9551 & n24877 ) | ( ~n23537 & n24877 ) ;
  assign n24879 = ( n3183 & n6895 ) | ( n3183 & ~n7604 ) | ( n6895 & ~n7604 ) ;
  assign n24880 = n24879 ^ n19112 ^ 1'b0 ;
  assign n24889 = ( n776 & n3753 ) | ( n776 & n5981 ) | ( n3753 & n5981 ) ;
  assign n24884 = n18721 ^ n11106 ^ n7592 ;
  assign n24885 = n10194 | n13796 ;
  assign n24886 = n24885 ^ n5740 ^ 1'b0 ;
  assign n24887 = n24886 ^ n13340 ^ n6434 ;
  assign n24888 = ( ~n12337 & n24884 ) | ( ~n12337 & n24887 ) | ( n24884 & n24887 ) ;
  assign n24881 = ( n5242 & n8492 ) | ( n5242 & n23509 ) | ( n8492 & n23509 ) ;
  assign n24882 = n24881 ^ n14968 ^ n14052 ;
  assign n24883 = ( n6326 & ~n19244 ) | ( n6326 & n24882 ) | ( ~n19244 & n24882 ) ;
  assign n24890 = n24889 ^ n24888 ^ n24883 ;
  assign n24891 = n22075 ^ n7990 ^ n6105 ;
  assign n24892 = ( n8445 & n11279 ) | ( n8445 & n24891 ) | ( n11279 & n24891 ) ;
  assign n24893 = n24892 ^ n21458 ^ 1'b0 ;
  assign n24894 = n17562 ^ n12104 ^ 1'b0 ;
  assign n24895 = ( n855 & ~n3703 ) | ( n855 & n8050 ) | ( ~n3703 & n8050 ) ;
  assign n24896 = ( ~n4156 & n21187 ) | ( ~n4156 & n24895 ) | ( n21187 & n24895 ) ;
  assign n24897 = n24896 ^ n16670 ^ n4618 ;
  assign n24898 = n11242 & n13377 ;
  assign n24899 = n24897 & n24898 ;
  assign n24900 = ( n2612 & n3578 ) | ( n2612 & ~n10918 ) | ( n3578 & ~n10918 ) ;
  assign n24901 = n24900 ^ n4735 ^ n2364 ;
  assign n24902 = n24901 ^ n4995 ^ n1450 ;
  assign n24903 = n24902 ^ n15275 ^ n4188 ;
  assign n24904 = n652 | n7557 ;
  assign n24905 = ( ~n319 & n3380 ) | ( ~n319 & n24904 ) | ( n3380 & n24904 ) ;
  assign n24906 = ( n3069 & n9214 ) | ( n3069 & n24905 ) | ( n9214 & n24905 ) ;
  assign n24907 = n12363 | n24906 ;
  assign n24908 = n24907 ^ n1246 ^ 1'b0 ;
  assign n24909 = ~n23326 & n24908 ;
  assign n24910 = ~n12661 & n24909 ;
  assign n24911 = ( ~n3155 & n21136 ) | ( ~n3155 & n21913 ) | ( n21136 & n21913 ) ;
  assign n24912 = ( n11773 & n12671 ) | ( n11773 & ~n19496 ) | ( n12671 & ~n19496 ) ;
  assign n24913 = ~n970 & n15469 ;
  assign n24914 = n24913 ^ n4192 ^ 1'b0 ;
  assign n24915 = n24914 ^ n16169 ^ n827 ;
  assign n24916 = n4839 & n15040 ;
  assign n24917 = n24916 ^ n17583 ^ 1'b0 ;
  assign n24918 = ~n5570 & n22595 ;
  assign n24919 = ( n5912 & n19623 ) | ( n5912 & ~n21081 ) | ( n19623 & ~n21081 ) ;
  assign n24920 = ( n2437 & ~n24918 ) | ( n2437 & n24919 ) | ( ~n24918 & n24919 ) ;
  assign n24921 = ( n1833 & ~n15774 ) | ( n1833 & n19464 ) | ( ~n15774 & n19464 ) ;
  assign n24922 = n24921 ^ n11965 ^ n4097 ;
  assign n24923 = n990 & ~n24922 ;
  assign n24924 = ~n6195 & n24923 ;
  assign n24925 = n21989 ^ n2117 ^ 1'b0 ;
  assign n24926 = n24925 ^ n22756 ^ x224 ;
  assign n24929 = n20848 ^ n4160 ^ 1'b0 ;
  assign n24927 = n7736 & ~n10396 ;
  assign n24928 = n24927 ^ n4853 ^ 1'b0 ;
  assign n24930 = n24929 ^ n24928 ^ n12533 ;
  assign n24931 = n20405 ^ n2287 ^ n721 ;
  assign n24932 = ( n4684 & n10500 ) | ( n4684 & ~n13481 ) | ( n10500 & ~n13481 ) ;
  assign n24933 = ( ~n962 & n24931 ) | ( ~n962 & n24932 ) | ( n24931 & n24932 ) ;
  assign n24934 = ( ~n16039 & n21543 ) | ( ~n16039 & n24933 ) | ( n21543 & n24933 ) ;
  assign n24941 = n12407 ^ n6043 ^ n6031 ;
  assign n24942 = n24941 ^ n19625 ^ n5337 ;
  assign n24937 = n15231 ^ n1608 ^ 1'b0 ;
  assign n24938 = n24937 ^ n12887 ^ n9937 ;
  assign n24939 = n24938 ^ n8333 ^ n4858 ;
  assign n24940 = n24939 ^ n11109 ^ n6036 ;
  assign n24935 = n9117 & n9519 ;
  assign n24936 = ~n17146 & n24935 ;
  assign n24943 = n24942 ^ n24940 ^ n24936 ;
  assign n24944 = n1527 & n7341 ;
  assign n24945 = ( x60 & ~n4698 ) | ( x60 & n5526 ) | ( ~n4698 & n5526 ) ;
  assign n24946 = n24945 ^ n12395 ^ 1'b0 ;
  assign n24947 = n23346 ^ n17618 ^ n2604 ;
  assign n24948 = ~n772 & n8595 ;
  assign n24949 = ~n24947 & n24948 ;
  assign n24950 = n1087 & n1774 ;
  assign n24951 = n24949 | n24950 ;
  assign n24952 = n11926 | n24951 ;
  assign n24953 = ( n11977 & n24946 ) | ( n11977 & ~n24952 ) | ( n24946 & ~n24952 ) ;
  assign n24954 = n13767 ^ n302 ^ 1'b0 ;
  assign n24955 = n14519 & n24954 ;
  assign n24956 = n24159 ^ n23450 ^ n10745 ;
  assign n24957 = n24956 ^ n8747 ^ 1'b0 ;
  assign n24958 = ~n22466 & n24957 ;
  assign n24959 = ~n24955 & n24958 ;
  assign n24960 = n24959 ^ n14998 ^ n4132 ;
  assign n24961 = n17937 ^ n3049 ^ 1'b0 ;
  assign n24962 = n21719 & n24961 ;
  assign n24963 = ( n16164 & n17536 ) | ( n16164 & n24642 ) | ( n17536 & n24642 ) ;
  assign n24964 = n24963 ^ n10291 ^ 1'b0 ;
  assign n24965 = n16520 | n24964 ;
  assign n24967 = ( x66 & n6610 ) | ( x66 & ~n10210 ) | ( n6610 & ~n10210 ) ;
  assign n24966 = ~n5312 & n10461 ;
  assign n24968 = n24967 ^ n24966 ^ 1'b0 ;
  assign n24969 = ( n6671 & n7139 ) | ( n6671 & n12516 ) | ( n7139 & n12516 ) ;
  assign n24970 = ( ~n6047 & n15268 ) | ( ~n6047 & n24969 ) | ( n15268 & n24969 ) ;
  assign n24971 = ( ~n4395 & n24968 ) | ( ~n4395 & n24970 ) | ( n24968 & n24970 ) ;
  assign n24972 = ( n269 & ~n6762 ) | ( n269 & n7804 ) | ( ~n6762 & n7804 ) ;
  assign n24973 = n8153 & ~n24972 ;
  assign n24974 = ( n536 & n10158 ) | ( n536 & n17322 ) | ( n10158 & n17322 ) ;
  assign n24975 = n24974 ^ n14631 ^ n380 ;
  assign n24976 = ( n2362 & n2820 ) | ( n2362 & ~n23695 ) | ( n2820 & ~n23695 ) ;
  assign n24977 = n24976 ^ n11348 ^ n330 ;
  assign n24978 = ( ~n4213 & n12948 ) | ( ~n4213 & n23171 ) | ( n12948 & n23171 ) ;
  assign n24979 = n16829 & n24978 ;
  assign n24980 = n24979 ^ n13630 ^ 1'b0 ;
  assign n24983 = ( n2582 & n8703 ) | ( n2582 & n13132 ) | ( n8703 & n13132 ) ;
  assign n24984 = ( n5542 & ~n20607 ) | ( n5542 & n23199 ) | ( ~n20607 & n23199 ) ;
  assign n24985 = ( ~n4350 & n24983 ) | ( ~n4350 & n24984 ) | ( n24983 & n24984 ) ;
  assign n24986 = n24985 ^ n7217 ^ n5189 ;
  assign n24981 = ( ~n1694 & n2226 ) | ( ~n1694 & n10035 ) | ( n2226 & n10035 ) ;
  assign n24982 = n23860 | n24981 ;
  assign n24987 = n24986 ^ n24982 ^ 1'b0 ;
  assign n24988 = ( n8881 & ~n14495 ) | ( n8881 & n18472 ) | ( ~n14495 & n18472 ) ;
  assign n24989 = n24988 ^ n15725 ^ n4060 ;
  assign n24993 = n12588 ^ n4935 ^ n1077 ;
  assign n24990 = n17954 ^ n13987 ^ n1551 ;
  assign n24991 = n24990 ^ n7497 ^ 1'b0 ;
  assign n24992 = n9958 & ~n24991 ;
  assign n24994 = n24993 ^ n24992 ^ 1'b0 ;
  assign n24995 = ( ~n4508 & n10284 ) | ( ~n4508 & n24994 ) | ( n10284 & n24994 ) ;
  assign n24996 = ~n5271 & n6308 ;
  assign n24997 = n24996 ^ n19172 ^ 1'b0 ;
  assign n24998 = n11051 ^ n5115 ^ n3720 ;
  assign n24999 = n11280 & ~n24998 ;
  assign n25000 = n10118 ^ n4914 ^ 1'b0 ;
  assign n25001 = n14730 & n25000 ;
  assign n25002 = ( n4735 & n17180 ) | ( n4735 & ~n25001 ) | ( n17180 & ~n25001 ) ;
  assign n25003 = n4688 & ~n5071 ;
  assign n25004 = ( ~n3691 & n23673 ) | ( ~n3691 & n25003 ) | ( n23673 & n25003 ) ;
  assign n25005 = ( n2318 & ~n12580 ) | ( n2318 & n25004 ) | ( ~n12580 & n25004 ) ;
  assign n25006 = n17879 ^ n6603 ^ n1909 ;
  assign n25007 = n25006 ^ n16025 ^ n3034 ;
  assign n25008 = ( n3942 & n9369 ) | ( n3942 & n23353 ) | ( n9369 & n23353 ) ;
  assign n25013 = n19752 & ~n21537 ;
  assign n25011 = n23331 ^ n13780 ^ 1'b0 ;
  assign n25012 = n8400 | n25011 ;
  assign n25009 = n17290 ^ n12670 ^ n6426 ;
  assign n25010 = n25009 ^ n11961 ^ n1471 ;
  assign n25014 = n25013 ^ n25012 ^ n25010 ;
  assign n25016 = ( n651 & n6360 ) | ( n651 & n7707 ) | ( n6360 & n7707 ) ;
  assign n25015 = ( n3421 & n6027 ) | ( n3421 & n11359 ) | ( n6027 & n11359 ) ;
  assign n25017 = n25016 ^ n25015 ^ n14135 ;
  assign n25018 = n15656 ^ n15271 ^ n9216 ;
  assign n25019 = n493 | n4847 ;
  assign n25020 = n25019 ^ n15848 ^ n582 ;
  assign n25021 = n2569 & n16473 ;
  assign n25022 = ( ~n3859 & n25020 ) | ( ~n3859 & n25021 ) | ( n25020 & n25021 ) ;
  assign n25023 = n25022 ^ n20349 ^ n15648 ;
  assign n25024 = ( n17022 & n18461 ) | ( n17022 & ~n25023 ) | ( n18461 & ~n25023 ) ;
  assign n25025 = ( n3862 & ~n7114 ) | ( n3862 & n8369 ) | ( ~n7114 & n8369 ) ;
  assign n25026 = ( n1828 & ~n9013 ) | ( n1828 & n25025 ) | ( ~n9013 & n25025 ) ;
  assign n25027 = n265 & ~n1190 ;
  assign n25028 = n25026 & n25027 ;
  assign n25029 = n21528 ^ n5328 ^ 1'b0 ;
  assign n25030 = n17229 & n25029 ;
  assign n25031 = ( n278 & ~n2514 ) | ( n278 & n5178 ) | ( ~n2514 & n5178 ) ;
  assign n25032 = n25031 ^ n11083 ^ 1'b0 ;
  assign n25033 = ( ~n1698 & n8057 ) | ( ~n1698 & n25032 ) | ( n8057 & n25032 ) ;
  assign n25034 = ( n4145 & n13772 ) | ( n4145 & n19894 ) | ( n13772 & n19894 ) ;
  assign n25035 = n25034 ^ n7082 ^ n5136 ;
  assign n25036 = ( n4677 & n7374 ) | ( n4677 & ~n9624 ) | ( n7374 & ~n9624 ) ;
  assign n25037 = ( n4294 & n7320 ) | ( n4294 & n8642 ) | ( n7320 & n8642 ) ;
  assign n25038 = n25037 ^ n23157 ^ n11750 ;
  assign n25039 = n10927 | n25038 ;
  assign n25040 = n25039 ^ n7517 ^ 1'b0 ;
  assign n25041 = ( n10607 & ~n25036 ) | ( n10607 & n25040 ) | ( ~n25036 & n25040 ) ;
  assign n25042 = n3946 & n25041 ;
  assign n25043 = n25042 ^ x89 ^ 1'b0 ;
  assign n25044 = ( ~n6540 & n25035 ) | ( ~n6540 & n25043 ) | ( n25035 & n25043 ) ;
  assign n25045 = ( ~n25030 & n25033 ) | ( ~n25030 & n25044 ) | ( n25033 & n25044 ) ;
  assign n25046 = n8475 ^ n5257 ^ n2379 ;
  assign n25047 = n22200 ^ n4541 ^ 1'b0 ;
  assign n25048 = n25047 ^ n23096 ^ n5466 ;
  assign n25049 = ( n310 & ~n1919 ) | ( n310 & n13644 ) | ( ~n1919 & n13644 ) ;
  assign n25050 = n4781 & n14571 ;
  assign n25051 = ~n3467 & n25050 ;
  assign n25052 = ( n1659 & n25049 ) | ( n1659 & n25051 ) | ( n25049 & n25051 ) ;
  assign n25053 = ( n10291 & ~n16170 ) | ( n10291 & n25052 ) | ( ~n16170 & n25052 ) ;
  assign n25054 = n25053 ^ n7727 ^ n7526 ;
  assign n25055 = ~n3717 & n18431 ;
  assign n25056 = n12183 & n25055 ;
  assign n25058 = n21960 ^ n18253 ^ n9428 ;
  assign n25057 = ( n2629 & ~n14382 ) | ( n2629 & n17559 ) | ( ~n14382 & n17559 ) ;
  assign n25059 = n25058 ^ n25057 ^ n716 ;
  assign n25060 = n16220 ^ n1402 ^ 1'b0 ;
  assign n25061 = n25060 ^ n9467 ^ n7473 ;
  assign n25062 = n25061 ^ n24244 ^ n16836 ;
  assign n25063 = n20413 ^ n9732 ^ n3498 ;
  assign n25064 = ( n9132 & n14972 ) | ( n9132 & ~n22793 ) | ( n14972 & ~n22793 ) ;
  assign n25065 = ~n8513 & n25064 ;
  assign n25069 = n13006 & n23618 ;
  assign n25070 = n13364 | n25069 ;
  assign n25066 = n20917 ^ n10184 ^ n3906 ;
  assign n25067 = n25066 ^ n16774 ^ n12477 ;
  assign n25068 = n25067 ^ n24337 ^ n23465 ;
  assign n25071 = n25070 ^ n25068 ^ 1'b0 ;
  assign n25072 = n25071 ^ n23695 ^ n19526 ;
  assign n25073 = n16024 ^ n10394 ^ n3989 ;
  assign n25074 = n25073 ^ n23839 ^ n10139 ;
  assign n25075 = n25074 ^ n13809 ^ n13564 ;
  assign n25076 = n7806 & ~n7946 ;
  assign n25077 = n25075 & n25076 ;
  assign n25078 = ( n977 & n22778 ) | ( n977 & ~n24682 ) | ( n22778 & ~n24682 ) ;
  assign n25079 = ( ~n6232 & n9243 ) | ( ~n6232 & n14104 ) | ( n9243 & n14104 ) ;
  assign n25080 = ( ~n11168 & n19430 ) | ( ~n11168 & n25079 ) | ( n19430 & n25079 ) ;
  assign n25081 = ( n24230 & n25078 ) | ( n24230 & n25080 ) | ( n25078 & n25080 ) ;
  assign n25082 = n23471 ^ x2 ^ 1'b0 ;
  assign n25083 = n19717 | n25082 ;
  assign n25084 = n13132 ^ n1686 ^ 1'b0 ;
  assign n25086 = n6669 ^ n4746 ^ n3486 ;
  assign n25085 = ~n2903 & n6612 ;
  assign n25087 = n25086 ^ n25085 ^ 1'b0 ;
  assign n25088 = n25087 ^ n24978 ^ n725 ;
  assign n25089 = ( n7994 & ~n10518 ) | ( n7994 & n10755 ) | ( ~n10518 & n10755 ) ;
  assign n25090 = ( n7639 & n13063 ) | ( n7639 & ~n25089 ) | ( n13063 & ~n25089 ) ;
  assign n25091 = n7236 ^ n1272 ^ 1'b0 ;
  assign n25092 = n25091 ^ n6811 ^ 1'b0 ;
  assign n25093 = n8935 & ~n20430 ;
  assign n25094 = n25093 ^ n17703 ^ n11295 ;
  assign n25095 = n12200 & ~n12600 ;
  assign n25096 = ~n13681 & n25095 ;
  assign n25097 = ( n1533 & n16852 ) | ( n1533 & n25096 ) | ( n16852 & n25096 ) ;
  assign n25098 = ( n20665 & n25094 ) | ( n20665 & n25097 ) | ( n25094 & n25097 ) ;
  assign n25099 = n7906 & n9654 ;
  assign n25100 = n5053 ^ n1842 ^ n1587 ;
  assign n25101 = n4658 | n8805 ;
  assign n25102 = ( ~n7644 & n12668 ) | ( ~n7644 & n25101 ) | ( n12668 & n25101 ) ;
  assign n25103 = ~n3073 & n12852 ;
  assign n25104 = n24675 & n25103 ;
  assign n25105 = n25104 ^ n8825 ^ n8806 ;
  assign n25106 = ( n25100 & n25102 ) | ( n25100 & ~n25105 ) | ( n25102 & ~n25105 ) ;
  assign n25107 = ( n9368 & n10015 ) | ( n9368 & n17913 ) | ( n10015 & n17913 ) ;
  assign n25108 = ( ~n2615 & n6925 ) | ( ~n2615 & n13753 ) | ( n6925 & n13753 ) ;
  assign n25109 = n14238 ^ n1635 ^ 1'b0 ;
  assign n25110 = ~n19459 & n25109 ;
  assign n25111 = ( n14824 & n25108 ) | ( n14824 & n25110 ) | ( n25108 & n25110 ) ;
  assign n25116 = n1202 & ~n14026 ;
  assign n25117 = n25116 ^ n12397 ^ 1'b0 ;
  assign n25115 = n11231 ^ n7517 ^ n1758 ;
  assign n25118 = n25117 ^ n25115 ^ n12739 ;
  assign n25112 = ( n11159 & ~n15576 ) | ( n11159 & n20519 ) | ( ~n15576 & n20519 ) ;
  assign n25113 = ( ~n13108 & n23476 ) | ( ~n13108 & n25112 ) | ( n23476 & n25112 ) ;
  assign n25114 = ~n15351 & n25113 ;
  assign n25119 = n25118 ^ n25114 ^ 1'b0 ;
  assign n25120 = ( ~n1667 & n2769 ) | ( ~n1667 & n24931 ) | ( n2769 & n24931 ) ;
  assign n25121 = ~n2864 & n25120 ;
  assign n25122 = n25121 ^ n7634 ^ 1'b0 ;
  assign n25123 = ( x23 & ~n7338 ) | ( x23 & n10573 ) | ( ~n7338 & n10573 ) ;
  assign n25124 = n19910 ^ n4217 ^ n2215 ;
  assign n25125 = ( n742 & n15025 ) | ( n742 & ~n25124 ) | ( n15025 & ~n25124 ) ;
  assign n25126 = ( n17556 & n23940 ) | ( n17556 & n25125 ) | ( n23940 & n25125 ) ;
  assign n25127 = n21835 & ~n25126 ;
  assign n25128 = ( n15064 & ~n19962 ) | ( n15064 & n21955 ) | ( ~n19962 & n21955 ) ;
  assign n25129 = n25128 ^ n3661 ^ n3523 ;
  assign n25130 = ( n3637 & n6210 ) | ( n3637 & ~n10999 ) | ( n6210 & ~n10999 ) ;
  assign n25131 = n25130 ^ n3918 ^ n2665 ;
  assign n25132 = n23633 ^ n12045 ^ 1'b0 ;
  assign n25133 = n8998 | n25132 ;
  assign n25134 = n10341 & n12012 ;
  assign n25135 = n25134 ^ n21912 ^ n13745 ;
  assign n25136 = n879 & n25135 ;
  assign n25137 = n25133 & n25136 ;
  assign n25138 = ( n4578 & n17162 ) | ( n4578 & ~n25137 ) | ( n17162 & ~n25137 ) ;
  assign n25139 = n4161 & ~n9984 ;
  assign n25140 = n25139 ^ n3010 ^ 1'b0 ;
  assign n25141 = n25140 ^ n22665 ^ n19305 ;
  assign n25142 = ( n9763 & n11567 ) | ( n9763 & ~n16029 ) | ( n11567 & ~n16029 ) ;
  assign n25143 = ( n6846 & n19821 ) | ( n6846 & n23667 ) | ( n19821 & n23667 ) ;
  assign n25144 = ( n25141 & n25142 ) | ( n25141 & n25143 ) | ( n25142 & n25143 ) ;
  assign n25145 = ( n13694 & n15952 ) | ( n13694 & n16147 ) | ( n15952 & n16147 ) ;
  assign n25146 = n10631 ^ n5539 ^ 1'b0 ;
  assign n25147 = n9619 & n22441 ;
  assign n25148 = n25147 ^ n23505 ^ 1'b0 ;
  assign n25149 = n22622 ^ n21141 ^ 1'b0 ;
  assign n25150 = n25148 & n25149 ;
  assign n25151 = n22108 ^ n480 ^ 1'b0 ;
  assign n25152 = n21737 | n25151 ;
  assign n25153 = n25152 ^ n22515 ^ 1'b0 ;
  assign n25154 = n1826 | n8686 ;
  assign n25155 = n25154 ^ n3706 ^ 1'b0 ;
  assign n25157 = n1818 & n14322 ;
  assign n25156 = n7553 ^ n382 ^ 1'b0 ;
  assign n25158 = n25157 ^ n25156 ^ n15206 ;
  assign n25159 = n25158 ^ n4760 ^ 1'b0 ;
  assign n25160 = ~n5233 & n25159 ;
  assign n25161 = ( n20689 & n25155 ) | ( n20689 & ~n25160 ) | ( n25155 & ~n25160 ) ;
  assign n25162 = n5615 & ~n7104 ;
  assign n25163 = n25162 ^ n10191 ^ n9435 ;
  assign n25164 = n10350 & ~n21019 ;
  assign n25165 = n25164 ^ n8722 ^ 1'b0 ;
  assign n25166 = n19342 ^ n19099 ^ n16838 ;
  assign n25167 = ( n7232 & n25165 ) | ( n7232 & ~n25166 ) | ( n25165 & ~n25166 ) ;
  assign n25168 = n10011 ^ n4222 ^ n3547 ;
  assign n25169 = ~n18461 & n25168 ;
  assign n25170 = n4816 & n25169 ;
  assign n25171 = ( n2608 & ~n7896 ) | ( n2608 & n15646 ) | ( ~n7896 & n15646 ) ;
  assign n25172 = ( ~n4037 & n6119 ) | ( ~n4037 & n25171 ) | ( n6119 & n25171 ) ;
  assign n25173 = n1860 | n25172 ;
  assign n25174 = ( n680 & n3803 ) | ( n680 & n25173 ) | ( n3803 & n25173 ) ;
  assign n25175 = n20420 ^ n7377 ^ 1'b0 ;
  assign n25176 = n13593 ^ n10232 ^ x48 ;
  assign n25177 = ( ~n10031 & n14705 ) | ( ~n10031 & n25176 ) | ( n14705 & n25176 ) ;
  assign n25178 = ( n1238 & n18957 ) | ( n1238 & ~n20264 ) | ( n18957 & ~n20264 ) ;
  assign n25179 = n25178 ^ n16079 ^ n10843 ;
  assign n25180 = n25179 ^ n21050 ^ n2569 ;
  assign n25181 = ( ~n12842 & n14836 ) | ( ~n12842 & n25180 ) | ( n14836 & n25180 ) ;
  assign n25182 = n18393 & n21065 ;
  assign n25183 = n498 | n937 ;
  assign n25184 = n25183 ^ n13687 ^ 1'b0 ;
  assign n25185 = n4712 ^ n2646 ^ n1904 ;
  assign n25186 = ( n410 & ~n8684 ) | ( n410 & n25185 ) | ( ~n8684 & n25185 ) ;
  assign n25187 = n25186 ^ n24493 ^ n1973 ;
  assign n25188 = ~n4988 & n14463 ;
  assign n25189 = n25188 ^ x86 ^ 1'b0 ;
  assign n25190 = n18005 ^ n10444 ^ 1'b0 ;
  assign n25191 = n22620 ^ n3939 ^ n3679 ;
  assign n25192 = n25191 ^ n22232 ^ 1'b0 ;
  assign n25193 = ( n2050 & ~n18451 ) | ( n2050 & n25192 ) | ( ~n18451 & n25192 ) ;
  assign n25194 = n20337 | n25193 ;
  assign n25195 = ( ~n12438 & n19500 ) | ( ~n12438 & n24332 ) | ( n19500 & n24332 ) ;
  assign n25199 = n18053 ^ n17843 ^ n4100 ;
  assign n25196 = n1971 & n10304 ;
  assign n25197 = n3051 & n25196 ;
  assign n25198 = n25197 ^ n1937 ^ n1278 ;
  assign n25200 = n25199 ^ n25198 ^ n4877 ;
  assign n25201 = n25200 ^ n22095 ^ n2985 ;
  assign n25202 = n9518 ^ n1243 ^ n842 ;
  assign n25203 = n25202 ^ n24094 ^ n5408 ;
  assign n25204 = ( n4059 & ~n4629 ) | ( n4059 & n14888 ) | ( ~n4629 & n14888 ) ;
  assign n25205 = ( n3935 & ~n17109 ) | ( n3935 & n25204 ) | ( ~n17109 & n25204 ) ;
  assign n25206 = ( n8503 & n25203 ) | ( n8503 & n25205 ) | ( n25203 & n25205 ) ;
  assign n25208 = n4721 & n18123 ;
  assign n25209 = n25208 ^ n4173 ^ 1'b0 ;
  assign n25210 = n25209 ^ n23049 ^ n21662 ;
  assign n25207 = ~n502 & n7537 ;
  assign n25211 = n25210 ^ n25207 ^ 1'b0 ;
  assign n25212 = n25211 ^ n2059 ^ n1459 ;
  assign n25213 = n15621 ^ n6160 ^ n4049 ;
  assign n25214 = n17173 ^ n13851 ^ n1227 ;
  assign n25215 = n3004 & n25214 ;
  assign n25216 = ( n15296 & ~n25213 ) | ( n15296 & n25215 ) | ( ~n25213 & n25215 ) ;
  assign n25221 = n17727 ^ n13928 ^ n2874 ;
  assign n25220 = n1291 & n4266 ;
  assign n25222 = n25221 ^ n25220 ^ 1'b0 ;
  assign n25217 = n5775 | n15993 ;
  assign n25218 = n25217 ^ n17805 ^ n2125 ;
  assign n25219 = n17052 & n25218 ;
  assign n25223 = n25222 ^ n25219 ^ 1'b0 ;
  assign n25224 = ( ~n14481 & n24827 ) | ( ~n14481 & n25223 ) | ( n24827 & n25223 ) ;
  assign n25225 = n313 & ~n14701 ;
  assign n25226 = n4630 ^ n3771 ^ 1'b0 ;
  assign n25227 = n13948 ^ n6652 ^ n614 ;
  assign n25228 = ( n9217 & ~n13788 ) | ( n9217 & n25227 ) | ( ~n13788 & n25227 ) ;
  assign n25229 = n10735 | n25228 ;
  assign n25230 = ( n6178 & ~n25226 ) | ( n6178 & n25229 ) | ( ~n25226 & n25229 ) ;
  assign n25231 = ( n9543 & n21250 ) | ( n9543 & ~n25230 ) | ( n21250 & ~n25230 ) ;
  assign n25232 = ( n12243 & ~n23955 ) | ( n12243 & n25231 ) | ( ~n23955 & n25231 ) ;
  assign n25233 = ( ~n24021 & n25225 ) | ( ~n24021 & n25232 ) | ( n25225 & n25232 ) ;
  assign n25234 = n17841 ^ n8846 ^ 1'b0 ;
  assign n25235 = ( ~n16905 & n17556 ) | ( ~n16905 & n18589 ) | ( n17556 & n18589 ) ;
  assign n25236 = n15969 ^ x171 ^ 1'b0 ;
  assign n25237 = n25235 & ~n25236 ;
  assign n25238 = ( n1481 & n8384 ) | ( n1481 & ~n9665 ) | ( n8384 & ~n9665 ) ;
  assign n25239 = n18585 ^ n6724 ^ 1'b0 ;
  assign n25240 = n24694 | n25239 ;
  assign n25241 = n8990 | n15604 ;
  assign n25242 = n1161 | n25241 ;
  assign n25243 = n2027 | n24217 ;
  assign n25244 = n2919 & ~n24206 ;
  assign n25245 = ( n25242 & n25243 ) | ( n25242 & ~n25244 ) | ( n25243 & ~n25244 ) ;
  assign n25246 = n21109 ^ n12679 ^ 1'b0 ;
  assign n25247 = n14966 | n25246 ;
  assign n25248 = n25247 ^ n25168 ^ 1'b0 ;
  assign n25249 = n24896 ^ n18906 ^ n17633 ;
  assign n25250 = ( ~n4471 & n21450 ) | ( ~n4471 & n25249 ) | ( n21450 & n25249 ) ;
  assign n25251 = ( n14685 & n21117 ) | ( n14685 & ~n25250 ) | ( n21117 & ~n25250 ) ;
  assign n25254 = n680 | n2806 ;
  assign n25255 = n25254 ^ n17672 ^ 1'b0 ;
  assign n25252 = ( n14161 & n15411 ) | ( n14161 & ~n16469 ) | ( n15411 & ~n16469 ) ;
  assign n25253 = n2498 & ~n25252 ;
  assign n25256 = n25255 ^ n25253 ^ n7966 ;
  assign n25257 = n17802 ^ n5536 ^ n2477 ;
  assign n25258 = n13681 ^ n9374 ^ n7865 ;
  assign n25259 = ( n1561 & ~n4467 ) | ( n1561 & n9144 ) | ( ~n4467 & n9144 ) ;
  assign n25260 = ( n3894 & n5950 ) | ( n3894 & n25259 ) | ( n5950 & n25259 ) ;
  assign n25266 = n24076 ^ n21628 ^ n9231 ;
  assign n25261 = x103 & ~n468 ;
  assign n25262 = ~n1344 & n25261 ;
  assign n25263 = n24646 ^ n14903 ^ n10079 ;
  assign n25264 = n25262 | n25263 ;
  assign n25265 = n25264 ^ n22615 ^ 1'b0 ;
  assign n25267 = n25266 ^ n25265 ^ n10469 ;
  assign n25268 = ( ~n301 & n25260 ) | ( ~n301 & n25267 ) | ( n25260 & n25267 ) ;
  assign n25269 = ( ~n7483 & n11278 ) | ( ~n7483 & n18912 ) | ( n11278 & n18912 ) ;
  assign n25270 = ( n803 & n11484 ) | ( n803 & n25269 ) | ( n11484 & n25269 ) ;
  assign n25271 = ( ~n3223 & n6029 ) | ( ~n3223 & n9840 ) | ( n6029 & n9840 ) ;
  assign n25276 = n12737 | n20447 ;
  assign n25277 = n25276 ^ n21951 ^ n20180 ;
  assign n25275 = n16171 ^ n10253 ^ 1'b0 ;
  assign n25272 = n12025 ^ n11349 ^ n3739 ;
  assign n25273 = n25272 ^ n10067 ^ n7225 ;
  assign n25274 = n7787 & ~n25273 ;
  assign n25278 = n25277 ^ n25275 ^ n25274 ;
  assign n25279 = n7366 ^ n6696 ^ n2658 ;
  assign n25280 = n25279 ^ n375 ^ 1'b0 ;
  assign n25281 = n6928 & n25280 ;
  assign n25282 = ( n3724 & n12899 ) | ( n3724 & n16664 ) | ( n12899 & n16664 ) ;
  assign n25283 = n25244 ^ n14147 ^ n2003 ;
  assign n25284 = ( ~n4745 & n25282 ) | ( ~n4745 & n25283 ) | ( n25282 & n25283 ) ;
  assign n25287 = ( n2447 & n3685 ) | ( n2447 & ~n5463 ) | ( n3685 & ~n5463 ) ;
  assign n25285 = n2146 & n4784 ;
  assign n25286 = n25285 ^ n11263 ^ 1'b0 ;
  assign n25288 = n25287 ^ n25286 ^ n714 ;
  assign n25289 = ( ~x61 & n293 ) | ( ~x61 & n3855 ) | ( n293 & n3855 ) ;
  assign n25290 = ( n2954 & ~n10749 ) | ( n2954 & n25289 ) | ( ~n10749 & n25289 ) ;
  assign n25291 = n23848 ^ n5792 ^ x40 ;
  assign n25292 = n7589 ^ n2072 ^ 1'b0 ;
  assign n25293 = n2275 | n9708 ;
  assign n25294 = n25292 & ~n25293 ;
  assign n25295 = n25294 ^ n16836 ^ n7388 ;
  assign n25296 = ( ~n469 & n2405 ) | ( ~n469 & n6954 ) | ( n2405 & n6954 ) ;
  assign n25297 = n20049 ^ n9801 ^ n8945 ;
  assign n25298 = n25297 ^ n2492 ^ n875 ;
  assign n25299 = n13929 ^ n12304 ^ n5710 ;
  assign n25300 = n25299 ^ n21597 ^ n19647 ;
  assign n25301 = ~n25298 & n25300 ;
  assign n25302 = n25296 & n25301 ;
  assign n25303 = ( n1507 & n8588 ) | ( n1507 & n15227 ) | ( n8588 & n15227 ) ;
  assign n25304 = ( ~n602 & n4614 ) | ( ~n602 & n9164 ) | ( n4614 & n9164 ) ;
  assign n25305 = n25304 ^ n16102 ^ n5037 ;
  assign n25306 = n5946 & ~n18023 ;
  assign n25314 = n20295 ^ n10575 ^ n1830 ;
  assign n25307 = n12466 ^ n11356 ^ n6301 ;
  assign n25308 = n4396 & n25307 ;
  assign n25309 = n25308 ^ n1609 ^ 1'b0 ;
  assign n25310 = ~n13958 & n25309 ;
  assign n25311 = n9579 ^ n2501 ^ 1'b0 ;
  assign n25312 = n25310 & n25311 ;
  assign n25313 = ( n3592 & n9020 ) | ( n3592 & n25312 ) | ( n9020 & n25312 ) ;
  assign n25315 = n25314 ^ n25313 ^ 1'b0 ;
  assign n25316 = ( n1865 & n25306 ) | ( n1865 & ~n25315 ) | ( n25306 & ~n25315 ) ;
  assign n25317 = n25316 ^ n20034 ^ n17518 ;
  assign n25318 = ( n8473 & ~n25305 ) | ( n8473 & n25317 ) | ( ~n25305 & n25317 ) ;
  assign n25319 = ~n1376 & n5184 ;
  assign n25320 = ~n2154 & n25319 ;
  assign n25321 = n14573 ^ n9933 ^ 1'b0 ;
  assign n25322 = n25320 | n25321 ;
  assign n25329 = n24649 ^ n13680 ^ n12287 ;
  assign n25323 = n16634 ^ n4835 ^ n3388 ;
  assign n25324 = n7401 ^ n1939 ^ 1'b0 ;
  assign n25325 = n6345 & ~n25324 ;
  assign n25326 = ( n7986 & ~n9797 ) | ( n7986 & n25325 ) | ( ~n9797 & n25325 ) ;
  assign n25327 = ( n8500 & n21335 ) | ( n8500 & ~n25326 ) | ( n21335 & ~n25326 ) ;
  assign n25328 = n25323 & n25327 ;
  assign n25330 = n25329 ^ n25328 ^ 1'b0 ;
  assign n25331 = ( n5645 & ~n11665 ) | ( n5645 & n25330 ) | ( ~n11665 & n25330 ) ;
  assign n25332 = n1752 & ~n1822 ;
  assign n25333 = ~n7011 & n25332 ;
  assign n25334 = ~n6779 & n15342 ;
  assign n25335 = ~n17234 & n25334 ;
  assign n25336 = n7404 | n15199 ;
  assign n25337 = n23593 | n25336 ;
  assign n25338 = n25337 ^ n18680 ^ 1'b0 ;
  assign n25339 = n25338 ^ n1551 ^ 1'b0 ;
  assign n25345 = n9402 & ~n24243 ;
  assign n25346 = ~n1487 & n25345 ;
  assign n25344 = n21858 ^ n3443 ^ n3268 ;
  assign n25347 = n25346 ^ n25344 ^ n24619 ;
  assign n25348 = ( n8895 & ~n12624 ) | ( n8895 & n20085 ) | ( ~n12624 & n20085 ) ;
  assign n25349 = n25348 ^ n1712 ^ 1'b0 ;
  assign n25350 = ( ~n742 & n25347 ) | ( ~n742 & n25349 ) | ( n25347 & n25349 ) ;
  assign n25342 = n23962 ^ n18716 ^ n3898 ;
  assign n25341 = n8746 ^ n8188 ^ n4230 ;
  assign n25340 = n1172 ^ n1002 ^ 1'b0 ;
  assign n25343 = n25342 ^ n25341 ^ n25340 ;
  assign n25351 = n25350 ^ n25343 ^ n4223 ;
  assign n25352 = ( n707 & n14568 ) | ( n707 & n17404 ) | ( n14568 & n17404 ) ;
  assign n25353 = ( n1682 & n6844 ) | ( n1682 & n7394 ) | ( n6844 & n7394 ) ;
  assign n25354 = n25353 ^ n10368 ^ n1258 ;
  assign n25355 = n25354 ^ n7722 ^ n2457 ;
  assign n25356 = ( n20149 & n23194 ) | ( n20149 & n25355 ) | ( n23194 & n25355 ) ;
  assign n25357 = n11264 & n25356 ;
  assign n25358 = n25352 & n25357 ;
  assign n25359 = n25358 ^ n25118 ^ n8453 ;
  assign n25360 = ( n790 & n13250 ) | ( n790 & n14288 ) | ( n13250 & n14288 ) ;
  assign n25361 = ( n14694 & n22320 ) | ( n14694 & ~n25360 ) | ( n22320 & ~n25360 ) ;
  assign n25362 = ( n9404 & n13230 ) | ( n9404 & n14509 ) | ( n13230 & n14509 ) ;
  assign n25363 = n10134 ^ n5884 ^ n1703 ;
  assign n25364 = ( n1482 & ~n19729 ) | ( n1482 & n20826 ) | ( ~n19729 & n20826 ) ;
  assign n25365 = ( n1531 & n3922 ) | ( n1531 & ~n23871 ) | ( n3922 & ~n23871 ) ;
  assign n25366 = n25365 ^ n25168 ^ n10267 ;
  assign n25367 = ( n6396 & n7232 ) | ( n6396 & ~n23142 ) | ( n7232 & ~n23142 ) ;
  assign n25368 = n25367 ^ n7145 ^ n5463 ;
  assign n25369 = ( n5019 & ~n14221 ) | ( n5019 & n21867 ) | ( ~n14221 & n21867 ) ;
  assign n25370 = ~n25368 & n25369 ;
  assign n25371 = n23948 ^ n13109 ^ n10998 ;
  assign n25372 = ( n16988 & n21202 ) | ( n16988 & n25371 ) | ( n21202 & n25371 ) ;
  assign n25373 = n1635 & n6162 ;
  assign n25374 = ( n2331 & ~n15353 ) | ( n2331 & n25373 ) | ( ~n15353 & n25373 ) ;
  assign n25375 = n10688 ^ n7100 ^ 1'b0 ;
  assign n25376 = ~n4405 & n8778 ;
  assign n25377 = n25376 ^ n9121 ^ 1'b0 ;
  assign n25378 = n2303 ^ n1576 ^ n1410 ;
  assign n25379 = n4066 & n25378 ;
  assign n25380 = ( n4191 & ~n12652 ) | ( n4191 & n25379 ) | ( ~n12652 & n25379 ) ;
  assign n25381 = ( n25375 & n25377 ) | ( n25375 & n25380 ) | ( n25377 & n25380 ) ;
  assign n25382 = ( n511 & n18802 ) | ( n511 & ~n25381 ) | ( n18802 & ~n25381 ) ;
  assign n25383 = ( ~x245 & n299 ) | ( ~x245 & n7340 ) | ( n299 & n7340 ) ;
  assign n25384 = ( n2886 & ~n6771 ) | ( n2886 & n10957 ) | ( ~n6771 & n10957 ) ;
  assign n25385 = n25384 ^ n21161 ^ n771 ;
  assign n25386 = n10823 ^ n8210 ^ x213 ;
  assign n25387 = ( n2622 & n6512 ) | ( n2622 & ~n8426 ) | ( n6512 & ~n8426 ) ;
  assign n25388 = ( n430 & n2089 ) | ( n430 & n8713 ) | ( n2089 & n8713 ) ;
  assign n25389 = n5527 & n11895 ;
  assign n25390 = ~n25388 & n25389 ;
  assign n25391 = n25390 ^ n17449 ^ n16323 ;
  assign n25392 = n25391 ^ n11647 ^ n4938 ;
  assign n25393 = n21868 ^ n9561 ^ n2764 ;
  assign n25394 = x2 & ~n25393 ;
  assign n25395 = n25394 ^ n610 ^ 1'b0 ;
  assign n25396 = n25395 ^ n19133 ^ 1'b0 ;
  assign n25397 = n12749 | n25396 ;
  assign n25398 = n17097 ^ n15274 ^ n3236 ;
  assign n25399 = ( n567 & n2444 ) | ( n567 & n13924 ) | ( n2444 & n13924 ) ;
  assign n25400 = n25399 ^ n18029 ^ n4338 ;
  assign n25401 = ( n2917 & n3145 ) | ( n2917 & n25400 ) | ( n3145 & n25400 ) ;
  assign n25402 = ~n24137 & n25401 ;
  assign n25403 = ~n8617 & n25402 ;
  assign n25404 = ( n1410 & n3380 ) | ( n1410 & ~n25403 ) | ( n3380 & ~n25403 ) ;
  assign n25405 = ~n2974 & n4414 ;
  assign n25406 = n972 & n25405 ;
  assign n25407 = n23553 ^ n9829 ^ n749 ;
  assign n25408 = ( n4028 & ~n10548 ) | ( n4028 & n14698 ) | ( ~n10548 & n14698 ) ;
  assign n25409 = ( ~n25406 & n25407 ) | ( ~n25406 & n25408 ) | ( n25407 & n25408 ) ;
  assign n25410 = n20517 ^ n11391 ^ n4770 ;
  assign n25417 = n8223 ^ n4223 ^ n3428 ;
  assign n25416 = n19851 ^ n11056 ^ n3329 ;
  assign n25411 = n7463 | n16306 ;
  assign n25412 = n8191 & ~n10198 ;
  assign n25413 = n3941 & ~n5807 ;
  assign n25414 = ~n25412 & n25413 ;
  assign n25415 = ( n24319 & n25411 ) | ( n24319 & n25414 ) | ( n25411 & n25414 ) ;
  assign n25418 = n25417 ^ n25416 ^ n25415 ;
  assign n25419 = n11302 ^ n9914 ^ n9581 ;
  assign n25420 = ( ~x232 & n11920 ) | ( ~x232 & n25419 ) | ( n11920 & n25419 ) ;
  assign n25421 = n702 & n9763 ;
  assign n25422 = ( n11090 & n25348 ) | ( n11090 & ~n25421 ) | ( n25348 & ~n25421 ) ;
  assign n25423 = x56 & ~n25422 ;
  assign n25424 = n25420 & n25423 ;
  assign n25425 = n7793 ^ n7054 ^ 1'b0 ;
  assign n25426 = n25425 ^ n13627 ^ n2596 ;
  assign n25427 = n25426 ^ n7922 ^ n7716 ;
  assign n25428 = ( n667 & n6833 ) | ( n667 & ~n8364 ) | ( n6833 & ~n8364 ) ;
  assign n25429 = ( n1597 & n2779 ) | ( n1597 & n25428 ) | ( n2779 & n25428 ) ;
  assign n25430 = n25429 ^ n11182 ^ n475 ;
  assign n25432 = ~n3297 & n14411 ;
  assign n25433 = n25432 ^ n24492 ^ 1'b0 ;
  assign n25431 = n2324 & n17787 ;
  assign n25434 = n25433 ^ n25431 ^ 1'b0 ;
  assign n25435 = ( n4109 & n9454 ) | ( n4109 & n19226 ) | ( n9454 & n19226 ) ;
  assign n25436 = n25435 ^ n22587 ^ n3451 ;
  assign n25437 = n8100 ^ n282 ^ x23 ;
  assign n25438 = n25437 ^ n9758 ^ n3188 ;
  assign n25439 = n25438 ^ n14378 ^ n5273 ;
  assign n25440 = n25439 ^ n18086 ^ n1545 ;
  assign n25441 = ( n10845 & n11961 ) | ( n10845 & n19625 ) | ( n11961 & n19625 ) ;
  assign n25442 = n25441 ^ n12675 ^ n9950 ;
  assign n25443 = ( n4412 & n10437 ) | ( n4412 & ~n25442 ) | ( n10437 & ~n25442 ) ;
  assign n25444 = n25443 ^ n20902 ^ n4864 ;
  assign n25445 = ( n803 & ~n3604 ) | ( n803 & n15587 ) | ( ~n3604 & n15587 ) ;
  assign n25446 = n10225 & n16089 ;
  assign n25447 = n15811 & n25446 ;
  assign n25448 = n25447 ^ n10335 ^ 1'b0 ;
  assign n25449 = ( ~n19390 & n25445 ) | ( ~n19390 & n25448 ) | ( n25445 & n25448 ) ;
  assign n25450 = n13114 ^ n6762 ^ n5337 ;
  assign n25451 = n4158 & n13385 ;
  assign n25452 = n25450 & n25451 ;
  assign n25453 = n14041 ^ n7385 ^ n3058 ;
  assign n25454 = ~n13724 & n25453 ;
  assign n25455 = n629 & ~n18671 ;
  assign n25456 = n25455 ^ n19118 ^ 1'b0 ;
  assign n25457 = ( n25452 & ~n25454 ) | ( n25452 & n25456 ) | ( ~n25454 & n25456 ) ;
  assign n25458 = n25239 ^ n1779 ^ 1'b0 ;
  assign n25459 = n21188 & n25458 ;
  assign n25460 = ( ~n1371 & n7447 ) | ( ~n1371 & n25459 ) | ( n7447 & n25459 ) ;
  assign n25461 = ~n10572 & n18963 ;
  assign n25462 = ( ~n572 & n6609 ) | ( ~n572 & n25461 ) | ( n6609 & n25461 ) ;
  assign n25467 = ( ~n2865 & n3902 ) | ( ~n2865 & n4898 ) | ( n3902 & n4898 ) ;
  assign n25468 = n25467 ^ n11414 ^ n9697 ;
  assign n25466 = n24388 ^ n6324 ^ n2946 ;
  assign n25463 = n4190 ^ n3055 ^ n2223 ;
  assign n25464 = ( n2440 & n15159 ) | ( n2440 & n25463 ) | ( n15159 & n25463 ) ;
  assign n25465 = n25464 ^ n16738 ^ n13592 ;
  assign n25469 = n25468 ^ n25466 ^ n25465 ;
  assign n25470 = ( n24555 & n25462 ) | ( n24555 & ~n25469 ) | ( n25462 & ~n25469 ) ;
  assign n25473 = n11899 ^ n4011 ^ n824 ;
  assign n25472 = ( n2153 & n11427 ) | ( n2153 & n12643 ) | ( n11427 & n12643 ) ;
  assign n25471 = ( ~n1557 & n21746 ) | ( ~n1557 & n23600 ) | ( n21746 & n23600 ) ;
  assign n25474 = n25473 ^ n25472 ^ n25471 ;
  assign n25475 = ( n390 & ~n11593 ) | ( n390 & n25474 ) | ( ~n11593 & n25474 ) ;
  assign n25476 = n25475 ^ n22932 ^ n2140 ;
  assign n25477 = n4309 & ~n4459 ;
  assign n25478 = n3581 & n25477 ;
  assign n25479 = n10202 | n24096 ;
  assign n25480 = n25478 & ~n25479 ;
  assign n25481 = n635 | n16336 ;
  assign n25482 = n25481 ^ n5721 ^ 1'b0 ;
  assign n25483 = n6936 ^ n2836 ^ n907 ;
  assign n25484 = n21899 ^ n18841 ^ n10626 ;
  assign n25485 = n12207 & ~n17370 ;
  assign n25486 = n17021 & n25485 ;
  assign n25487 = n17253 | n24212 ;
  assign n25488 = ( ~n4281 & n25486 ) | ( ~n4281 & n25487 ) | ( n25486 & n25487 ) ;
  assign n25489 = n23087 ^ n9773 ^ n8796 ;
  assign n25490 = ( n9549 & ~n10316 ) | ( n9549 & n18730 ) | ( ~n10316 & n18730 ) ;
  assign n25491 = n2403 & n11849 ;
  assign n25492 = ( ~n13548 & n25490 ) | ( ~n13548 & n25491 ) | ( n25490 & n25491 ) ;
  assign n25493 = n9970 ^ n5880 ^ n1571 ;
  assign n25494 = n25493 ^ n24806 ^ n16225 ;
  assign n25495 = n21213 ^ n16044 ^ n7849 ;
  assign n25496 = n25495 ^ n8282 ^ n3177 ;
  assign n25497 = n25496 ^ n1131 ^ 1'b0 ;
  assign n25498 = n10697 | n18113 ;
  assign n25499 = ( ~n2202 & n22319 ) | ( ~n2202 & n25498 ) | ( n22319 & n25498 ) ;
  assign n25500 = ( ~n4395 & n17028 ) | ( ~n4395 & n25499 ) | ( n17028 & n25499 ) ;
  assign n25501 = n23730 | n25500 ;
  assign n25502 = n25501 ^ n635 ^ 1'b0 ;
  assign n25503 = n9135 ^ n6564 ^ 1'b0 ;
  assign n25504 = n11134 ^ n6523 ^ n4877 ;
  assign n25505 = ( ~n9220 & n13391 ) | ( ~n9220 & n25504 ) | ( n13391 & n25504 ) ;
  assign n25512 = n23340 ^ n21455 ^ 1'b0 ;
  assign n25506 = n1186 | n5110 ;
  assign n25507 = n25506 ^ n4853 ^ 1'b0 ;
  assign n25508 = n15407 & ~n25507 ;
  assign n25509 = n21941 ^ n12232 ^ 1'b0 ;
  assign n25510 = n25508 & ~n25509 ;
  assign n25511 = n12181 & n25510 ;
  assign n25513 = n25512 ^ n25511 ^ 1'b0 ;
  assign n25516 = n13266 ^ n8882 ^ n1723 ;
  assign n25514 = ( n5997 & n8881 ) | ( n5997 & ~n9676 ) | ( n8881 & ~n9676 ) ;
  assign n25515 = ( n14494 & ~n18026 ) | ( n14494 & n25514 ) | ( ~n18026 & n25514 ) ;
  assign n25517 = n25516 ^ n25515 ^ x202 ;
  assign n25518 = n14669 ^ n2046 ^ 1'b0 ;
  assign n25519 = n25518 ^ n21606 ^ n14752 ;
  assign n25520 = ( ~n6204 & n13017 ) | ( ~n6204 & n21146 ) | ( n13017 & n21146 ) ;
  assign n25521 = ( n8240 & n10212 ) | ( n8240 & n14113 ) | ( n10212 & n14113 ) ;
  assign n25522 = n23669 ^ n4132 ^ 1'b0 ;
  assign n25523 = n25521 & n25522 ;
  assign n25525 = ( n3105 & n3281 ) | ( n3105 & ~n6842 ) | ( n3281 & ~n6842 ) ;
  assign n25524 = n14209 ^ n2405 ^ 1'b0 ;
  assign n25526 = n25525 ^ n25524 ^ n12619 ;
  assign n25534 = n24078 ^ n12309 ^ n5048 ;
  assign n25532 = ( ~n2575 & n3102 ) | ( ~n2575 & n9270 ) | ( n3102 & n9270 ) ;
  assign n25528 = n1773 & ~n10744 ;
  assign n25529 = n21455 & n25528 ;
  assign n25527 = n19511 ^ n9416 ^ n721 ;
  assign n25530 = n25529 ^ n25527 ^ n5185 ;
  assign n25531 = ~n23290 & n25530 ;
  assign n25533 = n25532 ^ n25531 ^ 1'b0 ;
  assign n25535 = n25534 ^ n25533 ^ n5284 ;
  assign n25536 = ~n16907 & n22637 ;
  assign n25537 = ( n1597 & n23162 ) | ( n1597 & ~n23785 ) | ( n23162 & ~n23785 ) ;
  assign n25538 = n25537 ^ n12760 ^ n1338 ;
  assign n25539 = n25538 ^ n11922 ^ 1'b0 ;
  assign n25540 = n12153 ^ n7708 ^ n1616 ;
  assign n25541 = ( n10737 & n12628 ) | ( n10737 & n25540 ) | ( n12628 & n25540 ) ;
  assign n25542 = n16308 ^ n648 ^ 1'b0 ;
  assign n25543 = ~n14722 & n25542 ;
  assign n25544 = ( ~n12468 & n25541 ) | ( ~n12468 & n25543 ) | ( n25541 & n25543 ) ;
  assign n25551 = n1202 ^ x239 ^ 1'b0 ;
  assign n25552 = n402 & n25551 ;
  assign n25547 = x38 & ~n3588 ;
  assign n25548 = n3487 | n25547 ;
  assign n25549 = n25548 ^ n1958 ^ 1'b0 ;
  assign n25550 = n1361 & ~n25549 ;
  assign n25553 = n25552 ^ n25550 ^ 1'b0 ;
  assign n25546 = ( n1390 & n2492 ) | ( n1390 & n8678 ) | ( n2492 & n8678 ) ;
  assign n25545 = ( n2698 & n13297 ) | ( n2698 & n22895 ) | ( n13297 & n22895 ) ;
  assign n25554 = n25553 ^ n25546 ^ n25545 ;
  assign n25555 = ( ~n6832 & n6971 ) | ( ~n6832 & n17513 ) | ( n6971 & n17513 ) ;
  assign n25556 = ( n2553 & ~n10663 ) | ( n2553 & n25555 ) | ( ~n10663 & n25555 ) ;
  assign n25557 = ( ~n2557 & n13344 ) | ( ~n2557 & n25556 ) | ( n13344 & n25556 ) ;
  assign n25558 = n25557 ^ n21919 ^ n3160 ;
  assign n25559 = n10215 ^ n7272 ^ n6630 ;
  assign n25560 = n5862 & ~n25559 ;
  assign n25561 = ~n14863 & n25560 ;
  assign n25565 = n18697 ^ n1382 ^ 1'b0 ;
  assign n25562 = n8657 ^ n5283 ^ 1'b0 ;
  assign n25563 = n19336 & n25562 ;
  assign n25564 = ~n16382 & n25563 ;
  assign n25566 = n25565 ^ n25564 ^ 1'b0 ;
  assign n25567 = ( n2074 & ~n4488 ) | ( n2074 & n13312 ) | ( ~n4488 & n13312 ) ;
  assign n25568 = ( n25561 & ~n25566 ) | ( n25561 & n25567 ) | ( ~n25566 & n25567 ) ;
  assign n25569 = n7240 ^ n4726 ^ n710 ;
  assign n25570 = ( n16634 & ~n19297 ) | ( n16634 & n25569 ) | ( ~n19297 & n25569 ) ;
  assign n25571 = n2362 & ~n13452 ;
  assign n25572 = n1180 & n25571 ;
  assign n25573 = ( n4529 & n6975 ) | ( n4529 & ~n15923 ) | ( n6975 & ~n15923 ) ;
  assign n25574 = ( ~n5012 & n5353 ) | ( ~n5012 & n25573 ) | ( n5353 & n25573 ) ;
  assign n25575 = ~n25572 & n25574 ;
  assign n25576 = ( n2445 & n6113 ) | ( n2445 & ~n15749 ) | ( n6113 & ~n15749 ) ;
  assign n25577 = n25576 ^ n5346 ^ n3369 ;
  assign n25578 = n8985 ^ n3990 ^ n1765 ;
  assign n25579 = ( n5625 & ~n25577 ) | ( n5625 & n25578 ) | ( ~n25577 & n25578 ) ;
  assign n25580 = ~n4219 & n15900 ;
  assign n25581 = ~n25579 & n25580 ;
  assign n25582 = n5336 | n25581 ;
  assign n25583 = n25575 | n25582 ;
  assign n25584 = ( ~n4868 & n11050 ) | ( ~n4868 & n23750 ) | ( n11050 & n23750 ) ;
  assign n25585 = n6342 ^ n348 ^ 1'b0 ;
  assign n25586 = n713 & ~n25585 ;
  assign n25587 = ( n6503 & ~n8350 ) | ( n6503 & n25586 ) | ( ~n8350 & n25586 ) ;
  assign n25588 = ( ~n12907 & n18753 ) | ( ~n12907 & n25587 ) | ( n18753 & n25587 ) ;
  assign n25589 = n25588 ^ n10209 ^ n7681 ;
  assign n25592 = ( n14325 & n15344 ) | ( n14325 & n18672 ) | ( n15344 & n18672 ) ;
  assign n25590 = ( n18026 & ~n20505 ) | ( n18026 & n22744 ) | ( ~n20505 & n22744 ) ;
  assign n25591 = n25590 ^ n10384 ^ 1'b0 ;
  assign n25593 = n25592 ^ n25591 ^ n20997 ;
  assign n25594 = n21541 ^ n11382 ^ n10595 ;
  assign n25595 = n17863 ^ n2258 ^ 1'b0 ;
  assign n25596 = n25595 ^ n12589 ^ n7319 ;
  assign n25597 = ( ~n14478 & n14513 ) | ( ~n14478 & n18263 ) | ( n14513 & n18263 ) ;
  assign n25598 = ( n18335 & ~n25596 ) | ( n18335 & n25597 ) | ( ~n25596 & n25597 ) ;
  assign n25599 = n10556 ^ n4728 ^ n2671 ;
  assign n25600 = n25599 ^ n16082 ^ n1504 ;
  assign n25601 = n25600 ^ n17851 ^ n12490 ;
  assign n25602 = n25601 ^ n16699 ^ 1'b0 ;
  assign n25603 = n4164 ^ n2839 ^ 1'b0 ;
  assign n25604 = n11371 | n25603 ;
  assign n25605 = n25604 ^ n13826 ^ n2433 ;
  assign n25606 = n17044 & n18738 ;
  assign n25607 = ~n17333 & n25606 ;
  assign n25608 = ~n301 & n5312 ;
  assign n25609 = n25608 ^ n11033 ^ n901 ;
  assign n25610 = n25609 ^ n12506 ^ 1'b0 ;
  assign n25611 = n14257 ^ n7983 ^ 1'b0 ;
  assign n25612 = n25611 ^ n12694 ^ 1'b0 ;
  assign n25613 = n10705 & n25612 ;
  assign n25614 = ( ~n4732 & n17018 ) | ( ~n4732 & n25613 ) | ( n17018 & n25613 ) ;
  assign n25615 = ( n13847 & n13848 ) | ( n13847 & ~n25614 ) | ( n13848 & ~n25614 ) ;
  assign n25616 = ( n1372 & n10487 ) | ( n1372 & n14125 ) | ( n10487 & n14125 ) ;
  assign n25617 = n16125 ^ n9581 ^ 1'b0 ;
  assign n25618 = ( ~n814 & n16466 ) | ( ~n814 & n25617 ) | ( n16466 & n25617 ) ;
  assign n25619 = ( n14763 & n25616 ) | ( n14763 & ~n25618 ) | ( n25616 & ~n25618 ) ;
  assign n25620 = n25619 ^ n2100 ^ 1'b0 ;
  assign n25621 = ( n9881 & ~n19019 ) | ( n9881 & n19062 ) | ( ~n19019 & n19062 ) ;
  assign n25622 = n8617 & ~n15741 ;
  assign n25623 = n10175 & n25622 ;
  assign n25625 = n12135 ^ n7086 ^ n1308 ;
  assign n25624 = n4075 ^ n339 ^ x165 ;
  assign n25626 = n25625 ^ n25624 ^ n11362 ;
  assign n25627 = ( n10064 & n25623 ) | ( n10064 & ~n25626 ) | ( n25623 & ~n25626 ) ;
  assign n25628 = n25627 ^ n19544 ^ n17843 ;
  assign n25629 = ( ~n7331 & n17778 ) | ( ~n7331 & n25628 ) | ( n17778 & n25628 ) ;
  assign n25630 = n8166 ^ n6031 ^ n1136 ;
  assign n25631 = n25630 ^ n2744 ^ n1532 ;
  assign n25632 = n6800 | n21765 ;
  assign n25633 = n12523 & ~n19549 ;
  assign n25634 = ( n9133 & n25632 ) | ( n9133 & ~n25633 ) | ( n25632 & ~n25633 ) ;
  assign n25635 = ( n334 & ~n15122 ) | ( n334 & n18539 ) | ( ~n15122 & n18539 ) ;
  assign n25636 = ( n8704 & ~n19713 ) | ( n8704 & n25635 ) | ( ~n19713 & n25635 ) ;
  assign n25637 = ( ~n7396 & n15248 ) | ( ~n7396 & n16048 ) | ( n15248 & n16048 ) ;
  assign n25638 = n25637 ^ n24689 ^ n5962 ;
  assign n25639 = ( n3363 & ~n11993 ) | ( n3363 & n16367 ) | ( ~n11993 & n16367 ) ;
  assign n25640 = ( ~n1652 & n10002 ) | ( ~n1652 & n25639 ) | ( n10002 & n25639 ) ;
  assign n25641 = ( n6723 & ~n10816 ) | ( n6723 & n19774 ) | ( ~n10816 & n19774 ) ;
  assign n25642 = n260 | n5516 ;
  assign n25643 = n15007 | n25642 ;
  assign n25644 = n25643 ^ n10341 ^ n4597 ;
  assign n25645 = n25644 ^ n9890 ^ 1'b0 ;
  assign n25646 = n941 & ~n12056 ;
  assign n25647 = n11698 ^ n8901 ^ 1'b0 ;
  assign n25648 = ( n9619 & ~n25646 ) | ( n9619 & n25647 ) | ( ~n25646 & n25647 ) ;
  assign n25649 = n25648 ^ n7182 ^ 1'b0 ;
  assign n25650 = n4018 ^ n2026 ^ n651 ;
  assign n25651 = ( n18828 & n24243 ) | ( n18828 & ~n25650 ) | ( n24243 & ~n25650 ) ;
  assign n25652 = ( n347 & ~n20435 ) | ( n347 & n25651 ) | ( ~n20435 & n25651 ) ;
  assign n25653 = ( ~n17984 & n25649 ) | ( ~n17984 & n25652 ) | ( n25649 & n25652 ) ;
  assign n25654 = ( n2681 & n7550 ) | ( n2681 & ~n19486 ) | ( n7550 & ~n19486 ) ;
  assign n25655 = n25654 ^ n8773 ^ 1'b0 ;
  assign n25656 = ~x23 & n25655 ;
  assign n25657 = n19454 ^ n15565 ^ n8348 ;
  assign n25658 = n25657 ^ n2194 ^ n1562 ;
  assign n25659 = n10252 ^ n9081 ^ n6473 ;
  assign n25660 = n17568 ^ n7819 ^ 1'b0 ;
  assign n25661 = ( ~n2323 & n5757 ) | ( ~n2323 & n25660 ) | ( n5757 & n25660 ) ;
  assign n25662 = n25661 ^ n24846 ^ n16225 ;
  assign n25663 = ( n16326 & ~n19332 ) | ( n16326 & n25662 ) | ( ~n19332 & n25662 ) ;
  assign n25667 = ( n15505 & n20472 ) | ( n15505 & n23115 ) | ( n20472 & n23115 ) ;
  assign n25664 = n1188 & ~n20383 ;
  assign n25665 = n25664 ^ n14066 ^ 1'b0 ;
  assign n25666 = n7571 | n25665 ;
  assign n25668 = n25667 ^ n25666 ^ 1'b0 ;
  assign n25674 = ( n7109 & n7775 ) | ( n7109 & ~n25031 ) | ( n7775 & ~n25031 ) ;
  assign n25669 = ~n3172 & n23927 ;
  assign n25670 = n25669 ^ n10249 ^ 1'b0 ;
  assign n25671 = n19181 ^ n8408 ^ 1'b0 ;
  assign n25672 = n25670 & n25671 ;
  assign n25673 = n25672 ^ n956 ^ n918 ;
  assign n25675 = n25674 ^ n25673 ^ n3687 ;
  assign n25676 = n19152 ^ n17074 ^ 1'b0 ;
  assign n25677 = ( n16131 & n19417 ) | ( n16131 & ~n25676 ) | ( n19417 & ~n25676 ) ;
  assign n25678 = ( n3390 & ~n3727 ) | ( n3390 & n3835 ) | ( ~n3727 & n3835 ) ;
  assign n25679 = ( n3290 & ~n4005 ) | ( n3290 & n19306 ) | ( ~n4005 & n19306 ) ;
  assign n25680 = ( n737 & n905 ) | ( n737 & ~n4252 ) | ( n905 & ~n4252 ) ;
  assign n25681 = ( ~n14239 & n17232 ) | ( ~n14239 & n25680 ) | ( n17232 & n25680 ) ;
  assign n25682 = n25679 & ~n25681 ;
  assign n25683 = n6064 | n9414 ;
  assign n25684 = n25683 ^ n5787 ^ 1'b0 ;
  assign n25685 = ( n6214 & n11191 ) | ( n6214 & ~n25684 ) | ( n11191 & ~n25684 ) ;
  assign n25686 = ~n25682 & n25685 ;
  assign n25687 = n25686 ^ n16995 ^ 1'b0 ;
  assign n25688 = ( n2063 & ~n8684 ) | ( n2063 & n17841 ) | ( ~n8684 & n17841 ) ;
  assign n25689 = n25688 ^ n4340 ^ 1'b0 ;
  assign n25691 = n11885 ^ n11348 ^ n7408 ;
  assign n25690 = n15784 & ~n18129 ;
  assign n25692 = n25691 ^ n25690 ^ n3470 ;
  assign n25693 = n18802 ^ n11769 ^ n6706 ;
  assign n25694 = n25693 ^ n15711 ^ n9310 ;
  assign n25695 = ( ~n7103 & n23066 ) | ( ~n7103 & n25694 ) | ( n23066 & n25694 ) ;
  assign n25696 = n4590 & ~n10082 ;
  assign n25697 = n25696 ^ n11135 ^ n6260 ;
  assign n25704 = n12449 ^ n11832 ^ n11059 ;
  assign n25705 = n25704 ^ n15255 ^ n8867 ;
  assign n25698 = n24124 ^ n10007 ^ n3913 ;
  assign n25699 = ( n1384 & n15370 ) | ( n1384 & n25698 ) | ( n15370 & n25698 ) ;
  assign n25700 = n11679 & n25699 ;
  assign n25701 = n25700 ^ n16714 ^ n6061 ;
  assign n25702 = ( n3157 & n17627 ) | ( n3157 & n25701 ) | ( n17627 & n25701 ) ;
  assign n25703 = n8223 | n25702 ;
  assign n25706 = n25705 ^ n25703 ^ 1'b0 ;
  assign n25707 = ( ~n4071 & n5697 ) | ( ~n4071 & n8935 ) | ( n5697 & n8935 ) ;
  assign n25708 = n25707 ^ n8167 ^ n3428 ;
  assign n25709 = n1738 & n25708 ;
  assign n25710 = ( n1569 & n3962 ) | ( n1569 & ~n25709 ) | ( n3962 & ~n25709 ) ;
  assign n25711 = ( n8519 & n11612 ) | ( n8519 & ~n24140 ) | ( n11612 & ~n24140 ) ;
  assign n25713 = n5752 ^ n593 ^ 1'b0 ;
  assign n25716 = ( n1581 & n3266 ) | ( n1581 & ~n6330 ) | ( n3266 & ~n6330 ) ;
  assign n25714 = n5963 ^ n3557 ^ n559 ;
  assign n25715 = n25714 ^ n14004 ^ n2887 ;
  assign n25717 = n25716 ^ n25715 ^ 1'b0 ;
  assign n25718 = n25713 | n25717 ;
  assign n25712 = n4677 & ~n15896 ;
  assign n25719 = n25718 ^ n25712 ^ 1'b0 ;
  assign n25720 = ~n24507 & n25719 ;
  assign n25721 = n15253 & n25720 ;
  assign n25722 = n25711 & n25721 ;
  assign n25723 = n18499 & ~n21469 ;
  assign n25724 = n18863 ^ n13960 ^ n2499 ;
  assign n25725 = n15122 ^ n6970 ^ n3176 ;
  assign n25726 = n25725 ^ n7965 ^ 1'b0 ;
  assign n25727 = ( n4753 & ~n12531 ) | ( n4753 & n25726 ) | ( ~n12531 & n25726 ) ;
  assign n25728 = ( n1864 & n25724 ) | ( n1864 & ~n25727 ) | ( n25724 & ~n25727 ) ;
  assign n25729 = n17153 ^ n10835 ^ n10123 ;
  assign n25730 = n25729 ^ n19656 ^ n7124 ;
  assign n25731 = ( ~n21319 & n23875 ) | ( ~n21319 & n25730 ) | ( n23875 & n25730 ) ;
  assign n25732 = n21310 ^ n14752 ^ 1'b0 ;
  assign n25733 = ~n16178 & n25732 ;
  assign n25734 = ( n4836 & n15242 ) | ( n4836 & ~n21086 ) | ( n15242 & ~n21086 ) ;
  assign n25735 = n25734 ^ n20287 ^ n5578 ;
  assign n25736 = ( n5861 & n22590 ) | ( n5861 & ~n25735 ) | ( n22590 & ~n25735 ) ;
  assign n25739 = n10977 ^ n5542 ^ n4932 ;
  assign n25738 = n2206 | n20811 ;
  assign n25740 = n25739 ^ n25738 ^ 1'b0 ;
  assign n25737 = ( n2688 & ~n2840 ) | ( n2688 & n16611 ) | ( ~n2840 & n16611 ) ;
  assign n25741 = n25740 ^ n25737 ^ n10755 ;
  assign n25742 = n18029 ^ n9029 ^ 1'b0 ;
  assign n25743 = ( n2191 & n11338 ) | ( n2191 & n12071 ) | ( n11338 & n12071 ) ;
  assign n25744 = x77 & ~n24805 ;
  assign n25745 = n2883 & n25744 ;
  assign n25746 = n25745 ^ n13694 ^ n4809 ;
  assign n25747 = ~n5933 & n20810 ;
  assign n25748 = ( ~n23183 & n25746 ) | ( ~n23183 & n25747 ) | ( n25746 & n25747 ) ;
  assign n25749 = ( n3593 & n5103 ) | ( n3593 & ~n9372 ) | ( n5103 & ~n9372 ) ;
  assign n25750 = ( x113 & n16928 ) | ( x113 & ~n25749 ) | ( n16928 & ~n25749 ) ;
  assign n25751 = ~n12787 & n18346 ;
  assign n25752 = ~n25750 & n25751 ;
  assign n25753 = n12076 ^ n8316 ^ n6747 ;
  assign n25754 = ( n7979 & n9473 ) | ( n7979 & n21215 ) | ( n9473 & n21215 ) ;
  assign n25755 = n20811 ^ n11210 ^ n4195 ;
  assign n25756 = n12412 ^ n5675 ^ 1'b0 ;
  assign n25757 = n9148 | n25756 ;
  assign n25758 = ( ~n17166 & n25755 ) | ( ~n17166 & n25757 ) | ( n25755 & n25757 ) ;
  assign n25760 = ( n3624 & ~n19783 ) | ( n3624 & n22077 ) | ( ~n19783 & n22077 ) ;
  assign n25759 = ( n5332 & n5369 ) | ( n5332 & ~n11909 ) | ( n5369 & ~n11909 ) ;
  assign n25761 = n25760 ^ n25759 ^ n11270 ;
  assign n25762 = n25761 ^ n24929 ^ n21649 ;
  assign n25763 = ( ~n2052 & n15164 ) | ( ~n2052 & n25762 ) | ( n15164 & n25762 ) ;
  assign n25766 = n536 & n1886 ;
  assign n25765 = n2393 | n13595 ;
  assign n25764 = ( ~n5685 & n10494 ) | ( ~n5685 & n13939 ) | ( n10494 & n13939 ) ;
  assign n25767 = n25766 ^ n25765 ^ n25764 ;
  assign n25769 = n4747 ^ n2171 ^ 1'b0 ;
  assign n25768 = ~n4681 & n11825 ;
  assign n25770 = n25769 ^ n25768 ^ 1'b0 ;
  assign n25771 = n19226 ^ n13580 ^ n1686 ;
  assign n25772 = n25771 ^ n13403 ^ n12965 ;
  assign n25773 = n25772 ^ n16411 ^ 1'b0 ;
  assign n25774 = n25770 | n25773 ;
  assign n25775 = n25774 ^ n7711 ^ n7662 ;
  assign n25776 = ( n4281 & ~n18265 ) | ( n4281 & n21691 ) | ( ~n18265 & n21691 ) ;
  assign n25777 = ( n5648 & n5834 ) | ( n5648 & ~n17723 ) | ( n5834 & ~n17723 ) ;
  assign n25778 = n1756 & n8948 ;
  assign n25779 = ( n10417 & n25777 ) | ( n10417 & ~n25778 ) | ( n25777 & ~n25778 ) ;
  assign n25780 = n25779 ^ n17631 ^ n576 ;
  assign n25781 = ( n761 & ~n5098 ) | ( n761 & n13833 ) | ( ~n5098 & n13833 ) ;
  assign n25782 = ( n7393 & n9347 ) | ( n7393 & n25781 ) | ( n9347 & n25781 ) ;
  assign n25783 = n16984 ^ n1056 ^ 1'b0 ;
  assign n25784 = ( n7578 & n11324 ) | ( n7578 & ~n25783 ) | ( n11324 & ~n25783 ) ;
  assign n25786 = n12363 ^ n5975 ^ n5691 ;
  assign n25785 = n25305 ^ n13904 ^ x174 ;
  assign n25787 = n25786 ^ n25785 ^ n4582 ;
  assign n25788 = n20254 ^ n5590 ^ n2425 ;
  assign n25789 = ( n11098 & ~n25787 ) | ( n11098 & n25788 ) | ( ~n25787 & n25788 ) ;
  assign n25790 = ( n25782 & n25784 ) | ( n25782 & n25789 ) | ( n25784 & n25789 ) ;
  assign n25800 = ( n2922 & n4647 ) | ( n2922 & n16901 ) | ( n4647 & n16901 ) ;
  assign n25801 = n25800 ^ n19604 ^ n18316 ;
  assign n25794 = n11400 ^ x200 ^ 1'b0 ;
  assign n25793 = n8219 ^ n5441 ^ n3790 ;
  assign n25795 = n25794 ^ n25793 ^ n7585 ;
  assign n25791 = n8517 & ~n18368 ;
  assign n25792 = n25791 ^ n11872 ^ 1'b0 ;
  assign n25796 = n25795 ^ n25792 ^ n23775 ;
  assign n25797 = ( n9311 & n19259 ) | ( n9311 & n21858 ) | ( n19259 & n21858 ) ;
  assign n25798 = n25797 ^ n24723 ^ n14754 ;
  assign n25799 = n25796 | n25798 ;
  assign n25802 = n25801 ^ n25799 ^ n7907 ;
  assign n25803 = n708 & ~n3083 ;
  assign n25804 = ( n1172 & n8509 ) | ( n1172 & n20426 ) | ( n8509 & n20426 ) ;
  assign n25805 = ~n12023 & n25804 ;
  assign n25806 = ( n4828 & n25803 ) | ( n4828 & n25805 ) | ( n25803 & n25805 ) ;
  assign n25809 = ( ~n3047 & n4540 ) | ( ~n3047 & n10361 ) | ( n4540 & n10361 ) ;
  assign n25810 = n7719 & ~n25809 ;
  assign n25807 = n9041 ^ n8970 ^ n7344 ;
  assign n25808 = ~n23305 & n25807 ;
  assign n25811 = n25810 ^ n25808 ^ 1'b0 ;
  assign n25812 = n3319 & n25811 ;
  assign n25813 = n8223 ^ n6842 ^ n2493 ;
  assign n25814 = ( ~n8172 & n9286 ) | ( ~n8172 & n25813 ) | ( n9286 & n25813 ) ;
  assign n25815 = n8182 & ~n25814 ;
  assign n25816 = ( n6044 & ~n20275 ) | ( n6044 & n25815 ) | ( ~n20275 & n25815 ) ;
  assign n25817 = ( n6336 & n15054 ) | ( n6336 & n25325 ) | ( n15054 & n25325 ) ;
  assign n25818 = n19044 ^ n8382 ^ 1'b0 ;
  assign n25819 = n25817 & ~n25818 ;
  assign n25821 = n18275 ^ n15506 ^ n8704 ;
  assign n25820 = n19950 | n22892 ;
  assign n25822 = n25821 ^ n25820 ^ 1'b0 ;
  assign n25823 = ~n15776 & n21451 ;
  assign n25824 = n19984 & n25823 ;
  assign n25825 = ~n9472 & n15879 ;
  assign n25826 = n3149 & n13189 ;
  assign n25827 = n7076 & n25826 ;
  assign n25828 = n8594 | n25827 ;
  assign n25829 = n25828 ^ n2588 ^ 1'b0 ;
  assign n25830 = ( n1407 & n13507 ) | ( n1407 & ~n19833 ) | ( n13507 & ~n19833 ) ;
  assign n25831 = ( x243 & n14941 ) | ( x243 & ~n25830 ) | ( n14941 & ~n25830 ) ;
  assign n25832 = ( n9551 & n25829 ) | ( n9551 & n25831 ) | ( n25829 & n25831 ) ;
  assign n25833 = n7515 | n9186 ;
  assign n25834 = ( n9131 & ~n23761 ) | ( n9131 & n25833 ) | ( ~n23761 & n25833 ) ;
  assign n25835 = n10000 | n10844 ;
  assign n25836 = n1609 & ~n25835 ;
  assign n25837 = n13505 ^ n12663 ^ n12466 ;
  assign n25838 = n25837 ^ n18659 ^ n8746 ;
  assign n25839 = n5517 ^ n3018 ^ n2922 ;
  assign n25843 = ( ~n8735 & n8773 ) | ( ~n8735 & n21441 ) | ( n8773 & n21441 ) ;
  assign n25844 = n9799 & ~n10594 ;
  assign n25845 = n10925 ^ n5982 ^ n2607 ;
  assign n25846 = ( n2515 & ~n8461 ) | ( n2515 & n25845 ) | ( ~n8461 & n25845 ) ;
  assign n25847 = ( n14999 & ~n25844 ) | ( n14999 & n25846 ) | ( ~n25844 & n25846 ) ;
  assign n25848 = ( n5832 & n25843 ) | ( n5832 & n25847 ) | ( n25843 & n25847 ) ;
  assign n25840 = n14554 ^ n11067 ^ n3155 ;
  assign n25841 = n25840 ^ n12067 ^ n2427 ;
  assign n25842 = n25841 ^ n22511 ^ n17180 ;
  assign n25849 = n25848 ^ n25842 ^ n19346 ;
  assign n25851 = n23268 ^ n14334 ^ n14042 ;
  assign n25850 = n10312 ^ n6975 ^ n1543 ;
  assign n25852 = n25851 ^ n25850 ^ n4905 ;
  assign n25853 = n25338 ^ n4505 ^ n929 ;
  assign n25854 = n1221 & ~n15664 ;
  assign n25855 = n9466 ^ n7979 ^ 1'b0 ;
  assign n25856 = ~n18895 & n25855 ;
  assign n25857 = n25856 ^ n25842 ^ 1'b0 ;
  assign n25858 = n14950 ^ n3167 ^ n1023 ;
  assign n25859 = n25858 ^ n8977 ^ 1'b0 ;
  assign n25860 = n19281 ^ n8133 ^ 1'b0 ;
  assign n25861 = n4543 | n25860 ;
  assign n25862 = n13771 | n25861 ;
  assign n25863 = n19157 | n25862 ;
  assign n25864 = ( n2551 & ~n5845 ) | ( n2551 & n15475 ) | ( ~n5845 & n15475 ) ;
  assign n25865 = n16733 ^ n15701 ^ 1'b0 ;
  assign n25866 = ~n25864 & n25865 ;
  assign n25867 = ( ~n11400 & n12146 ) | ( ~n11400 & n24223 ) | ( n12146 & n24223 ) ;
  assign n25868 = n25867 ^ n25353 ^ n2524 ;
  assign n25869 = n25868 ^ n20231 ^ n20090 ;
  assign n25870 = n3686 & n17114 ;
  assign n25871 = n25870 ^ n5676 ^ 1'b0 ;
  assign n25872 = n25871 ^ n25221 ^ n3563 ;
  assign n25873 = ( n8585 & n24625 ) | ( n8585 & n25872 ) | ( n24625 & n25872 ) ;
  assign n25874 = n23606 ^ n19236 ^ n11183 ;
  assign n25877 = n16195 ^ n7256 ^ 1'b0 ;
  assign n25875 = n23103 ^ n16066 ^ n9378 ;
  assign n25876 = n25875 ^ n25604 ^ n14427 ;
  assign n25878 = n25877 ^ n25876 ^ x194 ;
  assign n25879 = n17823 ^ n3205 ^ 1'b0 ;
  assign n25880 = ( n373 & n7471 ) | ( n373 & n25879 ) | ( n7471 & n25879 ) ;
  assign n25881 = n13795 & n25880 ;
  assign n25882 = ( n4639 & n11386 ) | ( n4639 & ~n13412 ) | ( n11386 & ~n13412 ) ;
  assign n25883 = ( n3254 & n8665 ) | ( n3254 & ~n25882 ) | ( n8665 & ~n25882 ) ;
  assign n25884 = ( n6226 & ~n10439 ) | ( n6226 & n19580 ) | ( ~n10439 & n19580 ) ;
  assign n25885 = ( ~n23133 & n23544 ) | ( ~n23133 & n25884 ) | ( n23544 & n25884 ) ;
  assign n25886 = ( n1370 & n4249 ) | ( n1370 & ~n5929 ) | ( n4249 & ~n5929 ) ;
  assign n25888 = ~x243 & n12441 ;
  assign n25887 = ~n612 & n8055 ;
  assign n25889 = n25888 ^ n25887 ^ n18884 ;
  assign n25890 = ( ~n9708 & n22701 ) | ( ~n9708 & n25889 ) | ( n22701 & n25889 ) ;
  assign n25896 = ( ~n2180 & n4100 ) | ( ~n2180 & n4370 ) | ( n4100 & n4370 ) ;
  assign n25897 = n25896 ^ n13000 ^ n5132 ;
  assign n25891 = ( n276 & ~n2289 ) | ( n276 & n20608 ) | ( ~n2289 & n20608 ) ;
  assign n25892 = n2566 ^ n2451 ^ n2168 ;
  assign n25893 = n4142 | n25892 ;
  assign n25894 = n13881 | n25893 ;
  assign n25895 = n25891 & n25894 ;
  assign n25898 = n25897 ^ n25895 ^ 1'b0 ;
  assign n25903 = n17261 ^ n5369 ^ n2197 ;
  assign n25899 = n327 & ~n5696 ;
  assign n25900 = n25899 ^ n6592 ^ 1'b0 ;
  assign n25901 = ~n17801 & n25900 ;
  assign n25902 = n25901 ^ n19057 ^ n5910 ;
  assign n25904 = n25903 ^ n25902 ^ n9808 ;
  assign n25905 = ( ~n286 & n7835 ) | ( ~n286 & n14269 ) | ( n7835 & n14269 ) ;
  assign n25906 = n25905 ^ n25067 ^ n8553 ;
  assign n25907 = ( n7442 & n14843 ) | ( n7442 & ~n21326 ) | ( n14843 & ~n21326 ) ;
  assign n25908 = ( n4552 & n6743 ) | ( n4552 & ~n12302 ) | ( n6743 & ~n12302 ) ;
  assign n25909 = ( n2317 & ~n6159 ) | ( n2317 & n25908 ) | ( ~n6159 & n25908 ) ;
  assign n25910 = n25909 ^ n20677 ^ 1'b0 ;
  assign n25911 = n25907 & n25910 ;
  assign n25912 = n5530 & n21038 ;
  assign n25913 = n25912 ^ n11026 ^ n7718 ;
  assign n25914 = n23196 ^ n22377 ^ n6814 ;
  assign n25915 = ( n9713 & n11835 ) | ( n9713 & n17617 ) | ( n11835 & n17617 ) ;
  assign n25916 = ( n544 & ~n8551 ) | ( n544 & n25915 ) | ( ~n8551 & n25915 ) ;
  assign n25917 = n12395 ^ n6899 ^ n2468 ;
  assign n25918 = ( n1692 & n14814 ) | ( n1692 & n18515 ) | ( n14814 & n18515 ) ;
  assign n25919 = n25918 ^ n23235 ^ n15675 ;
  assign n25920 = ~n25917 & n25919 ;
  assign n25921 = ~n16789 & n18583 ;
  assign n25922 = n25921 ^ n3675 ^ 1'b0 ;
  assign n25923 = n10579 ^ n7179 ^ n4266 ;
  assign n25924 = n9764 | n19663 ;
  assign n25925 = n25924 ^ n4079 ^ 1'b0 ;
  assign n25926 = n15827 & ~n25925 ;
  assign n25927 = ( n1722 & n4703 ) | ( n1722 & ~n9711 ) | ( n4703 & ~n9711 ) ;
  assign n25928 = n22405 ^ n11378 ^ x156 ;
  assign n25929 = n18603 ^ n15560 ^ n12357 ;
  assign n25930 = n25929 ^ n21457 ^ n13192 ;
  assign n25931 = x209 & n4114 ;
  assign n25932 = n15010 ^ n4904 ^ n3811 ;
  assign n25933 = ( n14338 & ~n25931 ) | ( n14338 & n25932 ) | ( ~n25931 & n25932 ) ;
  assign n25934 = ( n1739 & n24367 ) | ( n1739 & ~n25933 ) | ( n24367 & ~n25933 ) ;
  assign n25940 = ~n665 & n5448 ;
  assign n25941 = n5792 & ~n25940 ;
  assign n25942 = n19974 & n25941 ;
  assign n25943 = ~n6417 & n10163 ;
  assign n25944 = ( n3131 & n25942 ) | ( n3131 & ~n25943 ) | ( n25942 & ~n25943 ) ;
  assign n25936 = n4411 & ~n6365 ;
  assign n25937 = ~n287 & n25936 ;
  assign n25935 = n16714 ^ n14709 ^ 1'b0 ;
  assign n25938 = n25937 ^ n25935 ^ n9437 ;
  assign n25939 = n25938 ^ n24936 ^ n22697 ;
  assign n25945 = n25944 ^ n25939 ^ n16841 ;
  assign n25946 = ( n1380 & ~n9820 ) | ( n1380 & n10716 ) | ( ~n9820 & n10716 ) ;
  assign n25947 = ( n20746 & n21328 ) | ( n20746 & ~n25946 ) | ( n21328 & ~n25946 ) ;
  assign n25948 = n4328 & n25947 ;
  assign n25949 = n25948 ^ n23821 ^ 1'b0 ;
  assign n25950 = ~n20078 & n20118 ;
  assign n25951 = n25950 ^ n708 ^ 1'b0 ;
  assign n25952 = n16440 ^ n15789 ^ n7392 ;
  assign n25953 = n21701 ^ n1959 ^ 1'b0 ;
  assign n25954 = n25952 & ~n25953 ;
  assign n25955 = ~n25951 & n25954 ;
  assign n25956 = n25955 ^ n23799 ^ 1'b0 ;
  assign n25957 = ( x85 & n10330 ) | ( x85 & n24542 ) | ( n10330 & n24542 ) ;
  assign n25958 = n25061 ^ n22369 ^ 1'b0 ;
  assign n25959 = n2527 & ~n25958 ;
  assign n25960 = ~n3402 & n25959 ;
  assign n25968 = n5664 ^ n5108 ^ n1389 ;
  assign n25969 = n1381 & n25968 ;
  assign n25970 = n689 & n25969 ;
  assign n25967 = n1519 & ~n7192 ;
  assign n25971 = n25970 ^ n25967 ^ 1'b0 ;
  assign n25963 = n8543 & n11580 ;
  assign n25964 = n25963 ^ n10647 ^ 1'b0 ;
  assign n25965 = n25964 ^ n14972 ^ n9535 ;
  assign n25961 = ( x95 & ~n3760 ) | ( x95 & n8193 ) | ( ~n3760 & n8193 ) ;
  assign n25962 = n23582 | n25961 ;
  assign n25966 = n25965 ^ n25962 ^ 1'b0 ;
  assign n25972 = n25971 ^ n25966 ^ n1042 ;
  assign n25973 = n16792 ^ n7461 ^ 1'b0 ;
  assign n25974 = ( n15117 & n16765 ) | ( n15117 & n25973 ) | ( n16765 & n25973 ) ;
  assign n25975 = n24908 ^ n18001 ^ n3243 ;
  assign n25976 = n17479 ^ n4646 ^ 1'b0 ;
  assign n25977 = n25975 & ~n25976 ;
  assign n25978 = n8537 & ~n25977 ;
  assign n25979 = ( n6494 & ~n13150 ) | ( n6494 & n19436 ) | ( ~n13150 & n19436 ) ;
  assign n25980 = n9216 ^ n5511 ^ n5258 ;
  assign n25981 = n25980 ^ n11120 ^ n7519 ;
  assign n25982 = ( ~n6459 & n8179 ) | ( ~n6459 & n13737 ) | ( n8179 & n13737 ) ;
  assign n25983 = n9379 & ~n24788 ;
  assign n25984 = n844 & n25983 ;
  assign n25985 = ( n7794 & ~n21599 ) | ( n7794 & n25984 ) | ( ~n21599 & n25984 ) ;
  assign n25986 = n25985 ^ n13378 ^ n3610 ;
  assign n25987 = n4318 | n6204 ;
  assign n25988 = n18618 & ~n25987 ;
  assign n25989 = n21319 | n25988 ;
  assign n25990 = n25989 ^ n17797 ^ 1'b0 ;
  assign n25991 = n18325 | n25990 ;
  assign n25992 = ( n11335 & n13989 ) | ( n11335 & ~n25991 ) | ( n13989 & ~n25991 ) ;
  assign n25993 = ~n3742 & n6501 ;
  assign n25994 = ~n9455 & n25993 ;
  assign n25995 = ( n3318 & n17975 ) | ( n3318 & n25994 ) | ( n17975 & n25994 ) ;
  assign n25996 = n25995 ^ n16504 ^ 1'b0 ;
  assign n25997 = n16725 ^ n3373 ^ 1'b0 ;
  assign n25998 = n7329 & ~n25997 ;
  assign n25999 = n16902 ^ n15973 ^ n3860 ;
  assign n26000 = ~n3349 & n16568 ;
  assign n26001 = n2219 | n26000 ;
  assign n26002 = ( n1908 & ~n4701 ) | ( n1908 & n26001 ) | ( ~n4701 & n26001 ) ;
  assign n26003 = n26002 ^ n18419 ^ 1'b0 ;
  assign n26004 = n24704 ^ n21552 ^ n11427 ;
  assign n26005 = ( ~n3399 & n14728 ) | ( ~n3399 & n26004 ) | ( n14728 & n26004 ) ;
  assign n26006 = ( n14149 & ~n26003 ) | ( n14149 & n26005 ) | ( ~n26003 & n26005 ) ;
  assign n26007 = ( ~n2030 & n25999 ) | ( ~n2030 & n26006 ) | ( n25999 & n26006 ) ;
  assign n26008 = n21090 ^ n1957 ^ n1204 ;
  assign n26009 = n26008 ^ n25388 ^ n15195 ;
  assign n26010 = n26009 ^ n7037 ^ 1'b0 ;
  assign n26011 = ~n10649 & n26010 ;
  assign n26012 = n26011 ^ n25342 ^ 1'b0 ;
  assign n26013 = ( ~n17966 & n24991 ) | ( ~n17966 & n26012 ) | ( n24991 & n26012 ) ;
  assign n26014 = ~n5867 & n26013 ;
  assign n26015 = n2442 & n4056 ;
  assign n26016 = n26015 ^ n6037 ^ 1'b0 ;
  assign n26017 = n17149 ^ n6272 ^ n4869 ;
  assign n26018 = ( n24299 & ~n26016 ) | ( n24299 & n26017 ) | ( ~n26016 & n26017 ) ;
  assign n26019 = n26018 ^ n21986 ^ 1'b0 ;
  assign n26020 = n18972 ^ n2015 ^ 1'b0 ;
  assign n26021 = n17196 & n26020 ;
  assign n26022 = n1216 & ~n16731 ;
  assign n26023 = ( x148 & ~n10390 ) | ( x148 & n26022 ) | ( ~n10390 & n26022 ) ;
  assign n26024 = ( n15878 & n26021 ) | ( n15878 & ~n26023 ) | ( n26021 & ~n26023 ) ;
  assign n26025 = n3862 ^ n2493 ^ n442 ;
  assign n26026 = n26025 ^ n11398 ^ n3574 ;
  assign n26027 = n17041 ^ n3593 ^ 1'b0 ;
  assign n26028 = n10747 | n26027 ;
  assign n26029 = n26028 ^ n11886 ^ n6287 ;
  assign n26030 = n663 | n3102 ;
  assign n26031 = n4647 | n26030 ;
  assign n26032 = ( n852 & ~n1225 ) | ( n852 & n5724 ) | ( ~n1225 & n5724 ) ;
  assign n26033 = n4131 | n16817 ;
  assign n26034 = ~n26032 & n26033 ;
  assign n26035 = ~n26031 & n26034 ;
  assign n26036 = ( n10233 & n26029 ) | ( n10233 & n26035 ) | ( n26029 & n26035 ) ;
  assign n26037 = n8116 & ~n15916 ;
  assign n26038 = n26037 ^ n22872 ^ 1'b0 ;
  assign n26039 = n13694 | n26038 ;
  assign n26040 = ( n2483 & n11212 ) | ( n2483 & ~n26039 ) | ( n11212 & ~n26039 ) ;
  assign n26042 = n4327 & ~n14810 ;
  assign n26043 = n13645 & n26042 ;
  assign n26044 = n26043 ^ n15493 ^ n3636 ;
  assign n26041 = n6762 & ~n9995 ;
  assign n26045 = n26044 ^ n26041 ^ 1'b0 ;
  assign n26046 = ( n4294 & n12521 ) | ( n4294 & n22623 ) | ( n12521 & n22623 ) ;
  assign n26047 = n26046 ^ n15625 ^ n9494 ;
  assign n26048 = n26047 ^ n18117 ^ n12250 ;
  assign n26049 = ~n3838 & n26048 ;
  assign n26057 = n8862 ^ n2760 ^ 1'b0 ;
  assign n26055 = n11033 ^ n2455 ^ 1'b0 ;
  assign n26051 = n6721 ^ n6328 ^ n6108 ;
  assign n26050 = n21599 ^ n17242 ^ n2062 ;
  assign n26052 = n26051 ^ n26050 ^ n12230 ;
  assign n26053 = ( n2609 & n6259 ) | ( n2609 & n26052 ) | ( n6259 & n26052 ) ;
  assign n26054 = n17712 & ~n26053 ;
  assign n26056 = n26055 ^ n26054 ^ 1'b0 ;
  assign n26058 = n26057 ^ n26056 ^ n1757 ;
  assign n26059 = n10272 ^ n7619 ^ n1792 ;
  assign n26060 = ( ~n22411 & n26058 ) | ( ~n22411 & n26059 ) | ( n26058 & n26059 ) ;
  assign n26061 = n9058 & ~n21705 ;
  assign n26062 = n26061 ^ n10381 ^ 1'b0 ;
  assign n26063 = n12394 | n26062 ;
  assign n26064 = n26063 ^ n24805 ^ n5675 ;
  assign n26065 = n23244 & ~n26064 ;
  assign n26066 = ( ~n5230 & n11095 ) | ( ~n5230 & n24677 ) | ( n11095 & n24677 ) ;
  assign n26067 = ( ~n13284 & n26065 ) | ( ~n13284 & n26066 ) | ( n26065 & n26066 ) ;
  assign n26068 = n2680 ^ n2150 ^ 1'b0 ;
  assign n26069 = n25762 | n26068 ;
  assign n26070 = ( n12271 & n25527 ) | ( n12271 & ~n26069 ) | ( n25527 & ~n26069 ) ;
  assign n26073 = ( n2256 & ~n3654 ) | ( n2256 & n4173 ) | ( ~n3654 & n4173 ) ;
  assign n26074 = n26073 ^ n11412 ^ n2505 ;
  assign n26075 = n26074 ^ n20487 ^ n19559 ;
  assign n26071 = n12620 & ~n16616 ;
  assign n26072 = n26071 ^ n5623 ^ 1'b0 ;
  assign n26076 = n26075 ^ n26072 ^ n7395 ;
  assign n26077 = n21130 ^ n9916 ^ 1'b0 ;
  assign n26078 = ( x82 & n2081 ) | ( x82 & n26077 ) | ( n2081 & n26077 ) ;
  assign n26079 = n26078 ^ n24137 ^ 1'b0 ;
  assign n26080 = ( n4565 & n4941 ) | ( n4565 & n7210 ) | ( n4941 & n7210 ) ;
  assign n26082 = n10307 ^ n9207 ^ n8024 ;
  assign n26081 = n22328 ^ n5587 ^ 1'b0 ;
  assign n26083 = n26082 ^ n26081 ^ n10132 ;
  assign n26087 = ( ~n1022 & n1790 ) | ( ~n1022 & n25168 ) | ( n1790 & n25168 ) ;
  assign n26084 = n17548 ^ n17441 ^ n3900 ;
  assign n26085 = n13615 ^ n8374 ^ n768 ;
  assign n26086 = ( ~n14598 & n26084 ) | ( ~n14598 & n26085 ) | ( n26084 & n26085 ) ;
  assign n26088 = n26087 ^ n26086 ^ n8254 ;
  assign n26089 = n4464 & ~n12314 ;
  assign n26090 = n1604 & n26089 ;
  assign n26091 = n26090 ^ n18658 ^ n14190 ;
  assign n26092 = ( n9442 & n18477 ) | ( n9442 & n24234 ) | ( n18477 & n24234 ) ;
  assign n26093 = n1808 | n16343 ;
  assign n26094 = n22242 | n26093 ;
  assign n26095 = n26092 & n26094 ;
  assign n26096 = n12115 ^ n8837 ^ 1'b0 ;
  assign n26097 = ( n3633 & ~n25217 ) | ( n3633 & n26096 ) | ( ~n25217 & n26096 ) ;
  assign n26098 = n7619 & ~n26097 ;
  assign n26099 = ( n14571 & ~n15279 ) | ( n14571 & n24687 ) | ( ~n15279 & n24687 ) ;
  assign n26100 = ( n1207 & n2636 ) | ( n1207 & ~n26099 ) | ( n2636 & ~n26099 ) ;
  assign n26101 = n13461 | n26100 ;
  assign n26102 = n26101 ^ n18825 ^ 1'b0 ;
  assign n26103 = ~n597 & n23473 ;
  assign n26104 = n26103 ^ x243 ^ 1'b0 ;
  assign n26105 = n9029 & n23567 ;
  assign n26106 = ~n4558 & n26105 ;
  assign n26107 = ( n271 & n8541 ) | ( n271 & ~n26106 ) | ( n8541 & ~n26106 ) ;
  assign n26108 = ( n5612 & n19669 ) | ( n5612 & n26107 ) | ( n19669 & n26107 ) ;
  assign n26109 = n20535 ^ n12868 ^ n9166 ;
  assign n26110 = ( ~n796 & n14860 ) | ( ~n796 & n19436 ) | ( n14860 & n19436 ) ;
  assign n26111 = n2852 | n12394 ;
  assign n26112 = n18905 | n26111 ;
  assign n26113 = ~n16614 & n26112 ;
  assign n26114 = n26113 ^ n402 ^ 1'b0 ;
  assign n26115 = n26114 ^ n9944 ^ n7419 ;
  assign n26116 = ( n872 & n1411 ) | ( n872 & n3794 ) | ( n1411 & n3794 ) ;
  assign n26117 = n16023 | n26116 ;
  assign n26118 = ( n4053 & n8926 ) | ( n4053 & n23128 ) | ( n8926 & n23128 ) ;
  assign n26119 = ( n8713 & n21207 ) | ( n8713 & ~n26118 ) | ( n21207 & ~n26118 ) ;
  assign n26120 = n1664 & n16238 ;
  assign n26121 = n5691 | n17022 ;
  assign n26123 = n5648 & ~n12188 ;
  assign n26124 = n26123 ^ n5636 ^ 1'b0 ;
  assign n26122 = ~n5815 & n25279 ;
  assign n26125 = n26124 ^ n26122 ^ 1'b0 ;
  assign n26126 = n26121 | n26125 ;
  assign n26130 = ( ~n1918 & n3178 ) | ( ~n1918 & n5370 ) | ( n3178 & n5370 ) ;
  assign n26131 = n10055 & n26130 ;
  assign n26127 = ( n1257 & n8545 ) | ( n1257 & ~n10721 ) | ( n8545 & ~n10721 ) ;
  assign n26128 = n11388 & n26127 ;
  assign n26129 = n4114 & ~n26128 ;
  assign n26132 = n26131 ^ n26129 ^ 1'b0 ;
  assign n26133 = n26132 ^ n8408 ^ 1'b0 ;
  assign n26134 = n7940 & ~n19717 ;
  assign n26135 = n26134 ^ n18236 ^ n5908 ;
  assign n26136 = ( ~n23910 & n25650 ) | ( ~n23910 & n26135 ) | ( n25650 & n26135 ) ;
  assign n26137 = ( n3796 & ~n25569 ) | ( n3796 & n26136 ) | ( ~n25569 & n26136 ) ;
  assign n26138 = n26137 ^ n25553 ^ n21078 ;
  assign n26139 = n9227 ^ n7868 ^ x189 ;
  assign n26142 = n7693 ^ n6323 ^ 1'b0 ;
  assign n26140 = n10316 & n18893 ;
  assign n26141 = n26140 ^ n25980 ^ n6152 ;
  assign n26143 = n26142 ^ n26141 ^ 1'b0 ;
  assign n26144 = ( n4991 & n12100 ) | ( n4991 & ~n16845 ) | ( n12100 & ~n16845 ) ;
  assign n26145 = n13829 ^ n12117 ^ n12097 ;
  assign n26146 = n342 | n2241 ;
  assign n26147 = n7259 ^ n3538 ^ 1'b0 ;
  assign n26148 = ~n26146 & n26147 ;
  assign n26149 = ~n10903 & n26148 ;
  assign n26150 = ( ~n4982 & n16283 ) | ( ~n4982 & n26149 ) | ( n16283 & n26149 ) ;
  assign n26157 = n12303 ^ n10759 ^ n9168 ;
  assign n26158 = n26157 ^ n14156 ^ x145 ;
  assign n26154 = n21601 ^ x134 ^ 1'b0 ;
  assign n26155 = n8566 & n26154 ;
  assign n26151 = n1773 & ~n5125 ;
  assign n26152 = n2091 & n26151 ;
  assign n26153 = n751 | n26152 ;
  assign n26156 = n26155 ^ n26153 ^ 1'b0 ;
  assign n26159 = n26158 ^ n26156 ^ n23918 ;
  assign n26160 = n9125 ^ n3213 ^ n576 ;
  assign n26161 = n26160 ^ n15977 ^ n11415 ;
  assign n26162 = ( ~n1707 & n2459 ) | ( ~n1707 & n7649 ) | ( n2459 & n7649 ) ;
  assign n26163 = n16345 ^ n14789 ^ 1'b0 ;
  assign n26164 = ( n1582 & n17361 ) | ( n1582 & ~n26163 ) | ( n17361 & ~n26163 ) ;
  assign n26165 = ( n5243 & n26162 ) | ( n5243 & n26164 ) | ( n26162 & n26164 ) ;
  assign n26166 = n3456 & n5144 ;
  assign n26167 = n9224 & n26166 ;
  assign n26168 = n19429 ^ n16411 ^ n8757 ;
  assign n26169 = ( n14368 & ~n26167 ) | ( n14368 & n26168 ) | ( ~n26167 & n26168 ) ;
  assign n26170 = n26169 ^ n11716 ^ n6397 ;
  assign n26171 = ~n5127 & n22458 ;
  assign n26172 = n22074 ^ n13887 ^ n11351 ;
  assign n26173 = n11897 ^ n1197 ^ 1'b0 ;
  assign n26174 = n26173 ^ n15986 ^ 1'b0 ;
  assign n26175 = ( n2152 & ~n4176 ) | ( n2152 & n7094 ) | ( ~n4176 & n7094 ) ;
  assign n26176 = ( x142 & ~n275 ) | ( x142 & n10445 ) | ( ~n275 & n10445 ) ;
  assign n26177 = n26176 ^ n8604 ^ n771 ;
  assign n26178 = n26177 ^ n606 ^ n564 ;
  assign n26179 = ( ~n17735 & n22704 ) | ( ~n17735 & n26178 ) | ( n22704 & n26178 ) ;
  assign n26180 = ~n17037 & n18358 ;
  assign n26181 = n17474 & n26180 ;
  assign n26182 = n13564 ^ n6069 ^ 1'b0 ;
  assign n26183 = ( n8204 & n21495 ) | ( n8204 & n26182 ) | ( n21495 & n26182 ) ;
  assign n26184 = n19836 ^ n8096 ^ 1'b0 ;
  assign n26185 = n26183 & n26184 ;
  assign n26186 = ( n3568 & ~n5554 ) | ( n3568 & n11850 ) | ( ~n5554 & n11850 ) ;
  assign n26187 = n26186 ^ n4070 ^ n1955 ;
  assign n26188 = n26187 ^ n6265 ^ 1'b0 ;
  assign n26189 = n14712 ^ n7804 ^ 1'b0 ;
  assign n26190 = ( ~n12391 & n15635 ) | ( ~n12391 & n25647 ) | ( n15635 & n25647 ) ;
  assign n26191 = ( n7462 & ~n16363 ) | ( n7462 & n26190 ) | ( ~n16363 & n26190 ) ;
  assign n26192 = ( n1042 & n19251 ) | ( n1042 & n26191 ) | ( n19251 & n26191 ) ;
  assign n26193 = n26192 ^ n7780 ^ 1'b0 ;
  assign n26194 = n26189 | n26193 ;
  assign n26195 = ( x206 & ~n864 ) | ( x206 & n26194 ) | ( ~n864 & n26194 ) ;
  assign n26196 = n11414 ^ n10058 ^ n2706 ;
  assign n26197 = n12133 ^ n11268 ^ 1'b0 ;
  assign n26198 = ( n5035 & n5498 ) | ( n5035 & ~n7938 ) | ( n5498 & ~n7938 ) ;
  assign n26199 = n26198 ^ n6657 ^ n2210 ;
  assign n26200 = ( ~n11869 & n26197 ) | ( ~n11869 & n26199 ) | ( n26197 & n26199 ) ;
  assign n26201 = ( n1635 & n25388 ) | ( n1635 & n26200 ) | ( n25388 & n26200 ) ;
  assign n26210 = ( n356 & ~n5176 ) | ( n356 & n9966 ) | ( ~n5176 & n9966 ) ;
  assign n26206 = ( ~n8249 & n13110 ) | ( ~n8249 & n18107 ) | ( n13110 & n18107 ) ;
  assign n26207 = n4056 & n18698 ;
  assign n26208 = ~n26206 & n26207 ;
  assign n26202 = n3578 & ~n23620 ;
  assign n26203 = n10654 ^ n4491 ^ n2884 ;
  assign n26204 = n26203 ^ n22064 ^ n6126 ;
  assign n26205 = ( n9165 & n26202 ) | ( n9165 & ~n26204 ) | ( n26202 & ~n26204 ) ;
  assign n26209 = n26208 ^ n26205 ^ n14912 ;
  assign n26211 = n26210 ^ n26209 ^ n22650 ;
  assign n26212 = x208 & n2597 ;
  assign n26213 = n1825 | n14124 ;
  assign n26214 = n9803 & ~n26213 ;
  assign n26215 = ( ~n24795 & n26212 ) | ( ~n24795 & n26214 ) | ( n26212 & n26214 ) ;
  assign n26216 = ( n2871 & ~n4172 ) | ( n2871 & n7515 ) | ( ~n4172 & n7515 ) ;
  assign n26217 = n26216 ^ n20619 ^ n800 ;
  assign n26218 = n26217 ^ n6940 ^ 1'b0 ;
  assign n26219 = n26218 ^ n19342 ^ n6508 ;
  assign n26223 = n25968 ^ n2622 ^ n2349 ;
  assign n26220 = ( n8286 & ~n22637 ) | ( n8286 & n24476 ) | ( ~n22637 & n24476 ) ;
  assign n26221 = n17318 | n26220 ;
  assign n26222 = n26221 ^ n25437 ^ 1'b0 ;
  assign n26224 = n26223 ^ n26222 ^ n7445 ;
  assign n26225 = ( n17820 & n25205 ) | ( n17820 & n26224 ) | ( n25205 & n26224 ) ;
  assign n26226 = ( ~n462 & n4636 ) | ( ~n462 & n20464 ) | ( n4636 & n20464 ) ;
  assign n26227 = n26226 ^ n20864 ^ 1'b0 ;
  assign n26228 = x67 & ~n26227 ;
  assign n26229 = ( ~n5290 & n5564 ) | ( ~n5290 & n8856 ) | ( n5564 & n8856 ) ;
  assign n26230 = n1346 & ~n2140 ;
  assign n26231 = n14555 & n26230 ;
  assign n26232 = ( n15248 & n26229 ) | ( n15248 & n26231 ) | ( n26229 & n26231 ) ;
  assign n26233 = ~n8428 & n13482 ;
  assign n26234 = n5742 ^ n3519 ^ n1447 ;
  assign n26235 = ( n5078 & ~n18023 ) | ( n5078 & n26234 ) | ( ~n18023 & n26234 ) ;
  assign n26236 = n26235 ^ n14357 ^ n5102 ;
  assign n26239 = n18466 ^ n18281 ^ n14554 ;
  assign n26237 = n13844 ^ n13330 ^ 1'b0 ;
  assign n26238 = n6640 & ~n26237 ;
  assign n26240 = n26239 ^ n26238 ^ 1'b0 ;
  assign n26241 = n13717 | n25478 ;
  assign n26242 = n26241 ^ n6739 ^ 1'b0 ;
  assign n26243 = ( ~n498 & n1604 ) | ( ~n498 & n26242 ) | ( n1604 & n26242 ) ;
  assign n26244 = ( n2371 & ~n2688 ) | ( n2371 & n13349 ) | ( ~n2688 & n13349 ) ;
  assign n26245 = n5790 ^ n4719 ^ 1'b0 ;
  assign n26246 = ~n14164 & n26245 ;
  assign n26247 = n26246 ^ n5691 ^ n3641 ;
  assign n26248 = ( n26243 & n26244 ) | ( n26243 & n26247 ) | ( n26244 & n26247 ) ;
  assign n26252 = ( n1444 & ~n12827 ) | ( n1444 & n13288 ) | ( ~n12827 & n13288 ) ;
  assign n26250 = n20236 ^ n5871 ^ n2408 ;
  assign n26251 = ( ~n3846 & n16492 ) | ( ~n3846 & n26250 ) | ( n16492 & n26250 ) ;
  assign n26249 = n14882 ^ n3231 ^ n459 ;
  assign n26253 = n26252 ^ n26251 ^ n26249 ;
  assign n26254 = n20070 ^ n4953 ^ n1370 ;
  assign n26255 = ( n308 & n9026 ) | ( n308 & ~n13815 ) | ( n9026 & ~n13815 ) ;
  assign n26256 = n8042 ^ n3959 ^ n1129 ;
  assign n26257 = n26256 ^ n4689 ^ n306 ;
  assign n26258 = ( n16390 & n26255 ) | ( n16390 & ~n26257 ) | ( n26255 & ~n26257 ) ;
  assign n26259 = n4096 & n20617 ;
  assign n26260 = n26259 ^ n15054 ^ 1'b0 ;
  assign n26261 = n23104 ^ n18105 ^ n13769 ;
  assign n26262 = n8946 & ~n24756 ;
  assign n26263 = ( ~n2944 & n18426 ) | ( ~n2944 & n25156 ) | ( n18426 & n25156 ) ;
  assign n26264 = n21165 ^ n8032 ^ n4132 ;
  assign n26265 = n26264 ^ n24321 ^ n15496 ;
  assign n26266 = n26265 ^ n13788 ^ 1'b0 ;
  assign n26267 = ~n8989 & n26266 ;
  assign n26268 = ( n4911 & n26263 ) | ( n4911 & n26267 ) | ( n26263 & n26267 ) ;
  assign n26275 = ( n2159 & n9310 ) | ( n2159 & ~n16225 ) | ( n9310 & ~n16225 ) ;
  assign n26273 = n17751 ^ n9936 ^ n8333 ;
  assign n26274 = ( ~n4051 & n11470 ) | ( ~n4051 & n26273 ) | ( n11470 & n26273 ) ;
  assign n26269 = n18975 | n19762 ;
  assign n26270 = n26269 ^ n12529 ^ 1'b0 ;
  assign n26271 = n5054 & n26270 ;
  assign n26272 = ~n17557 & n26271 ;
  assign n26276 = n26275 ^ n26274 ^ n26272 ;
  assign n26277 = n24884 ^ n2625 ^ n1132 ;
  assign n26280 = ( n2586 & ~n8789 ) | ( n2586 & n13052 ) | ( ~n8789 & n13052 ) ;
  assign n26278 = ( n2016 & ~n3208 ) | ( n2016 & n13603 ) | ( ~n3208 & n13603 ) ;
  assign n26279 = n26278 ^ n10944 ^ n9435 ;
  assign n26281 = n26280 ^ n26279 ^ n13919 ;
  assign n26282 = n5962 & n11586 ;
  assign n26283 = ( n6785 & n26281 ) | ( n6785 & ~n26282 ) | ( n26281 & ~n26282 ) ;
  assign n26284 = ( n5103 & n14795 ) | ( n5103 & n16746 ) | ( n14795 & n16746 ) ;
  assign n26285 = ( n22393 & n26283 ) | ( n22393 & n26284 ) | ( n26283 & n26284 ) ;
  assign n26286 = ~n14608 & n18704 ;
  assign n26287 = ( n15046 & n15182 ) | ( n15046 & n19159 ) | ( n15182 & n19159 ) ;
  assign n26288 = n26286 & ~n26287 ;
  assign n26289 = ( n4253 & n12311 ) | ( n4253 & ~n12728 ) | ( n12311 & ~n12728 ) ;
  assign n26290 = ~n4403 & n12880 ;
  assign n26291 = n26290 ^ n16988 ^ 1'b0 ;
  assign n26292 = ( ~n1320 & n20243 ) | ( ~n1320 & n26291 ) | ( n20243 & n26291 ) ;
  assign n26293 = n13647 & ~n23131 ;
  assign n26294 = ( n8342 & ~n10205 ) | ( n8342 & n11657 ) | ( ~n10205 & n11657 ) ;
  assign n26295 = n26294 ^ n11025 ^ 1'b0 ;
  assign n26296 = n3798 & ~n26295 ;
  assign n26297 = ( n974 & n26293 ) | ( n974 & n26296 ) | ( n26293 & n26296 ) ;
  assign n26298 = ( n5623 & n20616 ) | ( n5623 & ~n24359 ) | ( n20616 & ~n24359 ) ;
  assign n26299 = n12372 & n26298 ;
  assign n26300 = n24485 & n26299 ;
  assign n26301 = ( n10822 & n25250 ) | ( n10822 & n26300 ) | ( n25250 & n26300 ) ;
  assign n26302 = n7225 ^ n5733 ^ 1'b0 ;
  assign n26303 = n1903 & ~n26302 ;
  assign n26304 = n20231 ^ n2581 ^ 1'b0 ;
  assign n26305 = n26303 & n26304 ;
  assign n26307 = ~n2612 & n17245 ;
  assign n26308 = n24529 & n26307 ;
  assign n26306 = ( n10309 & n10509 ) | ( n10309 & ~n15715 ) | ( n10509 & ~n15715 ) ;
  assign n26309 = n26308 ^ n26306 ^ n9670 ;
  assign n26310 = n2294 | n5480 ;
  assign n26311 = n5595 | n6825 ;
  assign n26312 = n21899 | n26311 ;
  assign n26313 = ~n9850 & n26312 ;
  assign n26314 = n21793 & n26313 ;
  assign n26319 = n5426 ^ n1911 ^ 1'b0 ;
  assign n26320 = n14254 ^ n6750 ^ 1'b0 ;
  assign n26321 = n26319 & n26320 ;
  assign n26315 = n16763 ^ n2164 ^ n949 ;
  assign n26316 = ( n4485 & n21222 ) | ( n4485 & n26315 ) | ( n21222 & n26315 ) ;
  assign n26317 = n22691 | n26316 ;
  assign n26318 = n26317 ^ n15597 ^ 1'b0 ;
  assign n26322 = n26321 ^ n26318 ^ n18736 ;
  assign n26324 = n16528 ^ n12244 ^ n9352 ;
  assign n26323 = n23074 & ~n24665 ;
  assign n26325 = n26324 ^ n26323 ^ n20483 ;
  assign n26326 = n10744 ^ n8492 ^ n8376 ;
  assign n26327 = ( n10900 & n24656 ) | ( n10900 & ~n26326 ) | ( n24656 & ~n26326 ) ;
  assign n26328 = n26327 ^ n7174 ^ n3083 ;
  assign n26329 = ( n19083 & ~n25091 ) | ( n19083 & n26328 ) | ( ~n25091 & n26328 ) ;
  assign n26330 = ~n13306 & n16922 ;
  assign n26331 = n26330 ^ n25005 ^ 1'b0 ;
  assign n26332 = ( n5881 & n9997 ) | ( n5881 & n11827 ) | ( n9997 & n11827 ) ;
  assign n26333 = ( n7446 & ~n10817 ) | ( n7446 & n19267 ) | ( ~n10817 & n19267 ) ;
  assign n26334 = n26333 ^ n22271 ^ n11056 ;
  assign n26335 = ( ~n4545 & n5684 ) | ( ~n4545 & n21418 ) | ( n5684 & n21418 ) ;
  assign n26336 = ( ~n7589 & n22271 ) | ( ~n7589 & n26335 ) | ( n22271 & n26335 ) ;
  assign n26337 = n26336 ^ n15615 ^ n4543 ;
  assign n26341 = ( ~n2585 & n7944 ) | ( ~n2585 & n20013 ) | ( n7944 & n20013 ) ;
  assign n26338 = ~n6886 & n19321 ;
  assign n26339 = n26338 ^ n10073 ^ 1'b0 ;
  assign n26340 = n26339 ^ n11921 ^ 1'b0 ;
  assign n26342 = n26341 ^ n26340 ^ 1'b0 ;
  assign n26343 = n5070 ^ n4063 ^ n974 ;
  assign n26344 = ( ~n1347 & n2713 ) | ( ~n1347 & n5283 ) | ( n2713 & n5283 ) ;
  assign n26345 = ( ~n1697 & n12588 ) | ( ~n1697 & n26344 ) | ( n12588 & n26344 ) ;
  assign n26346 = ( ~n2298 & n6110 ) | ( ~n2298 & n7983 ) | ( n6110 & n7983 ) ;
  assign n26347 = ( n26343 & n26345 ) | ( n26343 & n26346 ) | ( n26345 & n26346 ) ;
  assign n26348 = ( ~n3181 & n15515 ) | ( ~n3181 & n24970 ) | ( n15515 & n24970 ) ;
  assign n26349 = n6125 & ~n18126 ;
  assign n26350 = n24959 & n26349 ;
  assign n26351 = n15989 ^ n11978 ^ n10775 ;
  assign n26352 = ~n3757 & n26351 ;
  assign n26353 = n15122 & n26352 ;
  assign n26354 = n26353 ^ n5452 ^ x3 ;
  assign n26355 = n26354 ^ n18713 ^ n7885 ;
  assign n26356 = n9383 ^ n7913 ^ 1'b0 ;
  assign n26357 = ~n7910 & n26356 ;
  assign n26360 = ~n17500 & n18073 ;
  assign n26361 = n6472 & n26360 ;
  assign n26362 = n26361 ^ n5587 ^ n614 ;
  assign n26358 = n10155 ^ n7163 ^ 1'b0 ;
  assign n26359 = n6272 & ~n26358 ;
  assign n26363 = n26362 ^ n26359 ^ 1'b0 ;
  assign n26364 = ( n972 & n6382 ) | ( n972 & n6842 ) | ( n6382 & n6842 ) ;
  assign n26365 = ( ~x2 & n18787 ) | ( ~x2 & n26364 ) | ( n18787 & n26364 ) ;
  assign n26366 = ( n4239 & n8844 ) | ( n4239 & ~n26365 ) | ( n8844 & ~n26365 ) ;
  assign n26367 = ( n2142 & ~n22025 ) | ( n2142 & n26366 ) | ( ~n22025 & n26366 ) ;
  assign n26368 = n18255 ^ n9708 ^ n2519 ;
  assign n26369 = ( n7686 & n11006 ) | ( n7686 & n26368 ) | ( n11006 & n26368 ) ;
  assign n26370 = n9464 ^ n9401 ^ n9262 ;
  assign n26371 = n26370 ^ n12257 ^ 1'b0 ;
  assign n26372 = n4827 ^ n3848 ^ n1767 ;
  assign n26373 = n19155 ^ n7745 ^ 1'b0 ;
  assign n26374 = n26372 & ~n26373 ;
  assign n26375 = ( n1550 & n1879 ) | ( n1550 & n26374 ) | ( n1879 & n26374 ) ;
  assign n26376 = ~n7039 & n13329 ;
  assign n26377 = ( ~n14398 & n20873 ) | ( ~n14398 & n26376 ) | ( n20873 & n26376 ) ;
  assign n26378 = n5175 & n26377 ;
  assign n26379 = ~n10611 & n26378 ;
  assign n26380 = n25015 ^ n19148 ^ n7858 ;
  assign n26381 = n26380 ^ n13843 ^ 1'b0 ;
  assign n26382 = n2644 & n26381 ;
  assign n26383 = n24819 ^ x213 ^ 1'b0 ;
  assign n26384 = ( ~n966 & n2347 ) | ( ~n966 & n26383 ) | ( n2347 & n26383 ) ;
  assign n26385 = ( n19183 & n22050 ) | ( n19183 & n26384 ) | ( n22050 & n26384 ) ;
  assign n26386 = n20194 ^ n3945 ^ 1'b0 ;
  assign n26387 = n26386 ^ n14630 ^ n1795 ;
  assign n26391 = ( n1461 & ~n14721 ) | ( n1461 & n16388 ) | ( ~n14721 & n16388 ) ;
  assign n26392 = n26391 ^ n15489 ^ n15406 ;
  assign n26388 = ~n1635 & n7124 ;
  assign n26389 = n26388 ^ n6333 ^ n5401 ;
  assign n26390 = n26389 ^ n11995 ^ 1'b0 ;
  assign n26393 = n26392 ^ n26390 ^ n4073 ;
  assign n26394 = ~n11043 & n22392 ;
  assign n26395 = n7370 & ~n9144 ;
  assign n26396 = ( n2318 & ~n6137 ) | ( n2318 & n18423 ) | ( ~n6137 & n18423 ) ;
  assign n26397 = ~n26395 & n26396 ;
  assign n26398 = ~n26394 & n26397 ;
  assign n26399 = ~n5324 & n16268 ;
  assign n26400 = n26399 ^ n7872 ^ n2786 ;
  assign n26401 = n26400 ^ n16744 ^ 1'b0 ;
  assign n26404 = n5053 ^ n4734 ^ n394 ;
  assign n26402 = n14503 ^ n1983 ^ x69 ;
  assign n26403 = ( n22780 & n25411 ) | ( n22780 & ~n26402 ) | ( n25411 & ~n26402 ) ;
  assign n26405 = n26404 ^ n26403 ^ n14181 ;
  assign n26406 = n6412 ^ n364 ^ 1'b0 ;
  assign n26407 = n10997 & n26406 ;
  assign n26408 = ( ~n9649 & n12273 ) | ( ~n9649 & n26407 ) | ( n12273 & n26407 ) ;
  assign n26409 = ( n8169 & n9053 ) | ( n8169 & ~n17607 ) | ( n9053 & ~n17607 ) ;
  assign n26410 = ( n1258 & ~n17104 ) | ( n1258 & n26409 ) | ( ~n17104 & n26409 ) ;
  assign n26411 = ( n7519 & n18871 ) | ( n7519 & ~n26410 ) | ( n18871 & ~n26410 ) ;
  assign n26412 = n26411 ^ n18597 ^ n277 ;
  assign n26413 = ( ~n4096 & n13658 ) | ( ~n4096 & n15426 ) | ( n13658 & n15426 ) ;
  assign n26414 = ~n19325 & n25260 ;
  assign n26415 = n26414 ^ n2577 ^ 1'b0 ;
  assign n26416 = n17792 & ~n22926 ;
  assign n26417 = n26416 ^ n2446 ^ 1'b0 ;
  assign n26418 = n12068 ^ n2177 ^ 1'b0 ;
  assign n26419 = ( n8025 & ~n15927 ) | ( n8025 & n20092 ) | ( ~n15927 & n20092 ) ;
  assign n26420 = n26419 ^ n12918 ^ 1'b0 ;
  assign n26421 = n26420 ^ n20062 ^ x45 ;
  assign n26422 = n12581 & n26421 ;
  assign n26423 = n26422 ^ n13306 ^ 1'b0 ;
  assign n26424 = n14719 & n26423 ;
  assign n26426 = ( ~n10799 & n14950 ) | ( ~n10799 & n19378 ) | ( n14950 & n19378 ) ;
  assign n26425 = n11217 | n23937 ;
  assign n26427 = n26426 ^ n26425 ^ 1'b0 ;
  assign n26428 = ( n660 & n6028 ) | ( n660 & n8430 ) | ( n6028 & n8430 ) ;
  assign n26429 = n17436 ^ n16204 ^ n13100 ;
  assign n26430 = ( n11862 & n26428 ) | ( n11862 & ~n26429 ) | ( n26428 & ~n26429 ) ;
  assign n26431 = n24063 ^ n23840 ^ n17757 ;
  assign n26432 = n8139 ^ n3327 ^ 1'b0 ;
  assign n26433 = n21016 ^ n17890 ^ n6633 ;
  assign n26434 = ( ~n20912 & n26432 ) | ( ~n20912 & n26433 ) | ( n26432 & n26433 ) ;
  assign n26435 = n16597 ^ n4117 ^ 1'b0 ;
  assign n26436 = ( n12944 & ~n26434 ) | ( n12944 & n26435 ) | ( ~n26434 & n26435 ) ;
  assign n26437 = n17692 ^ n15254 ^ n4064 ;
  assign n26438 = ~n8997 & n26437 ;
  assign n26439 = n7953 ^ n5785 ^ 1'b0 ;
  assign n26440 = n24690 & n26439 ;
  assign n26442 = n13712 ^ n7273 ^ x28 ;
  assign n26441 = n10890 ^ n8953 ^ n3437 ;
  assign n26443 = n26442 ^ n26441 ^ n19730 ;
  assign n26444 = ( x112 & n4604 ) | ( x112 & n19397 ) | ( n4604 & n19397 ) ;
  assign n26445 = ( n14254 & n17467 ) | ( n14254 & n19840 ) | ( n17467 & n19840 ) ;
  assign n26446 = ( n7153 & n13636 ) | ( n7153 & n26445 ) | ( n13636 & n26445 ) ;
  assign n26447 = n13330 ^ n7262 ^ n6231 ;
  assign n26448 = n7485 ^ n7102 ^ 1'b0 ;
  assign n26449 = ( n4204 & n9623 ) | ( n4204 & ~n18117 ) | ( n9623 & ~n18117 ) ;
  assign n26450 = ( ~n3305 & n9929 ) | ( ~n3305 & n26449 ) | ( n9929 & n26449 ) ;
  assign n26451 = ( n7251 & n26448 ) | ( n7251 & n26450 ) | ( n26448 & n26450 ) ;
  assign n26452 = ( n20492 & ~n26447 ) | ( n20492 & n26451 ) | ( ~n26447 & n26451 ) ;
  assign n26453 = n26452 ^ n24893 ^ 1'b0 ;
  assign n26454 = ( n9917 & ~n17276 ) | ( n9917 & n18095 ) | ( ~n17276 & n18095 ) ;
  assign n26455 = n1405 & ~n6617 ;
  assign n26456 = ~n2475 & n26455 ;
  assign n26457 = ( ~n8695 & n11406 ) | ( ~n8695 & n17883 ) | ( n11406 & n17883 ) ;
  assign n26458 = ( ~n15106 & n19528 ) | ( ~n15106 & n26457 ) | ( n19528 & n26457 ) ;
  assign n26459 = ( n3249 & n10628 ) | ( n3249 & ~n16176 ) | ( n10628 & ~n16176 ) ;
  assign n26460 = ( n5017 & n13070 ) | ( n5017 & ~n26459 ) | ( n13070 & ~n26459 ) ;
  assign n26461 = ( n2646 & ~n4644 ) | ( n2646 & n26460 ) | ( ~n4644 & n26460 ) ;
  assign n26462 = n19101 ^ n6373 ^ 1'b0 ;
  assign n26463 = n14873 & ~n26462 ;
  assign n26464 = ~n13241 & n13806 ;
  assign n26468 = ( n4388 & n5020 ) | ( n4388 & n8933 ) | ( n5020 & n8933 ) ;
  assign n26467 = n14039 ^ n9903 ^ n5388 ;
  assign n26469 = n26468 ^ n26467 ^ n16309 ;
  assign n26465 = n16463 ^ n11839 ^ n2565 ;
  assign n26466 = n26465 ^ n14702 ^ 1'b0 ;
  assign n26470 = n26469 ^ n26466 ^ 1'b0 ;
  assign n26471 = n26464 | n26470 ;
  assign n26472 = ( n3933 & n7845 ) | ( n3933 & n9250 ) | ( n7845 & n9250 ) ;
  assign n26473 = ( ~x131 & n5172 ) | ( ~x131 & n26472 ) | ( n5172 & n26472 ) ;
  assign n26474 = n4685 & n8149 ;
  assign n26475 = ( n2741 & ~n15776 ) | ( n2741 & n16846 ) | ( ~n15776 & n16846 ) ;
  assign n26476 = n26474 & n26475 ;
  assign n26477 = n26473 & n26476 ;
  assign n26478 = n26477 ^ n17193 ^ n5981 ;
  assign n26479 = n26478 ^ n15645 ^ 1'b0 ;
  assign n26480 = n9979 & n26479 ;
  assign n26481 = ( n870 & n15506 ) | ( n870 & n26480 ) | ( n15506 & n26480 ) ;
  assign n26482 = ( n915 & ~n21705 ) | ( n915 & n25590 ) | ( ~n21705 & n25590 ) ;
  assign n26483 = ( n4665 & n9500 ) | ( n4665 & n9851 ) | ( n9500 & n9851 ) ;
  assign n26484 = n6048 ^ n1876 ^ 1'b0 ;
  assign n26485 = n24672 | n26484 ;
  assign n26486 = ( n7734 & n26483 ) | ( n7734 & ~n26485 ) | ( n26483 & ~n26485 ) ;
  assign n26487 = n8778 ^ n8400 ^ n6269 ;
  assign n26488 = ( n1091 & n5643 ) | ( n1091 & ~n15500 ) | ( n5643 & ~n15500 ) ;
  assign n26489 = n5357 & n7245 ;
  assign n26490 = n26489 ^ n9283 ^ 1'b0 ;
  assign n26491 = n3845 & ~n26490 ;
  assign n26492 = n11550 ^ n10790 ^ x201 ;
  assign n26493 = ( n10244 & n15098 ) | ( n10244 & n26492 ) | ( n15098 & n26492 ) ;
  assign n26494 = n21412 ^ n15093 ^ n13249 ;
  assign n26495 = ( n1440 & n11729 ) | ( n1440 & ~n26494 ) | ( n11729 & ~n26494 ) ;
  assign n26496 = n11224 ^ n11131 ^ n11127 ;
  assign n26497 = n15339 ^ n11137 ^ 1'b0 ;
  assign n26500 = n11160 | n18903 ;
  assign n26498 = n6621 & ~n13571 ;
  assign n26499 = ( ~n8850 & n19636 ) | ( ~n8850 & n26498 ) | ( n19636 & n26498 ) ;
  assign n26501 = n26500 ^ n26499 ^ n20204 ;
  assign n26502 = n6216 & n12413 ;
  assign n26504 = ( ~n1777 & n6555 ) | ( ~n1777 & n23150 ) | ( n6555 & n23150 ) ;
  assign n26503 = n20219 & ~n25466 ;
  assign n26505 = n26504 ^ n26503 ^ 1'b0 ;
  assign n26506 = ( ~n4892 & n6151 ) | ( ~n4892 & n12724 ) | ( n6151 & n12724 ) ;
  assign n26507 = n12590 ^ n9162 ^ n3074 ;
  assign n26508 = n4656 ^ n2636 ^ 1'b0 ;
  assign n26509 = n18529 ^ n4914 ^ 1'b0 ;
  assign n26510 = ( ~n8525 & n12998 ) | ( ~n8525 & n21724 ) | ( n12998 & n21724 ) ;
  assign n26511 = ~n4899 & n5401 ;
  assign n26512 = ( n9051 & n13985 ) | ( n9051 & ~n26511 ) | ( n13985 & ~n26511 ) ;
  assign n26513 = n26512 ^ n1636 ^ 1'b0 ;
  assign n26514 = n26510 & ~n26513 ;
  assign n26515 = ( n26508 & ~n26509 ) | ( n26508 & n26514 ) | ( ~n26509 & n26514 ) ;
  assign n26516 = n3145 | n15450 ;
  assign n26517 = n4630 | n26516 ;
  assign n26518 = n26517 ^ n18842 ^ n11183 ;
  assign n26521 = n15262 ^ n6001 ^ n4946 ;
  assign n26519 = n24114 ^ n5252 ^ 1'b0 ;
  assign n26520 = ~n8738 & n26519 ;
  assign n26522 = n26521 ^ n26520 ^ 1'b0 ;
  assign n26523 = n14156 | n26522 ;
  assign n26524 = ( ~n8448 & n12288 ) | ( ~n8448 & n26371 ) | ( n12288 & n26371 ) ;
  assign n26526 = n11796 ^ n11519 ^ n3999 ;
  assign n26527 = n26526 ^ n3496 ^ n2873 ;
  assign n26528 = x23 & ~n13156 ;
  assign n26529 = ~n26527 & n26528 ;
  assign n26525 = ( n13843 & ~n15457 ) | ( n13843 & n20845 ) | ( ~n15457 & n20845 ) ;
  assign n26530 = n26529 ^ n26525 ^ n8945 ;
  assign n26531 = n1442 ^ n1164 ^ 1'b0 ;
  assign n26533 = n2404 | n3816 ;
  assign n26532 = ~n14092 & n20258 ;
  assign n26534 = n26533 ^ n26532 ^ 1'b0 ;
  assign n26535 = n26534 ^ n25388 ^ n13468 ;
  assign n26536 = n26535 ^ n10589 ^ n7979 ;
  assign n26537 = ( n10558 & n26531 ) | ( n10558 & n26536 ) | ( n26531 & n26536 ) ;
  assign n26538 = ( n4810 & n11433 ) | ( n4810 & n11961 ) | ( n11433 & n11961 ) ;
  assign n26539 = n12813 ^ n12713 ^ n1777 ;
  assign n26540 = n26539 ^ n26274 ^ n6309 ;
  assign n26541 = n17084 ^ n12595 ^ n12370 ;
  assign n26542 = n26541 ^ n25512 ^ 1'b0 ;
  assign n26543 = n9834 & n26542 ;
  assign n26544 = n24900 ^ n9359 ^ n2859 ;
  assign n26545 = n26544 ^ n12358 ^ n8117 ;
  assign n26546 = n5461 | n26545 ;
  assign n26547 = n24825 & ~n26546 ;
  assign n26548 = n6187 & ~n7019 ;
  assign n26549 = n26548 ^ n1027 ^ 1'b0 ;
  assign n26550 = ( n3468 & n18104 ) | ( n3468 & n26549 ) | ( n18104 & n26549 ) ;
  assign n26551 = ( n2506 & n6151 ) | ( n2506 & ~n10743 ) | ( n6151 & ~n10743 ) ;
  assign n26552 = n14432 & ~n26308 ;
  assign n26553 = ( n20037 & n25087 ) | ( n20037 & n26552 ) | ( n25087 & n26552 ) ;
  assign n26554 = n774 | n4379 ;
  assign n26555 = ( ~n21292 & n23998 ) | ( ~n21292 & n26554 ) | ( n23998 & n26554 ) ;
  assign n26556 = n6684 ^ n2038 ^ 1'b0 ;
  assign n26557 = n14635 & ~n26556 ;
  assign n26558 = n26557 ^ n17725 ^ 1'b0 ;
  assign n26559 = n3812 & ~n20737 ;
  assign n26560 = ( n6963 & n8886 ) | ( n6963 & n13062 ) | ( n8886 & n13062 ) ;
  assign n26561 = ( n3909 & ~n4974 ) | ( n3909 & n6117 ) | ( ~n4974 & n6117 ) ;
  assign n26562 = n21573 ^ n21152 ^ n1482 ;
  assign n26563 = ( n21733 & ~n26561 ) | ( n21733 & n26562 ) | ( ~n26561 & n26562 ) ;
  assign n26564 = ( n1264 & ~n9717 ) | ( n1264 & n14133 ) | ( ~n9717 & n14133 ) ;
  assign n26565 = n26564 ^ n12616 ^ 1'b0 ;
  assign n26566 = ( n1832 & n4993 ) | ( n1832 & ~n6737 ) | ( n4993 & ~n6737 ) ;
  assign n26567 = n26566 ^ n10282 ^ n3658 ;
  assign n26568 = ( n304 & n3855 ) | ( n304 & n26567 ) | ( n3855 & n26567 ) ;
  assign n26569 = n16011 & n22482 ;
  assign n26570 = ~n1905 & n26569 ;
  assign n26571 = n12266 ^ n10840 ^ n7383 ;
  assign n26572 = ( ~n11915 & n26570 ) | ( ~n11915 & n26571 ) | ( n26570 & n26571 ) ;
  assign n26573 = n21564 ^ n1859 ^ 1'b0 ;
  assign n26574 = ~n22884 & n26573 ;
  assign n26575 = n17001 ^ n12113 ^ n9822 ;
  assign n26576 = ( ~n5691 & n6600 ) | ( ~n5691 & n14955 ) | ( n6600 & n14955 ) ;
  assign n26577 = n16603 ^ n12589 ^ x235 ;
  assign n26578 = n26577 ^ n24654 ^ n21583 ;
  assign n26579 = ( n15652 & n26576 ) | ( n15652 & n26578 ) | ( n26576 & n26578 ) ;
  assign n26580 = ( ~n24198 & n26575 ) | ( ~n24198 & n26579 ) | ( n26575 & n26579 ) ;
  assign n26581 = n21118 ^ n8309 ^ n1496 ;
  assign n26582 = ( n4031 & n14845 ) | ( n4031 & n16276 ) | ( n14845 & n16276 ) ;
  assign n26583 = n16467 ^ n13964 ^ 1'b0 ;
  assign n26584 = ~n13115 & n26583 ;
  assign n26585 = n19885 ^ n17254 ^ 1'b0 ;
  assign n26586 = n25968 ^ n17443 ^ n1444 ;
  assign n26587 = ( n18438 & ~n19729 ) | ( n18438 & n26586 ) | ( ~n19729 & n26586 ) ;
  assign n26588 = n26587 ^ n23839 ^ n20692 ;
  assign n26589 = n15734 & ~n26588 ;
  assign n26590 = n20372 ^ n7576 ^ n5219 ;
  assign n26591 = ( n8677 & n24502 ) | ( n8677 & n26590 ) | ( n24502 & n26590 ) ;
  assign n26592 = n23349 & n26591 ;
  assign n26593 = n5959 ^ n3144 ^ n1467 ;
  assign n26594 = ~n4698 & n17903 ;
  assign n26595 = n26593 & n26594 ;
  assign n26596 = ( x56 & n19549 ) | ( x56 & n26595 ) | ( n19549 & n26595 ) ;
  assign n26597 = n26596 ^ n20208 ^ n17008 ;
  assign n26598 = ( n3968 & n23073 ) | ( n3968 & ~n26597 ) | ( n23073 & ~n26597 ) ;
  assign n26599 = ( ~n11453 & n13008 ) | ( ~n11453 & n26598 ) | ( n13008 & n26598 ) ;
  assign n26600 = n4758 & n11183 ;
  assign n26601 = n26600 ^ n373 ^ 1'b0 ;
  assign n26602 = n10497 & n17677 ;
  assign n26603 = ~n22264 & n26602 ;
  assign n26604 = ( n5566 & ~n11275 ) | ( n5566 & n24337 ) | ( ~n11275 & n24337 ) ;
  assign n26605 = ( n5973 & n11433 ) | ( n5973 & ~n26604 ) | ( n11433 & ~n26604 ) ;
  assign n26606 = ( n5332 & n6178 ) | ( n5332 & ~n11408 ) | ( n6178 & ~n11408 ) ;
  assign n26607 = n24640 ^ n19507 ^ n8860 ;
  assign n26608 = n3370 & ~n26607 ;
  assign n26609 = n26606 & n26608 ;
  assign n26612 = n14839 ^ n3464 ^ n423 ;
  assign n26613 = n26612 ^ n7292 ^ 1'b0 ;
  assign n26610 = n1980 & n4045 ;
  assign n26611 = ( ~n3773 & n15455 ) | ( ~n3773 & n26610 ) | ( n15455 & n26610 ) ;
  assign n26614 = n26613 ^ n26611 ^ n6078 ;
  assign n26615 = ( ~n407 & n14880 ) | ( ~n407 & n25086 ) | ( n14880 & n25086 ) ;
  assign n26616 = ( ~n6903 & n13792 ) | ( ~n6903 & n26615 ) | ( n13792 & n26615 ) ;
  assign n26617 = ~n6184 & n6641 ;
  assign n26618 = ~n6087 & n20892 ;
  assign n26619 = n14727 & n26618 ;
  assign n26620 = ( n8701 & n26617 ) | ( n8701 & ~n26619 ) | ( n26617 & ~n26619 ) ;
  assign n26621 = ~n26066 & n26620 ;
  assign n26622 = n19166 & n20526 ;
  assign n26623 = ~n26366 & n26622 ;
  assign n26624 = ( n5093 & n5993 ) | ( n5093 & ~n26623 ) | ( n5993 & ~n26623 ) ;
  assign n26625 = n23553 ^ n6257 ^ n4565 ;
  assign n26626 = n26625 ^ n13358 ^ n10568 ;
  assign n26627 = ~n1981 & n21752 ;
  assign n26628 = ~n686 & n26627 ;
  assign n26629 = ( n11132 & n26626 ) | ( n11132 & ~n26628 ) | ( n26626 & ~n26628 ) ;
  assign n26630 = n17801 ^ n12588 ^ n4230 ;
  assign n26631 = n14913 ^ n8600 ^ 1'b0 ;
  assign n26632 = n7862 & ~n26631 ;
  assign n26633 = n26632 ^ n21698 ^ 1'b0 ;
  assign n26634 = n26633 ^ n5329 ^ 1'b0 ;
  assign n26635 = ( n5252 & n6680 ) | ( n5252 & n26634 ) | ( n6680 & n26634 ) ;
  assign n26637 = n12972 ^ n11925 ^ n1624 ;
  assign n26636 = n15808 & ~n20060 ;
  assign n26638 = n26637 ^ n26636 ^ 1'b0 ;
  assign n26641 = n6028 ^ n3987 ^ n3583 ;
  assign n26639 = ( n1289 & n15976 ) | ( n1289 & n17804 ) | ( n15976 & n17804 ) ;
  assign n26640 = n26639 ^ n15898 ^ n7716 ;
  assign n26642 = n26641 ^ n26640 ^ 1'b0 ;
  assign n26643 = n26638 & n26642 ;
  assign n26644 = n6629 & ~n26643 ;
  assign n26645 = n3353 & n18516 ;
  assign n26646 = n22064 & n26645 ;
  assign n26647 = n26646 ^ n15347 ^ n3360 ;
  assign n26648 = n26647 ^ n17699 ^ n13645 ;
  assign n26649 = n26648 ^ n23905 ^ n11603 ;
  assign n26650 = ~n18317 & n26649 ;
  assign n26651 = n1208 ^ n1049 ^ 1'b0 ;
  assign n26652 = ( n4358 & n25375 ) | ( n4358 & ~n26651 ) | ( n25375 & ~n26651 ) ;
  assign n26653 = ( ~n11252 & n19226 ) | ( ~n11252 & n26652 ) | ( n19226 & n26652 ) ;
  assign n26654 = ~n18644 & n26653 ;
  assign n26655 = n18422 & n26654 ;
  assign n26656 = n26655 ^ n24585 ^ n363 ;
  assign n26657 = n26656 ^ n19072 ^ n7150 ;
  assign n26658 = n13580 ^ n2519 ^ 1'b0 ;
  assign n26659 = n14480 & ~n26658 ;
  assign n26660 = ( n3509 & n22642 ) | ( n3509 & n26659 ) | ( n22642 & n26659 ) ;
  assign n26664 = n14155 ^ n5174 ^ n4345 ;
  assign n26661 = n13320 ^ n1700 ^ n464 ;
  assign n26662 = n26661 ^ n23751 ^ n11518 ;
  assign n26663 = n6121 & ~n26662 ;
  assign n26665 = n26664 ^ n26663 ^ 1'b0 ;
  assign n26666 = ( ~n989 & n5497 ) | ( ~n989 & n10444 ) | ( n5497 & n10444 ) ;
  assign n26667 = ( n7763 & n14637 ) | ( n7763 & n16785 ) | ( n14637 & n16785 ) ;
  assign n26668 = n26667 ^ n16161 ^ n10817 ;
  assign n26669 = n5045 & ~n15979 ;
  assign n26670 = n26669 ^ n12082 ^ n6324 ;
  assign n26671 = ( n8095 & n10731 ) | ( n8095 & ~n20426 ) | ( n10731 & ~n20426 ) ;
  assign n26672 = ( ~n11641 & n22788 ) | ( ~n11641 & n26671 ) | ( n22788 & n26671 ) ;
  assign n26673 = n5021 & ~n7582 ;
  assign n26674 = n26673 ^ n12462 ^ 1'b0 ;
  assign n26675 = ( n26670 & ~n26672 ) | ( n26670 & n26674 ) | ( ~n26672 & n26674 ) ;
  assign n26676 = n1575 & n13626 ;
  assign n26677 = ~n4047 & n26676 ;
  assign n26678 = ( n7860 & n11270 ) | ( n7860 & n15066 ) | ( n11270 & n15066 ) ;
  assign n26679 = n26678 ^ n22319 ^ n6405 ;
  assign n26680 = n9257 & ~n21913 ;
  assign n26681 = n9200 ^ n8167 ^ n5871 ;
  assign n26682 = n26681 ^ n17227 ^ n16097 ;
  assign n26688 = n1559 & n21899 ;
  assign n26689 = n26688 ^ n22218 ^ 1'b0 ;
  assign n26687 = n9811 ^ n5983 ^ 1'b0 ;
  assign n26683 = n1028 ^ n533 ^ n346 ;
  assign n26684 = ( ~n781 & n1386 ) | ( ~n781 & n26683 ) | ( n1386 & n26683 ) ;
  assign n26685 = ( n436 & n10499 ) | ( n436 & ~n24849 ) | ( n10499 & ~n24849 ) ;
  assign n26686 = ( ~n11074 & n26684 ) | ( ~n11074 & n26685 ) | ( n26684 & n26685 ) ;
  assign n26690 = n26689 ^ n26687 ^ n26686 ;
  assign n26691 = n26682 | n26690 ;
  assign n26692 = n26691 ^ n24604 ^ n15906 ;
  assign n26693 = n3668 | n7136 ;
  assign n26694 = ( n6505 & n19046 ) | ( n6505 & ~n26693 ) | ( n19046 & ~n26693 ) ;
  assign n26695 = ( n6195 & n7722 ) | ( n6195 & ~n11604 ) | ( n7722 & ~n11604 ) ;
  assign n26696 = ( n1423 & n26694 ) | ( n1423 & ~n26695 ) | ( n26694 & ~n26695 ) ;
  assign n26697 = ~n5461 & n8352 ;
  assign n26698 = n26697 ^ n262 ^ 1'b0 ;
  assign n26699 = n9702 & ~n12721 ;
  assign n26700 = ( ~n18564 & n26698 ) | ( ~n18564 & n26699 ) | ( n26698 & n26699 ) ;
  assign n26701 = ( x121 & n15412 ) | ( x121 & ~n26700 ) | ( n15412 & ~n26700 ) ;
  assign n26702 = n26701 ^ n4023 ^ 1'b0 ;
  assign n26703 = n26702 ^ n17420 ^ n546 ;
  assign n26704 = n26703 ^ n12523 ^ n1069 ;
  assign n26705 = n26282 ^ n9320 ^ n4710 ;
  assign n26706 = ( n3633 & n5081 ) | ( n3633 & ~n19953 ) | ( n5081 & ~n19953 ) ;
  assign n26712 = n16568 ^ n13083 ^ 1'b0 ;
  assign n26713 = ( n3884 & n17000 ) | ( n3884 & n26712 ) | ( n17000 & n26712 ) ;
  assign n26707 = n2635 & ~n3726 ;
  assign n26708 = n26707 ^ n6553 ^ 1'b0 ;
  assign n26709 = n26708 ^ n17651 ^ n8049 ;
  assign n26710 = ~n13440 & n26709 ;
  assign n26711 = n7681 & n26710 ;
  assign n26714 = n26713 ^ n26711 ^ 1'b0 ;
  assign n26721 = n3963 ^ n2613 ^ n1551 ;
  assign n26722 = n4296 & ~n26721 ;
  assign n26723 = n11867 | n13054 ;
  assign n26724 = n26722 | n26723 ;
  assign n26725 = n26724 ^ n6389 ^ n5233 ;
  assign n26719 = n7302 ^ n6915 ^ n3107 ;
  assign n26720 = n26719 ^ n15811 ^ n13817 ;
  assign n26715 = n13770 ^ n13236 ^ n6491 ;
  assign n26716 = n10559 & n25856 ;
  assign n26717 = n26716 ^ n11758 ^ 1'b0 ;
  assign n26718 = ( n17944 & ~n26715 ) | ( n17944 & n26717 ) | ( ~n26715 & n26717 ) ;
  assign n26726 = n26725 ^ n26720 ^ n26718 ;
  assign n26727 = n16467 & n17608 ;
  assign n26728 = n23468 ^ n21665 ^ n3326 ;
  assign n26730 = n14178 | n24896 ;
  assign n26731 = n23593 & ~n26730 ;
  assign n26729 = n7045 | n23248 ;
  assign n26732 = n26731 ^ n26729 ^ 1'b0 ;
  assign n26733 = n26732 ^ n12653 ^ x53 ;
  assign n26734 = n8732 ^ n259 ^ 1'b0 ;
  assign n26735 = n20692 & ~n26734 ;
  assign n26736 = n26735 ^ n23549 ^ n11292 ;
  assign n26744 = n10554 | n21098 ;
  assign n26745 = n6587 & ~n26744 ;
  assign n26737 = n18667 ^ n15921 ^ 1'b0 ;
  assign n26738 = n9257 & ~n26737 ;
  assign n26739 = n26738 ^ n10499 ^ n2773 ;
  assign n26740 = n26739 ^ n22770 ^ n3682 ;
  assign n26741 = n26740 ^ n21363 ^ n17864 ;
  assign n26742 = n22203 & ~n26741 ;
  assign n26743 = ~n3894 & n26742 ;
  assign n26746 = n26745 ^ n26743 ^ n14790 ;
  assign n26747 = ~n8053 & n23926 ;
  assign n26748 = ( n4701 & ~n5732 ) | ( n4701 & n10269 ) | ( ~n5732 & n10269 ) ;
  assign n26749 = n26748 ^ n21319 ^ n4850 ;
  assign n26750 = ~n17139 & n26749 ;
  assign n26751 = n22764 ^ n11269 ^ n3072 ;
  assign n26752 = n26751 ^ n4747 ^ n4732 ;
  assign n26753 = ( ~x243 & n263 ) | ( ~x243 & n26752 ) | ( n263 & n26752 ) ;
  assign n26754 = n23349 ^ n21781 ^ n18442 ;
  assign n26755 = ~n13608 & n19576 ;
  assign n26756 = n26755 ^ n24038 ^ 1'b0 ;
  assign n26760 = ( n9168 & n15094 ) | ( n9168 & n19313 ) | ( n15094 & n19313 ) ;
  assign n26757 = n3060 | n7609 ;
  assign n26758 = n1738 & ~n26757 ;
  assign n26759 = n26758 ^ n24906 ^ n20028 ;
  assign n26761 = n26760 ^ n26759 ^ n7803 ;
  assign n26765 = n20412 ^ n18026 ^ 1'b0 ;
  assign n26766 = ( n20032 & n22637 ) | ( n20032 & ~n26765 ) | ( n22637 & ~n26765 ) ;
  assign n26762 = n3826 & n8778 ;
  assign n26763 = n26762 ^ n8504 ^ 1'b0 ;
  assign n26764 = ( n13845 & n26380 ) | ( n13845 & ~n26763 ) | ( n26380 & ~n26763 ) ;
  assign n26767 = n26766 ^ n26764 ^ n21310 ;
  assign n26768 = n13614 ^ n7114 ^ n868 ;
  assign n26769 = n4489 & ~n9512 ;
  assign n26770 = ( n2467 & ~n9639 ) | ( n2467 & n17077 ) | ( ~n9639 & n17077 ) ;
  assign n26771 = ( ~n6936 & n13388 ) | ( ~n6936 & n23921 ) | ( n13388 & n23921 ) ;
  assign n26772 = n7983 ^ n4684 ^ 1'b0 ;
  assign n26773 = n14057 ^ n3942 ^ 1'b0 ;
  assign n26774 = n26773 ^ n15856 ^ 1'b0 ;
  assign n26775 = ~n26772 & n26774 ;
  assign n26776 = n2832 ^ n2167 ^ 1'b0 ;
  assign n26779 = n9010 ^ n5956 ^ 1'b0 ;
  assign n26777 = n24110 ^ n7128 ^ n2241 ;
  assign n26778 = ( n8194 & ~n23984 ) | ( n8194 & n26777 ) | ( ~n23984 & n26777 ) ;
  assign n26780 = n26779 ^ n26778 ^ 1'b0 ;
  assign n26781 = n3619 | n25603 ;
  assign n26782 = n26781 ^ n3660 ^ 1'b0 ;
  assign n26783 = n17804 ^ n5943 ^ 1'b0 ;
  assign n26784 = n26351 ^ n21348 ^ n14739 ;
  assign n26785 = n26784 ^ n17754 ^ n16836 ;
  assign n26786 = n26783 & ~n26785 ;
  assign n26787 = ( n13621 & n26782 ) | ( n13621 & n26786 ) | ( n26782 & n26786 ) ;
  assign n26788 = ( n11996 & ~n12992 ) | ( n11996 & n17513 ) | ( ~n12992 & n17513 ) ;
  assign n26789 = n4337 | n10800 ;
  assign n26790 = ( n8450 & n15615 ) | ( n8450 & n26789 ) | ( n15615 & n26789 ) ;
  assign n26791 = n12945 ^ n9849 ^ n538 ;
  assign n26792 = ( ~n1785 & n20508 ) | ( ~n1785 & n26791 ) | ( n20508 & n26791 ) ;
  assign n26793 = n7342 ^ n1616 ^ 1'b0 ;
  assign n26794 = n9042 & ~n26793 ;
  assign n26795 = n26794 ^ n16920 ^ n4164 ;
  assign n26796 = n26795 ^ n9352 ^ 1'b0 ;
  assign n26797 = n15306 ^ n10230 ^ 1'b0 ;
  assign n26806 = ~n3981 & n9695 ;
  assign n26800 = n6574 ^ n5208 ^ n3802 ;
  assign n26798 = n21373 ^ n5310 ^ n894 ;
  assign n26799 = ~n4915 & n26798 ;
  assign n26801 = n26800 ^ n26799 ^ 1'b0 ;
  assign n26802 = n26606 ^ n26576 ^ n2827 ;
  assign n26803 = ( n13041 & n26801 ) | ( n13041 & n26802 ) | ( n26801 & n26802 ) ;
  assign n26804 = n26803 ^ n21355 ^ n9091 ;
  assign n26805 = n26804 ^ n19300 ^ n13071 ;
  assign n26807 = n26806 ^ n26805 ^ 1'b0 ;
  assign n26808 = n25944 ^ n25452 ^ 1'b0 ;
  assign n26809 = ~n5276 & n26808 ;
  assign n26810 = n22261 ^ n13612 ^ n3936 ;
  assign n26811 = ( n862 & n16848 ) | ( n862 & ~n21562 ) | ( n16848 & ~n21562 ) ;
  assign n26812 = n24853 ^ n10276 ^ n2077 ;
  assign n26813 = n26812 ^ n16556 ^ 1'b0 ;
  assign n26814 = n15717 & n26813 ;
  assign n26815 = n26814 ^ n12327 ^ 1'b0 ;
  assign n26816 = n26811 & ~n26815 ;
  assign n26817 = n25166 ^ n9185 ^ 1'b0 ;
  assign n26818 = n25909 ^ n7343 ^ n2827 ;
  assign n26819 = ( n4432 & n8628 ) | ( n4432 & n26818 ) | ( n8628 & n26818 ) ;
  assign n26820 = n20120 ^ n19930 ^ n1678 ;
  assign n26821 = n26820 ^ n22853 ^ n13755 ;
  assign n26822 = n1594 & n1940 ;
  assign n26828 = n25766 ^ n16391 ^ n12315 ;
  assign n26825 = ( n5734 & ~n9828 ) | ( n5734 & n16933 ) | ( ~n9828 & n16933 ) ;
  assign n26824 = n17834 ^ n11081 ^ 1'b0 ;
  assign n26826 = n26825 ^ n26824 ^ n6153 ;
  assign n26827 = ( n7435 & ~n15383 ) | ( n7435 & n26826 ) | ( ~n15383 & n26826 ) ;
  assign n26829 = n26828 ^ n26827 ^ n6616 ;
  assign n26823 = n26759 ^ n19160 ^ n18453 ;
  assign n26830 = n26829 ^ n26823 ^ n18278 ;
  assign n26833 = ~n3296 & n8272 ;
  assign n26831 = n13070 & ~n19901 ;
  assign n26832 = n25140 & n26831 ;
  assign n26834 = n26833 ^ n26832 ^ n25771 ;
  assign n26835 = n20988 ^ n4816 ^ 1'b0 ;
  assign n26836 = n3168 | n5380 ;
  assign n26837 = n26836 ^ n7099 ^ 1'b0 ;
  assign n26838 = n4247 ^ n293 ^ 1'b0 ;
  assign n26839 = ( n5134 & ~n12897 ) | ( n5134 & n26838 ) | ( ~n12897 & n26838 ) ;
  assign n26840 = ~n1870 & n14279 ;
  assign n26841 = ~n11209 & n26840 ;
  assign n26848 = n14857 ^ n8341 ^ 1'b0 ;
  assign n26849 = n17392 & n26848 ;
  assign n26850 = n26849 ^ n5043 ^ 1'b0 ;
  assign n26842 = n2594 ^ x127 ^ 1'b0 ;
  assign n26843 = n21684 ^ n8298 ^ x83 ;
  assign n26844 = n26843 ^ n8616 ^ n6249 ;
  assign n26845 = n25995 ^ n13613 ^ n11955 ;
  assign n26846 = ( n6593 & n26844 ) | ( n6593 & n26845 ) | ( n26844 & n26845 ) ;
  assign n26847 = ( n23037 & n26842 ) | ( n23037 & n26846 ) | ( n26842 & n26846 ) ;
  assign n26851 = n26850 ^ n26847 ^ 1'b0 ;
  assign n26852 = n10685 ^ n7514 ^ 1'b0 ;
  assign n26853 = n3160 | n26852 ;
  assign n26854 = ( ~n3880 & n17917 ) | ( ~n3880 & n26853 ) | ( n17917 & n26853 ) ;
  assign n26860 = n15398 ^ n7900 ^ n7090 ;
  assign n26859 = ( n6301 & n11424 ) | ( n6301 & ~n20562 ) | ( n11424 & ~n20562 ) ;
  assign n26861 = n26860 ^ n26859 ^ n6218 ;
  assign n26857 = n14936 ^ n5464 ^ 1'b0 ;
  assign n26858 = ( n5905 & ~n24367 ) | ( n5905 & n26857 ) | ( ~n24367 & n26857 ) ;
  assign n26862 = n26861 ^ n26858 ^ n22131 ;
  assign n26863 = n26862 ^ n18849 ^ n2090 ;
  assign n26855 = ~n9466 & n26653 ;
  assign n26856 = ~n19442 & n26855 ;
  assign n26864 = n26863 ^ n26856 ^ n17992 ;
  assign n26865 = n17609 ^ n5024 ^ 1'b0 ;
  assign n26866 = n8773 & ~n26865 ;
  assign n26867 = n6560 & n14974 ;
  assign n26868 = n15888 & n26867 ;
  assign n26869 = n6333 ^ n2289 ^ 1'b0 ;
  assign n26870 = n26869 ^ n7732 ^ n1965 ;
  assign n26871 = ( n16799 & n24384 ) | ( n16799 & ~n26870 ) | ( n24384 & ~n26870 ) ;
  assign n26872 = ( n1048 & n3583 ) | ( n1048 & n11911 ) | ( n3583 & n11911 ) ;
  assign n26873 = n26872 ^ n8181 ^ n5276 ;
  assign n26874 = ~n14830 & n26873 ;
  assign n26875 = n12334 ^ n10292 ^ n2753 ;
  assign n26877 = n1597 ^ n982 ^ n810 ;
  assign n26878 = n26877 ^ n1427 ^ n276 ;
  assign n26876 = ( ~n3735 & n7121 ) | ( ~n3735 & n13853 ) | ( n7121 & n13853 ) ;
  assign n26879 = n26878 ^ n26876 ^ n6886 ;
  assign n26880 = n26879 ^ n11957 ^ n3834 ;
  assign n26881 = n5724 ^ n4862 ^ n3264 ;
  assign n26882 = ( n9129 & ~n10110 ) | ( n9129 & n18802 ) | ( ~n10110 & n18802 ) ;
  assign n26883 = n19376 ^ n8879 ^ 1'b0 ;
  assign n26884 = ( n11274 & n26882 ) | ( n11274 & n26883 ) | ( n26882 & n26883 ) ;
  assign n26885 = ( n7145 & n26881 ) | ( n7145 & n26884 ) | ( n26881 & n26884 ) ;
  assign n26886 = n26885 ^ n13438 ^ 1'b0 ;
  assign n26887 = ( n26377 & n26880 ) | ( n26377 & n26886 ) | ( n26880 & n26886 ) ;
  assign n26888 = n12115 ^ n8476 ^ n3791 ;
  assign n26889 = n7775 ^ n1813 ^ n548 ;
  assign n26890 = ( n14895 & n15979 ) | ( n14895 & ~n26889 ) | ( n15979 & ~n26889 ) ;
  assign n26891 = ( n13552 & n26888 ) | ( n13552 & ~n26890 ) | ( n26888 & ~n26890 ) ;
  assign n26892 = ( ~n15509 & n21087 ) | ( ~n15509 & n26891 ) | ( n21087 & n26891 ) ;
  assign n26893 = n12844 ^ n7736 ^ 1'b0 ;
  assign n26894 = n5943 & ~n26893 ;
  assign n26899 = ( n5490 & ~n14347 ) | ( n5490 & n19326 ) | ( ~n14347 & n19326 ) ;
  assign n26895 = n5822 & ~n9660 ;
  assign n26896 = n10327 & n26895 ;
  assign n26897 = n9422 | n26896 ;
  assign n26898 = n25467 | n26897 ;
  assign n26900 = n26899 ^ n26898 ^ 1'b0 ;
  assign n26901 = n20186 & ~n26900 ;
  assign n26902 = n26901 ^ n3390 ^ 1'b0 ;
  assign n26903 = ~n11887 & n18228 ;
  assign n26904 = ( n7368 & n23869 ) | ( n7368 & ~n26903 ) | ( n23869 & ~n26903 ) ;
  assign n26905 = ~n16934 & n25426 ;
  assign n26906 = n5198 ^ n691 ^ 1'b0 ;
  assign n26909 = ( ~n728 & n9933 ) | ( ~n728 & n24969 ) | ( n9933 & n24969 ) ;
  assign n26907 = ( ~n1160 & n1875 ) | ( ~n1160 & n10271 ) | ( n1875 & n10271 ) ;
  assign n26908 = ( ~n12063 & n20615 ) | ( ~n12063 & n26907 ) | ( n20615 & n26907 ) ;
  assign n26910 = n26909 ^ n26908 ^ n4806 ;
  assign n26911 = ( n16767 & ~n26906 ) | ( n16767 & n26910 ) | ( ~n26906 & n26910 ) ;
  assign n26912 = n5118 ^ n3427 ^ n3194 ;
  assign n26913 = ( n13865 & n23494 ) | ( n13865 & n26912 ) | ( n23494 & n26912 ) ;
  assign n26914 = n26913 ^ n24800 ^ n8745 ;
  assign n26916 = n6936 | n7177 ;
  assign n26917 = n8017 & ~n26916 ;
  assign n26918 = n2296 | n10144 ;
  assign n26919 = n9929 | n26918 ;
  assign n26920 = ( n3880 & n11996 ) | ( n3880 & ~n21134 ) | ( n11996 & ~n21134 ) ;
  assign n26921 = ( n26917 & n26919 ) | ( n26917 & ~n26920 ) | ( n26919 & ~n26920 ) ;
  assign n26922 = n26921 ^ n23498 ^ n21062 ;
  assign n26915 = n1365 & n2096 ;
  assign n26923 = n26922 ^ n26915 ^ 1'b0 ;
  assign n26924 = n12977 ^ n8933 ^ 1'b0 ;
  assign n26925 = n1711 | n26924 ;
  assign n26929 = n22134 ^ n5740 ^ n3691 ;
  assign n26926 = n9877 | n18324 ;
  assign n26927 = n26926 ^ n855 ^ 1'b0 ;
  assign n26928 = ( ~x242 & n1692 ) | ( ~x242 & n26927 ) | ( n1692 & n26927 ) ;
  assign n26930 = n26929 ^ n26928 ^ n9926 ;
  assign n26931 = ( n21023 & n26925 ) | ( n21023 & ~n26930 ) | ( n26925 & ~n26930 ) ;
  assign n26932 = n26931 ^ n9830 ^ 1'b0 ;
  assign n26933 = n2604 & n26932 ;
  assign n26934 = n1246 & n25186 ;
  assign n26935 = n26934 ^ n15953 ^ 1'b0 ;
  assign n26936 = ( n13599 & ~n15762 ) | ( n13599 & n21113 ) | ( ~n15762 & n21113 ) ;
  assign n26937 = ( n5153 & n10959 ) | ( n5153 & n26936 ) | ( n10959 & n26936 ) ;
  assign n26938 = n10651 ^ n3126 ^ n1252 ;
  assign n26939 = ~n15080 & n24054 ;
  assign n26940 = n26939 ^ n19113 ^ 1'b0 ;
  assign n26941 = ( n9486 & ~n26938 ) | ( n9486 & n26940 ) | ( ~n26938 & n26940 ) ;
  assign n26947 = n10374 ^ n2884 ^ n2535 ;
  assign n26948 = n26947 ^ n5085 ^ n1555 ;
  assign n26945 = n23770 ^ n16060 ^ n1805 ;
  assign n26942 = n13778 ^ n8154 ^ 1'b0 ;
  assign n26943 = n26942 ^ n19208 ^ n1407 ;
  assign n26944 = ( n2358 & ~n13167 ) | ( n2358 & n26943 ) | ( ~n13167 & n26943 ) ;
  assign n26946 = n26945 ^ n26944 ^ n22193 ;
  assign n26949 = n26948 ^ n26946 ^ n3819 ;
  assign n26951 = ( ~n1782 & n14431 ) | ( ~n1782 & n21791 ) | ( n14431 & n21791 ) ;
  assign n26950 = n25034 ^ n18148 ^ n16171 ;
  assign n26952 = n26951 ^ n26950 ^ n4779 ;
  assign n26953 = ( n4209 & ~n10867 ) | ( n4209 & n19646 ) | ( ~n10867 & n19646 ) ;
  assign n26954 = n26953 ^ n25597 ^ 1'b0 ;
  assign n26955 = ~n5718 & n18918 ;
  assign n26956 = ( n10435 & ~n16418 ) | ( n10435 & n26955 ) | ( ~n16418 & n26955 ) ;
  assign n26957 = x131 & ~n4882 ;
  assign n26958 = n21300 ^ n15159 ^ n7988 ;
  assign n26959 = ( ~n13245 & n26957 ) | ( ~n13245 & n26958 ) | ( n26957 & n26958 ) ;
  assign n26960 = ~n4489 & n26096 ;
  assign n26961 = n17675 & n26960 ;
  assign n26962 = ( n26956 & n26959 ) | ( n26956 & n26961 ) | ( n26959 & n26961 ) ;
  assign n26963 = n17449 ^ n5970 ^ 1'b0 ;
  assign n26964 = n2572 & ~n19952 ;
  assign n26965 = n26964 ^ n10564 ^ 1'b0 ;
  assign n26966 = ( ~n1445 & n2794 ) | ( ~n1445 & n26965 ) | ( n2794 & n26965 ) ;
  assign n26967 = ~n5709 & n21457 ;
  assign n26968 = ~n14196 & n26967 ;
  assign n26969 = ~n999 & n26968 ;
  assign n26970 = n667 | n7534 ;
  assign n26971 = n26970 ^ n3605 ^ 1'b0 ;
  assign n26972 = n8543 & n26971 ;
  assign n26973 = n26972 ^ n23922 ^ 1'b0 ;
  assign n26974 = ( ~n2516 & n4712 ) | ( ~n2516 & n19378 ) | ( n4712 & n19378 ) ;
  assign n26975 = n4520 & n5029 ;
  assign n26976 = ~n9611 & n26975 ;
  assign n26977 = n13976 ^ n11147 ^ n2023 ;
  assign n26978 = ~n9094 & n26977 ;
  assign n26979 = ~n9296 & n26978 ;
  assign n26980 = ( n17812 & n26976 ) | ( n17812 & ~n26979 ) | ( n26976 & ~n26979 ) ;
  assign n26981 = ( n1191 & ~n26974 ) | ( n1191 & n26980 ) | ( ~n26974 & n26980 ) ;
  assign n26982 = ( n15432 & n23524 ) | ( n15432 & n25486 ) | ( n23524 & n25486 ) ;
  assign n26983 = n12097 ^ n11525 ^ 1'b0 ;
  assign n26984 = n10554 | n26983 ;
  assign n26985 = n9126 & n18059 ;
  assign n26986 = n10865 & n26985 ;
  assign n26987 = n26986 ^ n19087 ^ n17889 ;
  assign n26988 = n973 | n26987 ;
  assign n26989 = n26988 ^ n25091 ^ 1'b0 ;
  assign n26990 = n21933 ^ n16933 ^ 1'b0 ;
  assign n26991 = ( n7193 & ~n8153 ) | ( n7193 & n17917 ) | ( ~n8153 & n17917 ) ;
  assign n26992 = n26408 | n26991 ;
  assign n26993 = n26992 ^ n3648 ^ 1'b0 ;
  assign n26994 = ( n4919 & n10846 ) | ( n4919 & ~n13458 ) | ( n10846 & ~n13458 ) ;
  assign n26995 = n21702 & ~n26994 ;
  assign n26996 = n26995 ^ n22226 ^ 1'b0 ;
  assign n26997 = ( ~n2077 & n7945 ) | ( ~n2077 & n18568 ) | ( n7945 & n18568 ) ;
  assign n26998 = ( ~n1885 & n13213 ) | ( ~n1885 & n17589 ) | ( n13213 & n17589 ) ;
  assign n26999 = n26998 ^ n22777 ^ n2783 ;
  assign n27000 = n26667 | n26999 ;
  assign n27001 = n18801 | n27000 ;
  assign n27002 = n4916 & n27001 ;
  assign n27003 = n14185 & n27002 ;
  assign n27004 = n27003 ^ n25173 ^ n24124 ;
  assign n27005 = ( n8975 & n10196 ) | ( n8975 & ~n22553 ) | ( n10196 & ~n22553 ) ;
  assign n27006 = ( ~n22913 & n23162 ) | ( ~n22913 & n27005 ) | ( n23162 & n27005 ) ;
  assign n27007 = ~n14762 & n21864 ;
  assign n27008 = n27007 ^ n2307 ^ 1'b0 ;
  assign n27009 = n6434 & n9462 ;
  assign n27011 = n22881 ^ n7832 ^ n5071 ;
  assign n27012 = n2587 | n27011 ;
  assign n27013 = n16768 & ~n27012 ;
  assign n27014 = ( n9278 & ~n9636 ) | ( n9278 & n27013 ) | ( ~n9636 & n27013 ) ;
  assign n27010 = n18659 ^ n17289 ^ n10795 ;
  assign n27015 = n27014 ^ n27010 ^ n9972 ;
  assign n27016 = n23115 ^ n9811 ^ n2190 ;
  assign n27017 = n20013 ^ n16459 ^ n11867 ;
  assign n27018 = ( n4847 & ~n27016 ) | ( n4847 & n27017 ) | ( ~n27016 & n27017 ) ;
  assign n27019 = ( n11902 & n15448 ) | ( n11902 & n26772 ) | ( n15448 & n26772 ) ;
  assign n27020 = ( n16705 & n21264 ) | ( n16705 & n27019 ) | ( n21264 & n27019 ) ;
  assign n27021 = ( n1877 & ~n20807 ) | ( n1877 & n27020 ) | ( ~n20807 & n27020 ) ;
  assign n27022 = n17137 ^ n11166 ^ n3695 ;
  assign n27023 = n27022 ^ n3486 ^ 1'b0 ;
  assign n27024 = n10339 & n27023 ;
  assign n27025 = n20764 ^ n14285 ^ n9147 ;
  assign n27026 = ( ~n9380 & n15894 ) | ( ~n9380 & n27025 ) | ( n15894 & n27025 ) ;
  assign n27027 = n840 & n2208 ;
  assign n27028 = n27027 ^ n15773 ^ 1'b0 ;
  assign n27029 = n27026 & n27028 ;
  assign n27030 = n19266 ^ n7898 ^ n4055 ;
  assign n27031 = n16951 ^ n10857 ^ n9633 ;
  assign n27032 = n27031 ^ n2545 ^ 1'b0 ;
  assign n27033 = ( n10496 & n27030 ) | ( n10496 & n27032 ) | ( n27030 & n27032 ) ;
  assign n27034 = n20368 ^ n3318 ^ 1'b0 ;
  assign n27035 = ~n13041 & n27034 ;
  assign n27036 = n2312 & n4920 ;
  assign n27037 = ~n27035 & n27036 ;
  assign n27038 = ( ~n9067 & n15437 ) | ( ~n9067 & n27037 ) | ( n15437 & n27037 ) ;
  assign n27045 = n1055 | n13670 ;
  assign n27046 = ( n1294 & n11349 ) | ( n1294 & ~n27045 ) | ( n11349 & ~n27045 ) ;
  assign n27040 = ( n5574 & n20956 ) | ( n5574 & n24230 ) | ( n20956 & n24230 ) ;
  assign n27041 = n19491 & n25867 ;
  assign n27042 = n27041 ^ n15557 ^ 1'b0 ;
  assign n27043 = ( n10042 & ~n27040 ) | ( n10042 & n27042 ) | ( ~n27040 & n27042 ) ;
  assign n27039 = n5909 ^ n4536 ^ n4213 ;
  assign n27044 = n27043 ^ n27039 ^ n18627 ;
  assign n27047 = n27046 ^ n27044 ^ n14390 ;
  assign n27048 = n19146 ^ n19124 ^ n3388 ;
  assign n27049 = n7224 & n8643 ;
  assign n27050 = n9662 ^ n1373 ^ n721 ;
  assign n27051 = ( ~n15450 & n21201 ) | ( ~n15450 & n27050 ) | ( n21201 & n27050 ) ;
  assign n27052 = ( ~n4272 & n6232 ) | ( ~n4272 & n27051 ) | ( n6232 & n27051 ) ;
  assign n27053 = ( n1796 & ~n2949 ) | ( n1796 & n16470 ) | ( ~n2949 & n16470 ) ;
  assign n27054 = n21447 & n24684 ;
  assign n27055 = ~n4239 & n27054 ;
  assign n27056 = n27055 ^ n24712 ^ 1'b0 ;
  assign n27057 = n5355 & ~n27056 ;
  assign n27058 = n27057 ^ n7581 ^ 1'b0 ;
  assign n27059 = ~n27053 & n27058 ;
  assign n27060 = n27059 ^ n16998 ^ x243 ;
  assign n27061 = n27060 ^ n16093 ^ n12073 ;
  assign n27062 = n7708 ^ n4567 ^ x134 ;
  assign n27063 = n12715 ^ n8797 ^ n6069 ;
  assign n27064 = ( ~n15987 & n27062 ) | ( ~n15987 & n27063 ) | ( n27062 & n27063 ) ;
  assign n27065 = ( n2687 & ~n5679 ) | ( n2687 & n10421 ) | ( ~n5679 & n10421 ) ;
  assign n27066 = n27065 ^ n2894 ^ 1'b0 ;
  assign n27067 = n8773 | n25051 ;
  assign n27068 = n14206 ^ n9090 ^ 1'b0 ;
  assign n27069 = n17663 | n27068 ;
  assign n27070 = n27069 ^ n6707 ^ n420 ;
  assign n27071 = ( n3335 & n19665 ) | ( n3335 & ~n27070 ) | ( n19665 & ~n27070 ) ;
  assign n27072 = ( ~n3612 & n7259 ) | ( ~n3612 & n16992 ) | ( n7259 & n16992 ) ;
  assign n27073 = ( n6913 & n25557 ) | ( n6913 & n27072 ) | ( n25557 & n27072 ) ;
  assign n27074 = n7578 | n16651 ;
  assign n27075 = n27074 ^ n23181 ^ n21649 ;
  assign n27076 = ~x33 & n7050 ;
  assign n27077 = ( n6430 & n6987 ) | ( n6430 & n20341 ) | ( n6987 & n20341 ) ;
  assign n27078 = n10473 & n20211 ;
  assign n27079 = n27078 ^ n4152 ^ 1'b0 ;
  assign n27080 = ( ~n12467 & n18513 ) | ( ~n12467 & n27079 ) | ( n18513 & n27079 ) ;
  assign n27081 = n17939 & n18908 ;
  assign n27082 = ~n26092 & n27081 ;
  assign n27083 = ( ~n27077 & n27080 ) | ( ~n27077 & n27082 ) | ( n27080 & n27082 ) ;
  assign n27084 = ( x206 & n1963 ) | ( x206 & n4256 ) | ( n1963 & n4256 ) ;
  assign n27085 = ~n8253 & n27084 ;
  assign n27086 = n27085 ^ n13392 ^ 1'b0 ;
  assign n27087 = ( n2595 & n5251 ) | ( n2595 & ~n17294 ) | ( n5251 & ~n17294 ) ;
  assign n27088 = n27087 ^ n18498 ^ 1'b0 ;
  assign n27089 = ~n18291 & n27088 ;
  assign n27090 = ( n23123 & n27086 ) | ( n23123 & ~n27089 ) | ( n27086 & ~n27089 ) ;
  assign n27092 = ( n2487 & n2740 ) | ( n2487 & n9185 ) | ( n2740 & n9185 ) ;
  assign n27091 = n20537 & ~n23553 ;
  assign n27093 = n27092 ^ n27091 ^ 1'b0 ;
  assign n27094 = ( n18409 & n27090 ) | ( n18409 & ~n27093 ) | ( n27090 & ~n27093 ) ;
  assign n27095 = n17380 ^ n16248 ^ n7447 ;
  assign n27096 = n12233 ^ n5045 ^ n1809 ;
  assign n27097 = n13605 ^ n11022 ^ 1'b0 ;
  assign n27098 = n18547 ^ n15807 ^ n11654 ;
  assign n27099 = n3531 ^ n1924 ^ n1840 ;
  assign n27100 = n27099 ^ n5448 ^ n1873 ;
  assign n27102 = n24325 ^ n10666 ^ 1'b0 ;
  assign n27103 = n27102 ^ n21557 ^ n15052 ;
  assign n27101 = n8983 ^ n1041 ^ 1'b0 ;
  assign n27104 = n27103 ^ n27101 ^ 1'b0 ;
  assign n27105 = n659 & n6372 ;
  assign n27106 = n17026 & n27105 ;
  assign n27107 = n27106 ^ n8312 ^ 1'b0 ;
  assign n27108 = n4418 & ~n12931 ;
  assign n27109 = ( n9969 & n19069 ) | ( n9969 & ~n26077 ) | ( n19069 & ~n26077 ) ;
  assign n27110 = ~n9217 & n9637 ;
  assign n27111 = ~n10276 & n27110 ;
  assign n27112 = ( n6946 & n20617 ) | ( n6946 & ~n27111 ) | ( n20617 & ~n27111 ) ;
  assign n27113 = n27112 ^ n24203 ^ n3930 ;
  assign n27114 = n13376 | n21427 ;
  assign n27115 = n14319 ^ n11438 ^ 1'b0 ;
  assign n27117 = ( n4194 & n16338 ) | ( n4194 & ~n24945 ) | ( n16338 & ~n24945 ) ;
  assign n27118 = n27117 ^ n17137 ^ n7822 ;
  assign n27116 = n22026 ^ n18116 ^ 1'b0 ;
  assign n27119 = n27118 ^ n27116 ^ n4990 ;
  assign n27120 = n12811 | n27119 ;
  assign n27121 = ( ~n2727 & n27115 ) | ( ~n2727 & n27120 ) | ( n27115 & n27120 ) ;
  assign n27122 = n12026 ^ n8007 ^ 1'b0 ;
  assign n27123 = n9833 & n27122 ;
  assign n27124 = ( ~n9243 & n19691 ) | ( ~n9243 & n27123 ) | ( n19691 & n27123 ) ;
  assign n27125 = ( n1418 & ~n6432 ) | ( n1418 & n7535 ) | ( ~n6432 & n7535 ) ;
  assign n27126 = ( n18572 & n22528 ) | ( n18572 & n27125 ) | ( n22528 & n27125 ) ;
  assign n27127 = n27126 ^ n9519 ^ n8831 ;
  assign n27128 = n2384 ^ n1062 ^ 1'b0 ;
  assign n27129 = n27127 & n27128 ;
  assign n27130 = n27129 ^ n16408 ^ n1370 ;
  assign n27131 = ( n1366 & ~n20349 ) | ( n1366 & n27130 ) | ( ~n20349 & n27130 ) ;
  assign n27132 = n24030 ^ n12224 ^ 1'b0 ;
  assign n27133 = n12079 & n21756 ;
  assign n27134 = ( n6820 & ~n10920 ) | ( n6820 & n15114 ) | ( ~n10920 & n15114 ) ;
  assign n27135 = n27134 ^ n1296 ^ 1'b0 ;
  assign n27136 = n12452 & ~n27135 ;
  assign n27137 = ~n27133 & n27136 ;
  assign n27138 = n27137 ^ n18156 ^ 1'b0 ;
  assign n27139 = n1492 | n14518 ;
  assign n27140 = n27139 ^ n8397 ^ 1'b0 ;
  assign n27141 = ( ~n10599 & n10932 ) | ( ~n10599 & n18314 ) | ( n10932 & n18314 ) ;
  assign n27142 = ( n11351 & n19463 ) | ( n11351 & n27141 ) | ( n19463 & n27141 ) ;
  assign n27143 = ( n12995 & n14830 ) | ( n12995 & n27142 ) | ( n14830 & n27142 ) ;
  assign n27144 = ( n8394 & n15455 ) | ( n8394 & n20154 ) | ( n15455 & n20154 ) ;
  assign n27145 = n27144 ^ n24089 ^ n7795 ;
  assign n27146 = ( ~n7078 & n21705 ) | ( ~n7078 & n27145 ) | ( n21705 & n27145 ) ;
  assign n27147 = ( n927 & n3801 ) | ( n927 & n11612 ) | ( n3801 & n11612 ) ;
  assign n27148 = ( n13022 & n21083 ) | ( n13022 & ~n27147 ) | ( n21083 & ~n27147 ) ;
  assign n27149 = n1020 & n7165 ;
  assign n27150 = n27149 ^ n2426 ^ 1'b0 ;
  assign n27151 = n22950 ^ n4177 ^ 1'b0 ;
  assign n27152 = ( n2869 & ~n2912 ) | ( n2869 & n27151 ) | ( ~n2912 & n27151 ) ;
  assign n27153 = ( ~n2824 & n27150 ) | ( ~n2824 & n27152 ) | ( n27150 & n27152 ) ;
  assign n27154 = n10843 & ~n27153 ;
  assign n27155 = n13708 & n27154 ;
  assign n27163 = n1796 | n2615 ;
  assign n27162 = n4688 & ~n21774 ;
  assign n27156 = n2860 | n14597 ;
  assign n27157 = n27156 ^ n7217 ^ 1'b0 ;
  assign n27158 = n17275 & n27157 ;
  assign n27159 = n27158 ^ n5297 ^ 1'b0 ;
  assign n27160 = n27159 ^ n7029 ^ n549 ;
  assign n27161 = ( n14426 & n27115 ) | ( n14426 & ~n27160 ) | ( n27115 & ~n27160 ) ;
  assign n27164 = n27163 ^ n27162 ^ n27161 ;
  assign n27167 = ( x235 & n4743 ) | ( x235 & ~n6004 ) | ( n4743 & ~n6004 ) ;
  assign n27168 = n27167 ^ n6248 ^ n1649 ;
  assign n27169 = ( n18123 & n23921 ) | ( n18123 & ~n27168 ) | ( n23921 & ~n27168 ) ;
  assign n27165 = ( n11749 & n14238 ) | ( n11749 & ~n16792 ) | ( n14238 & ~n16792 ) ;
  assign n27166 = ~n20550 & n27165 ;
  assign n27170 = n27169 ^ n27166 ^ 1'b0 ;
  assign n27171 = ( ~n4355 & n4840 ) | ( ~n4355 & n24752 ) | ( n4840 & n24752 ) ;
  assign n27172 = n16862 ^ n14903 ^ n13500 ;
  assign n27173 = n27172 ^ n20178 ^ n2910 ;
  assign n27174 = n26483 ^ n19302 ^ x120 ;
  assign n27179 = n3700 & n6899 ;
  assign n27180 = ~n11746 & n27179 ;
  assign n27181 = ( n1501 & ~n4765 ) | ( n1501 & n27180 ) | ( ~n4765 & n27180 ) ;
  assign n27178 = ( n8146 & n17035 ) | ( n8146 & n25959 ) | ( n17035 & n25959 ) ;
  assign n27176 = n17272 ^ n11988 ^ n1226 ;
  assign n27175 = x185 & n12451 ;
  assign n27177 = n27176 ^ n27175 ^ 1'b0 ;
  assign n27182 = n27181 ^ n27178 ^ n27177 ;
  assign n27183 = n21587 ^ n8543 ^ n6333 ;
  assign n27184 = n18200 ^ n4109 ^ n2495 ;
  assign n27185 = n27184 ^ n17194 ^ n3383 ;
  assign n27193 = n9035 ^ n3826 ^ n737 ;
  assign n27187 = ( n402 & ~n4178 ) | ( n402 & n6259 ) | ( ~n4178 & n6259 ) ;
  assign n27186 = n8652 ^ n6694 ^ 1'b0 ;
  assign n27188 = n27187 ^ n27186 ^ 1'b0 ;
  assign n27189 = n17640 | n27188 ;
  assign n27190 = n27189 ^ n3132 ^ 1'b0 ;
  assign n27191 = ~n16849 & n27190 ;
  assign n27192 = ( n20335 & n23171 ) | ( n20335 & ~n27191 ) | ( n23171 & ~n27191 ) ;
  assign n27194 = n27193 ^ n27192 ^ n22158 ;
  assign n27195 = n13898 ^ n10696 ^ n3209 ;
  assign n27196 = n27195 ^ n21841 ^ 1'b0 ;
  assign n27197 = n5283 | n7943 ;
  assign n27198 = n17024 ^ n8244 ^ 1'b0 ;
  assign n27199 = n27197 | n27198 ;
  assign n27208 = ( ~n1282 & n7183 ) | ( ~n1282 & n14564 ) | ( n7183 & n14564 ) ;
  assign n27204 = n18147 ^ n12605 ^ n8512 ;
  assign n27205 = n27204 ^ n8571 ^ 1'b0 ;
  assign n27206 = ~n10624 & n27205 ;
  assign n27200 = n7253 & n10367 ;
  assign n27201 = n27200 ^ n8289 ^ 1'b0 ;
  assign n27202 = ( x132 & ~n893 ) | ( x132 & n4823 ) | ( ~n893 & n4823 ) ;
  assign n27203 = n27201 | n27202 ;
  assign n27207 = n27206 ^ n27203 ^ 1'b0 ;
  assign n27209 = n27208 ^ n27207 ^ n2369 ;
  assign n27210 = n27209 ^ n17320 ^ n3321 ;
  assign n27211 = n11062 ^ n2593 ^ 1'b0 ;
  assign n27212 = ( n10372 & n12295 ) | ( n10372 & n27211 ) | ( n12295 & n27211 ) ;
  assign n27213 = n6411 ^ n2653 ^ 1'b0 ;
  assign n27214 = n27213 ^ n12670 ^ n5337 ;
  assign n27215 = n27214 ^ n21006 ^ n20704 ;
  assign n27216 = ( n6153 & n11295 ) | ( n6153 & ~n13032 ) | ( n11295 & ~n13032 ) ;
  assign n27217 = ( n4992 & n27215 ) | ( n4992 & ~n27216 ) | ( n27215 & ~n27216 ) ;
  assign n27218 = n26906 ^ n13765 ^ n11829 ;
  assign n27219 = ( x204 & ~n16685 ) | ( x204 & n27218 ) | ( ~n16685 & n27218 ) ;
  assign n27220 = ~n15101 & n27219 ;
  assign n27221 = n27220 ^ n14319 ^ 1'b0 ;
  assign n27222 = n20527 ^ n10452 ^ 1'b0 ;
  assign n27223 = ~n9851 & n27222 ;
  assign n27224 = ~n459 & n18725 ;
  assign n27225 = n27224 ^ n10461 ^ 1'b0 ;
  assign n27226 = n27225 ^ n23257 ^ n22098 ;
  assign n27227 = ( n27221 & ~n27223 ) | ( n27221 & n27226 ) | ( ~n27223 & n27226 ) ;
  assign n27228 = n14554 ^ n1508 ^ 1'b0 ;
  assign n27229 = n27228 ^ n25980 ^ n23311 ;
  assign n27231 = ( n3640 & n8702 ) | ( n3640 & n8873 ) | ( n8702 & n8873 ) ;
  assign n27232 = ( n14210 & n25490 ) | ( n14210 & n27231 ) | ( n25490 & n27231 ) ;
  assign n27230 = n15820 & ~n20303 ;
  assign n27233 = n27232 ^ n27230 ^ 1'b0 ;
  assign n27234 = n4039 & ~n27233 ;
  assign n27235 = n27229 & n27234 ;
  assign n27236 = ~n3973 & n6815 ;
  assign n27237 = n20801 & n27236 ;
  assign n27238 = ( ~n5010 & n6042 ) | ( ~n5010 & n6130 ) | ( n6042 & n6130 ) ;
  assign n27239 = ~n10438 & n27238 ;
  assign n27240 = n27239 ^ n14519 ^ 1'b0 ;
  assign n27241 = n27240 ^ n2699 ^ n869 ;
  assign n27242 = x144 & n27241 ;
  assign n27243 = n27237 & n27242 ;
  assign n27244 = n14598 | n27243 ;
  assign n27245 = n17622 | n27244 ;
  assign n27246 = ( n3421 & n10337 ) | ( n3421 & ~n23774 ) | ( n10337 & ~n23774 ) ;
  assign n27247 = n11537 ^ n10394 ^ 1'b0 ;
  assign n27248 = ~n18219 & n27247 ;
  assign n27249 = n27246 | n27248 ;
  assign n27250 = n17992 ^ n13394 ^ 1'b0 ;
  assign n27251 = n27250 ^ n10833 ^ 1'b0 ;
  assign n27252 = ( ~n1555 & n16399 ) | ( ~n1555 & n27251 ) | ( n16399 & n27251 ) ;
  assign n27253 = ( n3747 & ~n4078 ) | ( n3747 & n27252 ) | ( ~n4078 & n27252 ) ;
  assign n27254 = n26708 ^ n17955 ^ n17797 ;
  assign n27264 = ( n6724 & ~n12565 ) | ( n6724 & n13209 ) | ( ~n12565 & n13209 ) ;
  assign n27265 = n27264 ^ n13138 ^ n2576 ;
  assign n27259 = ( ~n16988 & n24449 ) | ( ~n16988 & n27246 ) | ( n24449 & n27246 ) ;
  assign n27260 = n26324 ^ n13849 ^ 1'b0 ;
  assign n27261 = n2318 & n27260 ;
  assign n27262 = ( n3897 & n27259 ) | ( n3897 & n27261 ) | ( n27259 & n27261 ) ;
  assign n27263 = n27262 ^ n21447 ^ n16950 ;
  assign n27255 = ( n1836 & n3414 ) | ( n1836 & n7557 ) | ( n3414 & n7557 ) ;
  assign n27256 = n2299 ^ n622 ^ 1'b0 ;
  assign n27257 = n523 & ~n27256 ;
  assign n27258 = ( n3534 & ~n27255 ) | ( n3534 & n27257 ) | ( ~n27255 & n27257 ) ;
  assign n27266 = n27265 ^ n27263 ^ n27258 ;
  assign n27267 = n6562 | n9327 ;
  assign n27268 = n27267 ^ n25597 ^ 1'b0 ;
  assign n27269 = n9396 & n27268 ;
  assign n27270 = ( ~n2940 & n26922 ) | ( ~n2940 & n27269 ) | ( n26922 & n27269 ) ;
  assign n27271 = n12508 ^ n6817 ^ x52 ;
  assign n27272 = n27271 ^ n13951 ^ 1'b0 ;
  assign n27273 = n10341 & ~n23527 ;
  assign n27274 = ~n27272 & n27273 ;
  assign n27275 = n27274 ^ n9998 ^ 1'b0 ;
  assign n27276 = n6434 & ~n27275 ;
  assign n27277 = n7848 & n25438 ;
  assign n27278 = ~n6018 & n27277 ;
  assign n27279 = n14357 ^ n2076 ^ 1'b0 ;
  assign n27280 = n4741 & n27279 ;
  assign n27281 = n19971 ^ n16411 ^ n4061 ;
  assign n27282 = n14915 ^ n12071 ^ n3372 ;
  assign n27283 = ~n10919 & n19880 ;
  assign n27284 = ( n898 & n27282 ) | ( n898 & n27283 ) | ( n27282 & n27283 ) ;
  assign n27285 = ( x23 & n27281 ) | ( x23 & ~n27284 ) | ( n27281 & ~n27284 ) ;
  assign n27286 = ( n7870 & ~n12180 ) | ( n7870 & n21552 ) | ( ~n12180 & n21552 ) ;
  assign n27287 = ( n27280 & ~n27285 ) | ( n27280 & n27286 ) | ( ~n27285 & n27286 ) ;
  assign n27288 = n8951 & n27287 ;
  assign n27289 = n9717 ^ n612 ^ 1'b0 ;
  assign n27290 = ~n16187 & n27289 ;
  assign n27291 = ( n11836 & n12148 ) | ( n11836 & n24793 ) | ( n12148 & n24793 ) ;
  assign n27292 = n12742 ^ n10993 ^ 1'b0 ;
  assign n27293 = ( n1331 & ~n3808 ) | ( n1331 & n27292 ) | ( ~n3808 & n27292 ) ;
  assign n27294 = ( n667 & n7102 ) | ( n667 & n10001 ) | ( n7102 & n10001 ) ;
  assign n27295 = n26336 & ~n27294 ;
  assign n27296 = n27293 & n27295 ;
  assign n27297 = ( x252 & ~n1481 ) | ( x252 & n8785 ) | ( ~n1481 & n8785 ) ;
  assign n27298 = n27297 ^ n3048 ^ 1'b0 ;
  assign n27299 = ( n1777 & n5507 ) | ( n1777 & ~n27298 ) | ( n5507 & ~n27298 ) ;
  assign n27300 = n27299 ^ n23530 ^ n286 ;
  assign n27301 = ( n12368 & n27296 ) | ( n12368 & ~n27300 ) | ( n27296 & ~n27300 ) ;
  assign n27302 = n17570 ^ n16166 ^ n11988 ;
  assign n27303 = n12835 ^ n9796 ^ n9121 ;
  assign n27304 = ( n15649 & n23317 ) | ( n15649 & n27303 ) | ( n23317 & n27303 ) ;
  assign n27305 = ( n4958 & ~n23598 ) | ( n4958 & n26319 ) | ( ~n23598 & n26319 ) ;
  assign n27306 = n27305 ^ n22539 ^ n2979 ;
  assign n27307 = n27306 ^ n22676 ^ n16561 ;
  assign n27308 = n8817 & n25521 ;
  assign n27309 = n27308 ^ n22185 ^ 1'b0 ;
  assign n27310 = n26319 ^ n20585 ^ n2899 ;
  assign n27311 = n27310 ^ n6647 ^ 1'b0 ;
  assign n27312 = n868 & ~n27311 ;
  assign n27313 = ( ~n4536 & n8727 ) | ( ~n4536 & n16707 ) | ( n8727 & n16707 ) ;
  assign n27314 = n27313 ^ n23596 ^ 1'b0 ;
  assign n27315 = n6044 ^ n2815 ^ 1'b0 ;
  assign n27316 = ( n7518 & n13396 ) | ( n7518 & ~n26021 ) | ( n13396 & ~n26021 ) ;
  assign n27317 = ( n12199 & ~n13639 ) | ( n12199 & n15376 ) | ( ~n13639 & n15376 ) ;
  assign n27318 = n25369 ^ n11920 ^ 1'b0 ;
  assign n27319 = ~n7777 & n27318 ;
  assign n27320 = n27319 ^ n25108 ^ n8686 ;
  assign n27321 = n27320 ^ n23715 ^ n2104 ;
  assign n27322 = ( ~n4039 & n12825 ) | ( ~n4039 & n21191 ) | ( n12825 & n21191 ) ;
  assign n27323 = n2002 & n2630 ;
  assign n27324 = n27323 ^ n6445 ^ 1'b0 ;
  assign n27325 = n20031 & n27324 ;
  assign n27326 = ~n19393 & n27325 ;
  assign n27327 = ( n23132 & n27322 ) | ( n23132 & ~n27326 ) | ( n27322 & ~n27326 ) ;
  assign n27328 = n12068 & ~n27327 ;
  assign n27329 = n27328 ^ n15110 ^ 1'b0 ;
  assign n27330 = ( ~x54 & n5573 ) | ( ~x54 & n10594 ) | ( n5573 & n10594 ) ;
  assign n27331 = n6972 & n18748 ;
  assign n27332 = n27330 & n27331 ;
  assign n27333 = ( n830 & n1575 ) | ( n830 & ~n10795 ) | ( n1575 & ~n10795 ) ;
  assign n27334 = n23102 ^ n10606 ^ n2027 ;
  assign n27335 = n12525 ^ n6256 ^ n6249 ;
  assign n27336 = n27335 ^ n16128 ^ n9698 ;
  assign n27338 = n6162 | n14407 ;
  assign n27337 = n15637 & ~n27022 ;
  assign n27339 = n27338 ^ n27337 ^ 1'b0 ;
  assign n27340 = n18280 ^ n2593 ^ n1873 ;
  assign n27341 = n27340 ^ n25186 ^ n17379 ;
  assign n27342 = n2774 | n27341 ;
  assign n27343 = n27342 ^ n7457 ^ 1'b0 ;
  assign n27344 = n27343 ^ n22458 ^ n4904 ;
  assign n27347 = n18412 ^ n8517 ^ n5975 ;
  assign n27345 = ( ~n5172 & n5962 ) | ( ~n5172 & n8191 ) | ( n5962 & n8191 ) ;
  assign n27346 = ( n17360 & ~n24955 ) | ( n17360 & n27345 ) | ( ~n24955 & n27345 ) ;
  assign n27348 = n27347 ^ n27346 ^ n10787 ;
  assign n27349 = ( ~n3315 & n3701 ) | ( ~n3315 & n13409 ) | ( n3701 & n13409 ) ;
  assign n27350 = ( n17069 & n23207 ) | ( n17069 & ~n27349 ) | ( n23207 & ~n27349 ) ;
  assign n27351 = ( n1138 & n17340 ) | ( n1138 & ~n27350 ) | ( n17340 & ~n27350 ) ;
  assign n27352 = n1826 ^ n1136 ^ n387 ;
  assign n27354 = ( ~x147 & n2185 ) | ( ~x147 & n22410 ) | ( n2185 & n22410 ) ;
  assign n27353 = ~n10438 & n17655 ;
  assign n27355 = n27354 ^ n27353 ^ 1'b0 ;
  assign n27356 = ( n18784 & n27352 ) | ( n18784 & ~n27355 ) | ( n27352 & ~n27355 ) ;
  assign n27357 = ( n4699 & ~n10015 ) | ( n4699 & n15265 ) | ( ~n10015 & n15265 ) ;
  assign n27358 = n27357 ^ n20207 ^ n10856 ;
  assign n27359 = ( n12105 & n13404 ) | ( n12105 & ~n13813 ) | ( n13404 & ~n13813 ) ;
  assign n27360 = n24370 ^ n14023 ^ 1'b0 ;
  assign n27361 = ~n27359 & n27360 ;
  assign n27362 = n23508 ^ n18517 ^ n3545 ;
  assign n27363 = ~n9880 & n25908 ;
  assign n27364 = n1460 & n27363 ;
  assign n27365 = n27364 ^ n16975 ^ 1'b0 ;
  assign n27366 = ( n7054 & ~n25596 ) | ( n7054 & n27365 ) | ( ~n25596 & n27365 ) ;
  assign n27367 = n14334 ^ n13025 ^ n7086 ;
  assign n27368 = n3379 ^ n3003 ^ n688 ;
  assign n27369 = n27368 ^ n13790 ^ 1'b0 ;
  assign n27370 = ~n14509 & n18951 ;
  assign n27371 = n27370 ^ n9197 ^ n7448 ;
  assign n27372 = ~n27369 & n27371 ;
  assign n27373 = n27372 ^ n23573 ^ 1'b0 ;
  assign n27374 = ( n1328 & ~n3488 ) | ( n1328 & n14860 ) | ( ~n3488 & n14860 ) ;
  assign n27375 = ( ~n3869 & n9620 ) | ( ~n3869 & n27374 ) | ( n9620 & n27374 ) ;
  assign n27376 = ( n2496 & ~n14529 ) | ( n2496 & n27375 ) | ( ~n14529 & n27375 ) ;
  assign n27377 = n8007 | n27376 ;
  assign n27378 = n27373 | n27377 ;
  assign n27379 = ( ~n9913 & n27367 ) | ( ~n9913 & n27378 ) | ( n27367 & n27378 ) ;
  assign n27381 = n4463 ^ n772 ^ 1'b0 ;
  assign n27380 = n3470 & n18835 ;
  assign n27382 = n27381 ^ n27380 ^ 1'b0 ;
  assign n27383 = ( n2102 & ~n2381 ) | ( n2102 & n5426 ) | ( ~n2381 & n5426 ) ;
  assign n27385 = n7197 & n11150 ;
  assign n27386 = n27385 ^ x171 ^ 1'b0 ;
  assign n27387 = n27386 ^ n7335 ^ n2332 ;
  assign n27384 = ( n6351 & n12754 ) | ( n6351 & n26186 ) | ( n12754 & n26186 ) ;
  assign n27388 = n27387 ^ n27384 ^ n16331 ;
  assign n27389 = ~n27383 & n27388 ;
  assign n27390 = n27389 ^ n3577 ^ 1'b0 ;
  assign n27392 = n19036 ^ n4758 ^ 1'b0 ;
  assign n27391 = n9539 & ~n17675 ;
  assign n27393 = n27392 ^ n27391 ^ 1'b0 ;
  assign n27394 = n14247 | n15153 ;
  assign n27395 = ( n14569 & ~n27393 ) | ( n14569 & n27394 ) | ( ~n27393 & n27394 ) ;
  assign n27396 = ( n2839 & n10611 ) | ( n2839 & n10956 ) | ( n10611 & n10956 ) ;
  assign n27397 = ( n3618 & n7786 ) | ( n3618 & n26051 ) | ( n7786 & n26051 ) ;
  assign n27398 = ( n22471 & ~n23477 ) | ( n22471 & n27397 ) | ( ~n23477 & n27397 ) ;
  assign n27399 = ( n7444 & n7934 ) | ( n7444 & ~n22774 ) | ( n7934 & ~n22774 ) ;
  assign n27400 = n17461 | n21236 ;
  assign n27401 = n15406 | n27400 ;
  assign n27403 = ~n17976 & n19836 ;
  assign n27404 = n16592 & n27403 ;
  assign n27402 = n6434 & n13900 ;
  assign n27405 = n27404 ^ n27402 ^ 1'b0 ;
  assign n27406 = ( n6862 & n10004 ) | ( n6862 & ~n24539 ) | ( n10004 & ~n24539 ) ;
  assign n27407 = ( n1425 & ~n13552 ) | ( n1425 & n27406 ) | ( ~n13552 & n27406 ) ;
  assign n27408 = n17619 ^ n15218 ^ n7097 ;
  assign n27409 = n1313 & ~n6092 ;
  assign n27410 = n1808 & n27409 ;
  assign n27411 = n27410 ^ n22357 ^ n19017 ;
  assign n27412 = ( ~n5385 & n27408 ) | ( ~n5385 & n27411 ) | ( n27408 & n27411 ) ;
  assign n27421 = n6710 ^ n2731 ^ 1'b0 ;
  assign n27420 = ( n16974 & n17313 ) | ( n16974 & n19448 ) | ( n17313 & n19448 ) ;
  assign n27415 = n784 & n5314 ;
  assign n27416 = n27415 ^ n1499 ^ 1'b0 ;
  assign n27417 = n27416 ^ n25493 ^ n1286 ;
  assign n27413 = ( x124 & n20243 ) | ( x124 & n22010 ) | ( n20243 & n22010 ) ;
  assign n27414 = ( n15401 & ~n15933 ) | ( n15401 & n27413 ) | ( ~n15933 & n27413 ) ;
  assign n27418 = n27417 ^ n27414 ^ 1'b0 ;
  assign n27419 = n25437 | n27418 ;
  assign n27422 = n27421 ^ n27420 ^ n27419 ;
  assign n27423 = ( n2133 & ~n10325 ) | ( n2133 & n14187 ) | ( ~n10325 & n14187 ) ;
  assign n27424 = n9160 & ~n27423 ;
  assign n27425 = n27424 ^ n19131 ^ 1'b0 ;
  assign n27426 = x239 & n8905 ;
  assign n27427 = n27426 ^ n4806 ^ n2618 ;
  assign n27428 = n27427 ^ n15788 ^ n10659 ;
  assign n27429 = n27428 ^ n24929 ^ n4536 ;
  assign n27438 = n3041 ^ n1324 ^ 1'b0 ;
  assign n27439 = n19514 | n27438 ;
  assign n27435 = n2014 | n19353 ;
  assign n27436 = n27435 ^ n1507 ^ 1'b0 ;
  assign n27437 = n1279 & ~n27436 ;
  assign n27440 = n27439 ^ n27437 ^ n5255 ;
  assign n27432 = ( ~n1792 & n11906 ) | ( ~n1792 & n15733 ) | ( n11906 & n15733 ) ;
  assign n27430 = n9189 ^ n2219 ^ n1834 ;
  assign n27431 = n27430 ^ n4661 ^ x145 ;
  assign n27433 = n27432 ^ n27431 ^ n20445 ;
  assign n27434 = n7971 & n27433 ;
  assign n27441 = n27440 ^ n27434 ^ 1'b0 ;
  assign n27442 = ( ~n2036 & n5545 ) | ( ~n2036 & n11242 ) | ( n5545 & n11242 ) ;
  assign n27443 = n13317 ^ n7930 ^ n7451 ;
  assign n27444 = ( n13642 & n22351 ) | ( n13642 & n27443 ) | ( n22351 & n27443 ) ;
  assign n27445 = n27444 ^ n13997 ^ n10064 ;
  assign n27446 = n6936 ^ n1891 ^ 1'b0 ;
  assign n27447 = ~n2413 & n27446 ;
  assign n27448 = ( n2923 & ~n2994 ) | ( n2923 & n4383 ) | ( ~n2994 & n4383 ) ;
  assign n27449 = ( n4200 & ~n27447 ) | ( n4200 & n27448 ) | ( ~n27447 & n27448 ) ;
  assign n27450 = n25193 | n27449 ;
  assign n27451 = n11512 & n13336 ;
  assign n27452 = n27451 ^ n8830 ^ 1'b0 ;
  assign n27453 = ( n1004 & n15445 ) | ( n1004 & ~n21505 ) | ( n15445 & ~n21505 ) ;
  assign n27454 = ( n7191 & ~n10404 ) | ( n7191 & n17205 ) | ( ~n10404 & n17205 ) ;
  assign n27455 = ~n2100 & n14380 ;
  assign n27456 = n27455 ^ n9054 ^ 1'b0 ;
  assign n27457 = n20349 ^ n12691 ^ n3377 ;
  assign n27458 = ( ~n6906 & n14239 ) | ( ~n6906 & n27457 ) | ( n14239 & n27457 ) ;
  assign n27459 = n27458 ^ n18622 ^ n4034 ;
  assign n27462 = n8543 ^ n7030 ^ x134 ;
  assign n27460 = ( n3451 & ~n11840 ) | ( n3451 & n12419 ) | ( ~n11840 & n12419 ) ;
  assign n27461 = n27460 ^ n6299 ^ n3421 ;
  assign n27463 = n27462 ^ n27461 ^ n24198 ;
  assign n27464 = ( ~n1781 & n27459 ) | ( ~n1781 & n27463 ) | ( n27459 & n27463 ) ;
  assign n27465 = ( n26389 & n27456 ) | ( n26389 & ~n27464 ) | ( n27456 & ~n27464 ) ;
  assign n27466 = ( n10064 & n14172 ) | ( n10064 & n17372 ) | ( n14172 & n17372 ) ;
  assign n27467 = ( n5081 & n7669 ) | ( n5081 & ~n7683 ) | ( n7669 & ~n7683 ) ;
  assign n27471 = n2586 | n5186 ;
  assign n27472 = n27471 ^ n14694 ^ 1'b0 ;
  assign n27469 = n9627 ^ n7376 ^ n3493 ;
  assign n27468 = n5160 & ~n7306 ;
  assign n27470 = n27469 ^ n27468 ^ n3746 ;
  assign n27473 = n27472 ^ n27470 ^ n18051 ;
  assign n27476 = ( ~n7398 & n12473 ) | ( ~n7398 & n14069 ) | ( n12473 & n14069 ) ;
  assign n27474 = ( ~n3451 & n15936 ) | ( ~n3451 & n21492 ) | ( n15936 & n21492 ) ;
  assign n27475 = x7 & n27474 ;
  assign n27477 = n27476 ^ n27475 ^ 1'b0 ;
  assign n27478 = ( n15076 & ~n27473 ) | ( n15076 & n27477 ) | ( ~n27473 & n27477 ) ;
  assign n27479 = ( n12911 & n27467 ) | ( n12911 & ~n27478 ) | ( n27467 & ~n27478 ) ;
  assign n27480 = n27479 ^ n16059 ^ 1'b0 ;
  assign n27481 = n22317 & ~n25472 ;
  assign n27482 = n27481 ^ n12526 ^ 1'b0 ;
  assign n27483 = n27482 ^ n13096 ^ n9033 ;
  assign n27484 = n785 & ~n9147 ;
  assign n27485 = n27484 ^ n7269 ^ 1'b0 ;
  assign n27486 = n16251 & ~n27485 ;
  assign n27487 = n23264 & ~n23997 ;
  assign n27488 = n27487 ^ n10816 ^ 1'b0 ;
  assign n27489 = n5330 & ~n10996 ;
  assign n27490 = n25086 ^ n1218 ^ 1'b0 ;
  assign n27493 = n7920 & ~n9819 ;
  assign n27494 = ~n24742 & n27493 ;
  assign n27491 = n13809 ^ n8120 ^ n472 ;
  assign n27492 = ( ~n22496 & n25755 ) | ( ~n22496 & n27491 ) | ( n25755 & n27491 ) ;
  assign n27495 = n27494 ^ n27492 ^ n13574 ;
  assign n27496 = ( ~n940 & n27490 ) | ( ~n940 & n27495 ) | ( n27490 & n27495 ) ;
  assign n27497 = n4581 ^ n3223 ^ n528 ;
  assign n27498 = n27497 ^ n13531 ^ 1'b0 ;
  assign n27499 = n5379 & n19930 ;
  assign n27500 = n12037 ^ n5793 ^ 1'b0 ;
  assign n27501 = n27500 ^ n18110 ^ n1645 ;
  assign n27502 = n17895 ^ n10963 ^ n575 ;
  assign n27503 = n27502 ^ n25134 ^ n21256 ;
  assign n27504 = ( n1553 & n15449 ) | ( n1553 & n27503 ) | ( n15449 & n27503 ) ;
  assign n27505 = n27504 ^ n21424 ^ n16764 ;
  assign n27509 = n17185 ^ n15548 ^ n8464 ;
  assign n27506 = x143 & n25388 ;
  assign n27507 = n27506 ^ n13297 ^ n9572 ;
  assign n27508 = ~n16442 & n27507 ;
  assign n27510 = n27509 ^ n27508 ^ 1'b0 ;
  assign n27511 = ( n8973 & n10166 ) | ( n8973 & n27510 ) | ( n10166 & n27510 ) ;
  assign n27512 = ( ~x147 & n6803 ) | ( ~x147 & n16308 ) | ( n6803 & n16308 ) ;
  assign n27513 = n25464 ^ n8279 ^ 1'b0 ;
  assign n27514 = n27513 ^ n5303 ^ 1'b0 ;
  assign n27515 = n27512 & n27514 ;
  assign n27516 = ( ~n2102 & n9133 ) | ( ~n2102 & n26607 ) | ( n9133 & n26607 ) ;
  assign n27517 = n26247 & n27516 ;
  assign n27518 = n17589 ^ n7497 ^ n4575 ;
  assign n27519 = n6094 ^ n5658 ^ n1752 ;
  assign n27520 = n27519 ^ n26860 ^ 1'b0 ;
  assign n27521 = n27518 | n27520 ;
  assign n27523 = ( ~n19876 & n22574 ) | ( ~n19876 & n25578 ) | ( n22574 & n25578 ) ;
  assign n27522 = ( x249 & ~n6703 ) | ( x249 & n13201 ) | ( ~n6703 & n13201 ) ;
  assign n27524 = n27523 ^ n27522 ^ n3337 ;
  assign n27525 = ( n2973 & n27521 ) | ( n2973 & ~n27524 ) | ( n27521 & ~n27524 ) ;
  assign n27526 = n3599 | n8477 ;
  assign n27527 = n27526 ^ n25412 ^ n22021 ;
  assign n27528 = ( n1852 & ~n6238 ) | ( n1852 & n18256 ) | ( ~n6238 & n18256 ) ;
  assign n27529 = ( n16671 & ~n18955 ) | ( n16671 & n27528 ) | ( ~n18955 & n27528 ) ;
  assign n27530 = n5121 | n8735 ;
  assign n27531 = n7538 & ~n27530 ;
  assign n27532 = n15078 & ~n27531 ;
  assign n27533 = n25608 ^ n4301 ^ n4176 ;
  assign n27534 = n5357 & ~n10512 ;
  assign n27535 = n27533 & n27534 ;
  assign n27536 = ( n6737 & n11677 ) | ( n6737 & n27535 ) | ( n11677 & n27535 ) ;
  assign n27537 = ( ~n2058 & n8743 ) | ( ~n2058 & n27536 ) | ( n8743 & n27536 ) ;
  assign n27539 = ( n413 & n523 ) | ( n413 & ~n1220 ) | ( n523 & ~n1220 ) ;
  assign n27538 = n16660 & n20158 ;
  assign n27540 = n27539 ^ n27538 ^ n24921 ;
  assign n27541 = ( n12295 & n14392 ) | ( n12295 & n27540 ) | ( n14392 & n27540 ) ;
  assign n27542 = n23882 ^ n12129 ^ n6780 ;
  assign n27543 = ~n388 & n27542 ;
  assign n27544 = n13428 & ~n24459 ;
  assign n27545 = n27544 ^ n24855 ^ 1'b0 ;
  assign n27546 = ( n9501 & ~n27543 ) | ( n9501 & n27545 ) | ( ~n27543 & n27545 ) ;
  assign n27547 = n7496 & n17562 ;
  assign n27548 = n5006 & n27547 ;
  assign n27549 = n27548 ^ n6579 ^ n2103 ;
  assign n27550 = ( ~n4777 & n17428 ) | ( ~n4777 & n27549 ) | ( n17428 & n27549 ) ;
  assign n27551 = n13452 & ~n18376 ;
  assign n27552 = n14083 & ~n27551 ;
  assign n27553 = n11991 ^ n5203 ^ n3628 ;
  assign n27554 = n4787 & ~n17077 ;
  assign n27555 = n27554 ^ n8316 ^ n5173 ;
  assign n27556 = ( ~n10855 & n15358 ) | ( ~n10855 & n27555 ) | ( n15358 & n27555 ) ;
  assign n27557 = n27553 & ~n27556 ;
  assign n27558 = n27552 & n27557 ;
  assign n27559 = ( n5358 & ~n9444 ) | ( n5358 & n15396 ) | ( ~n9444 & n15396 ) ;
  assign n27560 = ( n9606 & n11462 ) | ( n9606 & ~n16800 ) | ( n11462 & ~n16800 ) ;
  assign n27561 = ( n820 & ~n18033 ) | ( n820 & n27560 ) | ( ~n18033 & n27560 ) ;
  assign n27563 = n7729 | n10328 ;
  assign n27562 = n3095 & ~n16338 ;
  assign n27564 = n27563 ^ n27562 ^ n13812 ;
  assign n27565 = n27564 ^ n20446 ^ n13050 ;
  assign n27566 = n6143 & n23984 ;
  assign n27567 = n15618 & n27566 ;
  assign n27574 = ( n678 & n3258 ) | ( n678 & n4187 ) | ( n3258 & n4187 ) ;
  assign n27575 = n27574 ^ n17662 ^ n10515 ;
  assign n27568 = ~n10098 & n17424 ;
  assign n27569 = n2900 & n27568 ;
  assign n27570 = n9919 | n27569 ;
  assign n27571 = n5777 | n27570 ;
  assign n27572 = ( n1530 & ~n10657 ) | ( n1530 & n27571 ) | ( ~n10657 & n27571 ) ;
  assign n27573 = n27572 ^ n12233 ^ n8582 ;
  assign n27576 = n27575 ^ n27573 ^ n17777 ;
  assign n27577 = ~n16768 & n18261 ;
  assign n27580 = ( ~n2759 & n16701 ) | ( ~n2759 & n25416 ) | ( n16701 & n25416 ) ;
  assign n27581 = n2368 ^ n1863 ^ 1'b0 ;
  assign n27582 = ~n27580 & n27581 ;
  assign n27583 = ( ~n6461 & n9151 ) | ( ~n6461 & n27582 ) | ( n9151 & n27582 ) ;
  assign n27578 = n2141 ^ n416 ^ 1'b0 ;
  assign n27579 = n15027 | n27578 ;
  assign n27584 = n27583 ^ n27579 ^ 1'b0 ;
  assign n27590 = ( n822 & n5579 ) | ( n822 & ~n14789 ) | ( n5579 & ~n14789 ) ;
  assign n27585 = n11734 ^ n10136 ^ n6393 ;
  assign n27586 = n21733 ^ n6816 ^ n4761 ;
  assign n27587 = n27586 ^ n13351 ^ 1'b0 ;
  assign n27588 = n27585 & n27587 ;
  assign n27589 = ( n11548 & n22367 ) | ( n11548 & n27588 ) | ( n22367 & n27588 ) ;
  assign n27591 = n27590 ^ n27589 ^ 1'b0 ;
  assign n27592 = n10011 ^ n8813 ^ 1'b0 ;
  assign n27593 = n27591 | n27592 ;
  assign n27594 = n3133 ^ n941 ^ 1'b0 ;
  assign n27595 = ( n3673 & n23588 ) | ( n3673 & n24777 ) | ( n23588 & n24777 ) ;
  assign n27596 = ( n6736 & ~n19539 ) | ( n6736 & n26265 ) | ( ~n19539 & n26265 ) ;
  assign n27597 = ( n26064 & n27595 ) | ( n26064 & ~n27596 ) | ( n27595 & ~n27596 ) ;
  assign n27598 = ( n2426 & n10979 ) | ( n2426 & n27597 ) | ( n10979 & n27597 ) ;
  assign n27601 = ~n15811 & n23390 ;
  assign n27602 = n16940 & n27601 ;
  assign n27599 = n9209 | n16809 ;
  assign n27600 = n27599 ^ n10335 ^ 1'b0 ;
  assign n27603 = n27602 ^ n27600 ^ 1'b0 ;
  assign n27604 = n2006 | n27603 ;
  assign n27605 = n27604 ^ n27153 ^ 1'b0 ;
  assign n27606 = ( n2054 & n10214 ) | ( n2054 & ~n22218 ) | ( n10214 & ~n22218 ) ;
  assign n27607 = n27606 ^ n15897 ^ 1'b0 ;
  assign n27608 = n4777 | n27607 ;
  assign n27609 = ~n1644 & n18110 ;
  assign n27610 = ~n27608 & n27609 ;
  assign n27611 = ( n9422 & n13039 ) | ( n9422 & ~n15141 ) | ( n13039 & ~n15141 ) ;
  assign n27612 = ( n4485 & n21416 ) | ( n4485 & n27611 ) | ( n21416 & n27611 ) ;
  assign n27613 = ( n3592 & n4040 ) | ( n3592 & ~n21204 ) | ( n4040 & ~n21204 ) ;
  assign n27614 = n11516 | n27613 ;
  assign n27615 = ( n5713 & n27612 ) | ( n5713 & ~n27614 ) | ( n27612 & ~n27614 ) ;
  assign n27616 = n313 & n14839 ;
  assign n27617 = n27616 ^ n21755 ^ 1'b0 ;
  assign n27618 = n14510 ^ n6816 ^ n1560 ;
  assign n27619 = n27618 ^ n11497 ^ 1'b0 ;
  assign n27620 = n21191 ^ n3959 ^ 1'b0 ;
  assign n27621 = ( n4841 & n4968 ) | ( n4841 & ~n11201 ) | ( n4968 & ~n11201 ) ;
  assign n27622 = n27621 ^ n7648 ^ n6080 ;
  assign n27623 = n15899 ^ n14836 ^ 1'b0 ;
  assign n27624 = ~n27622 & n27623 ;
  assign n27625 = n27624 ^ n1700 ^ 1'b0 ;
  assign n27626 = n27620 & ~n27625 ;
  assign n27627 = ( n27617 & n27619 ) | ( n27617 & n27626 ) | ( n27619 & n27626 ) ;
  assign n27628 = ( ~n3983 & n11467 ) | ( ~n3983 & n24313 ) | ( n11467 & n24313 ) ;
  assign n27629 = ( ~n6517 & n27627 ) | ( ~n6517 & n27628 ) | ( n27627 & n27628 ) ;
  assign n27630 = n16081 ^ n9834 ^ n2903 ;
  assign n27631 = n3668 & n14069 ;
  assign n27632 = n27631 ^ n18915 ^ 1'b0 ;
  assign n27633 = ( n2998 & n10183 ) | ( n2998 & n11091 ) | ( n10183 & n11091 ) ;
  assign n27634 = n27633 ^ n8126 ^ n7659 ;
  assign n27635 = n7951 | n27634 ;
  assign n27636 = n27632 & ~n27635 ;
  assign n27637 = ( ~n4668 & n19338 ) | ( ~n4668 & n27636 ) | ( n19338 & n27636 ) ;
  assign n27640 = x48 & ~n9438 ;
  assign n27641 = n27640 ^ n16831 ^ 1'b0 ;
  assign n27638 = n8008 ^ n2801 ^ n270 ;
  assign n27639 = n17488 | n27638 ;
  assign n27642 = n27641 ^ n27639 ^ 1'b0 ;
  assign n27643 = n22226 ^ n5127 ^ n1215 ;
  assign n27644 = ( ~n1161 & n2738 ) | ( ~n1161 & n27643 ) | ( n2738 & n27643 ) ;
  assign n27645 = n7847 ^ n1500 ^ 1'b0 ;
  assign n27646 = n4196 & ~n6151 ;
  assign n27650 = n5983 & n8253 ;
  assign n27649 = n7737 & n12792 ;
  assign n27651 = n27650 ^ n27649 ^ n4219 ;
  assign n27647 = x32 & ~n16953 ;
  assign n27648 = n7976 & n27647 ;
  assign n27652 = n27651 ^ n27648 ^ 1'b0 ;
  assign n27653 = n4741 | n9653 ;
  assign n27656 = ( n548 & n3614 ) | ( n548 & ~n9587 ) | ( n3614 & ~n9587 ) ;
  assign n27654 = n10191 | n12124 ;
  assign n27655 = n19305 | n27654 ;
  assign n27657 = n27656 ^ n27655 ^ n10510 ;
  assign n27658 = n27657 ^ n6856 ^ n5486 ;
  assign n27659 = n13302 ^ n734 ^ 1'b0 ;
  assign n27660 = n9182 & ~n27659 ;
  assign n27661 = n23860 ^ n20881 ^ 1'b0 ;
  assign n27662 = n6559 ^ n1944 ^ x77 ;
  assign n27663 = n27662 ^ n6398 ^ n1349 ;
  assign n27664 = n11995 & n14767 ;
  assign n27665 = n27663 & n27664 ;
  assign n27666 = n14785 & n18772 ;
  assign n27667 = n27665 & n27666 ;
  assign n27668 = n16271 ^ n737 ^ 1'b0 ;
  assign n27669 = n5103 ^ n1356 ^ x64 ;
  assign n27670 = ( n14579 & ~n19017 ) | ( n14579 & n27669 ) | ( ~n19017 & n27669 ) ;
  assign n27671 = ( n9904 & n17393 ) | ( n9904 & ~n27670 ) | ( n17393 & ~n27670 ) ;
  assign n27672 = ( n4371 & n21835 ) | ( n4371 & ~n24066 ) | ( n21835 & ~n24066 ) ;
  assign n27673 = n17402 & n17901 ;
  assign n27674 = n20410 ^ n18736 ^ n18350 ;
  assign n27675 = n25943 | n27674 ;
  assign n27676 = n27675 ^ n11267 ^ 1'b0 ;
  assign n27684 = n14510 ^ n8595 ^ n2968 ;
  assign n27685 = ( n14958 & ~n25040 ) | ( n14958 & n27684 ) | ( ~n25040 & n27684 ) ;
  assign n27681 = n17728 ^ n12266 ^ n368 ;
  assign n27677 = n790 | n8688 ;
  assign n27678 = n27677 ^ n11588 ^ 1'b0 ;
  assign n27679 = n27678 ^ n13070 ^ n3213 ;
  assign n27680 = ( n706 & n4729 ) | ( n706 & n27679 ) | ( n4729 & n27679 ) ;
  assign n27682 = n27681 ^ n27680 ^ n4191 ;
  assign n27683 = n12791 & ~n27682 ;
  assign n27686 = n27685 ^ n27683 ^ 1'b0 ;
  assign n27689 = n21416 ^ n10437 ^ n354 ;
  assign n27687 = n20984 ^ n12896 ^ n10989 ;
  assign n27688 = n27687 ^ n8397 ^ n1616 ;
  assign n27690 = n27689 ^ n27688 ^ x201 ;
  assign n27691 = ( n911 & ~n15796 ) | ( n911 & n27690 ) | ( ~n15796 & n27690 ) ;
  assign n27692 = n10222 & n19464 ;
  assign n27693 = n27692 ^ n8341 ^ 1'b0 ;
  assign n27694 = n27693 ^ n25115 ^ n19869 ;
  assign n27695 = n5519 ^ n2860 ^ n2763 ;
  assign n27696 = n4757 | n27695 ;
  assign n27697 = ( x17 & n8686 ) | ( x17 & ~n12423 ) | ( n8686 & ~n12423 ) ;
  assign n27698 = ( ~n1879 & n9615 ) | ( ~n1879 & n15514 ) | ( n9615 & n15514 ) ;
  assign n27699 = ( n27696 & ~n27697 ) | ( n27696 & n27698 ) | ( ~n27697 & n27698 ) ;
  assign n27700 = ~n16390 & n23896 ;
  assign n27701 = ~n8950 & n27700 ;
  assign n27702 = ( n2012 & ~n4837 ) | ( n2012 & n10514 ) | ( ~n4837 & n10514 ) ;
  assign n27703 = ( ~n730 & n6452 ) | ( ~n730 & n27702 ) | ( n6452 & n27702 ) ;
  assign n27704 = n27703 ^ n9075 ^ 1'b0 ;
  assign n27705 = n9621 & n10551 ;
  assign n27706 = n26167 & n27705 ;
  assign n27707 = n27706 ^ n18403 ^ 1'b0 ;
  assign n27708 = ~n7957 & n27707 ;
  assign n27709 = ~n10022 & n27708 ;
  assign n27710 = n26204 ^ n23477 ^ n3570 ;
  assign n27711 = n564 | n2623 ;
  assign n27712 = n25718 | n27711 ;
  assign n27713 = n27710 | n27712 ;
  assign n27714 = ( n1344 & n11001 ) | ( n1344 & ~n21567 ) | ( n11001 & ~n21567 ) ;
  assign n27715 = ( n11017 & ~n27713 ) | ( n11017 & n27714 ) | ( ~n27713 & n27714 ) ;
  assign n27716 = n11201 ^ n11074 ^ 1'b0 ;
  assign n27717 = n12412 | n27716 ;
  assign n27718 = n27717 ^ n8123 ^ n3120 ;
  assign n27719 = ( n4556 & ~n4830 ) | ( n4556 & n8708 ) | ( ~n4830 & n8708 ) ;
  assign n27720 = n27719 ^ n16867 ^ n16079 ;
  assign n27721 = n27720 ^ n24877 ^ n8689 ;
  assign n27722 = ( n3939 & n12647 ) | ( n3939 & n14795 ) | ( n12647 & n14795 ) ;
  assign n27725 = n22097 ^ n20337 ^ n18973 ;
  assign n27726 = ( n6546 & n25630 ) | ( n6546 & ~n27725 ) | ( n25630 & ~n27725 ) ;
  assign n27727 = n27726 ^ n6128 ^ n6001 ;
  assign n27728 = n27727 ^ n27638 ^ n5209 ;
  assign n27723 = ( ~n7563 & n13989 ) | ( ~n7563 & n24472 ) | ( n13989 & n24472 ) ;
  assign n27724 = ~n944 & n27723 ;
  assign n27729 = n27728 ^ n27724 ^ 1'b0 ;
  assign n27730 = ( n27595 & n27722 ) | ( n27595 & ~n27729 ) | ( n27722 & ~n27729 ) ;
  assign n27731 = n17218 ^ n8043 ^ n874 ;
  assign n27732 = n27731 ^ n5915 ^ 1'b0 ;
  assign n27733 = n1938 & n9214 ;
  assign n27734 = ( n7253 & n25784 ) | ( n7253 & ~n27733 ) | ( n25784 & ~n27733 ) ;
  assign n27735 = n23236 ^ n4101 ^ 1'b0 ;
  assign n27736 = n6477 | n10838 ;
  assign n27737 = n27736 ^ n18987 ^ n4612 ;
  assign n27738 = ( n2883 & n15575 ) | ( n2883 & ~n17784 ) | ( n15575 & ~n17784 ) ;
  assign n27739 = ~n21957 & n27738 ;
  assign n27740 = n27739 ^ n10416 ^ n8150 ;
  assign n27741 = n27740 ^ n14182 ^ n3768 ;
  assign n27742 = ~n2464 & n6189 ;
  assign n27743 = n27742 ^ n3872 ^ 1'b0 ;
  assign n27744 = ( n4487 & n9598 ) | ( n4487 & ~n27743 ) | ( n9598 & ~n27743 ) ;
  assign n27745 = n8084 | n9453 ;
  assign n27746 = n27745 ^ n9898 ^ 1'b0 ;
  assign n27747 = ( n19557 & ~n27744 ) | ( n19557 & n27746 ) | ( ~n27744 & n27746 ) ;
  assign n27758 = ( x250 & ~n4651 ) | ( x250 & n21191 ) | ( ~n4651 & n21191 ) ;
  assign n27752 = n12963 ^ n11429 ^ n1047 ;
  assign n27750 = n4761 ^ n1313 ^ 1'b0 ;
  assign n27751 = n27750 ^ n24881 ^ x139 ;
  assign n27748 = ( n10140 & n19593 ) | ( n10140 & ~n26198 ) | ( n19593 & ~n26198 ) ;
  assign n27749 = ( n19233 & n24941 ) | ( n19233 & n27748 ) | ( n24941 & n27748 ) ;
  assign n27753 = n27752 ^ n27751 ^ n27749 ;
  assign n27754 = n25942 ^ n12125 ^ n2509 ;
  assign n27755 = n27754 ^ n16616 ^ n11345 ;
  assign n27756 = n27755 ^ n18650 ^ 1'b0 ;
  assign n27757 = n27753 & ~n27756 ;
  assign n27759 = n27758 ^ n27757 ^ n8964 ;
  assign n27760 = n27759 ^ n20239 ^ n2577 ;
  assign n27761 = ( ~n4512 & n11534 ) | ( ~n4512 & n11576 ) | ( n11534 & n11576 ) ;
  assign n27762 = ( n1137 & n7141 ) | ( n1137 & n11905 ) | ( n7141 & n11905 ) ;
  assign n27763 = n27762 ^ n25766 ^ n7883 ;
  assign n27764 = n27763 ^ n7551 ^ n839 ;
  assign n27768 = ( ~n5727 & n7906 ) | ( ~n5727 & n11165 ) | ( n7906 & n11165 ) ;
  assign n27765 = n7639 ^ n5621 ^ n3396 ;
  assign n27766 = ( n9600 & n16244 ) | ( n9600 & n27765 ) | ( n16244 & n27765 ) ;
  assign n27767 = ( n6991 & n7896 ) | ( n6991 & ~n27766 ) | ( n7896 & ~n27766 ) ;
  assign n27769 = n27768 ^ n27767 ^ 1'b0 ;
  assign n27770 = ~n17987 & n27769 ;
  assign n27773 = n7646 | n17134 ;
  assign n27774 = n27773 ^ n11767 ^ 1'b0 ;
  assign n27771 = n14473 ^ n12456 ^ 1'b0 ;
  assign n27772 = n27771 ^ n25320 ^ n7504 ;
  assign n27775 = n27774 ^ n27772 ^ 1'b0 ;
  assign n27776 = ~n13984 & n17471 ;
  assign n27777 = ( n447 & n10777 ) | ( n447 & n10785 ) | ( n10777 & n10785 ) ;
  assign n27778 = n27777 ^ n7128 ^ n5426 ;
  assign n27779 = n27778 ^ n17113 ^ 1'b0 ;
  assign n27780 = n23924 ^ n18397 ^ n3848 ;
  assign n27781 = ~n1693 & n7612 ;
  assign n27782 = n27781 ^ n7624 ^ n4109 ;
  assign n27783 = n5541 & n27782 ;
  assign n27784 = n27783 ^ n23156 ^ 1'b0 ;
  assign n27785 = n27345 ^ n13334 ^ n3117 ;
  assign n27786 = n6625 & n27785 ;
  assign n27794 = n321 & n4547 ;
  assign n27795 = n27794 ^ n2114 ^ n1044 ;
  assign n27793 = ( n6477 & n10672 ) | ( n6477 & n21030 ) | ( n10672 & n21030 ) ;
  assign n27789 = ( n4965 & ~n7979 ) | ( n4965 & n12648 ) | ( ~n7979 & n12648 ) ;
  assign n27788 = ( n3077 & ~n5125 ) | ( n3077 & n14286 ) | ( ~n5125 & n14286 ) ;
  assign n27790 = n27789 ^ n27788 ^ n1027 ;
  assign n27791 = n27790 ^ n12398 ^ n6270 ;
  assign n27787 = ~n2574 & n17764 ;
  assign n27792 = n27791 ^ n27787 ^ 1'b0 ;
  assign n27796 = n27795 ^ n27793 ^ n27792 ;
  assign n27797 = ( n8620 & n14637 ) | ( n8620 & n25965 ) | ( n14637 & n25965 ) ;
  assign n27798 = n27797 ^ n6789 ^ 1'b0 ;
  assign n27799 = ~n27796 & n27798 ;
  assign n27800 = ( n5560 & n10943 ) | ( n5560 & n14759 ) | ( n10943 & n14759 ) ;
  assign n27801 = n800 & n27800 ;
  assign n27802 = n27801 ^ n3715 ^ 1'b0 ;
  assign n27803 = ( n623 & n25750 ) | ( n623 & ~n27802 ) | ( n25750 & ~n27802 ) ;
  assign n27804 = ( n3144 & ~n9657 ) | ( n3144 & n15811 ) | ( ~n9657 & n15811 ) ;
  assign n27805 = n27804 ^ n19024 ^ n3638 ;
  assign n27806 = n27805 ^ n21829 ^ n16238 ;
  assign n27807 = ( ~n7710 & n8784 ) | ( ~n7710 & n22187 ) | ( n8784 & n22187 ) ;
  assign n27808 = n27807 ^ n19118 ^ n1729 ;
  assign n27809 = n5419 ^ n828 ^ 1'b0 ;
  assign n27810 = n12543 & ~n27809 ;
  assign n27811 = ( ~x140 & n27808 ) | ( ~x140 & n27810 ) | ( n27808 & n27810 ) ;
  assign n27812 = n24657 ^ n20931 ^ n17257 ;
  assign n27813 = n12316 ^ n2299 ^ 1'b0 ;
  assign n27819 = ( n1261 & ~n14865 ) | ( n1261 & n22941 ) | ( ~n14865 & n22941 ) ;
  assign n27820 = n7240 | n27819 ;
  assign n27821 = n27820 ^ n16807 ^ 1'b0 ;
  assign n27822 = ~n1045 & n27821 ;
  assign n27814 = n2974 & ~n12690 ;
  assign n27815 = ( n665 & n3803 ) | ( n665 & ~n4241 ) | ( n3803 & ~n4241 ) ;
  assign n27816 = n27815 ^ n19315 ^ 1'b0 ;
  assign n27817 = ( n6171 & n27814 ) | ( n6171 & ~n27816 ) | ( n27814 & ~n27816 ) ;
  assign n27818 = n16269 | n27817 ;
  assign n27823 = n27822 ^ n27818 ^ 1'b0 ;
  assign n27824 = ( n15987 & n22432 ) | ( n15987 & n27823 ) | ( n22432 & n27823 ) ;
  assign n27825 = n27824 ^ n2102 ^ 1'b0 ;
  assign n27826 = n4258 ^ n3405 ^ n3124 ;
  assign n27827 = n27826 ^ n21044 ^ n7312 ;
  assign n27828 = ( n9556 & ~n15496 ) | ( n9556 & n27827 ) | ( ~n15496 & n27827 ) ;
  assign n27829 = ( n21448 & ~n22781 ) | ( n21448 & n27828 ) | ( ~n22781 & n27828 ) ;
  assign n27830 = n16069 ^ n1863 ^ 1'b0 ;
  assign n27831 = n26539 | n27830 ;
  assign n27832 = n8949 ^ x75 ^ 1'b0 ;
  assign n27833 = ~n11043 & n27832 ;
  assign n27834 = ( ~n15845 & n16000 ) | ( ~n15845 & n27833 ) | ( n16000 & n27833 ) ;
  assign n27835 = ( x217 & ~n10946 ) | ( x217 & n12909 ) | ( ~n10946 & n12909 ) ;
  assign n27836 = n27834 & n27835 ;
  assign n27837 = ~n2677 & n27836 ;
  assign n27838 = n12134 | n27837 ;
  assign n27839 = n27838 ^ n9527 ^ 1'b0 ;
  assign n27840 = ( n11961 & ~n14006 ) | ( n11961 & n27839 ) | ( ~n14006 & n27839 ) ;
  assign n27841 = n3849 ^ n2049 ^ n1813 ;
  assign n27842 = ~n782 & n18228 ;
  assign n27843 = ~n11481 & n27842 ;
  assign n27844 = ( n2178 & n6164 ) | ( n2178 & ~n27843 ) | ( n6164 & ~n27843 ) ;
  assign n27845 = n27844 ^ n14999 ^ n484 ;
  assign n27846 = ( n10908 & n27841 ) | ( n10908 & ~n27845 ) | ( n27841 & ~n27845 ) ;
  assign n27847 = x117 & ~n23543 ;
  assign n27848 = x85 & n7181 ;
  assign n27849 = ( n4375 & n8865 ) | ( n4375 & ~n14572 ) | ( n8865 & ~n14572 ) ;
  assign n27850 = n27849 ^ n12451 ^ n8207 ;
  assign n27851 = n9882 ^ n7370 ^ n4968 ;
  assign n27852 = ( n897 & n17901 ) | ( n897 & ~n27851 ) | ( n17901 & ~n27851 ) ;
  assign n27853 = ( n2873 & n4650 ) | ( n2873 & ~n24667 ) | ( n4650 & ~n24667 ) ;
  assign n27854 = ( ~n709 & n8461 ) | ( ~n709 & n26198 ) | ( n8461 & n26198 ) ;
  assign n27855 = n1482 & ~n9660 ;
  assign n27856 = ~n3363 & n27855 ;
  assign n27857 = n4221 & ~n9717 ;
  assign n27858 = n4647 ^ n3750 ^ n1930 ;
  assign n27859 = ( n8698 & n16548 ) | ( n8698 & ~n27858 ) | ( n16548 & ~n27858 ) ;
  assign n27860 = ( n3565 & ~n27857 ) | ( n3565 & n27859 ) | ( ~n27857 & n27859 ) ;
  assign n27861 = ( n16593 & n23474 ) | ( n16593 & ~n27860 ) | ( n23474 & ~n27860 ) ;
  assign n27862 = ( n4081 & ~n27856 ) | ( n4081 & n27861 ) | ( ~n27856 & n27861 ) ;
  assign n27863 = n18061 | n27862 ;
  assign n27864 = n27863 ^ n9368 ^ 1'b0 ;
  assign n27865 = ( n7634 & ~n10381 ) | ( n7634 & n27864 ) | ( ~n10381 & n27864 ) ;
  assign n27866 = ( n6520 & n27854 ) | ( n6520 & ~n27865 ) | ( n27854 & ~n27865 ) ;
  assign n27867 = n12398 ^ n4128 ^ n848 ;
  assign n27868 = ( ~n7754 & n12429 ) | ( ~n7754 & n27867 ) | ( n12429 & n27867 ) ;
  assign n27869 = n6899 & n27193 ;
  assign n27870 = n27869 ^ n2307 ^ 1'b0 ;
  assign n27871 = ( n23032 & n24142 ) | ( n23032 & n27870 ) | ( n24142 & n27870 ) ;
  assign n27872 = n27871 ^ n6309 ^ 1'b0 ;
  assign n27873 = ( n10618 & ~n14084 ) | ( n10618 & n22450 ) | ( ~n14084 & n22450 ) ;
  assign n27874 = n15669 ^ n12543 ^ n12318 ;
  assign n27875 = n12743 ^ n3978 ^ n1013 ;
  assign n27876 = n27875 ^ n24179 ^ n7830 ;
  assign n27877 = ( n2524 & n22510 ) | ( n2524 & n27876 ) | ( n22510 & n27876 ) ;
  assign n27878 = ( n1794 & ~n6082 ) | ( n1794 & n11623 ) | ( ~n6082 & n11623 ) ;
  assign n27879 = n27878 ^ n18271 ^ n14886 ;
  assign n27880 = ( n829 & n2234 ) | ( n829 & n27879 ) | ( n2234 & n27879 ) ;
  assign n27881 = n6508 ^ n3642 ^ n280 ;
  assign n27882 = n27881 ^ n4063 ^ 1'b0 ;
  assign n27883 = n8028 & ~n27882 ;
  assign n27884 = n27883 ^ n13235 ^ n3799 ;
  assign n27885 = ( n2763 & n14430 ) | ( n2763 & ~n19496 ) | ( n14430 & ~n19496 ) ;
  assign n27886 = ( n722 & n10755 ) | ( n722 & ~n20250 ) | ( n10755 & ~n20250 ) ;
  assign n27887 = ( n27796 & ~n27885 ) | ( n27796 & n27886 ) | ( ~n27885 & n27886 ) ;
  assign n27888 = ( n1942 & ~n4385 ) | ( n1942 & n16158 ) | ( ~n4385 & n16158 ) ;
  assign n27889 = ( n6395 & ~n19045 ) | ( n6395 & n19771 ) | ( ~n19045 & n19771 ) ;
  assign n27890 = n27889 ^ n17909 ^ n10580 ;
  assign n27891 = ( n19816 & ~n27888 ) | ( n19816 & n27890 ) | ( ~n27888 & n27890 ) ;
  assign n27892 = ( ~n5266 & n5941 ) | ( ~n5266 & n18026 ) | ( n5941 & n18026 ) ;
  assign n27893 = n27892 ^ n766 ^ n600 ;
  assign n27894 = n27893 ^ n11369 ^ 1'b0 ;
  assign n27895 = n26700 | n27894 ;
  assign n27896 = ( n4153 & n9958 ) | ( n4153 & ~n20911 ) | ( n9958 & ~n20911 ) ;
  assign n27897 = n22179 ^ n17081 ^ n1629 ;
  assign n27898 = n6616 & ~n18548 ;
  assign n27899 = n27898 ^ n3978 ^ 1'b0 ;
  assign n27900 = ( ~n8548 & n17742 ) | ( ~n8548 & n27208 ) | ( n17742 & n27208 ) ;
  assign n27901 = n27900 ^ n18308 ^ 1'b0 ;
  assign n27902 = ( ~n385 & n26237 ) | ( ~n385 & n27901 ) | ( n26237 & n27901 ) ;
  assign n27903 = ( n7009 & ~n8325 ) | ( n7009 & n24620 ) | ( ~n8325 & n24620 ) ;
  assign n27905 = ( n9075 & n11531 ) | ( n9075 & n15594 ) | ( n11531 & n15594 ) ;
  assign n27904 = ( n9431 & ~n9833 ) | ( n9431 & n19507 ) | ( ~n9833 & n19507 ) ;
  assign n27906 = n27905 ^ n27904 ^ n10186 ;
  assign n27912 = n9820 ^ n1144 ^ 1'b0 ;
  assign n27910 = n4534 & ~n12390 ;
  assign n27907 = ( n7509 & n8191 ) | ( n7509 & n17750 ) | ( n8191 & n17750 ) ;
  assign n27908 = ( n7457 & n8428 ) | ( n7457 & n27907 ) | ( n8428 & n27907 ) ;
  assign n27909 = n23395 & ~n27908 ;
  assign n27911 = n27910 ^ n27909 ^ n20370 ;
  assign n27913 = n27912 ^ n27911 ^ n9722 ;
  assign n27914 = ~n6844 & n22297 ;
  assign n27915 = ( n13522 & ~n15256 ) | ( n13522 & n27914 ) | ( ~n15256 & n27914 ) ;
  assign n27916 = ( n10289 & ~n20183 ) | ( n10289 & n20890 ) | ( ~n20183 & n20890 ) ;
  assign n27917 = n27916 ^ n23128 ^ 1'b0 ;
  assign n27919 = n6612 ^ n2115 ^ n617 ;
  assign n27918 = ( ~n2218 & n8632 ) | ( ~n2218 & n13711 ) | ( n8632 & n13711 ) ;
  assign n27920 = n27919 ^ n27918 ^ x225 ;
  assign n27921 = n11548 ^ n7816 ^ n1205 ;
  assign n27922 = n27921 ^ n10579 ^ n5790 ;
  assign n27923 = n18909 & ~n27922 ;
  assign n27925 = ( n10339 & ~n11412 ) | ( n10339 & n13054 ) | ( ~n11412 & n13054 ) ;
  assign n27924 = n2525 & ~n4791 ;
  assign n27926 = n27925 ^ n27924 ^ 1'b0 ;
  assign n27927 = n27886 ^ n14257 ^ n13142 ;
  assign n27928 = ( ~n1364 & n6296 ) | ( ~n1364 & n17213 ) | ( n6296 & n17213 ) ;
  assign n27929 = n9431 & ~n24555 ;
  assign n27930 = ( ~n8631 & n27928 ) | ( ~n8631 & n27929 ) | ( n27928 & n27929 ) ;
  assign n27931 = n22249 | n24858 ;
  assign n27932 = ( n1383 & n10567 ) | ( n1383 & ~n27410 ) | ( n10567 & ~n27410 ) ;
  assign n27933 = n27932 ^ n4841 ^ n2740 ;
  assign n27934 = n27933 ^ n3455 ^ 1'b0 ;
  assign n27935 = ( n973 & n10106 ) | ( n973 & ~n15811 ) | ( n10106 & ~n15811 ) ;
  assign n27936 = n17282 | n27935 ;
  assign n27937 = n27936 ^ n16123 ^ 1'b0 ;
  assign n27938 = n27937 ^ n19640 ^ 1'b0 ;
  assign n27939 = ~n27934 & n27938 ;
  assign n27940 = n20972 ^ n19551 ^ n8408 ;
  assign n27941 = ( n5159 & n8151 ) | ( n5159 & ~n27940 ) | ( n8151 & ~n27940 ) ;
  assign n27942 = ( n1299 & n10062 ) | ( n1299 & ~n27941 ) | ( n10062 & ~n27941 ) ;
  assign n27943 = ~n822 & n13021 ;
  assign n27944 = ( n8334 & ~n22450 ) | ( n8334 & n27943 ) | ( ~n22450 & n27943 ) ;
  assign n27947 = n21589 ^ n8671 ^ n5408 ;
  assign n27948 = n15357 | n27947 ;
  assign n27949 = n20545 & ~n27948 ;
  assign n27945 = n13201 ^ n3079 ^ 1'b0 ;
  assign n27946 = n27945 ^ n15264 ^ n8182 ;
  assign n27950 = n27949 ^ n27946 ^ n4726 ;
  assign n27951 = n27950 ^ n1581 ^ n1144 ;
  assign n27952 = n27951 ^ n16011 ^ n6559 ;
  assign n27957 = ~n9144 & n15987 ;
  assign n27958 = n27957 ^ n3525 ^ 1'b0 ;
  assign n27953 = n27634 ^ n5439 ^ n861 ;
  assign n27954 = n2828 & n27953 ;
  assign n27955 = n27954 ^ n18083 ^ 1'b0 ;
  assign n27956 = ( n3096 & n23115 ) | ( n3096 & ~n27955 ) | ( n23115 & ~n27955 ) ;
  assign n27959 = n27958 ^ n27956 ^ n7768 ;
  assign n27960 = ( ~n2299 & n8506 ) | ( ~n2299 & n9659 ) | ( n8506 & n9659 ) ;
  assign n27961 = n21358 & n24882 ;
  assign n27962 = n6980 & n27961 ;
  assign n27963 = n27960 & ~n27962 ;
  assign n27964 = ~n27005 & n27405 ;
  assign n27965 = n27964 ^ n18593 ^ 1'b0 ;
  assign n27966 = n10645 & n22495 ;
  assign n27967 = n27966 ^ n15781 ^ 1'b0 ;
  assign n27968 = ~n9265 & n13516 ;
  assign n27969 = n27968 ^ n11986 ^ n1697 ;
  assign n27970 = n6056 & n12808 ;
  assign n27971 = n24076 ^ n20360 ^ n8830 ;
  assign n27972 = ~n8181 & n27971 ;
  assign n27973 = n764 | n4938 ;
  assign n27974 = n19006 & ~n27973 ;
  assign n27975 = n24021 ^ n15923 ^ n5430 ;
  assign n27989 = ~n3100 & n3679 ;
  assign n27990 = n10277 | n27989 ;
  assign n27991 = n5660 & ~n27990 ;
  assign n27976 = n18022 ^ n3913 ^ n3328 ;
  assign n27977 = ( n5820 & ~n17138 ) | ( n5820 & n27976 ) | ( ~n17138 & n27976 ) ;
  assign n27979 = n23620 ^ n13411 ^ n10911 ;
  assign n27980 = ( n3243 & ~n13800 ) | ( n3243 & n27979 ) | ( ~n13800 & n27979 ) ;
  assign n27978 = n17471 ^ n8394 ^ n5882 ;
  assign n27981 = n27980 ^ n27978 ^ 1'b0 ;
  assign n27982 = n13748 & n27981 ;
  assign n27983 = n8504 ^ n7562 ^ n7412 ;
  assign n27984 = n19268 & ~n26442 ;
  assign n27985 = ~n11687 & n27984 ;
  assign n27986 = n7027 & ~n27985 ;
  assign n27987 = n27983 & n27986 ;
  assign n27988 = ( ~n27977 & n27982 ) | ( ~n27977 & n27987 ) | ( n27982 & n27987 ) ;
  assign n27992 = n27991 ^ n27988 ^ n9578 ;
  assign n27993 = ( n5703 & ~n20530 ) | ( n5703 & n27992 ) | ( ~n20530 & n27992 ) ;
  assign n27994 = ( n2558 & n7046 ) | ( n2558 & ~n16251 ) | ( n7046 & ~n16251 ) ;
  assign n27995 = n4910 | n13301 ;
  assign n27996 = n27995 ^ n15379 ^ 1'b0 ;
  assign n27997 = ( n9069 & ~n10513 ) | ( n9069 & n27996 ) | ( ~n10513 & n27996 ) ;
  assign n27998 = ( n8228 & ~n13154 ) | ( n8228 & n27997 ) | ( ~n13154 & n27997 ) ;
  assign n27999 = n27998 ^ n15374 ^ n5899 ;
  assign n28000 = n5577 ^ n3253 ^ n2978 ;
  assign n28001 = ( n12420 & n21707 ) | ( n12420 & ~n28000 ) | ( n21707 & ~n28000 ) ;
  assign n28002 = n12369 ^ n9980 ^ n9443 ;
  assign n28003 = ~n12938 & n28002 ;
  assign n28004 = n5138 ^ n494 ^ 1'b0 ;
  assign n28005 = n25915 & n28004 ;
  assign n28006 = n9055 ^ n4610 ^ x180 ;
  assign n28007 = n28006 ^ n12218 ^ 1'b0 ;
  assign n28008 = n14023 & ~n28007 ;
  assign n28009 = ( n12502 & ~n14622 ) | ( n12502 & n18667 ) | ( ~n14622 & n18667 ) ;
  assign n28010 = n28009 ^ n1013 ^ 1'b0 ;
  assign n28021 = ( n1093 & n8441 ) | ( n1093 & n16357 ) | ( n8441 & n16357 ) ;
  assign n28020 = ~n5707 & n9012 ;
  assign n28022 = n28021 ^ n28020 ^ n1039 ;
  assign n28023 = n28022 ^ n21496 ^ n8095 ;
  assign n28011 = n4403 | n20761 ;
  assign n28012 = n28011 ^ n8570 ^ 1'b0 ;
  assign n28013 = n18507 & n18963 ;
  assign n28014 = n28013 ^ n5272 ^ 1'b0 ;
  assign n28015 = n28014 ^ n17044 ^ n8728 ;
  assign n28016 = n28015 ^ n27298 ^ n6373 ;
  assign n28017 = n28016 ^ n19750 ^ n10443 ;
  assign n28018 = ~n23979 & n28017 ;
  assign n28019 = ( n5598 & n28012 ) | ( n5598 & n28018 ) | ( n28012 & n28018 ) ;
  assign n28024 = n28023 ^ n28019 ^ n26135 ;
  assign n28025 = n2787 & ~n11978 ;
  assign n28026 = n28025 ^ n13098 ^ 1'b0 ;
  assign n28027 = ( n7246 & ~n15315 ) | ( n7246 & n28026 ) | ( ~n15315 & n28026 ) ;
  assign n28028 = ~n9683 & n9838 ;
  assign n28029 = n28028 ^ n7290 ^ 1'b0 ;
  assign n28030 = ( n2631 & ~n12132 ) | ( n2631 & n24466 ) | ( ~n12132 & n24466 ) ;
  assign n28031 = ~n3867 & n10048 ;
  assign n28032 = ( ~n1495 & n17275 ) | ( ~n1495 & n28031 ) | ( n17275 & n28031 ) ;
  assign n28034 = ( ~n5657 & n13877 ) | ( ~n5657 & n16354 ) | ( n13877 & n16354 ) ;
  assign n28033 = n19880 | n24555 ;
  assign n28035 = n28034 ^ n28033 ^ 1'b0 ;
  assign n28036 = ( ~n7043 & n25666 ) | ( ~n7043 & n28035 ) | ( n25666 & n28035 ) ;
  assign n28037 = n1254 | n27192 ;
  assign n28038 = n28037 ^ n7455 ^ 1'b0 ;
  assign n28039 = n27619 ^ n16779 ^ n13804 ;
  assign n28040 = ( n5570 & n12196 ) | ( n5570 & ~n28039 ) | ( n12196 & ~n28039 ) ;
  assign n28041 = n28040 ^ n21269 ^ n11391 ;
  assign n28042 = ( n11044 & ~n28038 ) | ( n11044 & n28041 ) | ( ~n28038 & n28041 ) ;
  assign n28043 = n13936 ^ n9197 ^ n9132 ;
  assign n28044 = n8315 & ~n28043 ;
  assign n28045 = ( ~n28036 & n28042 ) | ( ~n28036 & n28044 ) | ( n28042 & n28044 ) ;
  assign n28046 = n19435 ^ n14368 ^ n7314 ;
  assign n28048 = n1834 ^ n1424 ^ n1036 ;
  assign n28047 = ( n311 & n1423 ) | ( n311 & ~n15152 ) | ( n1423 & ~n15152 ) ;
  assign n28049 = n28048 ^ n28047 ^ n11069 ;
  assign n28051 = n4837 & n20058 ;
  assign n28050 = n25611 ^ n6181 ^ n1191 ;
  assign n28052 = n28051 ^ n28050 ^ n1870 ;
  assign n28053 = ( n804 & n3548 ) | ( n804 & n18296 ) | ( n3548 & n18296 ) ;
  assign n28054 = ( n9052 & ~n16473 ) | ( n9052 & n17632 ) | ( ~n16473 & n17632 ) ;
  assign n28055 = n11475 ^ n6975 ^ n1627 ;
  assign n28056 = n28055 ^ n6214 ^ n4849 ;
  assign n28057 = ( n4631 & n26125 ) | ( n4631 & n28056 ) | ( n26125 & n28056 ) ;
  assign n28064 = n9189 | n15586 ;
  assign n28065 = n28064 ^ n1168 ^ 1'b0 ;
  assign n28067 = ( n3182 & ~n10089 ) | ( n3182 & n20139 ) | ( ~n10089 & n20139 ) ;
  assign n28066 = n15602 & ~n18046 ;
  assign n28068 = n28067 ^ n28066 ^ 1'b0 ;
  assign n28069 = ( n15691 & ~n23634 ) | ( n15691 & n28068 ) | ( ~n23634 & n28068 ) ;
  assign n28070 = ( n17382 & n28065 ) | ( n17382 & n28069 ) | ( n28065 & n28069 ) ;
  assign n28058 = n18866 ^ n12020 ^ x205 ;
  assign n28059 = n10812 ^ n2805 ^ 1'b0 ;
  assign n28060 = n1610 | n28059 ;
  assign n28061 = n28060 ^ n6938 ^ 1'b0 ;
  assign n28062 = ( n6196 & n10407 ) | ( n6196 & ~n15460 ) | ( n10407 & ~n15460 ) ;
  assign n28063 = ( ~n28058 & n28061 ) | ( ~n28058 & n28062 ) | ( n28061 & n28062 ) ;
  assign n28071 = n28070 ^ n28063 ^ 1'b0 ;
  assign n28072 = n22012 & ~n28071 ;
  assign n28073 = ( n28054 & n28057 ) | ( n28054 & n28072 ) | ( n28057 & n28072 ) ;
  assign n28074 = ( n10431 & n28053 ) | ( n10431 & ~n28073 ) | ( n28053 & ~n28073 ) ;
  assign n28075 = n15376 ^ n7673 ^ n2107 ;
  assign n28076 = n24030 ^ n19346 ^ 1'b0 ;
  assign n28077 = ( n1601 & n9776 ) | ( n1601 & n25765 ) | ( n9776 & n25765 ) ;
  assign n28078 = n4604 ^ n1427 ^ 1'b0 ;
  assign n28079 = ( n3433 & ~n28077 ) | ( n3433 & n28078 ) | ( ~n28077 & n28078 ) ;
  assign n28080 = ( ~n22732 & n28076 ) | ( ~n22732 & n28079 ) | ( n28076 & n28079 ) ;
  assign n28081 = ~n1026 & n8294 ;
  assign n28082 = n28081 ^ n8315 ^ 1'b0 ;
  assign n28083 = n28082 ^ n15715 ^ 1'b0 ;
  assign n28084 = n3361 & n15864 ;
  assign n28085 = n28084 ^ n7253 ^ 1'b0 ;
  assign n28086 = n28083 & ~n28085 ;
  assign n28087 = ( n3026 & n8377 ) | ( n3026 & ~n18933 ) | ( n8377 & ~n18933 ) ;
  assign n28088 = ( n7174 & n7429 ) | ( n7174 & n7516 ) | ( n7429 & n7516 ) ;
  assign n28089 = ( n27339 & n28087 ) | ( n27339 & ~n28088 ) | ( n28087 & ~n28088 ) ;
  assign n28090 = ( n10828 & ~n14777 ) | ( n10828 & n25608 ) | ( ~n14777 & n25608 ) ;
  assign n28091 = n28090 ^ n19285 ^ n4011 ;
  assign n28092 = ( n4028 & n20243 ) | ( n4028 & ~n28091 ) | ( n20243 & ~n28091 ) ;
  assign n28093 = n28092 ^ n26022 ^ n21930 ;
  assign n28094 = n5266 | n6368 ;
  assign n28095 = n28094 ^ n1252 ^ 1'b0 ;
  assign n28096 = ( ~n6899 & n16741 ) | ( ~n6899 & n21180 ) | ( n16741 & n21180 ) ;
  assign n28097 = n14719 ^ n3146 ^ n2590 ;
  assign n28098 = ( n16463 & n18138 ) | ( n16463 & n28097 ) | ( n18138 & n28097 ) ;
  assign n28099 = n23130 ^ n7986 ^ 1'b0 ;
  assign n28100 = ( n9767 & n28098 ) | ( n9767 & n28099 ) | ( n28098 & n28099 ) ;
  assign n28101 = ( ~n1469 & n13639 ) | ( ~n1469 & n15630 ) | ( n13639 & n15630 ) ;
  assign n28102 = n28101 ^ n21694 ^ n5566 ;
  assign n28103 = n27867 ^ n25708 ^ n25486 ;
  assign n28104 = n28103 ^ n17299 ^ n12014 ;
  assign n28105 = n8436 | n25157 ;
  assign n28106 = n14114 | n28105 ;
  assign n28107 = n28106 ^ n15153 ^ n11711 ;
  assign n28108 = ( n15141 & n26086 ) | ( n15141 & n28107 ) | ( n26086 & n28107 ) ;
  assign n28109 = ( n9079 & n13400 ) | ( n9079 & ~n28108 ) | ( n13400 & ~n28108 ) ;
  assign n28110 = ( n4359 & ~n20416 ) | ( n4359 & n20447 ) | ( ~n20416 & n20447 ) ;
  assign n28111 = n28110 ^ n27459 ^ 1'b0 ;
  assign n28112 = ~n4241 & n9723 ;
  assign n28113 = ~n5833 & n28112 ;
  assign n28114 = n14425 ^ n6851 ^ n6024 ;
  assign n28115 = ( ~n3661 & n28113 ) | ( ~n3661 & n28114 ) | ( n28113 & n28114 ) ;
  assign n28116 = n622 & ~n10814 ;
  assign n28117 = ~n17233 & n28116 ;
  assign n28118 = ( n2421 & n25989 ) | ( n2421 & ~n28117 ) | ( n25989 & ~n28117 ) ;
  assign n28120 = x181 & n23573 ;
  assign n28119 = ~n14456 & n19021 ;
  assign n28121 = n28120 ^ n28119 ^ 1'b0 ;
  assign n28123 = ~n7314 & n17478 ;
  assign n28124 = ( n18727 & n25377 ) | ( n18727 & n28123 ) | ( n25377 & n28123 ) ;
  assign n28122 = ( n3435 & n5966 ) | ( n3435 & n20538 ) | ( n5966 & n20538 ) ;
  assign n28125 = n28124 ^ n28122 ^ n9217 ;
  assign n28126 = ~n660 & n28125 ;
  assign n28127 = n28126 ^ n22275 ^ n5885 ;
  assign n28128 = n21658 ^ n6931 ^ n2824 ;
  assign n28129 = n28128 ^ n25365 ^ n551 ;
  assign n28136 = ~n1656 & n1922 ;
  assign n28130 = n10617 ^ n4991 ^ x27 ;
  assign n28131 = ( n11318 & n22083 ) | ( n11318 & n28130 ) | ( n22083 & n28130 ) ;
  assign n28132 = n27925 ^ n16010 ^ n10944 ;
  assign n28133 = ( n22445 & n22628 ) | ( n22445 & ~n28132 ) | ( n22628 & ~n28132 ) ;
  assign n28134 = ( n8345 & n28131 ) | ( n8345 & n28133 ) | ( n28131 & n28133 ) ;
  assign n28135 = n28134 ^ n20264 ^ n5255 ;
  assign n28137 = n28136 ^ n28135 ^ n8124 ;
  assign n28140 = ~n8673 & n16762 ;
  assign n28138 = n6544 ^ n5118 ^ n1551 ;
  assign n28139 = n28138 ^ n5884 ^ n1343 ;
  assign n28141 = n28140 ^ n28139 ^ n14329 ;
  assign n28142 = ( n2265 & n4133 ) | ( n2265 & n4729 ) | ( n4133 & n4729 ) ;
  assign n28143 = n28142 ^ n11882 ^ n7857 ;
  assign n28144 = ( ~n11829 & n20767 ) | ( ~n11829 & n28143 ) | ( n20767 & n28143 ) ;
  assign n28145 = n28144 ^ n28084 ^ n13151 ;
  assign n28146 = ( x173 & ~n12926 ) | ( x173 & n17242 ) | ( ~n12926 & n17242 ) ;
  assign n28147 = n11427 | n28146 ;
  assign n28148 = n9411 & ~n28147 ;
  assign n28149 = ( ~n17683 & n21151 ) | ( ~n17683 & n21965 ) | ( n21151 & n21965 ) ;
  assign n28150 = n28149 ^ n846 ^ 1'b0 ;
  assign n28151 = ( n16787 & ~n23786 ) | ( n16787 & n28150 ) | ( ~n23786 & n28150 ) ;
  assign n28152 = ( n13444 & n28148 ) | ( n13444 & n28151 ) | ( n28148 & n28151 ) ;
  assign n28153 = n21692 & n28152 ;
  assign n28154 = n8989 ^ n2389 ^ 1'b0 ;
  assign n28155 = ( n2170 & n22704 ) | ( n2170 & ~n22984 ) | ( n22704 & ~n22984 ) ;
  assign n28156 = ( ~n20965 & n28154 ) | ( ~n20965 & n28155 ) | ( n28154 & n28155 ) ;
  assign n28157 = ~n8395 & n16663 ;
  assign n28158 = ( ~n1935 & n3628 ) | ( ~n1935 & n12035 ) | ( n3628 & n12035 ) ;
  assign n28159 = n28158 ^ n18084 ^ n5024 ;
  assign n28160 = n15236 ^ n10209 ^ n9106 ;
  assign n28161 = ( n10048 & n22945 ) | ( n10048 & ~n24771 ) | ( n22945 & ~n24771 ) ;
  assign n28162 = ( n14353 & n17716 ) | ( n14353 & n28161 ) | ( n17716 & n28161 ) ;
  assign n28163 = ( n7060 & ~n19932 ) | ( n7060 & n28162 ) | ( ~n19932 & n28162 ) ;
  assign n28164 = ( n417 & n3685 ) | ( n417 & ~n5531 ) | ( n3685 & ~n5531 ) ;
  assign n28165 = n5614 | n7660 ;
  assign n28166 = n21419 & ~n28165 ;
  assign n28167 = ( n22594 & ~n28164 ) | ( n22594 & n28166 ) | ( ~n28164 & n28166 ) ;
  assign n28168 = n21436 ^ n16033 ^ n11209 ;
  assign n28169 = n12498 & n13304 ;
  assign n28170 = n22577 ^ n10389 ^ n2316 ;
  assign n28171 = ~n11464 & n28170 ;
  assign n28172 = n10363 & n28171 ;
  assign n28173 = n6714 ^ n3322 ^ 1'b0 ;
  assign n28174 = n2731 & ~n28173 ;
  assign n28175 = n19857 ^ n19181 ^ 1'b0 ;
  assign n28176 = ~n23553 & n28175 ;
  assign n28177 = ( n939 & n12693 ) | ( n939 & ~n28176 ) | ( n12693 & ~n28176 ) ;
  assign n28178 = n19558 ^ n11948 ^ n10073 ;
  assign n28179 = n11068 & ~n28178 ;
  assign n28180 = n11223 | n28179 ;
  assign n28181 = ( n28174 & n28177 ) | ( n28174 & n28180 ) | ( n28177 & n28180 ) ;
  assign n28182 = n28181 ^ n22478 ^ n13904 ;
  assign n28184 = ( n5565 & n6970 ) | ( n5565 & n13803 ) | ( n6970 & n13803 ) ;
  assign n28185 = ~n1626 & n28184 ;
  assign n28186 = ~n7401 & n28185 ;
  assign n28183 = ( n13430 & n13750 ) | ( n13430 & n22559 ) | ( n13750 & n22559 ) ;
  assign n28187 = n28186 ^ n28183 ^ n9128 ;
  assign n28188 = ~n4014 & n12166 ;
  assign n28189 = n25283 ^ n14220 ^ n13976 ;
  assign n28190 = n28188 | n28189 ;
  assign n28197 = ( n697 & n2732 ) | ( n697 & n11004 ) | ( n2732 & n11004 ) ;
  assign n28198 = n6890 ^ n5015 ^ 1'b0 ;
  assign n28199 = ~n28197 & n28198 ;
  assign n28200 = ( n4633 & n23867 ) | ( n4633 & n28199 ) | ( n23867 & n28199 ) ;
  assign n28196 = n10320 ^ n3979 ^ n3040 ;
  assign n28194 = ( ~n4021 & n8582 ) | ( ~n4021 & n15941 ) | ( n8582 & n15941 ) ;
  assign n28192 = n19375 ^ n14468 ^ 1'b0 ;
  assign n28193 = n815 & ~n28192 ;
  assign n28191 = n11695 ^ n4807 ^ 1'b0 ;
  assign n28195 = n28194 ^ n28193 ^ n28191 ;
  assign n28201 = n28200 ^ n28196 ^ n28195 ;
  assign n28202 = n24352 ^ n19967 ^ n3123 ;
  assign n28203 = ( ~n8784 & n10923 ) | ( ~n8784 & n24179 ) | ( n10923 & n24179 ) ;
  assign n28204 = n28202 & n28203 ;
  assign n28212 = n15542 ^ n7607 ^ n4143 ;
  assign n28210 = ( n3629 & ~n7989 ) | ( n3629 & n14231 ) | ( ~n7989 & n14231 ) ;
  assign n28209 = n2208 | n21382 ;
  assign n28211 = n28210 ^ n28209 ^ 1'b0 ;
  assign n28213 = n28212 ^ n28211 ^ n5907 ;
  assign n28205 = ~n455 & n10165 ;
  assign n28206 = n28205 ^ n7329 ^ 1'b0 ;
  assign n28207 = ( n20234 & n27524 ) | ( n20234 & n28206 ) | ( n27524 & n28206 ) ;
  assign n28208 = ~n18630 & n28207 ;
  assign n28214 = n28213 ^ n28208 ^ 1'b0 ;
  assign n28215 = n7689 ^ n6390 ^ 1'b0 ;
  assign n28216 = n12689 & n28215 ;
  assign n28217 = n21500 & ~n21529 ;
  assign n28218 = n21211 ^ n15129 ^ n12785 ;
  assign n28219 = n23101 ^ n16575 ^ 1'b0 ;
  assign n28220 = n20971 & ~n28219 ;
  assign n28221 = n28220 ^ n7172 ^ n1153 ;
  assign n28222 = ~n1669 & n22058 ;
  assign n28223 = n28222 ^ n3772 ^ 1'b0 ;
  assign n28224 = n21457 ^ n4978 ^ 1'b0 ;
  assign n28225 = ~n28223 & n28224 ;
  assign n28226 = n22998 ^ n13313 ^ n4395 ;
  assign n28227 = n11835 & ~n12995 ;
  assign n28228 = n4172 & n28227 ;
  assign n28229 = ( ~n4497 & n7572 ) | ( ~n4497 & n28228 ) | ( n7572 & n28228 ) ;
  assign n28230 = ( ~n9236 & n28226 ) | ( ~n9236 & n28229 ) | ( n28226 & n28229 ) ;
  assign n28231 = ~n11983 & n28230 ;
  assign n28232 = n623 & n28231 ;
  assign n28233 = ( ~n9141 & n9764 ) | ( ~n9141 & n22642 ) | ( n9764 & n22642 ) ;
  assign n28234 = ~n17030 & n28233 ;
  assign n28235 = n28232 & n28234 ;
  assign n28243 = n7612 & ~n21081 ;
  assign n28244 = n28243 ^ n25051 ^ 1'b0 ;
  assign n28241 = n24874 ^ n22189 ^ 1'b0 ;
  assign n28242 = n28241 ^ n1535 ^ n551 ;
  assign n28236 = n22946 ^ n1138 ^ 1'b0 ;
  assign n28237 = ~n1922 & n28236 ;
  assign n28238 = n20805 ^ n10319 ^ n623 ;
  assign n28239 = ( n5399 & n17050 ) | ( n5399 & ~n28238 ) | ( n17050 & ~n28238 ) ;
  assign n28240 = ( n11446 & n28237 ) | ( n11446 & ~n28239 ) | ( n28237 & ~n28239 ) ;
  assign n28245 = n28244 ^ n28242 ^ n28240 ;
  assign n28246 = ( n2524 & n7293 ) | ( n2524 & ~n13352 ) | ( n7293 & ~n13352 ) ;
  assign n28248 = ( n4254 & n8145 ) | ( n4254 & n20335 ) | ( n8145 & n20335 ) ;
  assign n28249 = n17126 & ~n28248 ;
  assign n28247 = n569 | n24274 ;
  assign n28250 = n28249 ^ n28247 ^ 1'b0 ;
  assign n28251 = n6590 & ~n28250 ;
  assign n28252 = ( n4048 & ~n5900 ) | ( n4048 & n14659 ) | ( ~n5900 & n14659 ) ;
  assign n28256 = n18326 ^ n6439 ^ n1731 ;
  assign n28253 = n6293 & ~n23332 ;
  assign n28254 = ~n10226 & n28253 ;
  assign n28255 = n23903 | n28254 ;
  assign n28257 = n28256 ^ n28255 ^ 1'b0 ;
  assign n28258 = ( ~n1447 & n4804 ) | ( ~n1447 & n20852 ) | ( n4804 & n20852 ) ;
  assign n28259 = n1753 | n24901 ;
  assign n28260 = n28259 ^ n10775 ^ 1'b0 ;
  assign n28261 = n1830 & n11641 ;
  assign n28262 = n28261 ^ n3212 ^ 1'b0 ;
  assign n28263 = n28262 ^ n20998 ^ n18665 ;
  assign n28264 = ( ~n12168 & n28260 ) | ( ~n12168 & n28263 ) | ( n28260 & n28263 ) ;
  assign n28265 = ( ~n532 & n9886 ) | ( ~n532 & n13340 ) | ( n9886 & n13340 ) ;
  assign n28266 = ( ~x216 & n4719 ) | ( ~x216 & n28265 ) | ( n4719 & n28265 ) ;
  assign n28267 = ~n18840 & n28266 ;
  assign n28269 = n3906 | n6072 ;
  assign n28270 = n10837 ^ n10272 ^ n4741 ;
  assign n28271 = ( n8314 & n25603 ) | ( n8314 & ~n28270 ) | ( n25603 & ~n28270 ) ;
  assign n28272 = ( n3845 & n28269 ) | ( n3845 & n28271 ) | ( n28269 & n28271 ) ;
  assign n28268 = n16273 ^ n3341 ^ n1190 ;
  assign n28273 = n28272 ^ n28268 ^ n27221 ;
  assign n28274 = n23131 ^ n16364 ^ n6139 ;
  assign n28275 = n28274 ^ n8375 ^ n5941 ;
  assign n28276 = x123 & n10726 ;
  assign n28277 = n28276 ^ n6658 ^ 1'b0 ;
  assign n28278 = ( ~n5286 & n12994 ) | ( ~n5286 & n28277 ) | ( n12994 & n28277 ) ;
  assign n28279 = n28278 ^ n1806 ^ 1'b0 ;
  assign n28280 = ( n6694 & ~n13116 ) | ( n6694 & n25086 ) | ( ~n13116 & n25086 ) ;
  assign n28281 = ( n5151 & ~n25538 ) | ( n5151 & n28280 ) | ( ~n25538 & n28280 ) ;
  assign n28282 = n16712 ^ n6285 ^ 1'b0 ;
  assign n28284 = n2851 ^ n1325 ^ x10 ;
  assign n28283 = n600 & n12682 ;
  assign n28285 = n28284 ^ n28283 ^ 1'b0 ;
  assign n28286 = n28285 ^ n11929 ^ n10966 ;
  assign n28287 = n28286 ^ n15857 ^ 1'b0 ;
  assign n28288 = n14218 ^ n5805 ^ n2586 ;
  assign n28289 = ( n4399 & n12390 ) | ( n4399 & n28288 ) | ( n12390 & n28288 ) ;
  assign n28290 = n18419 | n28012 ;
  assign n28291 = ( n402 & n7199 ) | ( n402 & ~n28290 ) | ( n7199 & ~n28290 ) ;
  assign n28292 = n28291 ^ n18022 ^ n364 ;
  assign n28293 = n3776 ^ n3300 ^ 1'b0 ;
  assign n28294 = ( n5050 & n28292 ) | ( n5050 & ~n28293 ) | ( n28292 & ~n28293 ) ;
  assign n28295 = n24645 ^ n23511 ^ n5756 ;
  assign n28296 = n28295 ^ n18495 ^ 1'b0 ;
  assign n28297 = n8233 & n28296 ;
  assign n28298 = n14685 & n21578 ;
  assign n28299 = ~n11039 & n27883 ;
  assign n28300 = ( ~n5076 & n7392 ) | ( ~n5076 & n28299 ) | ( n7392 & n28299 ) ;
  assign n28301 = n28300 ^ n15568 ^ n1721 ;
  assign n28302 = n21348 ^ n4466 ^ 1'b0 ;
  assign n28303 = n4859 & ~n10292 ;
  assign n28304 = n28303 ^ n1812 ^ 1'b0 ;
  assign n28305 = n28304 ^ n17594 ^ n5189 ;
  assign n28306 = n24196 | n28305 ;
  assign n28307 = n28306 ^ n20936 ^ 1'b0 ;
  assign n28308 = n17515 ^ n11933 ^ n3417 ;
  assign n28309 = n28308 ^ n9955 ^ n5184 ;
  assign n28310 = ( n1282 & n5900 ) | ( n1282 & ~n11489 ) | ( n5900 & ~n11489 ) ;
  assign n28311 = ( ~n3288 & n16097 ) | ( ~n3288 & n28310 ) | ( n16097 & n28310 ) ;
  assign n28312 = n11962 ^ n11664 ^ n4580 ;
  assign n28313 = ( n4457 & ~n24443 ) | ( n4457 & n28312 ) | ( ~n24443 & n28312 ) ;
  assign n28314 = ( n17322 & n24768 ) | ( n17322 & ~n28313 ) | ( n24768 & ~n28313 ) ;
  assign n28315 = n18646 | n24299 ;
  assign n28316 = n22796 & ~n28315 ;
  assign n28317 = n28316 ^ n24555 ^ n16705 ;
  assign n28318 = ( ~n599 & n11348 ) | ( ~n599 & n19177 ) | ( n11348 & n19177 ) ;
  assign n28319 = n20524 & ~n28318 ;
  assign n28320 = n22847 ^ n9034 ^ n582 ;
  assign n28321 = n7272 | n21778 ;
  assign n28322 = n28320 & ~n28321 ;
  assign n28323 = n28322 ^ n708 ^ 1'b0 ;
  assign n28329 = n25336 ^ n16465 ^ n10668 ;
  assign n28324 = n4066 | n10478 ;
  assign n28325 = n11501 & ~n28324 ;
  assign n28326 = n17699 ^ n9771 ^ 1'b0 ;
  assign n28327 = n28326 ^ n21177 ^ n800 ;
  assign n28328 = ( ~n11300 & n28325 ) | ( ~n11300 & n28327 ) | ( n28325 & n28327 ) ;
  assign n28330 = n28329 ^ n28328 ^ n27042 ;
  assign n28331 = n11996 & ~n24197 ;
  assign n28332 = n28331 ^ n6614 ^ 1'b0 ;
  assign n28333 = n23227 ^ n13517 ^ 1'b0 ;
  assign n28334 = ( ~n9954 & n19699 ) | ( ~n9954 & n28333 ) | ( n19699 & n28333 ) ;
  assign n28335 = n2003 & n28334 ;
  assign n28336 = n28335 ^ n7731 ^ 1'b0 ;
  assign n28337 = n21166 ^ n19183 ^ 1'b0 ;
  assign n28338 = ~n28336 & n28337 ;
  assign n28339 = ( n1317 & n2285 ) | ( n1317 & n8120 ) | ( n2285 & n8120 ) ;
  assign n28340 = ( n1379 & ~n6585 ) | ( n1379 & n28339 ) | ( ~n6585 & n28339 ) ;
  assign n28341 = ( n1389 & ~n5036 ) | ( n1389 & n19297 ) | ( ~n5036 & n19297 ) ;
  assign n28342 = n1384 & ~n15058 ;
  assign n28343 = n4753 & ~n6995 ;
  assign n28344 = ( n28341 & n28342 ) | ( n28341 & n28343 ) | ( n28342 & n28343 ) ;
  assign n28345 = n10236 ^ n2879 ^ n1057 ;
  assign n28346 = ( n680 & n1944 ) | ( n680 & n28345 ) | ( n1944 & n28345 ) ;
  assign n28347 = ( n8358 & n10843 ) | ( n8358 & n28346 ) | ( n10843 & n28346 ) ;
  assign n28348 = ( n28340 & n28344 ) | ( n28340 & n28347 ) | ( n28344 & n28347 ) ;
  assign n28369 = ( ~n12248 & n22080 ) | ( ~n12248 & n23676 ) | ( n22080 & n23676 ) ;
  assign n28349 = n25049 ^ n3437 ^ 1'b0 ;
  assign n28350 = n3315 & n28349 ;
  assign n28351 = n21334 ^ n8231 ^ 1'b0 ;
  assign n28352 = n26279 & ~n28351 ;
  assign n28353 = n28350 & n28352 ;
  assign n28354 = n18558 & n28353 ;
  assign n28361 = n21460 ^ n1315 ^ 1'b0 ;
  assign n28362 = n10450 | n28361 ;
  assign n28363 = n28362 ^ n27983 ^ 1'b0 ;
  assign n28364 = ( ~n413 & n18469 ) | ( ~n413 & n28363 ) | ( n18469 & n28363 ) ;
  assign n28355 = ( n1614 & n18237 ) | ( n1614 & ~n22191 ) | ( n18237 & ~n22191 ) ;
  assign n28356 = x144 & n28355 ;
  assign n28357 = n28356 ^ n19777 ^ 1'b0 ;
  assign n28358 = n28357 ^ n14910 ^ n7792 ;
  assign n28359 = ( ~n14281 & n14606 ) | ( ~n14281 & n15288 ) | ( n14606 & n15288 ) ;
  assign n28360 = n28358 & n28359 ;
  assign n28365 = n28364 ^ n28360 ^ 1'b0 ;
  assign n28366 = ~n7176 & n28365 ;
  assign n28367 = n28366 ^ n16562 ^ 1'b0 ;
  assign n28368 = ( ~n6947 & n28354 ) | ( ~n6947 & n28367 ) | ( n28354 & n28367 ) ;
  assign n28370 = n28369 ^ n28368 ^ n14246 ;
  assign n28371 = n986 & ~n6364 ;
  assign n28372 = n1219 & n28371 ;
  assign n28373 = ( ~n11527 & n14561 ) | ( ~n11527 & n28372 ) | ( n14561 & n28372 ) ;
  assign n28374 = n24956 ^ n21048 ^ n13062 ;
  assign n28375 = n28374 ^ n24111 ^ 1'b0 ;
  assign n28376 = n19300 ^ n14488 ^ n5771 ;
  assign n28377 = n28376 ^ n10641 ^ 1'b0 ;
  assign n28378 = n9758 & n28377 ;
  assign n28379 = ( n13298 & ~n17237 ) | ( n13298 & n24074 ) | ( ~n17237 & n24074 ) ;
  assign n28380 = ( n5493 & n11371 ) | ( n5493 & ~n14967 ) | ( n11371 & ~n14967 ) ;
  assign n28381 = n28379 | n28380 ;
  assign n28386 = n25700 ^ n17618 ^ n15360 ;
  assign n28384 = n6834 ^ n2782 ^ n1975 ;
  assign n28385 = n28384 ^ n10014 ^ n5865 ;
  assign n28382 = ( n9728 & n12691 ) | ( n9728 & n13490 ) | ( n12691 & n13490 ) ;
  assign n28383 = n6630 & ~n28382 ;
  assign n28387 = n28386 ^ n28385 ^ n28383 ;
  assign n28388 = ~n4630 & n10709 ;
  assign n28389 = n28388 ^ n8436 ^ n7466 ;
  assign n28390 = ( n395 & n16166 ) | ( n395 & n18008 ) | ( n16166 & n18008 ) ;
  assign n28391 = x72 & n7850 ;
  assign n28392 = ( n2374 & ~n11647 ) | ( n2374 & n28391 ) | ( ~n11647 & n28391 ) ;
  assign n28393 = n28392 ^ n12462 ^ 1'b0 ;
  assign n28394 = ( x47 & n2850 ) | ( x47 & n7780 ) | ( n2850 & n7780 ) ;
  assign n28395 = n28394 ^ n19466 ^ n7799 ;
  assign n28396 = ( ~n7911 & n10682 ) | ( ~n7911 & n18917 ) | ( n10682 & n18917 ) ;
  assign n28399 = ( ~n5929 & n10917 ) | ( ~n5929 & n14360 ) | ( n10917 & n14360 ) ;
  assign n28397 = n12453 ^ n10061 ^ 1'b0 ;
  assign n28398 = n13039 | n28397 ;
  assign n28400 = n28399 ^ n28398 ^ n2472 ;
  assign n28401 = ( n1275 & ~n11583 ) | ( n1275 & n24741 ) | ( ~n11583 & n24741 ) ;
  assign n28402 = ~n15671 & n21450 ;
  assign n28403 = n22033 & n28402 ;
  assign n28404 = x22 & n18491 ;
  assign n28405 = n28403 & n28404 ;
  assign n28406 = n28405 ^ n22858 ^ x171 ;
  assign n28407 = n28401 & ~n28406 ;
  assign n28408 = n26539 ^ n19390 ^ n5653 ;
  assign n28409 = n28408 ^ n13420 ^ 1'b0 ;
  assign n28410 = n7295 & ~n28409 ;
  assign n28411 = n17958 & n28410 ;
  assign n28412 = n10393 & n16345 ;
  assign n28413 = ~n28411 & n28412 ;
  assign n28414 = n4269 ^ n1125 ^ x234 ;
  assign n28415 = n28414 ^ n15456 ^ n3866 ;
  assign n28416 = n1815 & ~n28415 ;
  assign n28417 = ( n3899 & n16717 ) | ( n3899 & ~n18223 ) | ( n16717 & ~n18223 ) ;
  assign n28418 = ~n19310 & n27465 ;
  assign n28419 = ( ~n4382 & n28417 ) | ( ~n4382 & n28418 ) | ( n28417 & n28418 ) ;
  assign n28420 = n16795 ^ n15309 ^ 1'b0 ;
  assign n28421 = n21533 ^ n680 ^ 1'b0 ;
  assign n28422 = ( ~n8466 & n20928 ) | ( ~n8466 & n23901 ) | ( n20928 & n23901 ) ;
  assign n28423 = ( n968 & ~n28421 ) | ( n968 & n28422 ) | ( ~n28421 & n28422 ) ;
  assign n28425 = n1438 & ~n9914 ;
  assign n28426 = n28425 ^ n342 ^ 1'b0 ;
  assign n28424 = n6426 & ~n18585 ;
  assign n28427 = n28426 ^ n28424 ^ 1'b0 ;
  assign n28428 = ( ~n9185 & n9694 ) | ( ~n9185 & n28427 ) | ( n9694 & n28427 ) ;
  assign n28429 = n28428 ^ n6183 ^ n5328 ;
  assign n28430 = n23638 ^ n8718 ^ n2328 ;
  assign n28431 = n28430 ^ n455 ^ x56 ;
  assign n28432 = n10149 | n28431 ;
  assign n28433 = n28429 | n28432 ;
  assign n28434 = ( ~n10455 & n20146 ) | ( ~n10455 & n28433 ) | ( n20146 & n28433 ) ;
  assign n28435 = n19894 ^ n17333 ^ 1'b0 ;
  assign n28436 = n5902 & n28435 ;
  assign n28437 = n28436 ^ n19626 ^ n12807 ;
  assign n28438 = ( n6955 & n14034 ) | ( n6955 & ~n24087 ) | ( n14034 & ~n24087 ) ;
  assign n28439 = n28438 ^ n20831 ^ 1'b0 ;
  assign n28440 = n12407 & n28439 ;
  assign n28442 = n6015 & ~n14372 ;
  assign n28441 = n21216 ^ n19975 ^ n12534 ;
  assign n28443 = n28442 ^ n28441 ^ n16117 ;
  assign n28444 = ( n13308 & ~n28440 ) | ( n13308 & n28443 ) | ( ~n28440 & n28443 ) ;
  assign n28445 = ( n2421 & ~n12834 ) | ( n2421 & n25380 ) | ( ~n12834 & n25380 ) ;
  assign n28446 = ( n13738 & n22485 ) | ( n13738 & ~n28445 ) | ( n22485 & ~n28445 ) ;
  assign n28447 = n19927 ^ n13754 ^ n9001 ;
  assign n28448 = ( ~n3104 & n6164 ) | ( ~n3104 & n26073 ) | ( n6164 & n26073 ) ;
  assign n28449 = ( n15304 & n25846 ) | ( n15304 & ~n28448 ) | ( n25846 & ~n28448 ) ;
  assign n28450 = ( n6231 & ~n10471 ) | ( n6231 & n20995 ) | ( ~n10471 & n20995 ) ;
  assign n28451 = ( n1604 & n6166 ) | ( n1604 & n7609 ) | ( n6166 & n7609 ) ;
  assign n28452 = n6037 ^ n5902 ^ 1'b0 ;
  assign n28453 = ( n4770 & ~n9452 ) | ( n4770 & n21846 ) | ( ~n9452 & n21846 ) ;
  assign n28454 = n1996 | n4485 ;
  assign n28455 = n28454 ^ n5793 ^ 1'b0 ;
  assign n28456 = n28455 ^ n25707 ^ n12869 ;
  assign n28457 = n20154 ^ n7352 ^ n6509 ;
  assign n28458 = ( n6536 & n28456 ) | ( n6536 & ~n28457 ) | ( n28456 & ~n28457 ) ;
  assign n28459 = ( n11212 & ~n11758 ) | ( n11212 & n24749 ) | ( ~n11758 & n24749 ) ;
  assign n28460 = n27322 ^ n18324 ^ n13455 ;
  assign n28461 = ( n5101 & ~n28459 ) | ( n5101 & n28460 ) | ( ~n28459 & n28460 ) ;
  assign n28462 = n8702 ^ n1908 ^ 1'b0 ;
  assign n28463 = ~n11390 & n28462 ;
  assign n28464 = ( n11364 & ~n17459 ) | ( n11364 & n26372 ) | ( ~n17459 & n26372 ) ;
  assign n28465 = ( ~n5130 & n7517 ) | ( ~n5130 & n23236 ) | ( n7517 & n23236 ) ;
  assign n28466 = n26882 & n28465 ;
  assign n28467 = ( ~n13283 & n14027 ) | ( ~n13283 & n20940 ) | ( n14027 & n20940 ) ;
  assign n28468 = ( n4614 & ~n5760 ) | ( n4614 & n26086 ) | ( ~n5760 & n26086 ) ;
  assign n28469 = n28468 ^ n5384 ^ n1555 ;
  assign n28470 = n6993 ^ n5954 ^ n4546 ;
  assign n28471 = ( ~n1455 & n13274 ) | ( ~n1455 & n14660 ) | ( n13274 & n14660 ) ;
  assign n28472 = ( n3421 & ~n27069 ) | ( n3421 & n28471 ) | ( ~n27069 & n28471 ) ;
  assign n28473 = ( n22713 & n28470 ) | ( n22713 & ~n28472 ) | ( n28470 & ~n28472 ) ;
  assign n28474 = ~n7390 & n28291 ;
  assign n28475 = n28473 & n28474 ;
  assign n28478 = ( n13449 & ~n17742 ) | ( n13449 & n19849 ) | ( ~n17742 & n19849 ) ;
  assign n28479 = ( n6430 & n10866 ) | ( n6430 & ~n28478 ) | ( n10866 & ~n28478 ) ;
  assign n28476 = n2208 & n7775 ;
  assign n28477 = ( n1392 & n20348 ) | ( n1392 & ~n28476 ) | ( n20348 & ~n28476 ) ;
  assign n28480 = n28479 ^ n28477 ^ 1'b0 ;
  assign n28481 = n8365 | n28480 ;
  assign n28482 = n28475 & ~n28481 ;
  assign n28483 = n17025 ^ n7062 ^ n3279 ;
  assign n28484 = n19846 ^ n5003 ^ 1'b0 ;
  assign n28485 = n11002 | n28484 ;
  assign n28488 = n7592 ^ n6837 ^ 1'b0 ;
  assign n28489 = n17853 & n28488 ;
  assign n28487 = n5965 & n6928 ;
  assign n28490 = n28489 ^ n28487 ^ n10269 ;
  assign n28486 = n4064 & n6701 ;
  assign n28491 = n28490 ^ n28486 ^ n22406 ;
  assign n28492 = n19477 ^ n14828 ^ n1658 ;
  assign n28493 = ( ~n525 & n21071 ) | ( ~n525 & n28492 ) | ( n21071 & n28492 ) ;
  assign n28494 = n10498 ^ n8937 ^ n2157 ;
  assign n28495 = ( n22419 & ~n28493 ) | ( n22419 & n28494 ) | ( ~n28493 & n28494 ) ;
  assign n28498 = n4103 ^ n3293 ^ n1062 ;
  assign n28496 = n16060 ^ n15443 ^ x69 ;
  assign n28497 = n28496 ^ n5998 ^ n2363 ;
  assign n28499 = n28498 ^ n28497 ^ n23370 ;
  assign n28500 = ( ~n3984 & n5858 ) | ( ~n3984 & n9944 ) | ( n5858 & n9944 ) ;
  assign n28501 = n9363 & ~n28500 ;
  assign n28505 = n16549 ^ n13925 ^ n4444 ;
  assign n28506 = n19296 ^ n3237 ^ 1'b0 ;
  assign n28507 = ~n19829 & n28506 ;
  assign n28508 = ( n15390 & ~n28505 ) | ( n15390 & n28507 ) | ( ~n28505 & n28507 ) ;
  assign n28509 = n28508 ^ n7226 ^ 1'b0 ;
  assign n28503 = ( n9170 & n9670 ) | ( n9170 & n18897 ) | ( n9670 & n18897 ) ;
  assign n28502 = n13514 ^ n2979 ^ n2900 ;
  assign n28504 = n28503 ^ n28502 ^ n12657 ;
  assign n28510 = n28509 ^ n28504 ^ n19605 ;
  assign n28511 = ( n3911 & ~n15085 ) | ( n3911 & n19169 ) | ( ~n15085 & n19169 ) ;
  assign n28512 = ~n3144 & n28511 ;
  assign n28513 = n13196 ^ n2035 ^ 1'b0 ;
  assign n28514 = ~n9840 & n28513 ;
  assign n28515 = n19313 ^ n15093 ^ 1'b0 ;
  assign n28516 = n17596 ^ n1133 ^ 1'b0 ;
  assign n28517 = n3365 & ~n28516 ;
  assign n28518 = n4361 ^ n1462 ^ 1'b0 ;
  assign n28519 = n28517 & ~n28518 ;
  assign n28520 = ~n1556 & n8725 ;
  assign n28521 = n24024 ^ n19506 ^ 1'b0 ;
  assign n28522 = ~n4795 & n28521 ;
  assign n28523 = ( n6425 & n12381 ) | ( n6425 & n28522 ) | ( n12381 & n28522 ) ;
  assign n28524 = ~n28520 & n28523 ;
  assign n28525 = n13474 & n28524 ;
  assign n28526 = n28525 ^ n10406 ^ n10046 ;
  assign n28527 = n27229 ^ n12555 ^ n2331 ;
  assign n28528 = ( n14794 & ~n22550 ) | ( n14794 & n28527 ) | ( ~n22550 & n28527 ) ;
  assign n28529 = ( n2610 & n6552 ) | ( n2610 & ~n28528 ) | ( n6552 & ~n28528 ) ;
  assign n28530 = n7549 | n15729 ;
  assign n28531 = n2694 & ~n28530 ;
  assign n28532 = n2608 | n28531 ;
  assign n28533 = n28532 ^ n7704 ^ 1'b0 ;
  assign n28534 = n28533 ^ n11243 ^ n9155 ;
  assign n28535 = ~n24610 & n28534 ;
  assign n28536 = ( n1952 & ~n8301 ) | ( n1952 & n8780 ) | ( ~n8301 & n8780 ) ;
  assign n28537 = ( ~n11252 & n16203 ) | ( ~n11252 & n28536 ) | ( n16203 & n28536 ) ;
  assign n28538 = ( n1061 & n6798 ) | ( n1061 & ~n28537 ) | ( n6798 & ~n28537 ) ;
  assign n28539 = ( n25208 & ~n28292 ) | ( n25208 & n28538 ) | ( ~n28292 & n28538 ) ;
  assign n28540 = n18534 ^ n16120 ^ n6229 ;
  assign n28541 = ( n16008 & n21425 ) | ( n16008 & n28540 ) | ( n21425 & n28540 ) ;
  assign n28542 = ~n9964 & n28541 ;
  assign n28543 = ( ~n20815 & n25135 ) | ( ~n20815 & n28542 ) | ( n25135 & n28542 ) ;
  assign n28544 = n3952 | n27243 ;
  assign n28545 = n28544 ^ n9022 ^ 1'b0 ;
  assign n28546 = n15810 ^ n3733 ^ 1'b0 ;
  assign n28547 = ~n1876 & n28546 ;
  assign n28548 = n15677 ^ n13960 ^ n7516 ;
  assign n28549 = n28547 & ~n28548 ;
  assign n28550 = ~n27084 & n28549 ;
  assign n28551 = ( n566 & n4642 ) | ( n566 & n17917 ) | ( n4642 & n17917 ) ;
  assign n28552 = n17280 ^ n5593 ^ 1'b0 ;
  assign n28553 = n20814 ^ n18116 ^ 1'b0 ;
  assign n28554 = n28553 ^ n14253 ^ n8379 ;
  assign n28555 = ( n28551 & n28552 ) | ( n28551 & ~n28554 ) | ( n28552 & ~n28554 ) ;
  assign n28556 = ( n562 & ~n1624 ) | ( n562 & n5418 ) | ( ~n1624 & n5418 ) ;
  assign n28557 = n462 & n17573 ;
  assign n28558 = ~n28556 & n28557 ;
  assign n28559 = ( n1116 & n8279 ) | ( n1116 & ~n28558 ) | ( n8279 & ~n28558 ) ;
  assign n28560 = ( n6610 & n7660 ) | ( n6610 & n23935 ) | ( n7660 & n23935 ) ;
  assign n28561 = ~n3229 & n6483 ;
  assign n28562 = n28561 ^ n2097 ^ 1'b0 ;
  assign n28563 = ( n16406 & n26494 ) | ( n16406 & n28562 ) | ( n26494 & n28562 ) ;
  assign n28569 = n14888 ^ n13100 ^ n1665 ;
  assign n28565 = n2703 & ~n26043 ;
  assign n28566 = n28565 ^ n2393 ^ 1'b0 ;
  assign n28567 = ~n1813 & n28566 ;
  assign n28564 = x81 & ~n3302 ;
  assign n28568 = n28567 ^ n28564 ^ 1'b0 ;
  assign n28570 = n28569 ^ n28568 ^ 1'b0 ;
  assign n28571 = n20826 | n23779 ;
  assign n28577 = n7023 ^ n5168 ^ n2433 ;
  assign n28578 = n9401 | n28577 ;
  assign n28572 = n3697 | n5669 ;
  assign n28573 = ( n1304 & n20455 ) | ( n1304 & ~n20853 ) | ( n20455 & ~n20853 ) ;
  assign n28574 = n10712 & ~n26056 ;
  assign n28575 = ~n28573 & n28574 ;
  assign n28576 = ( n15421 & ~n28572 ) | ( n15421 & n28575 ) | ( ~n28572 & n28575 ) ;
  assign n28579 = n28578 ^ n28576 ^ n10959 ;
  assign n28585 = ( n1601 & n4305 ) | ( n1601 & ~n4802 ) | ( n4305 & ~n4802 ) ;
  assign n28586 = n28585 ^ n2375 ^ n1067 ;
  assign n28584 = n18715 & ~n22583 ;
  assign n28587 = n28586 ^ n28584 ^ 1'b0 ;
  assign n28588 = n4175 | n28587 ;
  assign n28582 = ( n2631 & ~n7431 ) | ( n2631 & n16848 ) | ( ~n7431 & n16848 ) ;
  assign n28583 = n28582 ^ n17987 ^ n7706 ;
  assign n28589 = n28588 ^ n28583 ^ n13049 ;
  assign n28580 = n11929 | n27482 ;
  assign n28581 = n23411 & ~n28580 ;
  assign n28590 = n28589 ^ n28581 ^ n21232 ;
  assign n28595 = n3885 | n6904 ;
  assign n28596 = ( n1528 & ~n13258 ) | ( n1528 & n28595 ) | ( ~n13258 & n28595 ) ;
  assign n28597 = ( n2569 & ~n7051 ) | ( n2569 & n28596 ) | ( ~n7051 & n28596 ) ;
  assign n28598 = n23366 & n28597 ;
  assign n28599 = ~n24085 & n28598 ;
  assign n28591 = ( x236 & n985 ) | ( x236 & ~n5486 ) | ( n985 & ~n5486 ) ;
  assign n28592 = ( n5244 & n5587 ) | ( n5244 & n7056 ) | ( n5587 & n7056 ) ;
  assign n28593 = n5853 & n28592 ;
  assign n28594 = ~n28591 & n28593 ;
  assign n28600 = n28599 ^ n28594 ^ n411 ;
  assign n28602 = n6912 ^ n2933 ^ 1'b0 ;
  assign n28603 = n27905 & n28602 ;
  assign n28601 = ( n1505 & n10662 ) | ( n1505 & ~n18688 ) | ( n10662 & ~n18688 ) ;
  assign n28604 = n28603 ^ n28601 ^ 1'b0 ;
  assign n28605 = n28604 ^ n24058 ^ n2006 ;
  assign n28606 = n13115 ^ n10723 ^ n1001 ;
  assign n28607 = ( n12038 & n21798 ) | ( n12038 & n28606 ) | ( n21798 & n28606 ) ;
  assign n28608 = ~n1303 & n2094 ;
  assign n28609 = ( n11473 & n27370 ) | ( n11473 & n28608 ) | ( n27370 & n28608 ) ;
  assign n28610 = n24146 ^ n14480 ^ n1518 ;
  assign n28611 = n4681 | n23146 ;
  assign n28612 = n9437 | n28611 ;
  assign n28613 = ( n2525 & n8252 ) | ( n2525 & n24679 ) | ( n8252 & n24679 ) ;
  assign n28614 = ( ~n7046 & n17063 ) | ( ~n7046 & n20912 ) | ( n17063 & n20912 ) ;
  assign n28615 = n501 & n15445 ;
  assign n28616 = ~n27791 & n28615 ;
  assign n28617 = n28616 ^ n26725 ^ n3664 ;
  assign n28618 = ~n26327 & n28617 ;
  assign n28619 = n24592 ^ n4103 ^ n3990 ;
  assign n28620 = n27423 ^ n19164 ^ 1'b0 ;
  assign n28621 = n16446 ^ x20 ^ 1'b0 ;
  assign n28622 = n5885 | n28621 ;
  assign n28623 = n28622 ^ n27875 ^ n27518 ;
  assign n28624 = n27578 ^ n20012 ^ n6788 ;
  assign n28625 = ( n15731 & ~n27958 ) | ( n15731 & n28624 ) | ( ~n27958 & n28624 ) ;
  assign n28626 = ( n8209 & n19806 ) | ( n8209 & n28625 ) | ( n19806 & n28625 ) ;
  assign n28627 = ( n14828 & ~n23783 ) | ( n14828 & n25684 ) | ( ~n23783 & n25684 ) ;
  assign n28628 = n28627 ^ n17973 ^ n7377 ;
  assign n28629 = n22597 ^ n19934 ^ n3696 ;
  assign n28630 = n14034 ^ n7066 ^ 1'b0 ;
  assign n28631 = n28630 ^ n17723 ^ 1'b0 ;
  assign n28632 = ~n28629 & n28631 ;
  assign n28633 = ~n19544 & n28632 ;
  assign n28634 = ~n13244 & n20719 ;
  assign n28635 = ~n10050 & n28634 ;
  assign n28636 = ~n3168 & n3176 ;
  assign n28637 = n28635 & n28636 ;
  assign n28638 = n28637 ^ n2509 ^ 1'b0 ;
  assign n28639 = ( n7106 & n25381 ) | ( n7106 & n28638 ) | ( n25381 & n28638 ) ;
  assign n28640 = n27199 ^ n416 ^ 1'b0 ;
  assign n28641 = n297 & ~n17722 ;
  assign n28642 = ~n7875 & n28641 ;
  assign n28643 = n28642 ^ n24761 ^ n2336 ;
  assign n28644 = ~n14199 & n28643 ;
  assign n28645 = ( n1065 & n9958 ) | ( n1065 & ~n13254 ) | ( n9958 & ~n13254 ) ;
  assign n28646 = ( n6885 & n18438 ) | ( n6885 & n28645 ) | ( n18438 & n28645 ) ;
  assign n28648 = ( ~n1428 & n3359 ) | ( ~n1428 & n3910 ) | ( n3359 & n3910 ) ;
  assign n28647 = n1451 & n14419 ;
  assign n28649 = n28648 ^ n28647 ^ 1'b0 ;
  assign n28650 = n5017 ^ n4803 ^ 1'b0 ;
  assign n28651 = n3505 & n28650 ;
  assign n28652 = ( n3265 & n28649 ) | ( n3265 & ~n28651 ) | ( n28649 & ~n28651 ) ;
  assign n28653 = ( n3335 & ~n10671 ) | ( n3335 & n28652 ) | ( ~n10671 & n28652 ) ;
  assign n28654 = n425 & ~n7003 ;
  assign n28655 = n28654 ^ n3086 ^ 1'b0 ;
  assign n28656 = n8022 | n28655 ;
  assign n28657 = ( x243 & n28653 ) | ( x243 & ~n28656 ) | ( n28653 & ~n28656 ) ;
  assign n28658 = ( ~n1474 & n2058 ) | ( ~n1474 & n4087 ) | ( n2058 & n4087 ) ;
  assign n28659 = n28658 ^ n6262 ^ x216 ;
  assign n28660 = ~n2875 & n28659 ;
  assign n28661 = n28660 ^ n6127 ^ 1'b0 ;
  assign n28662 = ~n574 & n11794 ;
  assign n28663 = ~n953 & n28662 ;
  assign n28665 = n8703 ^ n1781 ^ 1'b0 ;
  assign n28664 = x105 & n9766 ;
  assign n28666 = n28665 ^ n28664 ^ 1'b0 ;
  assign n28667 = ~n28663 & n28666 ;
  assign n28668 = n11969 & n28667 ;
  assign n28669 = ( n1190 & n17613 ) | ( n1190 & n28578 ) | ( n17613 & n28578 ) ;
  assign n28670 = n28669 ^ n22462 ^ n6792 ;
  assign n28671 = ( n28661 & n28668 ) | ( n28661 & n28670 ) | ( n28668 & n28670 ) ;
  assign n28672 = n17843 & n25438 ;
  assign n28673 = n28672 ^ n11004 ^ 1'b0 ;
  assign n28674 = n28673 ^ n27165 ^ n13578 ;
  assign n28675 = n21005 ^ n17731 ^ n14411 ;
  assign n28676 = ( ~n25294 & n27951 ) | ( ~n25294 & n28675 ) | ( n27951 & n28675 ) ;
  assign n28677 = n19504 ^ n10570 ^ 1'b0 ;
  assign n28678 = n7607 & n28677 ;
  assign n28681 = ( ~n6006 & n12544 ) | ( ~n6006 & n24054 ) | ( n12544 & n24054 ) ;
  assign n28679 = ( n5623 & ~n10521 ) | ( n5623 & n25777 ) | ( ~n10521 & n25777 ) ;
  assign n28680 = n7417 & n28679 ;
  assign n28682 = n28681 ^ n28680 ^ 1'b0 ;
  assign n28683 = n28682 ^ n6971 ^ 1'b0 ;
  assign n28684 = ~n10554 & n28683 ;
  assign n28685 = ~n10468 & n25792 ;
  assign n28686 = n28685 ^ n7170 ^ 1'b0 ;
  assign n28687 = n12207 | n23185 ;
  assign n28688 = n13547 & ~n14789 ;
  assign n28689 = n25348 & n28688 ;
  assign n28690 = n28687 & ~n28689 ;
  assign n28691 = n18847 ^ n17146 ^ n8787 ;
  assign n28692 = n9001 ^ n3848 ^ n3837 ;
  assign n28693 = ( n2707 & n13469 ) | ( n2707 & ~n28692 ) | ( n13469 & ~n28692 ) ;
  assign n28694 = ( n11523 & n14295 ) | ( n11523 & n28693 ) | ( n14295 & n28693 ) ;
  assign n28695 = n28694 ^ n20672 ^ n8787 ;
  assign n28696 = n23903 ^ n21185 ^ n8776 ;
  assign n28697 = n26407 ^ n1627 ^ 1'b0 ;
  assign n28698 = n17226 | n28697 ;
  assign n28699 = n17381 ^ n10064 ^ 1'b0 ;
  assign n28700 = n25025 | n28699 ;
  assign n28701 = n28700 ^ n929 ^ 1'b0 ;
  assign n28702 = ( n2325 & n6588 ) | ( n2325 & ~n7795 ) | ( n6588 & ~n7795 ) ;
  assign n28703 = ( ~n25745 & n26354 ) | ( ~n25745 & n28702 ) | ( n26354 & n28702 ) ;
  assign n28704 = n28703 ^ n3679 ^ 1'b0 ;
  assign n28706 = ( n6276 & ~n24479 ) | ( n6276 & n28577 ) | ( ~n24479 & n28577 ) ;
  assign n28705 = n8345 & n13006 ;
  assign n28707 = n28706 ^ n28705 ^ 1'b0 ;
  assign n28708 = ~n19730 & n28707 ;
  assign n28709 = n18166 ^ n13623 ^ n9593 ;
  assign n28710 = n28709 ^ n20289 ^ n2636 ;
  assign n28711 = ( n5102 & n22324 ) | ( n5102 & ~n24152 ) | ( n22324 & ~n24152 ) ;
  assign n28712 = n10786 ^ n6712 ^ n6044 ;
  assign n28713 = ( n3524 & n20015 ) | ( n3524 & ~n28712 ) | ( n20015 & ~n28712 ) ;
  assign n28714 = ( n2136 & ~n2629 ) | ( n2136 & n3123 ) | ( ~n2629 & n3123 ) ;
  assign n28715 = ( n530 & n3047 ) | ( n530 & n28714 ) | ( n3047 & n28714 ) ;
  assign n28716 = n18797 ^ n14043 ^ 1'b0 ;
  assign n28717 = ~n9046 & n28716 ;
  assign n28718 = n28717 ^ n857 ^ 1'b0 ;
  assign n28719 = n21652 ^ n5786 ^ 1'b0 ;
  assign n28720 = n2593 & ~n28719 ;
  assign n28721 = ( n3528 & n10428 ) | ( n3528 & ~n28720 ) | ( n10428 & ~n28720 ) ;
  assign n28722 = n28721 ^ n15973 ^ 1'b0 ;
  assign n28723 = n16419 | n28722 ;
  assign n28724 = n9492 & ~n12840 ;
  assign n28725 = ( ~n16245 & n20499 ) | ( ~n16245 & n28724 ) | ( n20499 & n28724 ) ;
  assign n28726 = ( n2023 & ~n5325 ) | ( n2023 & n7455 ) | ( ~n5325 & n7455 ) ;
  assign n28727 = ( n4866 & ~n7709 ) | ( n4866 & n28726 ) | ( ~n7709 & n28726 ) ;
  assign n28728 = n6336 | n28727 ;
  assign n28729 = n12464 & ~n28728 ;
  assign n28730 = n28729 ^ n16919 ^ n14129 ;
  assign n28731 = ( n2525 & n14488 ) | ( n2525 & ~n28730 ) | ( n14488 & ~n28730 ) ;
  assign n28732 = n28731 ^ n15908 ^ n12300 ;
  assign n28733 = n3631 & ~n6852 ;
  assign n28734 = n28733 ^ n13098 ^ 1'b0 ;
  assign n28735 = n28734 ^ n7461 ^ 1'b0 ;
  assign n28736 = n13180 | n28735 ;
  assign n28737 = n14605 | n28736 ;
  assign n28738 = n28737 ^ n20285 ^ n3116 ;
  assign n28739 = n10452 ^ n5237 ^ x57 ;
  assign n28740 = n28739 ^ n12004 ^ n9604 ;
  assign n28741 = ( n793 & n2861 ) | ( n793 & n13977 ) | ( n2861 & n13977 ) ;
  assign n28742 = n9639 ^ n3917 ^ n3407 ;
  assign n28743 = n9893 & n28742 ;
  assign n28744 = n28743 ^ n4516 ^ n531 ;
  assign n28745 = n28744 ^ n22873 ^ 1'b0 ;
  assign n28746 = n27553 ^ n23924 ^ n7128 ;
  assign n28747 = n10829 | n28746 ;
  assign n28748 = n18635 & n19300 ;
  assign n28749 = n28748 ^ n11536 ^ 1'b0 ;
  assign n28750 = n12356 & ~n17674 ;
  assign n28751 = n6137 ^ n3163 ^ 1'b0 ;
  assign n28752 = ( ~n6983 & n11180 ) | ( ~n6983 & n28751 ) | ( n11180 & n28751 ) ;
  assign n28753 = ( n2396 & ~n13381 ) | ( n2396 & n28752 ) | ( ~n13381 & n28752 ) ;
  assign n28754 = ~n720 & n12239 ;
  assign n28755 = n28754 ^ n28652 ^ n18317 ;
  assign n28756 = n12303 ^ n9790 ^ 1'b0 ;
  assign n28757 = x16 & n28756 ;
  assign n28758 = ( n16813 & n28755 ) | ( n16813 & n28757 ) | ( n28755 & n28757 ) ;
  assign n28759 = n24832 ^ n7965 ^ n4249 ;
  assign n28760 = ( n9776 & ~n13173 ) | ( n9776 & n18437 ) | ( ~n13173 & n18437 ) ;
  assign n28761 = n19050 ^ n14458 ^ n12468 ;
  assign n28762 = ( ~n6204 & n7963 ) | ( ~n6204 & n28761 ) | ( n7963 & n28761 ) ;
  assign n28763 = n22907 ^ n12345 ^ 1'b0 ;
  assign n28764 = n28762 & n28763 ;
  assign n28765 = ( n5901 & ~n28760 ) | ( n5901 & n28764 ) | ( ~n28760 & n28764 ) ;
  assign n28766 = ( n2073 & n15541 ) | ( n2073 & n19174 ) | ( n15541 & n19174 ) ;
  assign n28767 = n28766 ^ n7033 ^ n3672 ;
  assign n28768 = n11611 ^ n2103 ^ 1'b0 ;
  assign n28769 = n1487 & n28768 ;
  assign n28770 = n28769 ^ n1186 ^ 1'b0 ;
  assign n28771 = ( n5650 & ~n5783 ) | ( n5650 & n5853 ) | ( ~n5783 & n5853 ) ;
  assign n28772 = n28771 ^ n7260 ^ n1958 ;
  assign n28773 = ( n6179 & n28770 ) | ( n6179 & n28772 ) | ( n28770 & n28772 ) ;
  assign n28774 = n8097 & ~n20483 ;
  assign n28777 = n15117 ^ n8547 ^ n5123 ;
  assign n28775 = ( n7554 & ~n27656 ) | ( n7554 & n27892 ) | ( ~n27656 & n27892 ) ;
  assign n28776 = n28775 ^ n27910 ^ 1'b0 ;
  assign n28778 = n28777 ^ n28776 ^ 1'b0 ;
  assign n28782 = n18805 ^ n2369 ^ n1370 ;
  assign n28780 = ( n5452 & ~n7088 ) | ( n5452 & n15849 ) | ( ~n7088 & n15849 ) ;
  assign n28779 = ~n2307 & n28734 ;
  assign n28781 = n28780 ^ n28779 ^ 1'b0 ;
  assign n28783 = n28782 ^ n28781 ^ x141 ;
  assign n28784 = n14619 ^ n8402 ^ n7605 ;
  assign n28785 = n28784 ^ n16867 ^ 1'b0 ;
  assign n28786 = n28785 ^ n26361 ^ n7172 ;
  assign n28787 = n12793 ^ n5090 ^ 1'b0 ;
  assign n28788 = n16580 ^ n15394 ^ 1'b0 ;
  assign n28789 = n28788 ^ n12594 ^ 1'b0 ;
  assign n28790 = n9559 | n28789 ;
  assign n28791 = n14075 ^ n6203 ^ 1'b0 ;
  assign n28792 = n17948 & ~n28791 ;
  assign n28793 = ( n23415 & n28790 ) | ( n23415 & ~n28792 ) | ( n28790 & ~n28792 ) ;
  assign n28794 = ( ~n6777 & n18621 ) | ( ~n6777 & n27655 ) | ( n18621 & n27655 ) ;
  assign n28795 = ~n13175 & n28794 ;
  assign n28796 = n28334 ^ n4647 ^ 1'b0 ;
  assign n28797 = n17112 | n23136 ;
  assign n28798 = n28797 ^ n5613 ^ 1'b0 ;
  assign n28799 = n28798 ^ n27214 ^ n24136 ;
  assign n28800 = n28799 ^ n17969 ^ 1'b0 ;
  assign n28801 = n926 & n28800 ;
  assign n28802 = n16287 ^ n15446 ^ n3196 ;
  assign n28803 = n28507 ^ n22602 ^ n7222 ;
  assign n28804 = n5674 ^ n666 ^ n288 ;
  assign n28805 = n28804 ^ n3844 ^ n2003 ;
  assign n28806 = n11500 ^ n4743 ^ 1'b0 ;
  assign n28807 = ~n28805 & n28806 ;
  assign n28808 = ( n1856 & n16008 ) | ( n1856 & ~n28807 ) | ( n16008 & ~n28807 ) ;
  assign n28809 = n28808 ^ n23478 ^ 1'b0 ;
  assign n28810 = n28520 ^ n25664 ^ n277 ;
  assign n28811 = n28810 ^ n20691 ^ n12320 ;
  assign n28812 = n15260 & n20169 ;
  assign n28813 = ( ~n25793 & n28679 ) | ( ~n25793 & n28812 ) | ( n28679 & n28812 ) ;
  assign n28814 = n4934 & ~n6086 ;
  assign n28815 = n28814 ^ n18066 ^ 1'b0 ;
  assign n28816 = ( n2491 & n4087 ) | ( n2491 & n8618 ) | ( n4087 & n8618 ) ;
  assign n28817 = n4688 ^ n4608 ^ x132 ;
  assign n28818 = ( x118 & n14888 ) | ( x118 & n24558 ) | ( n14888 & n24558 ) ;
  assign n28819 = n28818 ^ n9274 ^ 1'b0 ;
  assign n28820 = n18727 ^ n17734 ^ n3111 ;
  assign n28821 = n28820 ^ n23230 ^ n21384 ;
  assign n28822 = n26125 ^ n23073 ^ n18710 ;
  assign n28823 = n22734 ^ n3793 ^ 1'b0 ;
  assign n28824 = n4088 & ~n28823 ;
  assign n28825 = n2392 & ~n14722 ;
  assign n28826 = ~n5076 & n28825 ;
  assign n28827 = n11306 ^ n4989 ^ n2174 ;
  assign n28828 = n923 & n28827 ;
  assign n28829 = n28828 ^ n24770 ^ n9510 ;
  assign n28830 = n24371 ^ n14782 ^ n8455 ;
  assign n28831 = n7454 ^ n7086 ^ n2510 ;
  assign n28832 = n1481 & n28831 ;
  assign n28833 = n28832 ^ n10842 ^ 1'b0 ;
  assign n28834 = ( ~n28829 & n28830 ) | ( ~n28829 & n28833 ) | ( n28830 & n28833 ) ;
  assign n28835 = ( n6039 & n12358 ) | ( n6039 & n19310 ) | ( n12358 & n19310 ) ;
  assign n28836 = n28835 ^ n17743 ^ 1'b0 ;
  assign n28837 = n28836 ^ n19560 ^ n11521 ;
  assign n28838 = ( ~n9648 & n10925 ) | ( ~n9648 & n13679 ) | ( n10925 & n13679 ) ;
  assign n28839 = n743 & n11597 ;
  assign n28840 = n28839 ^ n4253 ^ 1'b0 ;
  assign n28841 = n13301 ^ n3002 ^ 1'b0 ;
  assign n28842 = ~n28840 & n28841 ;
  assign n28844 = n15208 ^ n12178 ^ n10981 ;
  assign n28843 = ( ~n20401 & n24460 ) | ( ~n20401 & n24756 ) | ( n24460 & n24756 ) ;
  assign n28845 = n28844 ^ n28843 ^ n1353 ;
  assign n28846 = ( n6968 & ~n27522 ) | ( n6968 & n28845 ) | ( ~n27522 & n28845 ) ;
  assign n28847 = ( n7269 & n10952 ) | ( n7269 & n11071 ) | ( n10952 & n11071 ) ;
  assign n28848 = n28847 ^ n15241 ^ n7688 ;
  assign n28849 = n5346 | n23656 ;
  assign n28850 = n28849 ^ n25064 ^ 1'b0 ;
  assign n28851 = ( n12566 & n28848 ) | ( n12566 & ~n28850 ) | ( n28848 & ~n28850 ) ;
  assign n28858 = n10187 ^ n3981 ^ 1'b0 ;
  assign n28854 = n12845 ^ n3926 ^ 1'b0 ;
  assign n28855 = ~n6898 & n28854 ;
  assign n28853 = n20332 ^ n19929 ^ n7378 ;
  assign n28852 = n23361 ^ n18785 ^ n12479 ;
  assign n28856 = n28855 ^ n28853 ^ n28852 ;
  assign n28857 = n28856 ^ n18931 ^ n8117 ;
  assign n28859 = n28858 ^ n28857 ^ n8487 ;
  assign n28860 = n7406 & n10145 ;
  assign n28861 = ~n12235 & n28860 ;
  assign n28862 = n22570 & ~n28861 ;
  assign n28863 = ( x68 & ~n823 ) | ( x68 & n1242 ) | ( ~n823 & n1242 ) ;
  assign n28864 = ~n3865 & n6317 ;
  assign n28865 = n10017 & n28864 ;
  assign n28866 = n26402 ^ n24969 ^ n10253 ;
  assign n28867 = ( n28863 & n28865 ) | ( n28863 & n28866 ) | ( n28865 & n28866 ) ;
  assign n28870 = ( n12059 & ~n16267 ) | ( n12059 & n16542 ) | ( ~n16267 & n16542 ) ;
  assign n28871 = n28870 ^ n24896 ^ n2950 ;
  assign n28868 = ( ~n528 & n2528 ) | ( ~n528 & n7863 ) | ( n2528 & n7863 ) ;
  assign n28869 = n5257 | n28868 ;
  assign n28872 = n28871 ^ n28869 ^ 1'b0 ;
  assign n28873 = n28872 ^ n18256 ^ x213 ;
  assign n28874 = n4352 & n28873 ;
  assign n28875 = ~n8932 & n28874 ;
  assign n28876 = n22633 | n28528 ;
  assign n28877 = ( n7625 & ~n13424 ) | ( n7625 & n14538 ) | ( ~n13424 & n14538 ) ;
  assign n28878 = n3991 | n9676 ;
  assign n28879 = n10778 | n28878 ;
  assign n28880 = ( n9310 & ~n28877 ) | ( n9310 & n28879 ) | ( ~n28877 & n28879 ) ;
  assign n28881 = ( n4894 & n12097 ) | ( n4894 & n28880 ) | ( n12097 & n28880 ) ;
  assign n28882 = ( n19677 & n28876 ) | ( n19677 & ~n28881 ) | ( n28876 & ~n28881 ) ;
  assign n28885 = n2302 & n17619 ;
  assign n28883 = n21063 ^ n15548 ^ n13184 ;
  assign n28884 = ( n9512 & n22170 ) | ( n9512 & n28883 ) | ( n22170 & n28883 ) ;
  assign n28886 = n28885 ^ n28884 ^ n2585 ;
  assign n28887 = n7692 & n11147 ;
  assign n28888 = n28798 ^ n18155 ^ n1666 ;
  assign n28889 = ~n4813 & n28888 ;
  assign n28890 = n14167 & ~n16209 ;
  assign n28891 = ( n9076 & n23143 ) | ( n9076 & ~n25782 ) | ( n23143 & ~n25782 ) ;
  assign n28892 = n28625 ^ n7177 ^ n3350 ;
  assign n28893 = ( n28890 & ~n28891 ) | ( n28890 & n28892 ) | ( ~n28891 & n28892 ) ;
  assign n28894 = n28893 ^ n28027 ^ n23104 ;
  assign n28895 = n10894 ^ n3296 ^ 1'b0 ;
  assign n28896 = ~n4910 & n28895 ;
  assign n28897 = n28896 ^ n19033 ^ 1'b0 ;
  assign n28900 = n27510 ^ n6875 ^ n3486 ;
  assign n28898 = n24566 ^ n19302 ^ n3195 ;
  assign n28899 = n28898 ^ n25215 ^ n3286 ;
  assign n28901 = n28900 ^ n28899 ^ n2734 ;
  assign n28902 = n24604 ^ n17313 ^ n6641 ;
  assign n28903 = n15594 & ~n28902 ;
  assign n28904 = ( n1706 & ~n13583 ) | ( n1706 & n28903 ) | ( ~n13583 & n28903 ) ;
  assign n28905 = n21983 ^ n17014 ^ n8473 ;
  assign n28906 = n26971 ^ n18953 ^ n305 ;
  assign n28907 = ( n6036 & ~n28905 ) | ( n6036 & n28906 ) | ( ~n28905 & n28906 ) ;
  assign n28908 = n25026 ^ n12709 ^ n4452 ;
  assign n28909 = n28908 ^ n24597 ^ n11433 ;
  assign n28914 = n1957 | n6839 ;
  assign n28915 = n7013 & ~n28914 ;
  assign n28916 = n15092 & ~n28915 ;
  assign n28917 = ~n9128 & n28916 ;
  assign n28918 = ( n12857 & n24093 ) | ( n12857 & ~n28917 ) | ( n24093 & ~n28917 ) ;
  assign n28910 = n12312 ^ n4947 ^ n451 ;
  assign n28911 = ~n965 & n28910 ;
  assign n28912 = n10749 & n28911 ;
  assign n28913 = n16958 & ~n28912 ;
  assign n28919 = n28918 ^ n28913 ^ 1'b0 ;
  assign n28920 = ( n5413 & n11945 ) | ( n5413 & ~n13236 ) | ( n11945 & ~n13236 ) ;
  assign n28921 = n28920 ^ n8168 ^ 1'b0 ;
  assign n28922 = n17048 & n28921 ;
  assign n28923 = n28922 ^ n10959 ^ n1914 ;
  assign n28924 = ~n17774 & n28923 ;
  assign n28925 = ( ~n16526 & n17975 ) | ( ~n16526 & n24420 ) | ( n17975 & n24420 ) ;
  assign n28926 = n28865 ^ n12247 ^ n7024 ;
  assign n28927 = n28851 ^ n6164 ^ 1'b0 ;
  assign n28928 = ( n13658 & n18001 ) | ( n13658 & n19979 ) | ( n18001 & n19979 ) ;
  assign n28931 = n14240 ^ n9276 ^ n5131 ;
  assign n28929 = ( n10485 & n13322 ) | ( n10485 & ~n22569 ) | ( n13322 & ~n22569 ) ;
  assign n28930 = ( x26 & n14261 ) | ( x26 & ~n28929 ) | ( n14261 & ~n28929 ) ;
  assign n28932 = n28931 ^ n28930 ^ n1116 ;
  assign n28933 = ( ~n13171 & n25830 ) | ( ~n13171 & n28932 ) | ( n25830 & n28932 ) ;
  assign n28934 = ( n6346 & ~n16926 ) | ( n6346 & n19677 ) | ( ~n16926 & n19677 ) ;
  assign n28935 = n2256 ^ n1564 ^ 1'b0 ;
  assign n28936 = ( ~n3372 & n28934 ) | ( ~n3372 & n28935 ) | ( n28934 & n28935 ) ;
  assign n28937 = n26965 & n27014 ;
  assign n28938 = ( n11062 & n11513 ) | ( n11062 & ~n12384 ) | ( n11513 & ~n12384 ) ;
  assign n28939 = n9000 & ~n28938 ;
  assign n28940 = n6177 & n28939 ;
  assign n28941 = n22938 ^ n13746 ^ n7183 ;
  assign n28942 = ( n2094 & n15484 ) | ( n2094 & n16348 ) | ( n15484 & n16348 ) ;
  assign n28944 = n12489 & ~n14238 ;
  assign n28943 = ( n10123 & n12141 ) | ( n10123 & ~n21348 ) | ( n12141 & ~n21348 ) ;
  assign n28945 = n28944 ^ n28943 ^ 1'b0 ;
  assign n28946 = ~n28942 & n28945 ;
  assign n28947 = ( n11014 & n16523 ) | ( n11014 & ~n28946 ) | ( n16523 & ~n28946 ) ;
  assign n28948 = n16988 ^ n6118 ^ 1'b0 ;
  assign n28949 = ~n7464 & n28948 ;
  assign n28950 = n28949 ^ n22981 ^ n21399 ;
  assign n28951 = n5212 ^ n1695 ^ n463 ;
  assign n28952 = ( n9995 & n28293 ) | ( n9995 & ~n28951 ) | ( n28293 & ~n28951 ) ;
  assign n28953 = n6813 & ~n28952 ;
  assign n28954 = n28953 ^ n17926 ^ 1'b0 ;
  assign n28955 = n6109 ^ n3263 ^ 1'b0 ;
  assign n28956 = ~n10428 & n28955 ;
  assign n28957 = ( ~n18481 & n20176 ) | ( ~n18481 & n28956 ) | ( n20176 & n28956 ) ;
  assign n28958 = n13290 ^ n12017 ^ n11267 ;
  assign n28959 = n12608 ^ n11671 ^ n3148 ;
  assign n28960 = n28959 ^ n6785 ^ n1834 ;
  assign n28961 = n28960 ^ n15115 ^ n4145 ;
  assign n28962 = n7561 | n21628 ;
  assign n28963 = n28962 ^ n13251 ^ 1'b0 ;
  assign n28964 = ( ~n10130 & n28961 ) | ( ~n10130 & n28963 ) | ( n28961 & n28963 ) ;
  assign n28965 = ( ~n17857 & n28958 ) | ( ~n17857 & n28964 ) | ( n28958 & n28964 ) ;
  assign n28966 = n26965 ^ n25579 ^ n21783 ;
  assign n28969 = n1778 | n15398 ;
  assign n28970 = n28969 ^ n3292 ^ 1'b0 ;
  assign n28967 = n14061 & n17449 ;
  assign n28968 = n24739 & n28967 ;
  assign n28971 = n28970 ^ n28968 ^ n12344 ;
  assign n28972 = n6676 | n15422 ;
  assign n28974 = n10099 ^ n8778 ^ 1'b0 ;
  assign n28975 = ~n14968 & n28974 ;
  assign n28976 = n27843 & n28975 ;
  assign n28973 = n11919 ^ n11588 ^ n9698 ;
  assign n28977 = n28976 ^ n28973 ^ n17864 ;
  assign n28978 = n28178 ^ n18475 ^ n6124 ;
  assign n28979 = n28978 ^ n4391 ^ 1'b0 ;
  assign n28983 = ( x107 & ~n2030 ) | ( x107 & n18079 ) | ( ~n2030 & n18079 ) ;
  assign n28984 = n28983 ^ n24344 ^ n9424 ;
  assign n28980 = n10407 ^ n4685 ^ n2739 ;
  assign n28981 = ( ~n954 & n5007 ) | ( ~n954 & n25968 ) | ( n5007 & n25968 ) ;
  assign n28982 = n28980 & n28981 ;
  assign n28985 = n28984 ^ n28982 ^ n9108 ;
  assign n28986 = ( n10295 & n28106 ) | ( n10295 & n28985 ) | ( n28106 & n28985 ) ;
  assign n28987 = n3163 & n17969 ;
  assign n28988 = ~n5462 & n28987 ;
  assign n28989 = ~n6353 & n24352 ;
  assign n28990 = n8455 & n28989 ;
  assign n28991 = n28990 ^ n9114 ^ 1'b0 ;
  assign n28992 = ~n11501 & n28991 ;
  assign n28993 = ( n5512 & ~n12662 ) | ( n5512 & n22466 ) | ( ~n12662 & n22466 ) ;
  assign n28994 = n5331 & n28993 ;
  assign n28995 = ~n28992 & n28994 ;
  assign n28996 = n8183 ^ n3915 ^ 1'b0 ;
  assign n28997 = ( ~n2672 & n4676 ) | ( ~n2672 & n18064 ) | ( n4676 & n18064 ) ;
  assign n28998 = n18841 | n28997 ;
  assign n28999 = n28996 | n28998 ;
  assign n29000 = n28999 ^ n25456 ^ 1'b0 ;
  assign n29001 = n2323 & ~n14319 ;
  assign n29002 = n29001 ^ n17123 ^ 1'b0 ;
  assign n29003 = ( n7545 & n15489 ) | ( n7545 & n29002 ) | ( n15489 & n29002 ) ;
  assign n29007 = n4579 & ~n22764 ;
  assign n29008 = n20959 & n29007 ;
  assign n29006 = ( n3366 & ~n7534 ) | ( n3366 & n14779 ) | ( ~n7534 & n14779 ) ;
  assign n29004 = n9209 ^ n8203 ^ n7092 ;
  assign n29005 = ( ~n3562 & n17566 ) | ( ~n3562 & n29004 ) | ( n17566 & n29004 ) ;
  assign n29009 = n29008 ^ n29006 ^ n29005 ;
  assign n29010 = n8199 | n8716 ;
  assign n29011 = n29010 ^ n13592 ^ 1'b0 ;
  assign n29012 = ( n16836 & n16905 ) | ( n16836 & ~n28134 ) | ( n16905 & ~n28134 ) ;
  assign n29013 = ( n24396 & n29011 ) | ( n24396 & ~n29012 ) | ( n29011 & ~n29012 ) ;
  assign n29014 = n24421 ^ n15144 ^ n13563 ;
  assign n29015 = n29014 ^ n1734 ^ x155 ;
  assign n29016 = n6325 ^ n478 ^ 1'b0 ;
  assign n29017 = ~n14021 & n29016 ;
  assign n29018 = n14702 ^ n10996 ^ n2219 ;
  assign n29019 = n23246 ^ n13053 ^ n9575 ;
  assign n29020 = n14735 & ~n26312 ;
  assign n29021 = n24117 & n29020 ;
  assign n29022 = ( n7388 & n16823 ) | ( n7388 & ~n17932 ) | ( n16823 & ~n17932 ) ;
  assign n29023 = n6624 ^ n2506 ^ 1'b0 ;
  assign n29024 = n16923 ^ n2527 ^ 1'b0 ;
  assign n29025 = n29023 | n29024 ;
  assign n29026 = ( n19582 & n29022 ) | ( n19582 & ~n29025 ) | ( n29022 & ~n29025 ) ;
  assign n29027 = ~n25924 & n26971 ;
  assign n29028 = n2992 & n18036 ;
  assign n29029 = n29027 & n29028 ;
  assign n29030 = ( ~n2569 & n8932 ) | ( ~n2569 & n16534 ) | ( n8932 & n16534 ) ;
  assign n29031 = n29030 ^ n20758 ^ n9492 ;
  assign n29032 = n29031 ^ n6792 ^ n5650 ;
  assign n29033 = ( n15198 & ~n15882 ) | ( n15198 & n29032 ) | ( ~n15882 & n29032 ) ;
  assign n29034 = ( ~n13001 & n16089 ) | ( ~n13001 & n29033 ) | ( n16089 & n29033 ) ;
  assign n29035 = n10194 ^ n2729 ^ n2548 ;
  assign n29036 = n29035 ^ n18277 ^ n17138 ;
  assign n29037 = ( n879 & n4783 ) | ( n879 & ~n29036 ) | ( n4783 & ~n29036 ) ;
  assign n29038 = n12250 ^ n2780 ^ n1084 ;
  assign n29039 = ( n7673 & n16518 ) | ( n7673 & n29038 ) | ( n16518 & n29038 ) ;
  assign n29040 = n9401 & ~n15293 ;
  assign n29041 = n3603 & n29040 ;
  assign n29042 = n11898 ^ n11877 ^ n9664 ;
  assign n29043 = ( n8344 & ~n15857 ) | ( n8344 & n29042 ) | ( ~n15857 & n29042 ) ;
  assign n29045 = n11098 ^ n2246 ^ n1023 ;
  assign n29046 = ( n425 & ~n5557 ) | ( n425 & n29045 ) | ( ~n5557 & n29045 ) ;
  assign n29044 = n11679 ^ n2909 ^ 1'b0 ;
  assign n29047 = n29046 ^ n29044 ^ n19549 ;
  assign n29048 = n6274 ^ n5541 ^ n1195 ;
  assign n29049 = n19933 ^ n12943 ^ 1'b0 ;
  assign n29050 = n6674 & n29049 ;
  assign n29051 = n11105 & n29050 ;
  assign n29052 = ( ~n979 & n12880 ) | ( ~n979 & n29051 ) | ( n12880 & n29051 ) ;
  assign n29053 = ( ~n11946 & n29048 ) | ( ~n11946 & n29052 ) | ( n29048 & n29052 ) ;
  assign n29054 = n4525 & ~n19105 ;
  assign n29055 = n546 & n29054 ;
  assign n29056 = ( n2193 & n5872 ) | ( n2193 & n29055 ) | ( n5872 & n29055 ) ;
  assign n29057 = n9852 ^ n1048 ^ n683 ;
  assign n29058 = ( n13982 & n28325 ) | ( n13982 & n29057 ) | ( n28325 & n29057 ) ;
  assign n29059 = n29058 ^ n22112 ^ n19953 ;
  assign n29060 = n29059 ^ n5769 ^ n555 ;
  assign n29061 = ( n2591 & ~n16126 ) | ( n2591 & n29060 ) | ( ~n16126 & n29060 ) ;
  assign n29067 = n2832 ^ n1376 ^ n937 ;
  assign n29068 = ( n1236 & ~n19313 ) | ( n1236 & n29067 ) | ( ~n19313 & n29067 ) ;
  assign n29069 = ( ~n6148 & n18062 ) | ( ~n6148 & n29068 ) | ( n18062 & n29068 ) ;
  assign n29070 = n9564 ^ n6128 ^ n1819 ;
  assign n29071 = ( n9104 & n12146 ) | ( n9104 & ~n29070 ) | ( n12146 & ~n29070 ) ;
  assign n29072 = n29071 ^ n7269 ^ n5848 ;
  assign n29073 = ( n19060 & n29069 ) | ( n19060 & n29072 ) | ( n29069 & n29072 ) ;
  assign n29062 = n19296 ^ n4407 ^ n929 ;
  assign n29063 = n29062 ^ n19790 ^ 1'b0 ;
  assign n29064 = n12050 & n29063 ;
  assign n29065 = n29064 ^ n19769 ^ n6160 ;
  assign n29066 = n15197 & n29065 ;
  assign n29074 = n29073 ^ n29066 ^ n26877 ;
  assign n29075 = n10044 & ~n15577 ;
  assign n29076 = ~n1485 & n29075 ;
  assign n29077 = n8014 ^ n3944 ^ n621 ;
  assign n29078 = ( n1837 & ~n6238 ) | ( n1837 & n29077 ) | ( ~n6238 & n29077 ) ;
  assign n29079 = ( n9615 & n19184 ) | ( n9615 & n21967 ) | ( n19184 & n21967 ) ;
  assign n29080 = n29079 ^ n27032 ^ n8890 ;
  assign n29081 = ( n8643 & n29078 ) | ( n8643 & n29080 ) | ( n29078 & n29080 ) ;
  assign n29084 = n15868 ^ n2786 ^ n2253 ;
  assign n29085 = ( n2032 & n4287 ) | ( n2032 & ~n29084 ) | ( n4287 & ~n29084 ) ;
  assign n29083 = n3556 | n21510 ;
  assign n29082 = n17371 ^ n15795 ^ n7289 ;
  assign n29086 = n29085 ^ n29083 ^ n29082 ;
  assign n29087 = n7215 ^ n4097 ^ n548 ;
  assign n29088 = ( n26478 & n28790 ) | ( n26478 & n29087 ) | ( n28790 & n29087 ) ;
  assign n29089 = ( n4000 & n9059 ) | ( n4000 & ~n29088 ) | ( n9059 & ~n29088 ) ;
  assign n29090 = n29089 ^ n20364 ^ n18864 ;
  assign n29091 = ( ~n6406 & n18678 ) | ( ~n6406 & n29090 ) | ( n18678 & n29090 ) ;
  assign n29092 = ( n1445 & n2643 ) | ( n1445 & ~n14518 ) | ( n2643 & ~n14518 ) ;
  assign n29093 = ( x142 & n12074 ) | ( x142 & ~n15893 ) | ( n12074 & ~n15893 ) ;
  assign n29094 = n29093 ^ n3724 ^ n3183 ;
  assign n29095 = ( ~n5582 & n7783 ) | ( ~n5582 & n29094 ) | ( n7783 & n29094 ) ;
  assign n29096 = n24502 ^ n19912 ^ n6502 ;
  assign n29097 = ( n5435 & n6405 ) | ( n5435 & ~n6658 ) | ( n6405 & ~n6658 ) ;
  assign n29098 = n29097 ^ n27285 ^ n870 ;
  assign n29108 = n11345 ^ n1994 ^ 1'b0 ;
  assign n29104 = n28146 ^ n7942 ^ 1'b0 ;
  assign n29105 = n671 | n29104 ;
  assign n29106 = ( n12673 & n18735 ) | ( n12673 & ~n28427 ) | ( n18735 & ~n28427 ) ;
  assign n29107 = ( n14689 & n29105 ) | ( n14689 & n29106 ) | ( n29105 & n29106 ) ;
  assign n29099 = n13929 ^ n4289 ^ n2720 ;
  assign n29100 = n469 & ~n29099 ;
  assign n29101 = n29100 ^ n5670 ^ 1'b0 ;
  assign n29102 = n18806 | n29101 ;
  assign n29103 = n25650 | n29102 ;
  assign n29109 = n29108 ^ n29107 ^ n29103 ;
  assign n29110 = n6139 & n27431 ;
  assign n29111 = n12722 & n29110 ;
  assign n29112 = n6295 | n29111 ;
  assign n29113 = ( n13989 & n14031 ) | ( n13989 & n18403 ) | ( n14031 & n18403 ) ;
  assign n29118 = ( n10185 & ~n18873 ) | ( n10185 & n22830 ) | ( ~n18873 & n22830 ) ;
  assign n29114 = n4920 & n21965 ;
  assign n29115 = n29114 ^ n590 ^ 1'b0 ;
  assign n29116 = ( ~n1763 & n2676 ) | ( ~n1763 & n29115 ) | ( n2676 & n29115 ) ;
  assign n29117 = n29116 ^ n2928 ^ n1380 ;
  assign n29119 = n29118 ^ n29117 ^ 1'b0 ;
  assign n29120 = n14529 & ~n29119 ;
  assign n29121 = n21979 ^ n13881 ^ n8190 ;
  assign n29122 = ( ~n2960 & n8787 ) | ( ~n2960 & n15042 ) | ( n8787 & n15042 ) ;
  assign n29123 = n29122 ^ x111 ^ 1'b0 ;
  assign n29124 = ( n3477 & n29121 ) | ( n3477 & n29123 ) | ( n29121 & n29123 ) ;
  assign n29125 = ~n11695 & n21861 ;
  assign n29126 = n7721 & n29125 ;
  assign n29127 = n29126 ^ n12785 ^ 1'b0 ;
  assign n29128 = n19602 | n29127 ;
  assign n29129 = n29128 ^ n7272 ^ 1'b0 ;
  assign n29130 = n23002 & n29129 ;
  assign n29131 = n29130 ^ n13431 ^ n11554 ;
  assign n29132 = n6116 & n18073 ;
  assign n29133 = ~n5050 & n29132 ;
  assign n29134 = n29133 ^ n6876 ^ n797 ;
  assign n29135 = x22 & ~n9614 ;
  assign n29136 = ~n2033 & n29135 ;
  assign n29137 = n1191 & ~n4591 ;
  assign n29138 = n29137 ^ n4145 ^ 1'b0 ;
  assign n29139 = ( n12678 & n29136 ) | ( n12678 & ~n29138 ) | ( n29136 & ~n29138 ) ;
  assign n29140 = n16411 ^ n9152 ^ n430 ;
  assign n29141 = n16486 ^ x231 ^ 1'b0 ;
  assign n29142 = n29140 & n29141 ;
  assign n29143 = n2688 & n29142 ;
  assign n29144 = n29143 ^ n28030 ^ 1'b0 ;
  assign n29145 = n18804 | n29144 ;
  assign n29146 = n14494 ^ n5696 ^ 1'b0 ;
  assign n29147 = n10310 | n29146 ;
  assign n29148 = ~n569 & n20810 ;
  assign n29149 = n29147 | n29148 ;
  assign n29150 = n19490 ^ n14482 ^ n12757 ;
  assign n29151 = n19088 ^ n4343 ^ 1'b0 ;
  assign n29152 = ( ~n623 & n15258 ) | ( ~n623 & n29151 ) | ( n15258 & n29151 ) ;
  assign n29153 = ( ~n9917 & n17573 ) | ( ~n9917 & n29152 ) | ( n17573 & n29152 ) ;
  assign n29154 = n29150 & n29153 ;
  assign n29156 = n16828 ^ n13476 ^ n3387 ;
  assign n29155 = n3340 & n25049 ;
  assign n29157 = n29156 ^ n29155 ^ 1'b0 ;
  assign n29158 = n29157 ^ n6661 ^ n1514 ;
  assign n29159 = n29154 & ~n29158 ;
  assign n29160 = n22902 ^ n16152 ^ 1'b0 ;
  assign n29161 = ~n2442 & n29160 ;
  assign n29162 = n24242 ^ n20274 ^ n6726 ;
  assign n29163 = n29162 ^ n12922 ^ n9131 ;
  assign n29164 = n25404 ^ n20117 ^ n4574 ;
  assign n29165 = n27657 ^ n24589 ^ n10514 ;
  assign n29166 = ( n283 & n708 ) | ( n283 & n8310 ) | ( n708 & n8310 ) ;
  assign n29167 = n29166 ^ n25864 ^ n14970 ;
  assign n29168 = n18396 & ~n29167 ;
  assign n29169 = n29168 ^ n20171 ^ n3920 ;
  assign n29170 = ~n7825 & n7873 ;
  assign n29171 = n29170 ^ n2216 ^ 1'b0 ;
  assign n29172 = n11572 & n12239 ;
  assign n29173 = ~n23541 & n29172 ;
  assign n29174 = n11772 & ~n23538 ;
  assign n29175 = n17516 & n29174 ;
  assign n29176 = n29175 ^ n14714 ^ 1'b0 ;
  assign n29177 = n11777 & n24004 ;
  assign n29178 = n29177 ^ n27521 ^ 1'b0 ;
  assign n29179 = ( n8394 & ~n15087 ) | ( n8394 & n29178 ) | ( ~n15087 & n29178 ) ;
  assign n29180 = n24433 ^ n20483 ^ 1'b0 ;
  assign n29181 = ( n3073 & ~n3105 ) | ( n3073 & n23250 ) | ( ~n3105 & n23250 ) ;
  assign n29182 = n29180 & ~n29181 ;
  assign n29183 = n16160 ^ n9798 ^ 1'b0 ;
  assign n29184 = n29183 ^ n27011 ^ n19432 ;
  assign n29185 = n6044 | n27016 ;
  assign n29186 = n25223 ^ n3035 ^ n2256 ;
  assign n29187 = ( n9763 & n17919 ) | ( n9763 & n19127 ) | ( n17919 & n19127 ) ;
  assign n29188 = ( ~n9347 & n15355 ) | ( ~n9347 & n25213 ) | ( n15355 & n25213 ) ;
  assign n29189 = n2039 | n23903 ;
  assign n29190 = n6537 | n29189 ;
  assign n29191 = ~n14551 & n29190 ;
  assign n29192 = n29191 ^ n19611 ^ n10453 ;
  assign n29193 = n21820 ^ n12021 ^ n11025 ;
  assign n29194 = ( n2877 & ~n8303 ) | ( n2877 & n29193 ) | ( ~n8303 & n29193 ) ;
  assign n29195 = n17682 ^ n2165 ^ 1'b0 ;
  assign n29196 = ( n9347 & ~n25836 ) | ( n9347 & n29195 ) | ( ~n25836 & n29195 ) ;
  assign n29197 = ( n585 & ~n5255 ) | ( n585 & n6737 ) | ( ~n5255 & n6737 ) ;
  assign n29198 = n29197 ^ n23783 ^ n13050 ;
  assign n29199 = ( n13150 & ~n26639 ) | ( n13150 & n29198 ) | ( ~n26639 & n29198 ) ;
  assign n29200 = ( n8163 & n10786 ) | ( n8163 & ~n13844 ) | ( n10786 & ~n13844 ) ;
  assign n29201 = n29200 ^ n21795 ^ n8115 ;
  assign n29202 = n3420 ^ n3407 ^ 1'b0 ;
  assign n29203 = n5927 & n29202 ;
  assign n29204 = ( n2384 & n15207 ) | ( n2384 & n29203 ) | ( n15207 & n29203 ) ;
  assign n29205 = ~n10507 & n29204 ;
  assign n29206 = ~n22984 & n29205 ;
  assign n29207 = n29206 ^ n24810 ^ n18911 ;
  assign n29208 = n8055 ^ n2014 ^ 1'b0 ;
  assign n29209 = n27943 & n29208 ;
  assign n29210 = ( n3949 & ~n8605 ) | ( n3949 & n29209 ) | ( ~n8605 & n29209 ) ;
  assign n29211 = n29210 ^ n24473 ^ n13847 ;
  assign n29212 = ( ~n4884 & n19035 ) | ( ~n4884 & n28910 ) | ( n19035 & n28910 ) ;
  assign n29213 = ( n2484 & n21570 ) | ( n2484 & n23626 ) | ( n21570 & n23626 ) ;
  assign n29214 = n29213 ^ n18752 ^ n10749 ;
  assign n29215 = ( n11256 & n22415 ) | ( n11256 & ~n29214 ) | ( n22415 & ~n29214 ) ;
  assign n29216 = n8336 & n19164 ;
  assign n29217 = n29216 ^ n8762 ^ 1'b0 ;
  assign n29218 = ~n1952 & n4568 ;
  assign n29219 = n29218 ^ n8638 ^ 1'b0 ;
  assign n29220 = n28655 ^ n4173 ^ n2319 ;
  assign n29221 = n11436 | n25314 ;
  assign n29222 = n26442 ^ n12332 ^ n2727 ;
  assign n29223 = n29222 ^ n14660 ^ n8668 ;
  assign n29224 = n22866 ^ n20585 ^ n2325 ;
  assign n29225 = ~n13250 & n29224 ;
  assign n29226 = n29225 ^ n8054 ^ 1'b0 ;
  assign n29227 = n18595 ^ n4061 ^ 1'b0 ;
  assign n29228 = n16967 ^ n16427 ^ 1'b0 ;
  assign n29229 = ( n2271 & ~n7083 ) | ( n2271 & n29228 ) | ( ~n7083 & n29228 ) ;
  assign n29230 = n4579 & n13886 ;
  assign n29231 = n14515 & n29230 ;
  assign n29232 = ( n2876 & ~n6435 ) | ( n2876 & n29231 ) | ( ~n6435 & n29231 ) ;
  assign n29233 = n19454 ^ n19386 ^ n10024 ;
  assign n29234 = ( n14794 & n15977 ) | ( n14794 & n29233 ) | ( n15977 & n29233 ) ;
  assign n29235 = n29234 ^ n28764 ^ 1'b0 ;
  assign n29236 = n29235 ^ n11484 ^ n5296 ;
  assign n29240 = ( ~n2527 & n2588 ) | ( ~n2527 & n16793 ) | ( n2588 & n16793 ) ;
  assign n29237 = n19757 ^ n19240 ^ n16320 ;
  assign n29238 = n27031 ^ n1888 ^ 1'b0 ;
  assign n29239 = n29237 | n29238 ;
  assign n29241 = n29240 ^ n29239 ^ n7602 ;
  assign n29248 = ( n11944 & n17905 ) | ( n11944 & n24377 ) | ( n17905 & n24377 ) ;
  assign n29245 = n21335 ^ n20586 ^ n954 ;
  assign n29246 = n29245 ^ n17668 ^ n6355 ;
  assign n29242 = n8229 & ~n9481 ;
  assign n29243 = n29242 ^ n3249 ^ 1'b0 ;
  assign n29244 = ( n2297 & ~n21829 ) | ( n2297 & n29243 ) | ( ~n21829 & n29243 ) ;
  assign n29247 = n29246 ^ n29244 ^ x234 ;
  assign n29249 = n29248 ^ n29247 ^ n22110 ;
  assign n29251 = n23766 ^ n939 ^ x97 ;
  assign n29250 = ( ~n10909 & n11561 ) | ( ~n10909 & n20498 ) | ( n11561 & n20498 ) ;
  assign n29252 = n29251 ^ n29250 ^ n14698 ;
  assign n29253 = n2666 | n24137 ;
  assign n29254 = n2925 | n29253 ;
  assign n29255 = n29254 ^ n7453 ^ n5140 ;
  assign n29256 = n4629 & ~n14185 ;
  assign n29257 = n29256 ^ n7046 ^ 1'b0 ;
  assign n29258 = n29257 ^ n15692 ^ n12931 ;
  assign n29259 = n18638 ^ n2385 ^ 1'b0 ;
  assign n29260 = n8412 | n29259 ;
  assign n29261 = ( n8767 & ~n29258 ) | ( n8767 & n29260 ) | ( ~n29258 & n29260 ) ;
  assign n29262 = ( n19922 & n29255 ) | ( n19922 & ~n29261 ) | ( n29255 & ~n29261 ) ;
  assign n29263 = ( n8603 & n17758 ) | ( n8603 & n27411 ) | ( n17758 & n27411 ) ;
  assign n29264 = ( n622 & n11845 ) | ( n622 & ~n16651 ) | ( n11845 & ~n16651 ) ;
  assign n29265 = n29264 ^ n11178 ^ n4585 ;
  assign n29266 = n18282 ^ n11453 ^ n3050 ;
  assign n29270 = n15533 ^ n12880 ^ 1'b0 ;
  assign n29267 = n5058 ^ n4764 ^ 1'b0 ;
  assign n29268 = n558 | n29267 ;
  assign n29269 = ( n1032 & n6313 ) | ( n1032 & ~n29268 ) | ( n6313 & ~n29268 ) ;
  assign n29271 = n29270 ^ n29269 ^ n5184 ;
  assign n29272 = n8334 ^ n5718 ^ 1'b0 ;
  assign n29273 = n29272 ^ n12444 ^ n7527 ;
  assign n29274 = n8914 & n10551 ;
  assign n29282 = n8690 ^ n3855 ^ n1093 ;
  assign n29276 = n3997 ^ n3453 ^ 1'b0 ;
  assign n29277 = n4989 & ~n29276 ;
  assign n29275 = n1036 | n14518 ;
  assign n29278 = n29277 ^ n29275 ^ 1'b0 ;
  assign n29279 = n29278 ^ n7897 ^ 1'b0 ;
  assign n29280 = ( n11573 & n15702 ) | ( n11573 & ~n29279 ) | ( n15702 & ~n29279 ) ;
  assign n29281 = ( ~n12624 & n19024 ) | ( ~n12624 & n29280 ) | ( n19024 & n29280 ) ;
  assign n29283 = n29282 ^ n29281 ^ n24091 ;
  assign n29284 = ( ~n1627 & n29274 ) | ( ~n1627 & n29283 ) | ( n29274 & n29283 ) ;
  assign n29285 = ( n1148 & n2959 ) | ( n1148 & n5090 ) | ( n2959 & n5090 ) ;
  assign n29286 = n29285 ^ n10660 ^ 1'b0 ;
  assign n29287 = ( n29273 & n29284 ) | ( n29273 & n29286 ) | ( n29284 & n29286 ) ;
  assign n29296 = n25003 ^ n5979 ^ n4285 ;
  assign n29297 = n29296 ^ n17576 ^ 1'b0 ;
  assign n29293 = n814 | n26051 ;
  assign n29294 = ~n21355 & n29293 ;
  assign n29288 = n12287 ^ n3191 ^ n3037 ;
  assign n29289 = ( ~n3823 & n8309 ) | ( ~n3823 & n8383 ) | ( n8309 & n8383 ) ;
  assign n29290 = n29289 ^ n6573 ^ n1453 ;
  assign n29291 = ( n14326 & ~n29288 ) | ( n14326 & n29290 ) | ( ~n29288 & n29290 ) ;
  assign n29292 = ~n19723 & n29291 ;
  assign n29295 = n29294 ^ n29292 ^ 1'b0 ;
  assign n29298 = n29297 ^ n29295 ^ n21814 ;
  assign n29302 = ( n8039 & n18509 ) | ( n8039 & n22317 ) | ( n18509 & n22317 ) ;
  assign n29299 = n23734 ^ n11062 ^ n2688 ;
  assign n29300 = ( n6842 & ~n20965 ) | ( n6842 & n29299 ) | ( ~n20965 & n29299 ) ;
  assign n29301 = n13831 & ~n29300 ;
  assign n29303 = n29302 ^ n29301 ^ 1'b0 ;
  assign n29304 = n29303 ^ n17274 ^ n12508 ;
  assign n29305 = n23374 ^ n12514 ^ n12358 ;
  assign n29306 = n29305 ^ n24806 ^ n292 ;
  assign n29307 = ( n1320 & n5153 ) | ( n1320 & n10885 ) | ( n5153 & n10885 ) ;
  assign n29308 = ~n14042 & n14153 ;
  assign n29309 = n11033 & n29308 ;
  assign n29310 = ( n2799 & n27092 ) | ( n2799 & ~n29309 ) | ( n27092 & ~n29309 ) ;
  assign n29311 = ~n13322 & n29310 ;
  assign n29312 = n29311 ^ x117 ^ 1'b0 ;
  assign n29313 = ( n10362 & n29307 ) | ( n10362 & n29312 ) | ( n29307 & n29312 ) ;
  assign n29314 = ( n1068 & n16492 ) | ( n1068 & n18472 ) | ( n16492 & n18472 ) ;
  assign n29315 = ( n7377 & n14135 ) | ( n7377 & ~n29314 ) | ( n14135 & ~n29314 ) ;
  assign n29316 = ( n4662 & n20741 ) | ( n4662 & n29315 ) | ( n20741 & n29315 ) ;
  assign n29317 = ( n29306 & ~n29313 ) | ( n29306 & n29316 ) | ( ~n29313 & n29316 ) ;
  assign n29318 = n4101 ^ n595 ^ 1'b0 ;
  assign n29319 = n4706 & n29318 ;
  assign n29320 = n25688 ^ n19460 ^ n17573 ;
  assign n29321 = ~n29319 & n29320 ;
  assign n29322 = n27374 ^ n2790 ^ n2527 ;
  assign n29323 = ( n19901 & ~n29321 ) | ( n19901 & n29322 ) | ( ~n29321 & n29322 ) ;
  assign n29324 = n6329 ^ n3969 ^ n2828 ;
  assign n29325 = ( ~n15697 & n15773 ) | ( ~n15697 & n29324 ) | ( n15773 & n29324 ) ;
  assign n29327 = n12671 ^ n10811 ^ n2100 ;
  assign n29326 = n9669 | n16960 ;
  assign n29328 = n29327 ^ n29326 ^ 1'b0 ;
  assign n29329 = n13503 & n29328 ;
  assign n29330 = n29329 ^ n5289 ^ 1'b0 ;
  assign n29332 = ~n746 & n4603 ;
  assign n29333 = n29332 ^ n13902 ^ n11812 ;
  assign n29334 = n29333 ^ n20533 ^ n17530 ;
  assign n29331 = n7479 & ~n14847 ;
  assign n29335 = n29334 ^ n29331 ^ 1'b0 ;
  assign n29336 = ( n370 & ~n532 ) | ( n370 & n827 ) | ( ~n532 & n827 ) ;
  assign n29337 = ( n2983 & n3582 ) | ( n2983 & n29336 ) | ( n3582 & n29336 ) ;
  assign n29338 = n29337 ^ n26526 ^ n845 ;
  assign n29339 = n7097 ^ n2524 ^ 1'b0 ;
  assign n29340 = ( n15391 & n17063 ) | ( n15391 & ~n22808 ) | ( n17063 & ~n22808 ) ;
  assign n29341 = n23987 ^ n7976 ^ n7837 ;
  assign n29342 = ( n29339 & ~n29340 ) | ( n29339 & n29341 ) | ( ~n29340 & n29341 ) ;
  assign n29344 = ( n1479 & n4533 ) | ( n1479 & n26521 ) | ( n4533 & n26521 ) ;
  assign n29343 = ( n7581 & n11083 ) | ( n7581 & ~n20945 ) | ( n11083 & ~n20945 ) ;
  assign n29345 = n29344 ^ n29343 ^ n25035 ;
  assign n29346 = n29345 ^ n22374 ^ n8994 ;
  assign n29347 = n9311 ^ n8971 ^ n2093 ;
  assign n29348 = n11446 & n28981 ;
  assign n29349 = ~n29347 & n29348 ;
  assign n29350 = n29349 ^ n5810 ^ n2535 ;
  assign n29351 = ( x118 & n4491 ) | ( x118 & ~n24928 ) | ( n4491 & ~n24928 ) ;
  assign n29352 = n29351 ^ n10023 ^ n8923 ;
  assign n29353 = n19626 ^ n10101 ^ 1'b0 ;
  assign n29354 = ( n9271 & ~n26698 ) | ( n9271 & n29353 ) | ( ~n26698 & n29353 ) ;
  assign n29355 = ( n4700 & ~n16930 ) | ( n4700 & n29354 ) | ( ~n16930 & n29354 ) ;
  assign n29356 = ( n13348 & n29352 ) | ( n13348 & n29355 ) | ( n29352 & n29355 ) ;
  assign n29357 = n21511 ^ n9328 ^ n739 ;
  assign n29358 = ( ~n13025 & n21878 ) | ( ~n13025 & n29357 ) | ( n21878 & n29357 ) ;
  assign n29359 = ( ~n10899 & n26889 ) | ( ~n10899 & n28146 ) | ( n26889 & n28146 ) ;
  assign n29360 = n9508 ^ n748 ^ n571 ;
  assign n29361 = n29360 ^ n22179 ^ n16982 ;
  assign n29362 = ( n18198 & n21142 ) | ( n18198 & ~n29361 ) | ( n21142 & ~n29361 ) ;
  assign n29364 = n4544 | n22094 ;
  assign n29365 = n323 & ~n29364 ;
  assign n29366 = n11140 | n29365 ;
  assign n29367 = n17022 | n29366 ;
  assign n29363 = n19883 ^ n12482 ^ n5246 ;
  assign n29368 = n29367 ^ n29363 ^ 1'b0 ;
  assign n29373 = n8492 & n10250 ;
  assign n29374 = n29373 ^ n3003 ^ n1832 ;
  assign n29369 = n20989 ^ n8896 ^ n2271 ;
  assign n29370 = n29369 ^ n8740 ^ n1572 ;
  assign n29371 = ( n4071 & ~n7991 ) | ( n4071 & n29370 ) | ( ~n7991 & n29370 ) ;
  assign n29372 = n29371 ^ n9614 ^ n3267 ;
  assign n29375 = n29374 ^ n29372 ^ 1'b0 ;
  assign n29376 = n13245 ^ n9571 ^ 1'b0 ;
  assign n29377 = n6302 ^ n5711 ^ 1'b0 ;
  assign n29378 = ( ~n9041 & n13556 ) | ( ~n9041 & n29377 ) | ( n13556 & n29377 ) ;
  assign n29379 = n27100 & n27893 ;
  assign n29380 = n29379 ^ n10611 ^ 1'b0 ;
  assign n29381 = n12254 ^ n4443 ^ 1'b0 ;
  assign n29382 = n27497 ^ n18237 ^ 1'b0 ;
  assign n29383 = n12529 & ~n29382 ;
  assign n29384 = ( n16731 & ~n29381 ) | ( n16731 & n29383 ) | ( ~n29381 & n29383 ) ;
  assign n29385 = n8977 | n15454 ;
  assign n29386 = ( n6092 & ~n25101 ) | ( n6092 & n25400 ) | ( ~n25101 & n25400 ) ;
  assign n29387 = ( n4799 & ~n6167 ) | ( n4799 & n20983 ) | ( ~n6167 & n20983 ) ;
  assign n29388 = n6952 | n29387 ;
  assign n29389 = n6563 | n29388 ;
  assign n29390 = n15833 ^ n12424 ^ n774 ;
  assign n29391 = n29390 ^ n13660 ^ 1'b0 ;
  assign n29392 = n1294 & ~n12698 ;
  assign n29393 = n29392 ^ n7727 ^ n3342 ;
  assign n29394 = n23815 ^ x120 ^ 1'b0 ;
  assign n29395 = ( n10441 & n11600 ) | ( n10441 & ~n22255 ) | ( n11600 & ~n22255 ) ;
  assign n29398 = ( n2666 & n5387 ) | ( n2666 & n12950 ) | ( n5387 & n12950 ) ;
  assign n29399 = ( ~n6034 & n16784 ) | ( ~n6034 & n19046 ) | ( n16784 & n19046 ) ;
  assign n29400 = n1915 | n29399 ;
  assign n29401 = ( n16960 & ~n29398 ) | ( n16960 & n29400 ) | ( ~n29398 & n29400 ) ;
  assign n29396 = n13145 | n29351 ;
  assign n29397 = ~n17090 & n29396 ;
  assign n29402 = n29401 ^ n29397 ^ 1'b0 ;
  assign n29403 = ( n6094 & n6591 ) | ( n6094 & ~n19781 ) | ( n6591 & ~n19781 ) ;
  assign n29404 = n29403 ^ n4537 ^ n2093 ;
  assign n29405 = n13788 | n29404 ;
  assign n29406 = ( n2846 & n29402 ) | ( n2846 & n29405 ) | ( n29402 & n29405 ) ;
  assign n29409 = ( n1279 & n2054 ) | ( n1279 & ~n3314 ) | ( n2054 & ~n3314 ) ;
  assign n29407 = ~n4189 & n11917 ;
  assign n29408 = n19383 & n29407 ;
  assign n29410 = n29409 ^ n29408 ^ n6185 ;
  assign n29411 = ( n1074 & n15074 ) | ( n1074 & n16740 ) | ( n15074 & n16740 ) ;
  assign n29412 = n22586 & n29411 ;
  assign n29413 = ~n6020 & n29412 ;
  assign n29414 = ( n8233 & ~n29410 ) | ( n8233 & n29413 ) | ( ~n29410 & n29413 ) ;
  assign n29415 = n25414 ^ n20219 ^ 1'b0 ;
  assign n29416 = n15207 & ~n29415 ;
  assign n29417 = n29416 ^ n13291 ^ 1'b0 ;
  assign n29418 = ( n14538 & n29414 ) | ( n14538 & n29417 ) | ( n29414 & n29417 ) ;
  assign n29419 = n13501 ^ n6891 ^ n2698 ;
  assign n29420 = n1074 & ~n23841 ;
  assign n29421 = ( ~n2587 & n13860 ) | ( ~n2587 & n20247 ) | ( n13860 & n20247 ) ;
  assign n29422 = ( n29419 & n29420 ) | ( n29419 & ~n29421 ) | ( n29420 & ~n29421 ) ;
  assign n29423 = ~n1499 & n12261 ;
  assign n29424 = n29423 ^ n10761 ^ 1'b0 ;
  assign n29425 = ( ~n12774 & n13544 ) | ( ~n12774 & n28784 ) | ( n13544 & n28784 ) ;
  assign n29426 = n25830 ^ n11569 ^ n545 ;
  assign n29427 = n29426 ^ n24009 ^ n12645 ;
  assign n29428 = ~n25430 & n29427 ;
  assign n29429 = n5543 & n29428 ;
  assign n29430 = n29429 ^ n15582 ^ n10538 ;
  assign n29431 = n6187 ^ n5871 ^ n2930 ;
  assign n29432 = ( n4270 & n6587 ) | ( n4270 & n13831 ) | ( n6587 & n13831 ) ;
  assign n29433 = n17792 & n29432 ;
  assign n29434 = n2169 & n29433 ;
  assign n29435 = n23701 ^ n22158 ^ n2830 ;
  assign n29436 = n29435 ^ n4160 ^ 1'b0 ;
  assign n29437 = n29004 | n29436 ;
  assign n29438 = n29437 ^ n19659 ^ 1'b0 ;
  assign n29439 = ( n6988 & n22564 ) | ( n6988 & n29438 ) | ( n22564 & n29438 ) ;
  assign n29440 = n29439 ^ n4574 ^ 1'b0 ;
  assign n29441 = n26595 ^ n11293 ^ x240 ;
  assign n29442 = ( x206 & ~n12770 ) | ( x206 & n29441 ) | ( ~n12770 & n29441 ) ;
  assign n29443 = n1352 | n23377 ;
  assign n29444 = n29443 ^ n3039 ^ 1'b0 ;
  assign n29445 = n11566 ^ n1295 ^ 1'b0 ;
  assign n29446 = n17880 ^ n15422 ^ n12830 ;
  assign n29447 = ( n29444 & n29445 ) | ( n29444 & n29446 ) | ( n29445 & n29446 ) ;
  assign n29448 = n10797 ^ n422 ^ 1'b0 ;
  assign n29449 = n14519 & n19053 ;
  assign n29450 = n10938 & n29449 ;
  assign n29451 = ( n7322 & n17677 ) | ( n7322 & n29450 ) | ( n17677 & n29450 ) ;
  assign n29452 = n17893 ^ n8013 ^ x211 ;
  assign n29453 = ( n13063 & n16952 ) | ( n13063 & n29452 ) | ( n16952 & n29452 ) ;
  assign n29454 = n18672 ^ n8346 ^ 1'b0 ;
  assign n29455 = n28540 ^ n19369 ^ 1'b0 ;
  assign n29456 = n29455 ^ n13122 ^ 1'b0 ;
  assign n29457 = n7523 | n29456 ;
  assign n29458 = n29454 | n29457 ;
  assign n29459 = n25253 ^ n23911 ^ 1'b0 ;
  assign n29460 = n6306 & ~n29459 ;
  assign n29461 = ( n1555 & n24888 ) | ( n1555 & ~n29460 ) | ( n24888 & ~n29460 ) ;
  assign n29462 = n29461 ^ n17528 ^ n10149 ;
  assign n29463 = ( n7313 & n11841 ) | ( n7313 & n21713 ) | ( n11841 & n21713 ) ;
  assign n29464 = n29463 ^ n5654 ^ n2983 ;
  assign n29465 = n29464 ^ n21711 ^ n3290 ;
  assign n29466 = n2107 | n5329 ;
  assign n29467 = n29466 ^ n17761 ^ 1'b0 ;
  assign n29468 = n19316 ^ n10139 ^ n9830 ;
  assign n29469 = ( ~n7485 & n29467 ) | ( ~n7485 & n29468 ) | ( n29467 & n29468 ) ;
  assign n29470 = ( n5061 & n9022 ) | ( n5061 & n29469 ) | ( n9022 & n29469 ) ;
  assign n29471 = ~n2344 & n15653 ;
  assign n29472 = n11360 & n29471 ;
  assign n29473 = n29472 ^ n26957 ^ n7466 ;
  assign n29474 = ( n8511 & n24000 ) | ( n8511 & n29473 ) | ( n24000 & n29473 ) ;
  assign n29475 = n29474 ^ n9620 ^ n8561 ;
  assign n29476 = n4216 ^ n1084 ^ 1'b0 ;
  assign n29477 = n3073 | n29476 ;
  assign n29481 = ( n12343 & n22623 ) | ( n12343 & ~n29351 ) | ( n22623 & ~n29351 ) ;
  assign n29478 = ( n8150 & ~n11930 ) | ( n8150 & n26124 ) | ( ~n11930 & n26124 ) ;
  assign n29479 = n2602 | n12867 ;
  assign n29480 = n29478 & ~n29479 ;
  assign n29482 = n29481 ^ n29480 ^ 1'b0 ;
  assign n29483 = n20084 ^ n9571 ^ 1'b0 ;
  assign n29484 = n29482 & n29483 ;
  assign n29485 = ( n4205 & n15506 ) | ( n4205 & n20851 ) | ( n15506 & n20851 ) ;
  assign n29486 = ( n9527 & n22764 ) | ( n9527 & ~n29485 ) | ( n22764 & ~n29485 ) ;
  assign n29495 = n2600 | n4887 ;
  assign n29492 = n9211 | n16450 ;
  assign n29493 = n29492 ^ n7177 ^ 1'b0 ;
  assign n29490 = ( ~n5411 & n12296 ) | ( ~n5411 & n14136 ) | ( n12296 & n14136 ) ;
  assign n29491 = ( n19348 & ~n19428 ) | ( n19348 & n29490 ) | ( ~n19428 & n29490 ) ;
  assign n29494 = n29493 ^ n29491 ^ n3860 ;
  assign n29496 = n29495 ^ n29494 ^ n13008 ;
  assign n29487 = x246 & n8332 ;
  assign n29488 = ~n10783 & n29487 ;
  assign n29489 = ( n7589 & n23104 ) | ( n7589 & ~n29488 ) | ( n23104 & ~n29488 ) ;
  assign n29497 = n29496 ^ n29489 ^ n13069 ;
  assign n29502 = ( n977 & ~n6636 ) | ( n977 & n8819 ) | ( ~n6636 & n8819 ) ;
  assign n29500 = ( n11137 & n16168 ) | ( n11137 & n19810 ) | ( n16168 & n19810 ) ;
  assign n29498 = ~n771 & n6961 ;
  assign n29499 = n29498 ^ n11969 ^ 1'b0 ;
  assign n29501 = n29500 ^ n29499 ^ n20818 ;
  assign n29503 = n29502 ^ n29501 ^ n7393 ;
  assign n29504 = ( n2491 & n7217 ) | ( n2491 & n20616 ) | ( n7217 & n20616 ) ;
  assign n29505 = n11979 ^ n8356 ^ n1485 ;
  assign n29506 = n29505 ^ n10803 ^ 1'b0 ;
  assign n29507 = ( n20133 & ~n29504 ) | ( n20133 & n29506 ) | ( ~n29504 & n29506 ) ;
  assign n29508 = ( ~n9908 & n15990 ) | ( ~n9908 & n26296 ) | ( n15990 & n26296 ) ;
  assign n29509 = n17060 ^ n12756 ^ 1'b0 ;
  assign n29510 = n4772 | n29509 ;
  assign n29511 = ( n3759 & ~n24183 ) | ( n3759 & n29510 ) | ( ~n24183 & n29510 ) ;
  assign n29512 = n9556 ^ n1102 ^ 1'b0 ;
  assign n29513 = n26648 ^ x166 ^ 1'b0 ;
  assign n29514 = n29513 ^ n29452 ^ n2941 ;
  assign n29515 = ( ~n3090 & n9885 ) | ( ~n3090 & n29514 ) | ( n9885 & n29514 ) ;
  assign n29522 = n17913 ^ n13583 ^ n8126 ;
  assign n29517 = ( n3671 & n6528 ) | ( n3671 & n9352 ) | ( n6528 & n9352 ) ;
  assign n29518 = n29517 ^ n24367 ^ n7793 ;
  assign n29519 = ( n1816 & n7006 ) | ( n1816 & ~n29518 ) | ( n7006 & ~n29518 ) ;
  assign n29520 = ( ~n8264 & n22171 ) | ( ~n8264 & n29519 ) | ( n22171 & n29519 ) ;
  assign n29521 = ( ~n496 & n25051 ) | ( ~n496 & n29520 ) | ( n25051 & n29520 ) ;
  assign n29516 = n22356 ^ n22120 ^ n3657 ;
  assign n29523 = n29522 ^ n29521 ^ n29516 ;
  assign n29524 = n2553 & ~n9082 ;
  assign n29525 = ~n5875 & n18663 ;
  assign n29526 = n29525 ^ n14641 ^ 1'b0 ;
  assign n29527 = ( n25679 & n25863 ) | ( n25679 & ~n28176 ) | ( n25863 & ~n28176 ) ;
  assign n29528 = ~n20957 & n21016 ;
  assign n29529 = ( n395 & ~n13587 ) | ( n395 & n15156 ) | ( ~n13587 & n15156 ) ;
  assign n29530 = ~n14490 & n29529 ;
  assign n29531 = ( n1543 & n2517 ) | ( n1543 & ~n16696 ) | ( n2517 & ~n16696 ) ;
  assign n29532 = n29531 ^ n8897 ^ n4299 ;
  assign n29533 = ( n5550 & ~n8656 ) | ( n5550 & n29532 ) | ( ~n8656 & n29532 ) ;
  assign n29535 = n22392 ^ n11715 ^ n9380 ;
  assign n29534 = ( n11198 & ~n12404 ) | ( n11198 & n19953 ) | ( ~n12404 & n19953 ) ;
  assign n29536 = n29535 ^ n29534 ^ n27583 ;
  assign n29537 = n29536 ^ n15255 ^ 1'b0 ;
  assign n29538 = n7337 & n29537 ;
  assign n29539 = ( n962 & n7794 ) | ( n962 & n21008 ) | ( n7794 & n21008 ) ;
  assign n29540 = n26380 ^ n6255 ^ n1817 ;
  assign n29541 = ( n10363 & n19460 ) | ( n10363 & n29540 ) | ( n19460 & n29540 ) ;
  assign n29542 = n21798 ^ n9642 ^ n6582 ;
  assign n29543 = n15011 & ~n29542 ;
  assign n29544 = n29543 ^ n11063 ^ n9610 ;
  assign n29545 = ( n847 & n14465 ) | ( n847 & ~n14687 ) | ( n14465 & ~n14687 ) ;
  assign n29546 = ( n3556 & n28355 ) | ( n3556 & ~n29545 ) | ( n28355 & ~n29545 ) ;
  assign n29547 = n8965 ^ n8036 ^ 1'b0 ;
  assign n29548 = n12780 | n29547 ;
  assign n29549 = n29548 ^ n10970 ^ n5689 ;
  assign n29550 = n29549 ^ n20642 ^ n13363 ;
  assign n29551 = n28364 ^ n11500 ^ n487 ;
  assign n29552 = n29551 ^ n20258 ^ n13069 ;
  assign n29553 = ( ~n642 & n4253 ) | ( ~n642 & n5736 ) | ( n4253 & n5736 ) ;
  assign n29554 = ~n25252 & n29553 ;
  assign n29555 = n29554 ^ n6730 ^ 1'b0 ;
  assign n29556 = n9758 & ~n29555 ;
  assign n29557 = ~n8967 & n29556 ;
  assign n29558 = ( n861 & n8408 ) | ( n861 & ~n12439 ) | ( n8408 & ~n12439 ) ;
  assign n29559 = n9686 & n29558 ;
  assign n29560 = ~n5953 & n29559 ;
  assign n29561 = ( n5506 & ~n29557 ) | ( n5506 & n29560 ) | ( ~n29557 & n29560 ) ;
  assign n29562 = n29561 ^ n24575 ^ n1042 ;
  assign n29563 = n25214 ^ n19200 ^ n4190 ;
  assign n29564 = n29563 ^ n1619 ^ 1'b0 ;
  assign n29566 = ( n10631 & n13297 ) | ( n10631 & ~n16081 ) | ( n13297 & ~n16081 ) ;
  assign n29565 = ( n2917 & n18278 ) | ( n2917 & ~n23555 ) | ( n18278 & ~n23555 ) ;
  assign n29567 = n29566 ^ n29565 ^ n23558 ;
  assign n29568 = ( n744 & ~n14162 ) | ( n744 & n17548 ) | ( ~n14162 & n17548 ) ;
  assign n29569 = n4024 & ~n20475 ;
  assign n29570 = ~n7378 & n29569 ;
  assign n29571 = ( n20226 & n23987 ) | ( n20226 & ~n29570 ) | ( n23987 & ~n29570 ) ;
  assign n29572 = n23667 ^ n7539 ^ n2408 ;
  assign n29573 = ( n414 & n5908 ) | ( n414 & n15078 ) | ( n5908 & n15078 ) ;
  assign n29574 = ~n9137 & n29573 ;
  assign n29575 = n29574 ^ n27996 ^ 1'b0 ;
  assign n29576 = ( ~n1881 & n29572 ) | ( ~n1881 & n29575 ) | ( n29572 & n29575 ) ;
  assign n29582 = ~n7869 & n11736 ;
  assign n29581 = n9289 & n29444 ;
  assign n29583 = n29582 ^ n29581 ^ 1'b0 ;
  assign n29578 = ( n3245 & ~n4142 ) | ( n3245 & n12042 ) | ( ~n4142 & n12042 ) ;
  assign n29577 = ( n1695 & n3069 ) | ( n1695 & ~n5867 ) | ( n3069 & ~n5867 ) ;
  assign n29579 = n29578 ^ n29577 ^ n7329 ;
  assign n29580 = n6409 & ~n29579 ;
  assign n29584 = n29583 ^ n29580 ^ n1325 ;
  assign n29587 = ~n3857 & n9253 ;
  assign n29588 = ~n5209 & n29587 ;
  assign n29585 = ( n418 & n1545 ) | ( n418 & ~n8182 ) | ( n1545 & ~n8182 ) ;
  assign n29586 = ( n20778 & n27436 ) | ( n20778 & ~n29585 ) | ( n27436 & ~n29585 ) ;
  assign n29589 = n29588 ^ n29586 ^ n19532 ;
  assign n29590 = n29589 ^ n29008 ^ 1'b0 ;
  assign n29591 = n29584 & n29590 ;
  assign n29592 = ( n1959 & n5337 ) | ( n1959 & ~n15346 ) | ( n5337 & ~n15346 ) ;
  assign n29593 = n29592 ^ n6788 ^ 1'b0 ;
  assign n29594 = n29593 ^ x5 ^ 1'b0 ;
  assign n29595 = n29594 ^ n18179 ^ 1'b0 ;
  assign n29596 = ( n283 & ~n4081 ) | ( n283 & n18894 ) | ( ~n4081 & n18894 ) ;
  assign n29597 = ( ~n7043 & n7576 ) | ( ~n7043 & n29596 ) | ( n7576 & n29596 ) ;
  assign n29598 = n9279 & n12374 ;
  assign n29599 = n29598 ^ n19527 ^ n16682 ;
  assign n29600 = ( n5312 & n29597 ) | ( n5312 & ~n29599 ) | ( n29597 & ~n29599 ) ;
  assign n29601 = n28196 ^ n9459 ^ 1'b0 ;
  assign n29602 = ( n2231 & ~n13515 ) | ( n2231 & n14762 ) | ( ~n13515 & n14762 ) ;
  assign n29603 = n29602 ^ n3029 ^ n916 ;
  assign n29604 = ~n631 & n29603 ;
  assign n29605 = n29604 ^ n7728 ^ 1'b0 ;
  assign n29609 = ~n5083 & n11989 ;
  assign n29610 = n29609 ^ n28760 ^ 1'b0 ;
  assign n29606 = n18383 ^ n12023 ^ n571 ;
  assign n29607 = n26718 ^ n25069 ^ n20593 ;
  assign n29608 = ~n29606 & n29607 ;
  assign n29611 = n29610 ^ n29608 ^ 1'b0 ;
  assign n29614 = n7110 ^ n6190 ^ n2823 ;
  assign n29612 = n15745 ^ n5231 ^ x189 ;
  assign n29613 = ( ~n3973 & n4692 ) | ( ~n3973 & n29612 ) | ( n4692 & n29612 ) ;
  assign n29615 = n29614 ^ n29613 ^ n14918 ;
  assign n29616 = n13241 ^ n2204 ^ 1'b0 ;
  assign n29617 = n29616 ^ n8471 ^ n1658 ;
  assign n29618 = n3018 ^ n2964 ^ x126 ;
  assign n29619 = ( n1882 & n10822 ) | ( n1882 & n29618 ) | ( n10822 & n29618 ) ;
  assign n29620 = ( ~n15324 & n19533 ) | ( ~n15324 & n29619 ) | ( n19533 & n29619 ) ;
  assign n29621 = n28539 ^ n22895 ^ n8546 ;
  assign n29622 = n7612 | n8110 ;
  assign n29623 = n17992 ^ n9692 ^ 1'b0 ;
  assign n29624 = n29623 ^ n12740 ^ 1'b0 ;
  assign n29625 = ( ~n17857 & n29622 ) | ( ~n17857 & n29624 ) | ( n29622 & n29624 ) ;
  assign n29627 = n3100 | n12067 ;
  assign n29628 = n16602 & ~n29627 ;
  assign n29629 = n15977 ^ n3701 ^ 1'b0 ;
  assign n29630 = n1886 & ~n29629 ;
  assign n29631 = ( n21806 & n29628 ) | ( n21806 & n29630 ) | ( n29628 & n29630 ) ;
  assign n29626 = n5019 ^ n2877 ^ 1'b0 ;
  assign n29632 = n29631 ^ n29626 ^ n29350 ;
  assign n29633 = ~n9999 & n10260 ;
  assign n29634 = ( ~n4096 & n13582 ) | ( ~n4096 & n20412 ) | ( n13582 & n20412 ) ;
  assign n29635 = ( n14770 & ~n17407 ) | ( n14770 & n29555 ) | ( ~n17407 & n29555 ) ;
  assign n29636 = ( n19373 & n24723 ) | ( n19373 & n29635 ) | ( n24723 & n29635 ) ;
  assign n29639 = ( n920 & n976 ) | ( n920 & ~n18044 ) | ( n976 & ~n18044 ) ;
  assign n29637 = ~n822 & n10897 ;
  assign n29638 = ~n8068 & n29637 ;
  assign n29640 = n29639 ^ n29638 ^ n17207 ;
  assign n29642 = n10803 ^ n5161 ^ n5133 ;
  assign n29643 = n13238 & n29642 ;
  assign n29641 = ( x8 & n15637 ) | ( x8 & ~n16496 ) | ( n15637 & ~n16496 ) ;
  assign n29644 = n29643 ^ n29641 ^ n936 ;
  assign n29645 = ( n3255 & n13505 ) | ( n3255 & n24082 ) | ( n13505 & n24082 ) ;
  assign n29646 = n9705 | n21256 ;
  assign n29647 = n29646 ^ n19877 ^ 1'b0 ;
  assign n29648 = n16646 ^ n13603 ^ n369 ;
  assign n29649 = ( n14746 & n17798 ) | ( n14746 & n29648 ) | ( n17798 & n29648 ) ;
  assign n29650 = ~n7388 & n18622 ;
  assign n29651 = ~n29649 & n29650 ;
  assign n29652 = ( ~n4375 & n11683 ) | ( ~n4375 & n29651 ) | ( n11683 & n29651 ) ;
  assign n29653 = n1696 & n9790 ;
  assign n29654 = ( ~n11490 & n23780 ) | ( ~n11490 & n27460 ) | ( n23780 & n27460 ) ;
  assign n29655 = ~n9737 & n10477 ;
  assign n29656 = n29655 ^ n3954 ^ 1'b0 ;
  assign n29657 = n29408 ^ n14976 ^ n5776 ;
  assign n29658 = n17343 ^ n16554 ^ 1'b0 ;
  assign n29659 = n29657 | n29658 ;
  assign n29660 = n29140 ^ n10631 ^ n2462 ;
  assign n29661 = ( n7966 & ~n19873 ) | ( n7966 & n26465 ) | ( ~n19873 & n26465 ) ;
  assign n29662 = n8619 & ~n29661 ;
  assign n29663 = n9579 ^ n8885 ^ n4221 ;
  assign n29664 = n29663 ^ n22516 ^ n7515 ;
  assign n29665 = ( n5935 & n6626 ) | ( n5935 & ~n29664 ) | ( n6626 & ~n29664 ) ;
  assign n29666 = ( n2028 & n20021 ) | ( n2028 & ~n26544 ) | ( n20021 & ~n26544 ) ;
  assign n29667 = n29666 ^ n22410 ^ n7909 ;
  assign n29668 = ( n3185 & n11348 ) | ( n3185 & ~n23685 ) | ( n11348 & ~n23685 ) ;
  assign n29669 = n29668 ^ n10918 ^ 1'b0 ;
  assign n29670 = n24539 & ~n29669 ;
  assign n29671 = ( x203 & ~n3154 ) | ( x203 & n29670 ) | ( ~n3154 & n29670 ) ;
  assign n29672 = n3132 & n29671 ;
  assign n29674 = n11545 | n28944 ;
  assign n29675 = n9507 | n29674 ;
  assign n29676 = ~n2107 & n29675 ;
  assign n29677 = n19880 & n29676 ;
  assign n29673 = n9255 & ~n17103 ;
  assign n29678 = n29677 ^ n29673 ^ 1'b0 ;
  assign n29679 = ( n15435 & ~n18440 ) | ( n15435 & n21506 ) | ( ~n18440 & n21506 ) ;
  assign n29680 = ( n6441 & ~n10779 ) | ( n6441 & n27070 ) | ( ~n10779 & n27070 ) ;
  assign n29682 = n23451 ^ n20906 ^ n3664 ;
  assign n29683 = ( n17099 & n24770 ) | ( n17099 & ~n29682 ) | ( n24770 & ~n29682 ) ;
  assign n29684 = n3742 | n29683 ;
  assign n29685 = n29684 ^ n12346 ^ 1'b0 ;
  assign n29681 = n20752 ^ n3190 ^ 1'b0 ;
  assign n29686 = n29685 ^ n29681 ^ n25066 ;
  assign n29687 = ( n4048 & n14727 ) | ( n4048 & ~n14945 ) | ( n14727 & ~n14945 ) ;
  assign n29688 = n10113 ^ n938 ^ 1'b0 ;
  assign n29689 = n29687 & ~n29688 ;
  assign n29693 = n25101 ^ n25006 ^ n17156 ;
  assign n29691 = ( ~n4834 & n6552 ) | ( ~n4834 & n16188 ) | ( n6552 & n16188 ) ;
  assign n29690 = n19184 ^ n3317 ^ 1'b0 ;
  assign n29692 = n29691 ^ n29690 ^ n14879 ;
  assign n29694 = n29693 ^ n29692 ^ n14380 ;
  assign n29695 = n16030 ^ n12290 ^ 1'b0 ;
  assign n29696 = n29694 & n29695 ;
  assign n29697 = ~n21530 & n29696 ;
  assign n29700 = n27250 ^ n16774 ^ n4075 ;
  assign n29698 = n8770 ^ n4205 ^ 1'b0 ;
  assign n29699 = ( n4830 & n28727 ) | ( n4830 & n29698 ) | ( n28727 & n29698 ) ;
  assign n29701 = n29700 ^ n29699 ^ n5253 ;
  assign n29702 = n20630 ^ n11758 ^ n3519 ;
  assign n29703 = n10131 & n29702 ;
  assign n29704 = n29703 ^ n16903 ^ 1'b0 ;
  assign n29705 = n2078 & n4446 ;
  assign n29706 = n29705 ^ n2257 ^ 1'b0 ;
  assign n29707 = n29706 ^ x94 ^ 1'b0 ;
  assign n29708 = n29707 ^ n17466 ^ 1'b0 ;
  assign n29709 = n851 & ~n29708 ;
  assign n29710 = n22581 ^ n6087 ^ 1'b0 ;
  assign n29711 = ( n1034 & n21533 ) | ( n1034 & ~n28840 ) | ( n21533 & ~n28840 ) ;
  assign n29717 = ( n11665 & n17191 ) | ( n11665 & n26889 ) | ( n17191 & n26889 ) ;
  assign n29712 = ( ~n3187 & n17549 ) | ( ~n3187 & n25272 ) | ( n17549 & n25272 ) ;
  assign n29713 = n29712 ^ n10356 ^ n622 ;
  assign n29714 = n19148 ^ n14998 ^ 1'b0 ;
  assign n29715 = ~n29713 & n29714 ;
  assign n29716 = ~n13890 & n29715 ;
  assign n29718 = n29717 ^ n29716 ^ 1'b0 ;
  assign n29719 = n23437 ^ n3892 ^ 1'b0 ;
  assign n29720 = ( n8369 & n24546 ) | ( n8369 & n29719 ) | ( n24546 & n29719 ) ;
  assign n29721 = ( n9859 & ~n11263 ) | ( n9859 & n23964 ) | ( ~n11263 & n23964 ) ;
  assign n29722 = ( n28884 & n29720 ) | ( n28884 & ~n29721 ) | ( n29720 & ~n29721 ) ;
  assign n29723 = n15501 ^ n6358 ^ n1781 ;
  assign n29724 = n29712 ^ n3430 ^ n651 ;
  assign n29725 = ( n589 & n16778 ) | ( n589 & n29724 ) | ( n16778 & n29724 ) ;
  assign n29726 = n18109 ^ n13526 ^ 1'b0 ;
  assign n29727 = n29726 ^ n9561 ^ 1'b0 ;
  assign n29728 = n10959 & ~n15983 ;
  assign n29729 = n29728 ^ n23511 ^ 1'b0 ;
  assign n29730 = n29729 ^ n473 ^ 1'b0 ;
  assign n29731 = n10718 ^ n2744 ^ n1832 ;
  assign n29732 = ( n4447 & n7627 ) | ( n4447 & ~n23091 ) | ( n7627 & ~n23091 ) ;
  assign n29733 = n29732 ^ n29372 ^ 1'b0 ;
  assign n29734 = ( n13999 & n15648 ) | ( n13999 & n29733 ) | ( n15648 & n29733 ) ;
  assign n29735 = ~n13008 & n29734 ;
  assign n29736 = ~n3565 & n29735 ;
  assign n29737 = ( n9510 & ~n29731 ) | ( n9510 & n29736 ) | ( ~n29731 & n29736 ) ;
  assign n29738 = n15713 ^ n5104 ^ 1'b0 ;
  assign n29739 = ~n7042 & n29738 ;
  assign n29743 = n25907 ^ n5049 ^ n2076 ;
  assign n29740 = x77 & ~n7792 ;
  assign n29741 = n29740 ^ n16390 ^ 1'b0 ;
  assign n29742 = n29741 ^ n22532 ^ n11782 ;
  assign n29744 = n29743 ^ n29742 ^ n20936 ;
  assign n29745 = n12026 | n19405 ;
  assign n29746 = ( n3837 & n7135 ) | ( n3837 & n13471 ) | ( n7135 & n13471 ) ;
  assign n29747 = ( n5114 & n29745 ) | ( n5114 & n29746 ) | ( n29745 & n29746 ) ;
  assign n29748 = ( n9833 & n20611 ) | ( n9833 & ~n25421 ) | ( n20611 & ~n25421 ) ;
  assign n29749 = n1734 | n3182 ;
  assign n29750 = n20572 | n29749 ;
  assign n29751 = n10728 ^ n10140 ^ n7606 ;
  assign n29752 = ( n6189 & n9046 ) | ( n6189 & ~n29751 ) | ( n9046 & ~n29751 ) ;
  assign n29753 = n29752 ^ n10975 ^ n8620 ;
  assign n29754 = ( n9109 & n9507 ) | ( n9109 & ~n13995 ) | ( n9507 & ~n13995 ) ;
  assign n29755 = ( n14135 & n25912 ) | ( n14135 & n29754 ) | ( n25912 & n29754 ) ;
  assign n29756 = ( x136 & ~n686 ) | ( x136 & n5090 ) | ( ~n686 & n5090 ) ;
  assign n29757 = x128 & ~n27436 ;
  assign n29758 = n3652 & n29757 ;
  assign n29759 = n29758 ^ n8468 ^ n1240 ;
  assign n29760 = ( n13138 & ~n29756 ) | ( n13138 & n29759 ) | ( ~n29756 & n29759 ) ;
  assign n29761 = n18799 ^ n8581 ^ 1'b0 ;
  assign n29762 = n28517 ^ n20595 ^ n16078 ;
  assign n29763 = ( ~n4512 & n5188 ) | ( ~n4512 & n10739 ) | ( n5188 & n10739 ) ;
  assign n29764 = n29763 ^ n9859 ^ n9542 ;
  assign n29765 = ( n11034 & n25189 ) | ( n11034 & n29764 ) | ( n25189 & n29764 ) ;
  assign n29766 = n9701 & n18680 ;
  assign n29767 = n29766 ^ n2465 ^ 1'b0 ;
  assign n29768 = n10184 & n25730 ;
  assign n29769 = n29767 & n29768 ;
  assign n29770 = n26441 & ~n29769 ;
  assign n29771 = n29770 ^ n26402 ^ 1'b0 ;
  assign n29772 = ( n281 & n3537 ) | ( n281 & ~n20718 ) | ( n3537 & ~n20718 ) ;
  assign n29773 = n892 & n29772 ;
  assign n29774 = n29773 ^ n20781 ^ 1'b0 ;
  assign n29775 = n5048 & ~n29774 ;
  assign n29779 = n5647 & n24900 ;
  assign n29780 = ~n4207 & n29779 ;
  assign n29781 = ( x156 & n4317 ) | ( x156 & ~n29780 ) | ( n4317 & ~n29780 ) ;
  assign n29776 = n5512 & n9816 ;
  assign n29777 = n11037 & n29776 ;
  assign n29778 = ( n11361 & ~n29064 ) | ( n11361 & n29777 ) | ( ~n29064 & n29777 ) ;
  assign n29782 = n29781 ^ n29778 ^ n12026 ;
  assign n29783 = ( n11360 & n17181 ) | ( n11360 & ~n24749 ) | ( n17181 & ~n24749 ) ;
  assign n29784 = ( ~n10828 & n20586 ) | ( ~n10828 & n28513 ) | ( n20586 & n28513 ) ;
  assign n29785 = n6480 ^ n4011 ^ 1'b0 ;
  assign n29786 = ( ~n5678 & n9937 ) | ( ~n5678 & n20576 ) | ( n9937 & n20576 ) ;
  assign n29787 = n29785 | n29786 ;
  assign n29788 = n29787 ^ n10607 ^ 1'b0 ;
  assign n29789 = ~n12507 & n24900 ;
  assign n29790 = ~n10813 & n29789 ;
  assign n29791 = n24969 ^ n2501 ^ n1079 ;
  assign n29792 = n29791 ^ n14131 ^ 1'b0 ;
  assign n29793 = n29790 | n29792 ;
  assign n29794 = n20580 & n26766 ;
  assign n29795 = ( n2172 & n14041 ) | ( n2172 & n25572 ) | ( n14041 & n25572 ) ;
  assign n29798 = n4785 & ~n11314 ;
  assign n29799 = n29798 ^ n12891 ^ 1'b0 ;
  assign n29796 = ( n13948 & n15219 ) | ( n13948 & n23962 ) | ( n15219 & n23962 ) ;
  assign n29797 = n9659 & ~n29796 ;
  assign n29800 = n29799 ^ n29797 ^ n12882 ;
  assign n29801 = n27162 ^ n5400 ^ 1'b0 ;
  assign n29802 = n931 | n29801 ;
  assign n29803 = n20044 ^ n15643 ^ n10563 ;
  assign n29804 = n29803 ^ n21399 ^ 1'b0 ;
  assign n29805 = n29804 ^ n13417 ^ n12370 ;
  assign n29806 = n13940 ^ n6294 ^ n2686 ;
  assign n29807 = ( n10859 & ~n21857 ) | ( n10859 & n29806 ) | ( ~n21857 & n29806 ) ;
  assign n29808 = ~n787 & n29807 ;
  assign n29811 = n3427 ^ n2014 ^ 1'b0 ;
  assign n29812 = n23568 | n29811 ;
  assign n29813 = n13142 | n29812 ;
  assign n29809 = n16292 | n23279 ;
  assign n29810 = n29809 ^ n17619 ^ 1'b0 ;
  assign n29814 = n29813 ^ n29810 ^ n24070 ;
  assign n29815 = n11281 ^ n643 ^ 1'b0 ;
  assign n29816 = n17278 & n29815 ;
  assign n29817 = ( n18594 & ~n20520 ) | ( n18594 & n22410 ) | ( ~n20520 & n22410 ) ;
  assign n29818 = ( n11827 & n29816 ) | ( n11827 & ~n29817 ) | ( n29816 & ~n29817 ) ;
  assign n29819 = ( n7838 & ~n29814 ) | ( n7838 & n29818 ) | ( ~n29814 & n29818 ) ;
  assign n29820 = n6000 & n18725 ;
  assign n29821 = ~n12881 & n29820 ;
  assign n29822 = ( n16418 & n25352 ) | ( n16418 & ~n29821 ) | ( n25352 & ~n29821 ) ;
  assign n29825 = ( n4825 & ~n8784 ) | ( n4825 & n18370 ) | ( ~n8784 & n18370 ) ;
  assign n29823 = ( n2199 & n3784 ) | ( n2199 & ~n5598 ) | ( n3784 & ~n5598 ) ;
  assign n29824 = n348 | n29823 ;
  assign n29826 = n29825 ^ n29824 ^ n15670 ;
  assign n29827 = ( ~n7627 & n7983 ) | ( ~n7627 & n25393 ) | ( n7983 & n25393 ) ;
  assign n29828 = n29827 ^ n3090 ^ 1'b0 ;
  assign n29829 = n29828 ^ n1986 ^ 1'b0 ;
  assign n29830 = n29829 ^ n18787 ^ n3864 ;
  assign n29831 = ( n784 & ~n10372 ) | ( n784 & n11414 ) | ( ~n10372 & n11414 ) ;
  assign n29832 = n29831 ^ n12630 ^ 1'b0 ;
  assign n29833 = n29830 | n29832 ;
  assign n29834 = n29833 ^ n1823 ^ 1'b0 ;
  assign n29835 = n4047 & n6468 ;
  assign n29836 = ~n4625 & n29835 ;
  assign n29844 = ~n1604 & n16887 ;
  assign n29837 = n17659 ^ n4503 ^ n3966 ;
  assign n29838 = ( x234 & ~n11535 ) | ( x234 & n29837 ) | ( ~n11535 & n29837 ) ;
  assign n29839 = ( n914 & n5174 ) | ( n914 & n14214 ) | ( n5174 & n14214 ) ;
  assign n29840 = n22064 & n29839 ;
  assign n29841 = n29840 ^ n15129 ^ n10425 ;
  assign n29842 = n29841 ^ n9794 ^ 1'b0 ;
  assign n29843 = n29838 & n29842 ;
  assign n29845 = n29844 ^ n29843 ^ 1'b0 ;
  assign n29846 = ~n13492 & n14729 ;
  assign n29847 = n16286 & n29846 ;
  assign n29848 = ~n2062 & n23174 ;
  assign n29849 = n22681 & n29848 ;
  assign n29850 = ( n21636 & n29847 ) | ( n21636 & ~n29849 ) | ( n29847 & ~n29849 ) ;
  assign n29851 = n5831 & ~n22568 ;
  assign n29855 = n21543 ^ n10508 ^ n5705 ;
  assign n29852 = n15617 ^ n4708 ^ n2877 ;
  assign n29853 = n6819 & ~n29852 ;
  assign n29854 = ~n6056 & n29853 ;
  assign n29856 = n29855 ^ n29854 ^ 1'b0 ;
  assign n29857 = ~n4887 & n29856 ;
  assign n29858 = n9931 ^ n1908 ^ 1'b0 ;
  assign n29859 = ~n1030 & n29858 ;
  assign n29860 = n23500 & n29859 ;
  assign n29861 = ( n752 & ~n7838 ) | ( n752 & n29860 ) | ( ~n7838 & n29860 ) ;
  assign n29862 = ( n16745 & ~n18161 ) | ( n16745 & n24532 ) | ( ~n18161 & n24532 ) ;
  assign n29863 = n29862 ^ n28372 ^ n8718 ;
  assign n29864 = n7210 & ~n29863 ;
  assign n29865 = n5704 & n29864 ;
  assign n29866 = ( n12652 & ~n27443 ) | ( n12652 & n29865 ) | ( ~n27443 & n29865 ) ;
  assign n29867 = n3418 & n6250 ;
  assign n29868 = n4175 & n29867 ;
  assign n29869 = n25657 ^ n6177 ^ 1'b0 ;
  assign n29870 = ~n9728 & n21768 ;
  assign n29871 = n29870 ^ n18261 ^ 1'b0 ;
  assign n29872 = ( n29868 & n29869 ) | ( n29868 & n29871 ) | ( n29869 & n29871 ) ;
  assign n29873 = n614 & ~n12983 ;
  assign n29874 = n28108 & n29873 ;
  assign n29875 = n17582 ^ n16214 ^ n3396 ;
  assign n29876 = n29875 ^ n21698 ^ n17629 ;
  assign n29877 = n1481 & n3951 ;
  assign n29878 = n29877 ^ n6487 ^ 1'b0 ;
  assign n29879 = n29878 ^ n3398 ^ n1972 ;
  assign n29880 = n29879 ^ n18049 ^ 1'b0 ;
  assign n29881 = ( n23173 & n23385 ) | ( n23173 & n29880 ) | ( n23385 & n29880 ) ;
  assign n29882 = ( n5260 & n18451 ) | ( n5260 & ~n24887 ) | ( n18451 & ~n24887 ) ;
  assign n29883 = ( n13286 & n29881 ) | ( n13286 & ~n29882 ) | ( n29881 & ~n29882 ) ;
  assign n29884 = ( n9717 & n18132 ) | ( n9717 & n27416 ) | ( n18132 & n27416 ) ;
  assign n29885 = n19380 & n29884 ;
  assign n29886 = n21215 ^ n7759 ^ 1'b0 ;
  assign n29887 = ~n8291 & n29886 ;
  assign n29888 = ( n5432 & n14165 ) | ( n5432 & n29887 ) | ( n14165 & n29887 ) ;
  assign n29889 = ( n6184 & n16492 ) | ( n6184 & ~n24646 ) | ( n16492 & ~n24646 ) ;
  assign n29890 = ( ~n23775 & n26725 ) | ( ~n23775 & n29889 ) | ( n26725 & n29889 ) ;
  assign n29891 = ( n3616 & n8930 ) | ( n3616 & n14414 ) | ( n8930 & n14414 ) ;
  assign n29892 = ~n8844 & n15047 ;
  assign n29893 = ~n29891 & n29892 ;
  assign n29894 = n29893 ^ n28178 ^ 1'b0 ;
  assign n29895 = n29890 & ~n29894 ;
  assign n29896 = n29888 & n29895 ;
  assign n29897 = n29896 ^ n3079 ^ 1'b0 ;
  assign n29898 = ( ~n2731 & n6284 ) | ( ~n2731 & n21408 ) | ( n6284 & n21408 ) ;
  assign n29899 = ( n3358 & n25183 ) | ( n3358 & ~n29898 ) | ( n25183 & ~n29898 ) ;
  assign n29900 = ( ~n3505 & n3514 ) | ( ~n3505 & n9760 ) | ( n3514 & n9760 ) ;
  assign n29901 = n11945 ^ n6592 ^ 1'b0 ;
  assign n29902 = ~n29900 & n29901 ;
  assign n29903 = ~n12403 & n29902 ;
  assign n29905 = ( n4582 & n14357 ) | ( n4582 & ~n16860 ) | ( n14357 & ~n16860 ) ;
  assign n29904 = ( n2993 & ~n13548 ) | ( n2993 & n25577 ) | ( ~n13548 & n25577 ) ;
  assign n29906 = n29905 ^ n29904 ^ n8036 ;
  assign n29907 = n2525 & ~n4992 ;
  assign n29908 = ~n4078 & n29907 ;
  assign n29909 = ~n5721 & n8346 ;
  assign n29910 = n29909 ^ n6609 ^ 1'b0 ;
  assign n29911 = ( n2251 & n29908 ) | ( n2251 & n29910 ) | ( n29908 & n29910 ) ;
  assign n29912 = n16842 | n27033 ;
  assign n29913 = n7312 & ~n29912 ;
  assign n29915 = n22057 ^ n20682 ^ 1'b0 ;
  assign n29916 = n4996 & n29915 ;
  assign n29914 = n6407 & ~n17282 ;
  assign n29917 = n29916 ^ n29914 ^ 1'b0 ;
  assign n29918 = n26751 ^ n1914 ^ x23 ;
  assign n29919 = ~n6096 & n29918 ;
  assign n29920 = n29919 ^ n28388 ^ n26222 ;
  assign n29921 = ( n4229 & n16324 ) | ( n4229 & ~n29291 ) | ( n16324 & ~n29291 ) ;
  assign n29922 = ( ~n1168 & n4466 ) | ( ~n1168 & n24649 ) | ( n4466 & n24649 ) ;
  assign n29923 = n24350 ^ n17583 ^ n12332 ;
  assign n29925 = n15371 | n25202 ;
  assign n29926 = ( n23474 & n28470 ) | ( n23474 & ~n29925 ) | ( n28470 & ~n29925 ) ;
  assign n29924 = n12544 ^ n287 ^ 1'b0 ;
  assign n29927 = n29926 ^ n29924 ^ 1'b0 ;
  assign n29928 = n29927 ^ n24670 ^ n19290 ;
  assign n29929 = n29928 ^ n11169 ^ n8917 ;
  assign n29930 = n11613 | n29929 ;
  assign n29931 = n20499 & ~n29930 ;
  assign n29932 = ( n29922 & n29923 ) | ( n29922 & n29931 ) | ( n29923 & n29931 ) ;
  assign n29934 = ( n337 & n5223 ) | ( n337 & n7760 ) | ( n5223 & n7760 ) ;
  assign n29935 = n29934 ^ n29409 ^ n494 ;
  assign n29936 = n29935 ^ n14253 ^ 1'b0 ;
  assign n29937 = n9144 ^ n5192 ^ 1'b0 ;
  assign n29938 = n22176 ^ n15856 ^ n10549 ;
  assign n29939 = n29938 ^ n26694 ^ n12256 ;
  assign n29940 = ( n29936 & n29937 ) | ( n29936 & n29939 ) | ( n29937 & n29939 ) ;
  assign n29933 = ( ~n5893 & n13612 ) | ( ~n5893 & n19308 ) | ( n13612 & n19308 ) ;
  assign n29941 = n29940 ^ n29933 ^ n19236 ;
  assign n29942 = ( n3207 & ~n18860 ) | ( n3207 & n20300 ) | ( ~n18860 & n20300 ) ;
  assign n29943 = n14584 | n29942 ;
  assign n29944 = ( n689 & n11915 ) | ( n689 & n26942 ) | ( n11915 & n26942 ) ;
  assign n29945 = n18704 ^ n18669 ^ 1'b0 ;
  assign n29946 = n1596 & n29945 ;
  assign n29947 = n12103 ^ n10987 ^ 1'b0 ;
  assign n29948 = ~n29852 & n29947 ;
  assign n29949 = n29948 ^ n25917 ^ n4281 ;
  assign n29950 = ( ~n15314 & n29946 ) | ( ~n15314 & n29949 ) | ( n29946 & n29949 ) ;
  assign n29951 = n3929 ^ n798 ^ 1'b0 ;
  assign n29952 = ( x18 & n15085 ) | ( x18 & n29951 ) | ( n15085 & n29951 ) ;
  assign n29953 = ( n3087 & n22510 ) | ( n3087 & ~n29952 ) | ( n22510 & ~n29952 ) ;
  assign n29954 = n29953 ^ n5634 ^ 1'b0 ;
  assign n29955 = ( n16977 & ~n22355 ) | ( n16977 & n29954 ) | ( ~n22355 & n29954 ) ;
  assign n29956 = ( n1250 & n13234 ) | ( n1250 & ~n13326 ) | ( n13234 & ~n13326 ) ;
  assign n29957 = n8547 | n22353 ;
  assign n29958 = n29956 & ~n29957 ;
  assign n29959 = n19436 ^ n17070 ^ n4347 ;
  assign n29960 = ( ~n6178 & n29958 ) | ( ~n6178 & n29959 ) | ( n29958 & n29959 ) ;
  assign n29961 = n27271 ^ n18334 ^ n17849 ;
  assign n29962 = ( ~n2425 & n19626 ) | ( ~n2425 & n21698 ) | ( n19626 & n21698 ) ;
  assign n29963 = n29962 ^ n4047 ^ n3355 ;
  assign n29964 = ( ~n272 & n3967 ) | ( ~n272 & n29963 ) | ( n3967 & n29963 ) ;
  assign n29965 = ( n2216 & n17637 ) | ( n2216 & n29964 ) | ( n17637 & n29964 ) ;
  assign n29966 = ( n2244 & ~n19050 ) | ( n2244 & n20858 ) | ( ~n19050 & n20858 ) ;
  assign n29967 = ~n315 & n8800 ;
  assign n29968 = ( n2869 & n16348 ) | ( n2869 & ~n29967 ) | ( n16348 & ~n29967 ) ;
  assign n29969 = ( n5164 & ~n25247 ) | ( n5164 & n26896 ) | ( ~n25247 & n26896 ) ;
  assign n29970 = ( n853 & n4537 ) | ( n853 & n9530 ) | ( n4537 & n9530 ) ;
  assign n29971 = n26112 ^ n20066 ^ n12263 ;
  assign n29972 = n29970 & ~n29971 ;
  assign n29973 = ~n16465 & n29972 ;
  assign n29974 = n5673 & ~n14266 ;
  assign n29975 = ~n21963 & n29974 ;
  assign n29976 = n1129 | n29975 ;
  assign n29977 = n29976 ^ n19409 ^ 1'b0 ;
  assign n29978 = n29977 ^ n13128 ^ n3721 ;
  assign n29979 = ( n1064 & n7086 ) | ( n1064 & ~n15339 ) | ( n7086 & ~n15339 ) ;
  assign n29980 = ( n19956 & ~n29936 ) | ( n19956 & n29979 ) | ( ~n29936 & n29979 ) ;
  assign n29981 = n5014 & n29980 ;
  assign n29982 = n23763 ^ n4239 ^ 1'b0 ;
  assign n29983 = n29982 ^ n18370 ^ n12725 ;
  assign n29985 = n26280 ^ n10718 ^ 1'b0 ;
  assign n29984 = ( n981 & n15729 ) | ( n981 & ~n21587 ) | ( n15729 & ~n21587 ) ;
  assign n29986 = n29985 ^ n29984 ^ 1'b0 ;
  assign n29990 = ( ~n7654 & n9393 ) | ( ~n7654 & n24016 ) | ( n9393 & n24016 ) ;
  assign n29989 = ( n3978 & n10129 ) | ( n3978 & ~n22174 ) | ( n10129 & ~n22174 ) ;
  assign n29987 = n993 | n14257 ;
  assign n29988 = n24161 & ~n29987 ;
  assign n29991 = n29990 ^ n29989 ^ n29988 ;
  assign n29992 = n10777 ^ n4408 ^ 1'b0 ;
  assign n29993 = n23346 ^ n5885 ^ n3807 ;
  assign n29994 = ( n2147 & ~n6341 ) | ( n2147 & n24137 ) | ( ~n6341 & n24137 ) ;
  assign n29995 = ( n21804 & n24771 ) | ( n21804 & n29994 ) | ( n24771 & n29994 ) ;
  assign n29996 = n1233 | n29995 ;
  assign n29997 = n28655 & ~n29996 ;
  assign n29998 = ( n29992 & n29993 ) | ( n29992 & ~n29997 ) | ( n29993 & ~n29997 ) ;
  assign n29999 = n10184 & ~n14645 ;
  assign n30000 = n29999 ^ n24711 ^ 1'b0 ;
  assign n30001 = n30000 ^ n25428 ^ n21086 ;
  assign n30002 = ( n3631 & n20501 ) | ( n3631 & ~n29062 ) | ( n20501 & ~n29062 ) ;
  assign n30003 = ( n9857 & n30001 ) | ( n9857 & ~n30002 ) | ( n30001 & ~n30002 ) ;
  assign n30004 = ( n5274 & n6410 ) | ( n5274 & n15198 ) | ( n6410 & n15198 ) ;
  assign n30005 = ( n1751 & ~n9306 ) | ( n1751 & n30004 ) | ( ~n9306 & n30004 ) ;
  assign n30006 = n10711 ^ n3174 ^ 1'b0 ;
  assign n30007 = ( ~n25298 & n30005 ) | ( ~n25298 & n30006 ) | ( n30005 & n30006 ) ;
  assign n30008 = n30007 ^ n1179 ^ 1'b0 ;
  assign n30009 = ( n10463 & ~n18913 ) | ( n10463 & n30008 ) | ( ~n18913 & n30008 ) ;
  assign n30010 = ( n8896 & n15902 ) | ( n8896 & ~n23453 ) | ( n15902 & ~n23453 ) ;
  assign n30011 = n24939 | n29373 ;
  assign n30012 = ( n1838 & n3902 ) | ( n1838 & ~n7710 ) | ( n3902 & ~n7710 ) ;
  assign n30013 = n30012 ^ n1926 ^ 1'b0 ;
  assign n30014 = ( ~n13374 & n18496 ) | ( ~n13374 & n23139 ) | ( n18496 & n23139 ) ;
  assign n30015 = n8457 ^ n2973 ^ 1'b0 ;
  assign n30016 = n3672 & ~n30015 ;
  assign n30017 = ( n8856 & ~n15568 ) | ( n8856 & n30016 ) | ( ~n15568 & n30016 ) ;
  assign n30018 = ( n7320 & n15762 ) | ( n7320 & n25793 ) | ( n15762 & n25793 ) ;
  assign n30019 = ( ~n30014 & n30017 ) | ( ~n30014 & n30018 ) | ( n30017 & n30018 ) ;
  assign n30020 = n10004 ^ n9786 ^ 1'b0 ;
  assign n30021 = ( n995 & n17423 ) | ( n995 & n30020 ) | ( n17423 & n30020 ) ;
  assign n30022 = ( n3547 & n13163 ) | ( n3547 & ~n30021 ) | ( n13163 & ~n30021 ) ;
  assign n30023 = ( n6408 & n26957 ) | ( n6408 & n29251 ) | ( n26957 & n29251 ) ;
  assign n30025 = n17478 ^ n2830 ^ 1'b0 ;
  assign n30026 = n11720 | n30025 ;
  assign n30024 = ( n8839 & n19078 ) | ( n8839 & n21895 ) | ( n19078 & n21895 ) ;
  assign n30027 = n30026 ^ n30024 ^ n10079 ;
  assign n30028 = ( n7125 & n8765 ) | ( n7125 & n30027 ) | ( n8765 & n30027 ) ;
  assign n30030 = n4168 & ~n20911 ;
  assign n30031 = n30030 ^ n6141 ^ 1'b0 ;
  assign n30029 = ( n7877 & n12774 ) | ( n7877 & n13856 ) | ( n12774 & n13856 ) ;
  assign n30032 = n30031 ^ n30029 ^ n19221 ;
  assign n30033 = n4526 ^ n2174 ^ x23 ;
  assign n30034 = ( n3477 & n22159 ) | ( n3477 & ~n30033 ) | ( n22159 & ~n30033 ) ;
  assign n30035 = ( ~n1903 & n22623 ) | ( ~n1903 & n30034 ) | ( n22623 & n30034 ) ;
  assign n30036 = ~n4783 & n30035 ;
  assign n30037 = n30036 ^ n23156 ^ 1'b0 ;
  assign n30040 = ( n5247 & n7376 ) | ( n5247 & ~n22242 ) | ( n7376 & ~n22242 ) ;
  assign n30041 = ( n14075 & n22411 ) | ( n14075 & n30040 ) | ( n22411 & n30040 ) ;
  assign n30038 = n26683 ^ n11822 ^ n5053 ;
  assign n30039 = ( n1046 & n7029 ) | ( n1046 & n30038 ) | ( n7029 & n30038 ) ;
  assign n30042 = n30041 ^ n30039 ^ n11609 ;
  assign n30043 = ( n7468 & ~n14310 ) | ( n7468 & n20668 ) | ( ~n14310 & n20668 ) ;
  assign n30044 = n30043 ^ n23210 ^ n6292 ;
  assign n30045 = n26160 ^ n22327 ^ n2892 ;
  assign n30046 = ( n593 & ~n7180 ) | ( n593 & n30045 ) | ( ~n7180 & n30045 ) ;
  assign n30047 = ( n25989 & ~n29462 ) | ( n25989 & n30046 ) | ( ~n29462 & n30046 ) ;
  assign n30048 = n14468 ^ n4062 ^ n1776 ;
  assign n30049 = n30048 ^ n23388 ^ n5157 ;
  assign n30050 = n30049 ^ n29752 ^ n4773 ;
  assign n30051 = n30050 ^ n16204 ^ n6582 ;
  assign n30052 = n15379 ^ n13516 ^ n3363 ;
  assign n30053 = n26756 & ~n30052 ;
  assign n30054 = n30053 ^ n13344 ^ 1'b0 ;
  assign n30055 = ( n1807 & n3587 ) | ( n1807 & n29336 ) | ( n3587 & n29336 ) ;
  assign n30056 = n30055 ^ n26326 ^ n3860 ;
  assign n30057 = ( n1263 & ~n10100 ) | ( n1263 & n20507 ) | ( ~n10100 & n20507 ) ;
  assign n30058 = n30057 ^ n14520 ^ n12111 ;
  assign n30059 = ( ~n18155 & n25532 ) | ( ~n18155 & n30058 ) | ( n25532 & n30058 ) ;
  assign n30060 = n30056 & n30059 ;
  assign n30061 = n22229 & n30060 ;
  assign n30062 = ( n494 & ~n3097 ) | ( n494 & n14368 ) | ( ~n3097 & n14368 ) ;
  assign n30063 = n26917 ^ n18576 ^ n4765 ;
  assign n30064 = ( n8338 & ~n23815 ) | ( n8338 & n30063 ) | ( ~n23815 & n30063 ) ;
  assign n30065 = ( x240 & n1112 ) | ( x240 & n11685 ) | ( n1112 & n11685 ) ;
  assign n30066 = ( n30062 & n30064 ) | ( n30062 & ~n30065 ) | ( n30064 & ~n30065 ) ;
  assign n30067 = ( ~n1847 & n12474 ) | ( ~n1847 & n29797 ) | ( n12474 & n29797 ) ;
  assign n30068 = n26472 ^ n10140 ^ n1142 ;
  assign n30069 = ( n12897 & ~n17805 ) | ( n12897 & n30068 ) | ( ~n17805 & n30068 ) ;
  assign n30070 = ( n10752 & n15475 ) | ( n10752 & n17636 ) | ( n15475 & n17636 ) ;
  assign n30071 = ( n11647 & n28981 ) | ( n11647 & n30070 ) | ( n28981 & n30070 ) ;
  assign n30072 = n30071 ^ n4921 ^ n2957 ;
  assign n30073 = ~n922 & n4540 ;
  assign n30074 = n30073 ^ n20512 ^ 1'b0 ;
  assign n30075 = ( n7527 & ~n18599 ) | ( n7527 & n26467 ) | ( ~n18599 & n26467 ) ;
  assign n30076 = n29847 ^ n12847 ^ n8158 ;
  assign n30078 = n1291 & ~n7071 ;
  assign n30077 = n6857 ^ n3667 ^ n409 ;
  assign n30079 = n30078 ^ n30077 ^ n1467 ;
  assign n30080 = ( n14113 & n16330 ) | ( n14113 & n26075 ) | ( n16330 & n26075 ) ;
  assign n30081 = n30080 ^ n6292 ^ x159 ;
  assign n30082 = ( n5500 & n30079 ) | ( n5500 & ~n30081 ) | ( n30079 & ~n30081 ) ;
  assign n30083 = n13605 ^ n8994 ^ n6351 ;
  assign n30084 = n30083 ^ n5322 ^ n1608 ;
  assign n30085 = n653 & ~n3714 ;
  assign n30086 = n30085 ^ n5497 ^ 1'b0 ;
  assign n30087 = n30086 ^ n6316 ^ x150 ;
  assign n30088 = n17753 ^ n16603 ^ 1'b0 ;
  assign n30089 = n30087 & ~n30088 ;
  assign n30090 = n5139 | n21362 ;
  assign n30091 = n23150 | n26601 ;
  assign n30092 = n30090 & ~n30091 ;
  assign n30093 = n8056 ^ n6399 ^ n464 ;
  assign n30094 = n14791 ^ n4166 ^ 1'b0 ;
  assign n30095 = n30093 & n30094 ;
  assign n30096 = n30095 ^ n29516 ^ n6407 ;
  assign n30097 = n3598 ^ n2444 ^ x9 ;
  assign n30098 = n8207 & n30097 ;
  assign n30099 = ( n9311 & n12506 ) | ( n9311 & ~n19075 ) | ( n12506 & ~n19075 ) ;
  assign n30100 = ~n11116 & n30099 ;
  assign n30101 = n11961 ^ n7570 ^ n1656 ;
  assign n30102 = ~n11811 & n20986 ;
  assign n30103 = n30102 ^ n10903 ^ 1'b0 ;
  assign n30104 = ( n3921 & n11348 ) | ( n3921 & ~n14810 ) | ( n11348 & ~n14810 ) ;
  assign n30105 = n12018 ^ n7163 ^ n6796 ;
  assign n30106 = ( ~n9593 & n26032 ) | ( ~n9593 & n30105 ) | ( n26032 & n30105 ) ;
  assign n30107 = n15301 ^ n9283 ^ n4710 ;
  assign n30108 = n4558 & ~n14518 ;
  assign n30109 = n30108 ^ n29691 ^ 1'b0 ;
  assign n30110 = n24540 | n30109 ;
  assign n30111 = n30107 & ~n30110 ;
  assign n30112 = ( ~n10131 & n22382 ) | ( ~n10131 & n30111 ) | ( n22382 & n30111 ) ;
  assign n30122 = n8689 ^ n898 ^ 1'b0 ;
  assign n30115 = ( x46 & n625 ) | ( x46 & n3785 ) | ( n625 & n3785 ) ;
  assign n30114 = n23670 ^ n13802 ^ n7104 ;
  assign n30116 = n30115 ^ n30114 ^ n10796 ;
  assign n30117 = n9890 & n11570 ;
  assign n30118 = n30116 & n30117 ;
  assign n30119 = n30118 ^ n25877 ^ n14913 ;
  assign n30113 = ( n4586 & ~n19502 ) | ( n4586 & n23982 ) | ( ~n19502 & n23982 ) ;
  assign n30120 = n30119 ^ n30113 ^ n3022 ;
  assign n30121 = n17720 & ~n30120 ;
  assign n30123 = n30122 ^ n30121 ^ 1'b0 ;
  assign n30124 = n5510 ^ n5394 ^ 1'b0 ;
  assign n30125 = n30124 ^ n11711 ^ n688 ;
  assign n30126 = n30125 ^ n26695 ^ n13428 ;
  assign n30127 = ( n10302 & n11183 ) | ( n10302 & n20796 ) | ( n11183 & n20796 ) ;
  assign n30128 = n18564 ^ n12569 ^ n2940 ;
  assign n30129 = ( ~n1259 & n3939 ) | ( ~n1259 & n30128 ) | ( n3939 & n30128 ) ;
  assign n30130 = ( n1009 & n2759 ) | ( n1009 & n30129 ) | ( n2759 & n30129 ) ;
  assign n30131 = n16865 ^ n11794 ^ n3674 ;
  assign n30132 = n30131 ^ n14273 ^ x114 ;
  assign n30133 = x134 & n26081 ;
  assign n30134 = n30133 ^ n22565 ^ 1'b0 ;
  assign n30135 = ( n8845 & n26351 ) | ( n8845 & n28194 ) | ( n26351 & n28194 ) ;
  assign n30136 = n30135 ^ n27327 ^ n14803 ;
  assign n30137 = n8663 ^ n8546 ^ n1618 ;
  assign n30138 = ( n262 & ~n4699 ) | ( n262 & n9795 ) | ( ~n4699 & n9795 ) ;
  assign n30139 = n11746 ^ n7165 ^ 1'b0 ;
  assign n30140 = ~n22249 & n30139 ;
  assign n30141 = n30140 ^ n9348 ^ 1'b0 ;
  assign n30142 = ( n2604 & n7573 ) | ( n2604 & ~n8734 ) | ( n7573 & ~n8734 ) ;
  assign n30143 = ( n3119 & n5799 ) | ( n3119 & n25681 ) | ( n5799 & n25681 ) ;
  assign n30144 = n30143 ^ n17865 ^ n2834 ;
  assign n30145 = ( n12776 & n30142 ) | ( n12776 & ~n30144 ) | ( n30142 & ~n30144 ) ;
  assign n30146 = ( n17436 & n30141 ) | ( n17436 & n30145 ) | ( n30141 & n30145 ) ;
  assign n30147 = n7141 | n28729 ;
  assign n30148 = ( n13320 & n20484 ) | ( n13320 & ~n26223 ) | ( n20484 & ~n26223 ) ;
  assign n30149 = ( n9648 & n24649 ) | ( n9648 & n30148 ) | ( n24649 & n30148 ) ;
  assign n30150 = ( ~n4760 & n7227 ) | ( ~n4760 & n9661 ) | ( n7227 & n9661 ) ;
  assign n30151 = n30150 ^ n24324 ^ n3592 ;
  assign n30152 = n14421 ^ n10797 ^ n5384 ;
  assign n30153 = ( ~n6295 & n22771 ) | ( ~n6295 & n30152 ) | ( n22771 & n30152 ) ;
  assign n30154 = ( n6750 & n10719 ) | ( n6750 & ~n22424 ) | ( n10719 & ~n22424 ) ;
  assign n30155 = ( ~n1208 & n20901 ) | ( ~n1208 & n29485 ) | ( n20901 & n29485 ) ;
  assign n30156 = ( n10598 & ~n14034 ) | ( n10598 & n30155 ) | ( ~n14034 & n30155 ) ;
  assign n30157 = n8727 & n18498 ;
  assign n30158 = n30157 ^ n5189 ^ 1'b0 ;
  assign n30159 = n30158 ^ n18480 ^ n4783 ;
  assign n30160 = n25764 ^ n1953 ^ 1'b0 ;
  assign n30161 = n6627 ^ n4759 ^ 1'b0 ;
  assign n30162 = ~n21705 & n30161 ;
  assign n30163 = n30162 ^ n22951 ^ n7224 ;
  assign n30164 = ~n14598 & n24330 ;
  assign n30165 = ~n18955 & n30164 ;
  assign n30166 = ( n26209 & n30163 ) | ( n26209 & n30165 ) | ( n30163 & n30165 ) ;
  assign n30167 = n3670 & n22970 ;
  assign n30168 = n30167 ^ n8348 ^ 1'b0 ;
  assign n30171 = n24076 ^ n2843 ^ n807 ;
  assign n30172 = ( n11314 & ~n16076 ) | ( n11314 & n30171 ) | ( ~n16076 & n30171 ) ;
  assign n30169 = n11918 ^ n4562 ^ n1314 ;
  assign n30170 = ( n2800 & n21452 ) | ( n2800 & n30169 ) | ( n21452 & n30169 ) ;
  assign n30173 = n30172 ^ n30170 ^ n1002 ;
  assign n30174 = n30173 ^ n29474 ^ n5384 ;
  assign n30175 = n1266 & n23382 ;
  assign n30176 = n30175 ^ n18583 ^ n9781 ;
  assign n30177 = n24904 ^ n3747 ^ 1'b0 ;
  assign n30178 = ~n1815 & n30177 ;
  assign n30179 = n29303 & n30178 ;
  assign n30180 = n29905 ^ n16086 ^ n14642 ;
  assign n30181 = n30180 ^ n29763 ^ n27405 ;
  assign n30182 = n13098 ^ n1189 ^ 1'b0 ;
  assign n30183 = n4865 | n30182 ;
  assign n30184 = ( n512 & n9283 ) | ( n512 & n30183 ) | ( n9283 & n30183 ) ;
  assign n30185 = n24087 | n29993 ;
  assign n30186 = n8408 ^ n446 ^ 1'b0 ;
  assign n30187 = n23283 | n30186 ;
  assign n30188 = n30185 | n30187 ;
  assign n30189 = ( ~n3993 & n5425 ) | ( ~n3993 & n25884 ) | ( n5425 & n25884 ) ;
  assign n30190 = n27472 ^ n15346 ^ n10978 ;
  assign n30191 = ~n17182 & n18148 ;
  assign n30192 = n30190 & n30191 ;
  assign n30193 = n30192 ^ n27914 ^ n17479 ;
  assign n30194 = n9975 | n27201 ;
  assign n30195 = n30194 ^ n12690 ^ 1'b0 ;
  assign n30196 = n17084 ^ n11487 ^ n7910 ;
  assign n30197 = n30196 ^ n28505 ^ n19271 ;
  assign n30198 = ( n6317 & n14813 ) | ( n6317 & n30197 ) | ( n14813 & n30197 ) ;
  assign n30199 = ( n13108 & n30195 ) | ( n13108 & n30198 ) | ( n30195 & n30198 ) ;
  assign n30200 = ~n851 & n7197 ;
  assign n30201 = n25681 ^ n11882 ^ n7919 ;
  assign n30202 = ~n30200 & n30201 ;
  assign n30203 = n30202 ^ n7819 ^ 1'b0 ;
  assign n30204 = n30203 ^ n8258 ^ 1'b0 ;
  assign n30205 = ( n1507 & n2197 ) | ( n1507 & n25325 ) | ( n2197 & n25325 ) ;
  assign n30206 = ( n15070 & n24400 ) | ( n15070 & n30205 ) | ( n24400 & n30205 ) ;
  assign n30207 = n22638 ^ n19527 ^ n17400 ;
  assign n30208 = ( n7686 & n13345 ) | ( n7686 & n30207 ) | ( n13345 & n30207 ) ;
  assign n30210 = ( n1724 & ~n7629 ) | ( n1724 & n12356 ) | ( ~n7629 & n12356 ) ;
  assign n30211 = n30210 ^ n24224 ^ n16365 ;
  assign n30209 = n29333 ^ n21865 ^ 1'b0 ;
  assign n30212 = n30211 ^ n30209 ^ n17237 ;
  assign n30218 = ( ~n3802 & n4581 ) | ( ~n3802 & n22256 ) | ( n4581 & n22256 ) ;
  assign n30213 = n11318 ^ n522 ^ 1'b0 ;
  assign n30214 = n5031 & n30213 ;
  assign n30215 = ( n542 & n17149 ) | ( n542 & n30214 ) | ( n17149 & n30214 ) ;
  assign n30216 = n20982 ^ n379 ^ 1'b0 ;
  assign n30217 = n30215 & n30216 ;
  assign n30219 = n30218 ^ n30217 ^ n258 ;
  assign n30220 = n15481 ^ n9877 ^ n6600 ;
  assign n30221 = ( n4560 & n8633 ) | ( n4560 & ~n30220 ) | ( n8633 & ~n30220 ) ;
  assign n30222 = ~n20524 & n30221 ;
  assign n30223 = n30222 ^ n9627 ^ 1'b0 ;
  assign n30224 = n14877 & ~n30223 ;
  assign n30225 = n30224 ^ n23329 ^ 1'b0 ;
  assign n30226 = ( n11325 & ~n18624 ) | ( n11325 & n28138 ) | ( ~n18624 & n28138 ) ;
  assign n30227 = ( ~n18663 & n19397 ) | ( ~n18663 & n30226 ) | ( n19397 & n30226 ) ;
  assign n30228 = n30227 ^ n15868 ^ 1'b0 ;
  assign n30229 = n24054 ^ n12377 ^ 1'b0 ;
  assign n30230 = ~n23466 & n30229 ;
  assign n30231 = n30230 ^ n24054 ^ n17054 ;
  assign n30232 = n2782 & ~n23349 ;
  assign n30233 = n30232 ^ n22540 ^ 1'b0 ;
  assign n30234 = ( n6751 & n12073 ) | ( n6751 & ~n19000 ) | ( n12073 & ~n19000 ) ;
  assign n30235 = ~n2833 & n15919 ;
  assign n30236 = n30235 ^ n19584 ^ 1'b0 ;
  assign n30237 = n792 | n18494 ;
  assign n30238 = n30237 ^ n1523 ^ 1'b0 ;
  assign n30239 = ( ~n12992 & n30236 ) | ( ~n12992 & n30238 ) | ( n30236 & n30238 ) ;
  assign n30240 = n30239 ^ n13407 ^ n1042 ;
  assign n30241 = n30240 ^ n13113 ^ n12822 ;
  assign n30242 = n15451 & ~n29281 ;
  assign n30243 = n17226 | n17491 ;
  assign n30244 = n2568 | n30243 ;
  assign n30245 = n28798 ^ n23520 ^ n21925 ;
  assign n30246 = ( n8810 & ~n24274 ) | ( n8810 & n25110 ) | ( ~n24274 & n25110 ) ;
  assign n30247 = n6820 & n22866 ;
  assign n30248 = ~n7659 & n30247 ;
  assign n30249 = ( ~n10238 & n26826 ) | ( ~n10238 & n30248 ) | ( n26826 & n30248 ) ;
  assign n30250 = ( n1541 & ~n7941 ) | ( n1541 & n10122 ) | ( ~n7941 & n10122 ) ;
  assign n30251 = n30250 ^ n22734 ^ n17121 ;
  assign n30252 = ( n6724 & n7671 ) | ( n6724 & ~n18010 ) | ( n7671 & ~n18010 ) ;
  assign n30253 = ( n10104 & ~n16196 ) | ( n10104 & n30252 ) | ( ~n16196 & n30252 ) ;
  assign n30254 = n2372 & n11402 ;
  assign n30255 = ( n6041 & ~n12448 ) | ( n6041 & n30254 ) | ( ~n12448 & n30254 ) ;
  assign n30256 = ~n16401 & n30255 ;
  assign n30257 = n30256 ^ n26485 ^ 1'b0 ;
  assign n30258 = n1811 & ~n17675 ;
  assign n30259 = n27265 & n30258 ;
  assign n30263 = n17079 ^ n10147 ^ n1231 ;
  assign n30260 = n20524 ^ n2935 ^ x224 ;
  assign n30261 = n30260 ^ n29520 ^ n2499 ;
  assign n30262 = ( n12254 & ~n14992 ) | ( n12254 & n30261 ) | ( ~n14992 & n30261 ) ;
  assign n30264 = n30263 ^ n30262 ^ 1'b0 ;
  assign n30265 = x94 & ~n19714 ;
  assign n30266 = ( n5020 & n27703 ) | ( n5020 & n30265 ) | ( n27703 & n30265 ) ;
  assign n30268 = n22522 ^ n4073 ^ n1285 ;
  assign n30267 = ~n9880 & n19062 ;
  assign n30269 = n30268 ^ n30267 ^ n18452 ;
  assign n30270 = n7015 ^ x149 ^ 1'b0 ;
  assign n30271 = n4077 & n29784 ;
  assign n30272 = n22638 ^ n5227 ^ n3066 ;
  assign n30273 = n24798 ^ n22975 ^ n4506 ;
  assign n30274 = n2586 ^ n1635 ^ 1'b0 ;
  assign n30275 = n2738 & n30274 ;
  assign n30276 = ~n8887 & n10576 ;
  assign n30277 = n30276 ^ n14187 ^ 1'b0 ;
  assign n30278 = n835 & n3039 ;
  assign n30279 = n30278 ^ n2046 ^ n556 ;
  assign n30280 = ( n3949 & ~n21302 ) | ( n3949 & n30279 ) | ( ~n21302 & n30279 ) ;
  assign n30281 = ( n27641 & n30277 ) | ( n27641 & n30280 ) | ( n30277 & n30280 ) ;
  assign n30282 = ( n3884 & ~n5462 ) | ( n3884 & n20175 ) | ( ~n5462 & n20175 ) ;
  assign n30283 = ( n22517 & n23290 ) | ( n22517 & ~n29401 ) | ( n23290 & ~n29401 ) ;
  assign n30284 = ( n9884 & ~n12986 ) | ( n9884 & n13003 ) | ( ~n12986 & n13003 ) ;
  assign n30285 = ( n7562 & n13430 ) | ( n7562 & ~n24675 ) | ( n13430 & ~n24675 ) ;
  assign n30286 = ( n3498 & n7362 ) | ( n3498 & ~n19391 ) | ( n7362 & ~n19391 ) ;
  assign n30287 = ( n30284 & n30285 ) | ( n30284 & ~n30286 ) | ( n30285 & ~n30286 ) ;
  assign n30288 = n22735 ^ n21775 ^ n15425 ;
  assign n30289 = ( ~n2629 & n30040 ) | ( ~n2629 & n30288 ) | ( n30040 & n30288 ) ;
  assign n30290 = ( n2992 & ~n11207 ) | ( n2992 & n27046 ) | ( ~n11207 & n27046 ) ;
  assign n30291 = n30290 ^ n6681 ^ 1'b0 ;
  assign n30292 = n8517 ^ n5998 ^ n5024 ;
  assign n30293 = n30292 ^ n7146 ^ n3636 ;
  assign n30294 = ( n2677 & n14509 ) | ( n2677 & n30293 ) | ( n14509 & n30293 ) ;
  assign n30295 = n30294 ^ n9988 ^ 1'b0 ;
  assign n30296 = n11924 | n12356 ;
  assign n30297 = n30296 ^ n2472 ^ 1'b0 ;
  assign n30298 = ~n26667 & n27352 ;
  assign n30299 = ~n15673 & n30298 ;
  assign n30300 = n30299 ^ n6024 ^ n2910 ;
  assign n30301 = n30300 ^ n18644 ^ n1926 ;
  assign n30302 = n5982 & n15187 ;
  assign n30303 = ( ~n3957 & n14455 ) | ( ~n3957 & n23150 ) | ( n14455 & n23150 ) ;
  assign n30304 = ( n3138 & n30302 ) | ( n3138 & ~n30303 ) | ( n30302 & ~n30303 ) ;
  assign n30305 = n28015 ^ n24355 ^ n1761 ;
  assign n30306 = n30305 ^ n25845 ^ 1'b0 ;
  assign n30307 = ( n9129 & n14755 ) | ( n9129 & ~n15925 ) | ( n14755 & ~n15925 ) ;
  assign n30308 = ~n14853 & n20172 ;
  assign n30309 = n30308 ^ n17916 ^ n14304 ;
  assign n30311 = ( ~n4437 & n7984 ) | ( ~n4437 & n12859 ) | ( n7984 & n12859 ) ;
  assign n30310 = n14088 ^ n13712 ^ n1537 ;
  assign n30312 = n30311 ^ n30310 ^ n15880 ;
  assign n30313 = n2865 | n30312 ;
  assign n30315 = n1332 & n6898 ;
  assign n30314 = n4395 | n9372 ;
  assign n30316 = n30315 ^ n30314 ^ 1'b0 ;
  assign n30317 = ( n11722 & n19896 ) | ( n11722 & n30316 ) | ( n19896 & n30316 ) ;
  assign n30318 = n9090 | n23283 ;
  assign n30319 = n30318 ^ n25487 ^ 1'b0 ;
  assign n30320 = n10166 | n18638 ;
  assign n30321 = n21479 ^ n19029 ^ n2408 ;
  assign n30322 = ( n12151 & n12966 ) | ( n12151 & ~n30321 ) | ( n12966 & ~n30321 ) ;
  assign n30323 = n11135 ^ n2692 ^ 1'b0 ;
  assign n30324 = n11484 | n30323 ;
  assign n30325 = n30324 ^ n17518 ^ x55 ;
  assign n30326 = ( ~n6111 & n30322 ) | ( ~n6111 & n30325 ) | ( n30322 & n30325 ) ;
  assign n30327 = ( n12151 & n26124 ) | ( n12151 & ~n30326 ) | ( n26124 & ~n30326 ) ;
  assign n30328 = n10656 & ~n18771 ;
  assign n30329 = ( n1780 & n2568 ) | ( n1780 & ~n8466 ) | ( n2568 & ~n8466 ) ;
  assign n30330 = n30329 ^ n13205 ^ n3231 ;
  assign n30331 = n16443 ^ n14470 ^ x159 ;
  assign n30333 = ( n8744 & n14307 ) | ( n8744 & ~n18813 ) | ( n14307 & ~n18813 ) ;
  assign n30332 = n15855 ^ n566 ^ 1'b0 ;
  assign n30334 = n30333 ^ n30332 ^ 1'b0 ;
  assign n30335 = ~n15325 & n30334 ;
  assign n30336 = ~n30331 & n30335 ;
  assign n30339 = n4960 ^ n3960 ^ n1822 ;
  assign n30340 = ( n5007 & n10260 ) | ( n5007 & n30339 ) | ( n10260 & n30339 ) ;
  assign n30341 = n30340 ^ n6177 ^ n1301 ;
  assign n30342 = ( ~n2568 & n27469 ) | ( ~n2568 & n30341 ) | ( n27469 & n30341 ) ;
  assign n30337 = n28762 ^ n10733 ^ n1249 ;
  assign n30338 = n30337 ^ n11666 ^ n1130 ;
  assign n30343 = n30342 ^ n30338 ^ n21973 ;
  assign n30344 = n22307 ^ n21930 ^ n1824 ;
  assign n30345 = n19625 ^ n15843 ^ 1'b0 ;
  assign n30346 = n20037 ^ n19494 ^ n6366 ;
  assign n30347 = ( n12254 & ~n30345 ) | ( n12254 & n30346 ) | ( ~n30345 & n30346 ) ;
  assign n30348 = n11361 ^ n3516 ^ 1'b0 ;
  assign n30349 = ~n27979 & n30348 ;
  assign n30356 = n28591 ^ n27788 ^ 1'b0 ;
  assign n30350 = ( n5015 & n23935 ) | ( n5015 & n27851 ) | ( n23935 & n27851 ) ;
  assign n30351 = ( n4036 & ~n10035 ) | ( n4036 & n12934 ) | ( ~n10035 & n12934 ) ;
  assign n30352 = n30351 ^ n8986 ^ 1'b0 ;
  assign n30353 = n19511 | n29731 ;
  assign n30354 = n30352 | n30353 ;
  assign n30355 = ( n8918 & n30350 ) | ( n8918 & n30354 ) | ( n30350 & n30354 ) ;
  assign n30357 = n30356 ^ n30355 ^ n4898 ;
  assign n30358 = n20748 ^ n18453 ^ 1'b0 ;
  assign n30359 = ( n9517 & n21038 ) | ( n9517 & n30358 ) | ( n21038 & n30358 ) ;
  assign n30360 = ~n10149 & n30359 ;
  assign n30361 = n6745 ^ n2599 ^ 1'b0 ;
  assign n30362 = n21457 & n30361 ;
  assign n30363 = ( ~n2759 & n16018 ) | ( ~n2759 & n30362 ) | ( n16018 & n30362 ) ;
  assign n30364 = n11193 ^ n6171 ^ 1'b0 ;
  assign n30365 = n30364 ^ n14437 ^ n4272 ;
  assign n30366 = n1905 & ~n20629 ;
  assign n30367 = n9401 & ~n30366 ;
  assign n30368 = n15981 ^ n4565 ^ 1'b0 ;
  assign n30369 = n5083 | n30368 ;
  assign n30370 = n422 & n6565 ;
  assign n30371 = n30370 ^ n4381 ^ 1'b0 ;
  assign n30372 = ~n30369 & n30371 ;
  assign n30373 = n22527 & ~n22562 ;
  assign n30374 = ~n30372 & n30373 ;
  assign n30375 = n8053 | n8876 ;
  assign n30377 = ~n5034 & n17874 ;
  assign n30376 = n12505 & n13441 ;
  assign n30378 = n30377 ^ n30376 ^ 1'b0 ;
  assign n30379 = ( ~n4851 & n6171 ) | ( ~n4851 & n17877 ) | ( n6171 & n17877 ) ;
  assign n30380 = ( n5890 & n23429 ) | ( n5890 & ~n30379 ) | ( n23429 & ~n30379 ) ;
  assign n30381 = n30378 | n30380 ;
  assign n30382 = n18644 & ~n30381 ;
  assign n30388 = ( n3872 & n9548 ) | ( n3872 & n19450 ) | ( n9548 & n19450 ) ;
  assign n30383 = n22603 ^ n9473 ^ 1'b0 ;
  assign n30384 = ( n4934 & n12306 ) | ( n4934 & n17513 ) | ( n12306 & n17513 ) ;
  assign n30385 = ( n10039 & n30383 ) | ( n10039 & n30384 ) | ( n30383 & n30384 ) ;
  assign n30386 = ( n5496 & ~n7881 ) | ( n5496 & n30385 ) | ( ~n7881 & n30385 ) ;
  assign n30387 = ( n937 & n19360 ) | ( n937 & n30386 ) | ( n19360 & n30386 ) ;
  assign n30389 = n30388 ^ n30387 ^ n2312 ;
  assign n30391 = n20026 ^ n11962 ^ n7338 ;
  assign n30392 = ( n3853 & n4179 ) | ( n3853 & n30391 ) | ( n4179 & n30391 ) ;
  assign n30390 = n6850 & n25021 ;
  assign n30393 = n30392 ^ n30390 ^ 1'b0 ;
  assign n30394 = n24109 ^ n23651 ^ n881 ;
  assign n30395 = ( n14902 & ~n30393 ) | ( n14902 & n30394 ) | ( ~n30393 & n30394 ) ;
  assign n30396 = n20210 & ~n28136 ;
  assign n30397 = n14257 | n16979 ;
  assign n30398 = ( n7596 & n20062 ) | ( n7596 & ~n27262 ) | ( n20062 & ~n27262 ) ;
  assign n30399 = n30398 ^ n19998 ^ 1'b0 ;
  assign n30400 = ~n18212 & n22630 ;
  assign n30401 = n16327 ^ n8399 ^ 1'b0 ;
  assign n30402 = ~n10790 & n30401 ;
  assign n30403 = ~n30400 & n30402 ;
  assign n30404 = n30403 ^ n22031 ^ n2775 ;
  assign n30405 = ( ~n2845 & n4571 ) | ( ~n2845 & n8160 ) | ( n4571 & n8160 ) ;
  assign n30406 = n30405 ^ n18917 ^ 1'b0 ;
  assign n30410 = ( n2858 & ~n3720 ) | ( n2858 & n6647 ) | ( ~n3720 & n6647 ) ;
  assign n30411 = n30410 ^ n12592 ^ 1'b0 ;
  assign n30412 = n9022 & ~n30411 ;
  assign n30407 = ( n7104 & ~n9907 ) | ( n7104 & n23305 ) | ( ~n9907 & n23305 ) ;
  assign n30408 = n30407 ^ n8285 ^ n2499 ;
  assign n30409 = n9102 & ~n30408 ;
  assign n30413 = n30412 ^ n30409 ^ 1'b0 ;
  assign n30414 = n425 & n5260 ;
  assign n30415 = n18271 & n30414 ;
  assign n30416 = n30415 ^ n29811 ^ n17879 ;
  assign n30419 = n26057 ^ n3562 ^ 1'b0 ;
  assign n30417 = ( n9598 & n16672 ) | ( n9598 & n24483 ) | ( n16672 & n24483 ) ;
  assign n30418 = n30417 ^ n28776 ^ n14309 ;
  assign n30420 = n30419 ^ n30418 ^ n28062 ;
  assign n30421 = n14423 ^ n4554 ^ n1236 ;
  assign n30422 = ~n20055 & n21213 ;
  assign n30423 = n2555 & n30422 ;
  assign n30424 = ( n11341 & ~n30421 ) | ( n11341 & n30423 ) | ( ~n30421 & n30423 ) ;
  assign n30425 = ~n14581 & n15472 ;
  assign n30426 = ~n12996 & n30425 ;
  assign n30427 = ( ~n6882 & n30424 ) | ( ~n6882 & n30426 ) | ( n30424 & n30426 ) ;
  assign n30428 = n14605 & n21002 ;
  assign n30429 = n3334 & n30428 ;
  assign n30430 = ( n1783 & n10357 ) | ( n1783 & ~n30429 ) | ( n10357 & ~n30429 ) ;
  assign n30434 = ( n5764 & n5893 ) | ( n5764 & n24723 ) | ( n5893 & n24723 ) ;
  assign n30435 = ( n9380 & n9813 ) | ( n9380 & n30434 ) | ( n9813 & n30434 ) ;
  assign n30432 = n20026 ^ n7956 ^ n396 ;
  assign n30433 = n30432 ^ n25794 ^ n8194 ;
  assign n30431 = n12882 ^ n3222 ^ n1088 ;
  assign n30436 = n30435 ^ n30433 ^ n30431 ;
  assign n30437 = ( n795 & n19749 ) | ( n795 & ~n30436 ) | ( n19749 & ~n30436 ) ;
  assign n30438 = n6965 & ~n30437 ;
  assign n30439 = ~n12308 & n30438 ;
  assign n30440 = ( ~n11572 & n15766 ) | ( ~n11572 & n19135 ) | ( n15766 & n19135 ) ;
  assign n30441 = n19888 ^ n8225 ^ n8102 ;
  assign n30442 = ( n13766 & ~n28022 ) | ( n13766 & n30441 ) | ( ~n28022 & n30441 ) ;
  assign n30443 = ( ~n623 & n11022 ) | ( ~n623 & n22226 ) | ( n11022 & n22226 ) ;
  assign n30444 = n30443 ^ n17703 ^ 1'b0 ;
  assign n30445 = ~n16377 & n30444 ;
  assign n30446 = n8107 & ~n30445 ;
  assign n30447 = ( n4016 & n30442 ) | ( n4016 & n30446 ) | ( n30442 & n30446 ) ;
  assign n30448 = n14337 & ~n21400 ;
  assign n30451 = ( n1363 & n8319 ) | ( n1363 & n8724 ) | ( n8319 & n8724 ) ;
  assign n30449 = ( n14130 & n16342 ) | ( n14130 & n25266 ) | ( n16342 & n25266 ) ;
  assign n30450 = n30449 ^ n19737 ^ n6346 ;
  assign n30452 = n30451 ^ n30450 ^ n24224 ;
  assign n30454 = n15710 ^ n8249 ^ n3413 ;
  assign n30455 = n30454 ^ n24521 ^ n16364 ;
  assign n30453 = n5340 & n13624 ;
  assign n30456 = n30455 ^ n30453 ^ 1'b0 ;
  assign n30457 = n8460 | n10077 ;
  assign n30458 = n1582 & ~n30457 ;
  assign n30459 = n28528 ^ n19299 ^ n15671 ;
  assign n30460 = ( n6021 & n12852 ) | ( n6021 & ~n30005 ) | ( n12852 & ~n30005 ) ;
  assign n30461 = ( n20122 & n30459 ) | ( n20122 & ~n30460 ) | ( n30459 & ~n30460 ) ;
  assign n30463 = ( x208 & ~n7938 ) | ( x208 & n23579 ) | ( ~n7938 & n23579 ) ;
  assign n30464 = n16326 | n18351 ;
  assign n30465 = n30463 & ~n30464 ;
  assign n30462 = n28124 ^ n17556 ^ n5997 ;
  assign n30466 = n30465 ^ n30462 ^ 1'b0 ;
  assign n30467 = n12851 & n15066 ;
  assign n30468 = ~n16209 & n30467 ;
  assign n30469 = n30308 & n30468 ;
  assign n30470 = ( n7856 & ~n14466 ) | ( n7856 & n30469 ) | ( ~n14466 & n30469 ) ;
  assign n30472 = n14967 ^ n5337 ^ n2539 ;
  assign n30473 = ~n6834 & n16951 ;
  assign n30474 = n30472 & n30473 ;
  assign n30471 = n5881 & n19783 ;
  assign n30475 = n30474 ^ n30471 ^ n3752 ;
  assign n30477 = n14776 | n14951 ;
  assign n30478 = n259 | n30477 ;
  assign n30476 = n9569 ^ n8180 ^ n7457 ;
  assign n30479 = n30478 ^ n30476 ^ n23765 ;
  assign n30480 = n13003 ^ n9539 ^ n7046 ;
  assign n30481 = n29278 ^ n24495 ^ 1'b0 ;
  assign n30483 = n1105 & n6926 ;
  assign n30482 = ( n3027 & n11758 ) | ( n3027 & n25404 ) | ( n11758 & n25404 ) ;
  assign n30484 = n30483 ^ n30482 ^ n23147 ;
  assign n30487 = ( n2566 & ~n12070 ) | ( n2566 & n24137 ) | ( ~n12070 & n24137 ) ;
  assign n30485 = x143 | n17283 ;
  assign n30486 = n30255 | n30485 ;
  assign n30488 = n30487 ^ n30486 ^ n14746 ;
  assign n30489 = ( n4504 & n5453 ) | ( n4504 & ~n9748 ) | ( n5453 & ~n9748 ) ;
  assign n30492 = ( ~n8386 & n20349 ) | ( ~n8386 & n25368 ) | ( n20349 & n25368 ) ;
  assign n30490 = n7516 ^ n1496 ^ n914 ;
  assign n30491 = ( ~n10668 & n24266 ) | ( ~n10668 & n30490 ) | ( n24266 & n30490 ) ;
  assign n30493 = n30492 ^ n30491 ^ n30465 ;
  assign n30494 = ~n21183 & n30493 ;
  assign n30495 = ( n5967 & n6302 ) | ( n5967 & ~n10381 ) | ( n6302 & ~n10381 ) ;
  assign n30496 = n18579 | n30495 ;
  assign n30497 = n30496 ^ n15574 ^ 1'b0 ;
  assign n30501 = ( n4704 & n9425 ) | ( n4704 & n17583 ) | ( n9425 & n17583 ) ;
  assign n30498 = n19894 ^ n14155 ^ n8442 ;
  assign n30499 = ( n3110 & n6958 ) | ( n3110 & ~n26272 ) | ( n6958 & ~n26272 ) ;
  assign n30500 = n30498 | n30499 ;
  assign n30502 = n30501 ^ n30500 ^ 1'b0 ;
  assign n30503 = n11676 & n29643 ;
  assign n30504 = ~n27184 & n30503 ;
  assign n30505 = n17468 ^ n9307 ^ n5924 ;
  assign n30506 = ( n16344 & n29309 ) | ( n16344 & n30505 ) | ( n29309 & n30505 ) ;
  assign n30507 = ( x204 & n2479 ) | ( x204 & ~n6304 ) | ( n2479 & ~n6304 ) ;
  assign n30508 = ( ~n1708 & n15813 ) | ( ~n1708 & n30507 ) | ( n15813 & n30507 ) ;
  assign n30509 = ( ~n8157 & n8316 ) | ( ~n8157 & n30508 ) | ( n8316 & n30508 ) ;
  assign n30510 = n3045 & ~n8205 ;
  assign n30511 = n30510 ^ n16634 ^ n4378 ;
  assign n30512 = n30511 ^ n11822 ^ n8760 ;
  assign n30513 = ( n5634 & ~n10182 ) | ( n5634 & n11385 ) | ( ~n10182 & n11385 ) ;
  assign n30514 = n30513 ^ n19883 ^ n436 ;
  assign n30515 = n13284 & n27461 ;
  assign n30516 = n15020 & n30515 ;
  assign n30517 = n12240 ^ n2404 ^ 1'b0 ;
  assign n30518 = n30517 ^ n29910 ^ n14124 ;
  assign n30519 = n11165 | n19640 ;
  assign n30520 = ( ~n7547 & n24095 ) | ( ~n7547 & n30519 ) | ( n24095 & n30519 ) ;
  assign n30521 = ( ~n3262 & n10504 ) | ( ~n3262 & n12101 ) | ( n10504 & n12101 ) ;
  assign n30522 = n30521 ^ n19677 ^ n7991 ;
  assign n30523 = n11591 ^ n8179 ^ 1'b0 ;
  assign n30524 = ~n7029 & n30523 ;
  assign n30525 = ( n8668 & n20166 ) | ( n8668 & ~n30524 ) | ( n20166 & ~n30524 ) ;
  assign n30526 = ( n5149 & n14968 ) | ( n5149 & ~n30525 ) | ( n14968 & ~n30525 ) ;
  assign n30527 = ( ~n11691 & n30522 ) | ( ~n11691 & n30526 ) | ( n30522 & n30526 ) ;
  assign n30528 = n25608 ^ n21552 ^ n757 ;
  assign n30529 = ( ~n9270 & n18583 ) | ( ~n9270 & n30528 ) | ( n18583 & n30528 ) ;
  assign n30530 = n24967 ^ n10979 ^ n6278 ;
  assign n30531 = ~n10747 & n10996 ;
  assign n30532 = ~n18879 & n30531 ;
  assign n30533 = n16442 ^ n4667 ^ n1954 ;
  assign n30534 = n22050 ^ n15550 ^ 1'b0 ;
  assign n30535 = ( ~n13783 & n30533 ) | ( ~n13783 & n30534 ) | ( n30533 & n30534 ) ;
  assign n30536 = ( n4246 & n10029 ) | ( n4246 & ~n24100 ) | ( n10029 & ~n24100 ) ;
  assign n30537 = n4718 & n30536 ;
  assign n30538 = n26198 ^ n23919 ^ n16708 ;
  assign n30539 = ~n2218 & n5684 ;
  assign n30540 = n30539 ^ n6497 ^ n947 ;
  assign n30541 = n27759 ^ n1489 ^ 1'b0 ;
  assign n30542 = n17099 | n30541 ;
  assign n30543 = n5452 & ~n17899 ;
  assign n30544 = ( n611 & n2032 ) | ( n611 & n7723 ) | ( n2032 & n7723 ) ;
  assign n30545 = ( n4906 & n13843 ) | ( n4906 & ~n30544 ) | ( n13843 & ~n30544 ) ;
  assign n30547 = n7640 & ~n29409 ;
  assign n30548 = n30547 ^ n12425 ^ 1'b0 ;
  assign n30546 = n23317 ^ n11838 ^ n10900 ;
  assign n30549 = n30548 ^ n30546 ^ n21780 ;
  assign n30550 = n15613 ^ n5221 ^ 1'b0 ;
  assign n30551 = ( n15649 & n18713 ) | ( n15649 & n30550 ) | ( n18713 & n30550 ) ;
  assign n30552 = n8408 & ~n13521 ;
  assign n30553 = n30552 ^ n12704 ^ 1'b0 ;
  assign n30554 = n6141 ^ n3669 ^ x172 ;
  assign n30555 = ( ~n11499 & n14401 ) | ( ~n11499 & n30554 ) | ( n14401 & n30554 ) ;
  assign n30556 = ( n1166 & n2970 ) | ( n1166 & ~n20029 ) | ( n2970 & ~n20029 ) ;
  assign n30557 = n30556 ^ n4233 ^ n1731 ;
  assign n30558 = ( n5066 & n30495 ) | ( n5066 & n30557 ) | ( n30495 & n30557 ) ;
  assign n30559 = n28265 ^ n8727 ^ n2768 ;
  assign n30560 = n30559 ^ n29683 ^ n15353 ;
  assign n30563 = ( n2561 & n10014 ) | ( n2561 & ~n13318 ) | ( n10014 & ~n13318 ) ;
  assign n30564 = n24386 | n30563 ;
  assign n30565 = n7856 | n30564 ;
  assign n30561 = ( n5241 & n11543 ) | ( n5241 & n25624 ) | ( n11543 & n25624 ) ;
  assign n30562 = ( ~n19177 & n25320 ) | ( ~n19177 & n30561 ) | ( n25320 & n30561 ) ;
  assign n30566 = n30565 ^ n30562 ^ n22323 ;
  assign n30568 = n12470 ^ n1334 ^ 1'b0 ;
  assign n30569 = n30568 ^ n5795 ^ n2174 ;
  assign n30567 = n2074 | n5977 ;
  assign n30570 = n30569 ^ n30567 ^ 1'b0 ;
  assign n30571 = n20215 ^ n6591 ^ 1'b0 ;
  assign n30572 = ~n19647 & n30571 ;
  assign n30573 = ( n10599 & n11230 ) | ( n10599 & ~n12089 ) | ( n11230 & ~n12089 ) ;
  assign n30574 = n28868 ^ n3873 ^ 1'b0 ;
  assign n30575 = n30574 ^ n20923 ^ n9005 ;
  assign n30576 = ( n23993 & ~n30573 ) | ( n23993 & n30575 ) | ( ~n30573 & n30575 ) ;
  assign n30577 = n14458 ^ n9392 ^ 1'b0 ;
  assign n30578 = n16123 & ~n30577 ;
  assign n30579 = n30578 ^ n7241 ^ n3822 ;
  assign n30580 = n12573 & ~n12821 ;
  assign n30581 = ( n22245 & n29062 ) | ( n22245 & ~n30400 ) | ( n29062 & ~n30400 ) ;
  assign n30582 = ( ~n623 & n4720 ) | ( ~n623 & n13967 ) | ( n4720 & n13967 ) ;
  assign n30583 = n30582 ^ n22036 ^ n6787 ;
  assign n30584 = n26250 & ~n30304 ;
  assign n30585 = n30584 ^ n10186 ^ 1'b0 ;
  assign n30586 = n12171 ^ n9519 ^ 1'b0 ;
  assign n30587 = n15274 & ~n30586 ;
  assign n30588 = ( n3380 & ~n7885 ) | ( n3380 & n15840 ) | ( ~n7885 & n15840 ) ;
  assign n30589 = n11796 & n30588 ;
  assign n30590 = ( n16025 & n30587 ) | ( n16025 & n30589 ) | ( n30587 & n30589 ) ;
  assign n30591 = ( n4121 & n25837 ) | ( n4121 & ~n27758 ) | ( n25837 & ~n27758 ) ;
  assign n30592 = n30591 ^ n19490 ^ n5942 ;
  assign n30596 = ( n2724 & n10171 ) | ( n2724 & n14240 ) | ( n10171 & n14240 ) ;
  assign n30595 = n26130 ^ n16846 ^ n9912 ;
  assign n30597 = n30596 ^ n30595 ^ n13599 ;
  assign n30593 = n19849 & ~n29156 ;
  assign n30594 = n30593 ^ n6485 ^ 1'b0 ;
  assign n30598 = n30597 ^ n30594 ^ 1'b0 ;
  assign n30599 = n12760 ^ n9753 ^ x50 ;
  assign n30600 = ( ~n15024 & n21871 ) | ( ~n15024 & n30599 ) | ( n21871 & n30599 ) ;
  assign n30601 = n2615 | n7387 ;
  assign n30602 = ~n889 & n30601 ;
  assign n30603 = n30602 ^ n25091 ^ 1'b0 ;
  assign n30604 = ( n1730 & n4187 ) | ( n1730 & ~n9174 ) | ( n4187 & ~n9174 ) ;
  assign n30605 = n30604 ^ n8872 ^ n5104 ;
  assign n30606 = n22873 ^ n6051 ^ n3950 ;
  assign n30607 = n30606 ^ n19559 ^ n18699 ;
  assign n30608 = n22527 ^ n18243 ^ 1'b0 ;
  assign n30609 = ( n15207 & ~n28132 ) | ( n15207 & n30608 ) | ( ~n28132 & n30608 ) ;
  assign n30610 = n30607 & ~n30609 ;
  assign n30611 = ( ~n12802 & n13113 ) | ( ~n12802 & n16972 ) | ( n13113 & n16972 ) ;
  assign n30612 = n12645 ^ n8205 ^ n1777 ;
  assign n30613 = n30612 ^ n9410 ^ n5971 ;
  assign n30614 = ( ~n3380 & n15714 ) | ( ~n3380 & n30613 ) | ( n15714 & n30613 ) ;
  assign n30615 = ( ~n12394 & n17304 ) | ( ~n12394 & n21044 ) | ( n17304 & n21044 ) ;
  assign n30616 = ( n10811 & n27283 ) | ( n10811 & n30615 ) | ( n27283 & n30615 ) ;
  assign n30617 = n5925 ^ n3204 ^ 1'b0 ;
  assign n30618 = ~n30616 & n30617 ;
  assign n30619 = n30618 ^ n16613 ^ n4581 ;
  assign n30620 = ( ~n10775 & n24205 ) | ( ~n10775 & n30619 ) | ( n24205 & n30619 ) ;
  assign n30621 = ( n9881 & ~n19114 ) | ( n9881 & n22069 ) | ( ~n19114 & n22069 ) ;
  assign n30623 = n25541 ^ n4547 ^ n1190 ;
  assign n30622 = ( ~n7141 & n13152 ) | ( ~n7141 & n16382 ) | ( n13152 & n16382 ) ;
  assign n30624 = n30623 ^ n30622 ^ 1'b0 ;
  assign n30625 = n1703 & ~n30624 ;
  assign n30626 = n8315 ^ n3333 ^ 1'b0 ;
  assign n30627 = ( n13291 & n30625 ) | ( n13291 & n30626 ) | ( n30625 & n30626 ) ;
  assign n30628 = n20223 ^ n14910 ^ n393 ;
  assign n30629 = n17380 ^ n1723 ^ 1'b0 ;
  assign n30630 = n30628 & ~n30629 ;
  assign n30631 = ( n12278 & n14361 ) | ( n12278 & n30630 ) | ( n14361 & n30630 ) ;
  assign n30632 = ~n30627 & n30631 ;
  assign n30633 = ~n30621 & n30632 ;
  assign n30634 = n2773 | n16597 ;
  assign n30635 = n21112 | n30634 ;
  assign n30636 = n26712 ^ n8339 ^ n2358 ;
  assign n30639 = ( n5844 & n9371 ) | ( n5844 & n22912 ) | ( n9371 & n22912 ) ;
  assign n30640 = ( ~n2615 & n24573 ) | ( ~n2615 & n30639 ) | ( n24573 & n30639 ) ;
  assign n30637 = ( n1787 & n8445 ) | ( n1787 & ~n15780 ) | ( n8445 & ~n15780 ) ;
  assign n30638 = ( n2927 & n30310 ) | ( n2927 & ~n30637 ) | ( n30310 & ~n30637 ) ;
  assign n30641 = n30640 ^ n30638 ^ n12141 ;
  assign n30642 = n995 | n17226 ;
  assign n30643 = ( n1734 & ~n1765 ) | ( n1734 & n4989 ) | ( ~n1765 & n4989 ) ;
  assign n30644 = n25514 ^ n21629 ^ 1'b0 ;
  assign n30645 = n30643 & ~n30644 ;
  assign n30646 = ( n14723 & ~n30642 ) | ( n14723 & n30645 ) | ( ~n30642 & n30645 ) ;
  assign n30647 = ( n746 & n18097 ) | ( n746 & ~n21649 ) | ( n18097 & ~n21649 ) ;
  assign n30649 = ( n414 & n4073 ) | ( n414 & ~n5056 ) | ( n4073 & ~n5056 ) ;
  assign n30650 = ( ~n487 & n4443 ) | ( ~n487 & n7034 ) | ( n4443 & n7034 ) ;
  assign n30651 = ( n19810 & n30649 ) | ( n19810 & n30650 ) | ( n30649 & n30650 ) ;
  assign n30652 = n30651 ^ n29840 ^ n19950 ;
  assign n30648 = n12480 ^ n10871 ^ n822 ;
  assign n30653 = n30652 ^ n30648 ^ n16990 ;
  assign n30654 = n18790 ^ n10250 ^ n8485 ;
  assign n30655 = n30654 ^ n21430 ^ n3001 ;
  assign n30656 = n30655 ^ n29206 ^ n17530 ;
  assign n30657 = n27390 ^ n17544 ^ n3224 ;
  assign n30659 = n10446 & n14595 ;
  assign n30660 = n30659 ^ n20380 ^ 1'b0 ;
  assign n30658 = n8820 ^ n7252 ^ n3085 ;
  assign n30661 = n30660 ^ n30658 ^ 1'b0 ;
  assign n30662 = n22833 ^ n14376 ^ n3176 ;
  assign n30663 = n30662 ^ n27177 ^ n6212 ;
  assign n30664 = ~n2344 & n29754 ;
  assign n30665 = n30664 ^ n4919 ^ 1'b0 ;
  assign n30666 = n30665 ^ n14159 ^ n7949 ;
  assign n30667 = n3262 ^ n2595 ^ 1'b0 ;
  assign n30668 = n30667 ^ n29432 ^ n18942 ;
  assign n30670 = n30421 ^ n15169 ^ n12610 ;
  assign n30669 = ( n3757 & n3959 ) | ( n3757 & ~n25439 ) | ( n3959 & ~n25439 ) ;
  assign n30671 = n30670 ^ n30669 ^ n10672 ;
  assign n30674 = n7903 & n9685 ;
  assign n30672 = n24291 | n26449 ;
  assign n30673 = n28249 & ~n30672 ;
  assign n30675 = n30674 ^ n30673 ^ n4322 ;
  assign n30676 = n7492 & n11391 ;
  assign n30677 = n11035 & n30676 ;
  assign n30678 = n19360 & ~n30677 ;
  assign n30679 = ~n7804 & n30678 ;
  assign n30680 = ( n3044 & ~n15829 ) | ( n3044 & n20743 ) | ( ~n15829 & n20743 ) ;
  assign n30681 = n30680 ^ n15936 ^ 1'b0 ;
  assign n30682 = n30681 ^ n24839 ^ n19756 ;
  assign n30683 = ( n17508 & n23469 ) | ( n17508 & n29123 ) | ( n23469 & n29123 ) ;
  assign n30685 = n7870 ^ n4158 ^ n1729 ;
  assign n30686 = ~n14596 & n30685 ;
  assign n30687 = n30686 ^ n12104 ^ 1'b0 ;
  assign n30684 = n22540 ^ n6784 ^ n3683 ;
  assign n30688 = n30687 ^ n30684 ^ n20464 ;
  assign n30693 = n11645 ^ n1207 ^ 1'b0 ;
  assign n30694 = ( n552 & n13951 ) | ( n552 & ~n30693 ) | ( n13951 & ~n30693 ) ;
  assign n30689 = n11977 & ~n13390 ;
  assign n30690 = ~n20359 & n30689 ;
  assign n30691 = n30690 ^ n23656 ^ n4651 ;
  assign n30692 = n18435 | n30691 ;
  assign n30695 = n30694 ^ n30692 ^ 1'b0 ;
  assign n30700 = n25155 ^ n13286 ^ n11463 ;
  assign n30696 = n12862 ^ n357 ^ 1'b0 ;
  assign n30697 = n30696 ^ n7576 ^ 1'b0 ;
  assign n30698 = n30697 ^ n16342 ^ n4143 ;
  assign n30699 = n5033 | n30698 ;
  assign n30701 = n30700 ^ n30699 ^ 1'b0 ;
  assign n30702 = n14104 ^ n8047 ^ 1'b0 ;
  assign n30703 = n10129 & n20493 ;
  assign n30704 = n8982 | n15705 ;
  assign n30705 = n30703 | n30704 ;
  assign n30706 = n30705 ^ n7403 ^ n2855 ;
  assign n30707 = ( n6961 & ~n8293 ) | ( n6961 & n27294 ) | ( ~n8293 & n27294 ) ;
  assign n30708 = ( n7909 & n21892 ) | ( n7909 & n30707 ) | ( n21892 & n30707 ) ;
  assign n30709 = ( n17218 & n29175 ) | ( n17218 & ~n30708 ) | ( n29175 & ~n30708 ) ;
  assign n30710 = ( n1936 & ~n6746 ) | ( n1936 & n15882 ) | ( ~n6746 & n15882 ) ;
  assign n30711 = n23185 ^ n21132 ^ n1904 ;
  assign n30712 = n1264 & ~n6138 ;
  assign n30713 = n13581 & n30712 ;
  assign n30714 = n15134 & ~n21028 ;
  assign n30715 = ~n12932 & n30714 ;
  assign n30716 = n2164 | n27789 ;
  assign n30717 = ( n313 & n15894 ) | ( n313 & n20569 ) | ( n15894 & n20569 ) ;
  assign n30718 = n30717 ^ n12990 ^ n1102 ;
  assign n30719 = n30718 ^ n26142 ^ n5436 ;
  assign n30720 = ( n4864 & ~n7862 ) | ( n4864 & n10444 ) | ( ~n7862 & n10444 ) ;
  assign n30721 = n30720 ^ n16000 ^ 1'b0 ;
  assign n30722 = n22547 ^ n1013 ^ 1'b0 ;
  assign n30723 = ( ~n3332 & n30721 ) | ( ~n3332 & n30722 ) | ( n30721 & n30722 ) ;
  assign n30724 = ( n836 & n3984 ) | ( n836 & ~n4565 ) | ( n3984 & ~n4565 ) ;
  assign n30725 = n30724 ^ n8505 ^ n4159 ;
  assign n30726 = n30725 ^ n28359 ^ n14424 ;
  assign n30741 = n25704 ^ n21222 ^ 1'b0 ;
  assign n30742 = ( n7245 & n26833 ) | ( n7245 & ~n30741 ) | ( n26833 & ~n30741 ) ;
  assign n30729 = n5708 ^ n2646 ^ 1'b0 ;
  assign n30730 = n7408 & ~n30729 ;
  assign n30731 = n23686 ^ n12760 ^ n8120 ;
  assign n30732 = ( n2134 & ~n8286 ) | ( n2134 & n12723 ) | ( ~n8286 & n12723 ) ;
  assign n30733 = n30732 ^ n8236 ^ 1'b0 ;
  assign n30734 = n12300 & ~n30733 ;
  assign n30735 = ( n2882 & n10802 ) | ( n2882 & ~n18552 ) | ( n10802 & ~n18552 ) ;
  assign n30736 = ( n6798 & n7434 ) | ( n6798 & n7822 ) | ( n7434 & n7822 ) ;
  assign n30737 = ( ~n6554 & n21682 ) | ( ~n6554 & n30736 ) | ( n21682 & n30736 ) ;
  assign n30738 = ( ~n17901 & n30735 ) | ( ~n17901 & n30737 ) | ( n30735 & n30737 ) ;
  assign n30739 = ( n19273 & n30734 ) | ( n19273 & n30738 ) | ( n30734 & n30738 ) ;
  assign n30740 = ( n30730 & ~n30731 ) | ( n30730 & n30739 ) | ( ~n30731 & n30739 ) ;
  assign n30727 = n28714 ^ n18475 ^ n1195 ;
  assign n30728 = n30727 ^ n9067 ^ n2345 ;
  assign n30743 = n30742 ^ n30740 ^ n30728 ;
  assign n30744 = ( n11593 & ~n18935 ) | ( n11593 & n21385 ) | ( ~n18935 & n21385 ) ;
  assign n30745 = n12346 ^ n3223 ^ 1'b0 ;
  assign n30746 = ~n30744 & n30745 ;
  assign n30747 = n30746 ^ n25074 ^ n9464 ;
  assign n30748 = n30747 ^ n26752 ^ 1'b0 ;
  assign n30749 = n16767 | n30748 ;
  assign n30750 = n15808 ^ n643 ^ 1'b0 ;
  assign n30751 = n27687 | n30750 ;
  assign n30752 = ( ~n3115 & n9758 ) | ( ~n3115 & n16354 ) | ( n9758 & n16354 ) ;
  assign n30753 = ( ~n2261 & n2283 ) | ( ~n2261 & n30752 ) | ( n2283 & n30752 ) ;
  assign n30754 = n30753 ^ n29209 ^ 1'b0 ;
  assign n30755 = n20958 ^ n2084 ^ 1'b0 ;
  assign n30756 = n30755 ^ n23721 ^ n16958 ;
  assign n30757 = ( n1808 & n5913 ) | ( n1808 & n8526 ) | ( n5913 & n8526 ) ;
  assign n30758 = ( n17126 & ~n28316 ) | ( n17126 & n30757 ) | ( ~n28316 & n30757 ) ;
  assign n30759 = ( ~n10516 & n12896 ) | ( ~n10516 & n30758 ) | ( n12896 & n30758 ) ;
  assign n30760 = n15943 ^ n11646 ^ n4313 ;
  assign n30761 = n20861 ^ n4908 ^ 1'b0 ;
  assign n30762 = ~n4269 & n30761 ;
  assign n30763 = n12391 & ~n18478 ;
  assign n30764 = n730 & n21349 ;
  assign n30765 = ~n1766 & n30764 ;
  assign n30766 = ( n21279 & ~n26498 ) | ( n21279 & n30765 ) | ( ~n26498 & n30765 ) ;
  assign n30767 = ( n2936 & n3309 ) | ( n2936 & n16797 ) | ( n3309 & n16797 ) ;
  assign n30768 = n16606 ^ n7593 ^ n2618 ;
  assign n30769 = ( ~n5504 & n8896 ) | ( ~n5504 & n10631 ) | ( n8896 & n10631 ) ;
  assign n30770 = n16764 | n28073 ;
  assign n30771 = n30770 ^ n18104 ^ 1'b0 ;
  assign n30772 = n22187 ^ n9370 ^ 1'b0 ;
  assign n30773 = n20983 | n30772 ;
  assign n30775 = ~n9005 & n16350 ;
  assign n30776 = ( ~n4231 & n23783 ) | ( ~n4231 & n30775 ) | ( n23783 & n30775 ) ;
  assign n30774 = ( n1891 & n7073 ) | ( n1891 & ~n16084 ) | ( n7073 & ~n16084 ) ;
  assign n30777 = n30776 ^ n30774 ^ n6559 ;
  assign n30778 = n5486 | n30777 ;
  assign n30779 = n19531 ^ n16327 ^ 1'b0 ;
  assign n30780 = n30779 ^ n25657 ^ 1'b0 ;
  assign n30781 = n7195 & ~n12279 ;
  assign n30782 = n30781 ^ n24139 ^ 1'b0 ;
  assign n30783 = n30782 ^ n4448 ^ n3067 ;
  assign n30784 = n1105 & n30783 ;
  assign n30785 = n21458 ^ n379 ^ 1'b0 ;
  assign n30786 = ( n7282 & n15839 ) | ( n7282 & ~n30785 ) | ( n15839 & ~n30785 ) ;
  assign n30787 = ( n582 & n24603 ) | ( n582 & n27246 ) | ( n24603 & n27246 ) ;
  assign n30788 = n895 & n8532 ;
  assign n30789 = n382 | n10660 ;
  assign n30790 = n30789 ^ n23643 ^ 1'b0 ;
  assign n30791 = n9085 ^ n2939 ^ 1'b0 ;
  assign n30794 = ( n2427 & n13249 ) | ( n2427 & ~n20965 ) | ( n13249 & ~n20965 ) ;
  assign n30792 = n10829 ^ n9913 ^ n2297 ;
  assign n30793 = n30792 ^ n16524 ^ n9168 ;
  assign n30795 = n30794 ^ n30793 ^ 1'b0 ;
  assign n30796 = n30601 ^ n8038 ^ n4425 ;
  assign n30797 = n30796 ^ n7363 ^ n5452 ;
  assign n30798 = n30797 ^ n7029 ^ 1'b0 ;
  assign n30799 = n14343 ^ n6037 ^ 1'b0 ;
  assign n30800 = n30799 ^ n10956 ^ n555 ;
  assign n30801 = n13492 ^ n7362 ^ x241 ;
  assign n30802 = n30801 ^ n16794 ^ n16189 ;
  assign n30803 = ( n13349 & n27960 ) | ( n13349 & n30802 ) | ( n27960 & n30802 ) ;
  assign n30804 = n11455 ^ n3368 ^ n2100 ;
  assign n30805 = ( n2154 & n5417 ) | ( n2154 & n20287 ) | ( n5417 & n20287 ) ;
  assign n30806 = ( n792 & n1491 ) | ( n792 & n7329 ) | ( n1491 & n7329 ) ;
  assign n30807 = n25729 ^ n16746 ^ n4624 ;
  assign n30808 = ( ~n1455 & n17686 ) | ( ~n1455 & n30807 ) | ( n17686 & n30807 ) ;
  assign n30809 = n30808 ^ n4512 ^ 1'b0 ;
  assign n30810 = ~n11527 & n30809 ;
  assign n30811 = n18772 ^ n4301 ^ n4188 ;
  assign n30812 = n30811 ^ n12795 ^ n6778 ;
  assign n30813 = n11926 & n30812 ;
  assign n30814 = ( n30806 & ~n30810 ) | ( n30806 & n30813 ) | ( ~n30810 & n30813 ) ;
  assign n30815 = ( n3215 & n6232 ) | ( n3215 & n7279 ) | ( n6232 & n7279 ) ;
  assign n30816 = n30815 ^ n19882 ^ n15394 ;
  assign n30817 = ~n3857 & n17992 ;
  assign n30818 = ~n2230 & n30817 ;
  assign n30819 = n30818 ^ n22066 ^ n13867 ;
  assign n30820 = n1896 & n10184 ;
  assign n30821 = n30820 ^ n1967 ^ 1'b0 ;
  assign n30822 = ~n30819 & n30821 ;
  assign n30823 = ~n4151 & n23390 ;
  assign n30824 = n8301 & n30823 ;
  assign n30825 = n30824 ^ n27055 ^ 1'b0 ;
  assign n30826 = ( n13074 & n14164 ) | ( n13074 & n15839 ) | ( n14164 & n15839 ) ;
  assign n30827 = n30826 ^ n10274 ^ 1'b0 ;
  assign n30828 = n30825 & n30827 ;
  assign n30829 = n6093 & ~n27862 ;
  assign n30830 = ( n5862 & ~n11656 ) | ( n5862 & n13266 ) | ( ~n11656 & n13266 ) ;
  assign n30831 = n30830 ^ n27237 ^ n11467 ;
  assign n30832 = ( n12215 & n14907 ) | ( n12215 & n30831 ) | ( n14907 & n30831 ) ;
  assign n30833 = ( n7810 & n10339 ) | ( n7810 & n12861 ) | ( n10339 & n12861 ) ;
  assign n30834 = ~n5575 & n23882 ;
  assign n30835 = n30833 & n30834 ;
  assign n30836 = n30835 ^ n24635 ^ 1'b0 ;
  assign n30837 = n3558 & n30836 ;
  assign n30838 = n4784 ^ n2927 ^ n785 ;
  assign n30839 = n30838 ^ n24227 ^ n7344 ;
  assign n30840 = n30839 ^ n29150 ^ 1'b0 ;
  assign n30841 = n19031 | n30840 ;
  assign n30842 = n4467 | n9803 ;
  assign n30843 = n30842 ^ n3536 ^ 1'b0 ;
  assign n30844 = n30843 ^ n22086 ^ 1'b0 ;
  assign n30845 = ( n8542 & ~n11993 ) | ( n8542 & n12350 ) | ( ~n11993 & n12350 ) ;
  assign n30846 = n30845 ^ n14340 ^ n914 ;
  assign n30847 = n30846 ^ n11948 ^ n7842 ;
  assign n30848 = n22428 ^ n17689 ^ n9676 ;
  assign n30849 = ( n2491 & ~n6933 ) | ( n2491 & n24733 ) | ( ~n6933 & n24733 ) ;
  assign n30850 = n15394 ^ n2080 ^ 1'b0 ;
  assign n30851 = ~n30849 & n30850 ;
  assign n30852 = n30851 ^ n20483 ^ 1'b0 ;
  assign n30853 = n30848 & ~n30852 ;
  assign n30854 = ( n2531 & n18840 ) | ( n2531 & n23356 ) | ( n18840 & n23356 ) ;
  assign n30855 = n16820 ^ n3689 ^ 1'b0 ;
  assign n30856 = n30854 & ~n30855 ;
  assign n30857 = n20445 ^ n19739 ^ n5898 ;
  assign n30858 = n30857 ^ n7162 ^ 1'b0 ;
  assign n30859 = n30856 & n30858 ;
  assign n30860 = n30859 ^ n13968 ^ n1233 ;
  assign n30863 = ( n1812 & n15416 ) | ( n1812 & ~n23591 ) | ( n15416 & ~n23591 ) ;
  assign n30861 = n20545 ^ n7019 ^ 1'b0 ;
  assign n30862 = n30574 & n30861 ;
  assign n30864 = n30863 ^ n30862 ^ n26392 ;
  assign n30865 = n12023 ^ n8285 ^ 1'b0 ;
  assign n30866 = n13574 | n30865 ;
  assign n30867 = n15378 ^ n9276 ^ 1'b0 ;
  assign n30868 = ~n30866 & n30867 ;
  assign n30869 = n21746 ^ n15241 ^ n10638 ;
  assign n30870 = n30869 ^ n30643 ^ n2486 ;
  assign n30871 = ( n8667 & n30868 ) | ( n8667 & ~n30870 ) | ( n30868 & ~n30870 ) ;
  assign n30872 = ( n3077 & n13879 ) | ( n3077 & n14743 ) | ( n13879 & n14743 ) ;
  assign n30873 = ( n6066 & n27062 ) | ( n6066 & ~n30872 ) | ( n27062 & ~n30872 ) ;
  assign n30874 = n1077 & ~n30873 ;
  assign n30875 = n21834 & ~n30874 ;
  assign n30882 = n11838 ^ n11037 ^ 1'b0 ;
  assign n30877 = ( n1461 & ~n5639 ) | ( n1461 & n18292 ) | ( ~n5639 & n18292 ) ;
  assign n30878 = ( n5166 & n5689 ) | ( n5166 & n20741 ) | ( n5689 & n20741 ) ;
  assign n30879 = ( ~n818 & n19477 ) | ( ~n818 & n23250 ) | ( n19477 & n23250 ) ;
  assign n30880 = ( n27447 & n30878 ) | ( n27447 & n30879 ) | ( n30878 & n30879 ) ;
  assign n30881 = ( n7807 & n30877 ) | ( n7807 & ~n30880 ) | ( n30877 & ~n30880 ) ;
  assign n30883 = n30882 ^ n30881 ^ n9454 ;
  assign n30876 = n9410 ^ n8039 ^ n2337 ;
  assign n30884 = n30883 ^ n30876 ^ n5650 ;
  assign n30885 = ( n3685 & ~n4765 ) | ( n3685 & n25015 ) | ( ~n4765 & n25015 ) ;
  assign n30886 = ( n407 & n3764 ) | ( n407 & ~n4993 ) | ( n3764 & ~n4993 ) ;
  assign n30887 = n2697 | n10845 ;
  assign n30888 = n30886 & ~n30887 ;
  assign n30889 = n30888 ^ n2138 ^ 1'b0 ;
  assign n30890 = ( n4916 & n17383 ) | ( n4916 & n30889 ) | ( n17383 & n30889 ) ;
  assign n30891 = ( ~n9912 & n13176 ) | ( ~n9912 & n30890 ) | ( n13176 & n30890 ) ;
  assign n30896 = n1326 | n7004 ;
  assign n30897 = n30896 ^ n24177 ^ n7198 ;
  assign n30892 = n3621 ^ n1889 ^ 1'b0 ;
  assign n30893 = n10941 | n30892 ;
  assign n30894 = n17378 | n30893 ;
  assign n30895 = n30894 ^ n6952 ^ 1'b0 ;
  assign n30898 = n30897 ^ n30895 ^ n20872 ;
  assign n30899 = ( n3288 & ~n4561 ) | ( n3288 & n21059 ) | ( ~n4561 & n21059 ) ;
  assign n30900 = ( n3767 & ~n3939 ) | ( n3767 & n23665 ) | ( ~n3939 & n23665 ) ;
  assign n30901 = n17577 ^ n15646 ^ 1'b0 ;
  assign n30902 = n30901 ^ n17949 ^ 1'b0 ;
  assign n30903 = n8261 & ~n30902 ;
  assign n30904 = ~n30900 & n30903 ;
  assign n30905 = n17559 ^ n15576 ^ n11099 ;
  assign n30906 = ( ~n6197 & n10998 ) | ( ~n6197 & n30905 ) | ( n10998 & n30905 ) ;
  assign n30907 = n30906 ^ n12191 ^ 1'b0 ;
  assign n30908 = n25286 ^ n23331 ^ 1'b0 ;
  assign n30909 = n30908 ^ n23503 ^ n10426 ;
  assign n30910 = n10049 ^ n7058 ^ n3491 ;
  assign n30911 = ( n3467 & n9831 ) | ( n3467 & n30910 ) | ( n9831 & n30910 ) ;
  assign n30913 = n7505 ^ n1656 ^ 1'b0 ;
  assign n30914 = n11046 & n30913 ;
  assign n30915 = n30914 ^ n21856 ^ n525 ;
  assign n30916 = ~n3132 & n3443 ;
  assign n30917 = n30916 ^ n9589 ^ 1'b0 ;
  assign n30918 = n30917 ^ n19857 ^ 1'b0 ;
  assign n30919 = ~n2443 & n30918 ;
  assign n30920 = n30915 & n30919 ;
  assign n30912 = n28635 ^ n28596 ^ n17576 ;
  assign n30921 = n30920 ^ n30912 ^ n6881 ;
  assign n30922 = ( n16790 & ~n30911 ) | ( n16790 & n30921 ) | ( ~n30911 & n30921 ) ;
  assign n30923 = n30922 ^ n6015 ^ n3380 ;
  assign n30924 = n24891 ^ n15552 ^ 1'b0 ;
  assign n30925 = ( n7417 & ~n16681 ) | ( n7417 & n27807 ) | ( ~n16681 & n27807 ) ;
  assign n30926 = ( n16610 & n19875 ) | ( n16610 & n30925 ) | ( n19875 & n30925 ) ;
  assign n30927 = ~n2723 & n4168 ;
  assign n30928 = n12846 ^ n6410 ^ 1'b0 ;
  assign n30929 = n30927 | n30928 ;
  assign n30930 = ( n4590 & n29521 ) | ( n4590 & n30929 ) | ( n29521 & n30929 ) ;
  assign n30931 = ( x177 & n1471 ) | ( x177 & ~n1824 ) | ( n1471 & ~n1824 ) ;
  assign n30932 = n1886 & n30931 ;
  assign n30933 = n30932 ^ n20041 ^ 1'b0 ;
  assign n30934 = n25630 ^ n7433 ^ n296 ;
  assign n30935 = n30934 ^ n3628 ^ 1'b0 ;
  assign n30936 = ( n10098 & n19435 ) | ( n10098 & ~n30935 ) | ( n19435 & ~n30935 ) ;
  assign n30937 = n30936 ^ n25937 ^ n2668 ;
  assign n30940 = n13163 ^ n12910 ^ n12668 ;
  assign n30938 = ( n4178 & n16068 ) | ( n4178 & ~n27548 ) | ( n16068 & ~n27548 ) ;
  assign n30939 = n30938 ^ n27655 ^ n8484 ;
  assign n30941 = n30940 ^ n30939 ^ n12269 ;
  assign n30942 = ( ~x119 & n8728 ) | ( ~x119 & n22393 ) | ( n8728 & n22393 ) ;
  assign n30943 = n15278 | n30942 ;
  assign n30944 = ( n4078 & n17371 ) | ( n4078 & ~n30943 ) | ( n17371 & ~n30943 ) ;
  assign n30945 = ( ~n6663 & n11022 ) | ( ~n6663 & n27284 ) | ( n11022 & n27284 ) ;
  assign n30946 = n5424 ^ n746 ^ 1'b0 ;
  assign n30947 = n8716 | n30946 ;
  assign n30948 = ( n1871 & n2476 ) | ( n1871 & n30947 ) | ( n2476 & n30947 ) ;
  assign n30949 = n26662 ^ n7290 ^ n577 ;
  assign n30950 = n30948 & ~n30949 ;
  assign n30951 = n16425 ^ n3269 ^ 1'b0 ;
  assign n30952 = n2939 ^ n1867 ^ n835 ;
  assign n30953 = ( ~n7590 & n11405 ) | ( ~n7590 & n30952 ) | ( n11405 & n30952 ) ;
  assign n30954 = ( ~n14130 & n23017 ) | ( ~n14130 & n30953 ) | ( n23017 & n30953 ) ;
  assign n30955 = n18593 ^ n16800 ^ n8751 ;
  assign n30956 = n30955 ^ n11218 ^ 1'b0 ;
  assign n30957 = ~n9162 & n30956 ;
  assign n30958 = n30957 ^ n11001 ^ 1'b0 ;
  assign n30959 = ~n28401 & n30958 ;
  assign n30960 = n20622 ^ n10111 ^ 1'b0 ;
  assign n30961 = n909 | n30960 ;
  assign n30963 = n13947 ^ n12857 ^ n8043 ;
  assign n30962 = n5694 | n23517 ;
  assign n30964 = n30963 ^ n30962 ^ 1'b0 ;
  assign n30965 = ( n19791 & n29142 ) | ( n19791 & n30964 ) | ( n29142 & n30964 ) ;
  assign n30966 = n30965 ^ n12470 ^ 1'b0 ;
  assign n30967 = ( n12758 & ~n15095 ) | ( n12758 & n30966 ) | ( ~n15095 & n30966 ) ;
  assign n30968 = ( ~n4697 & n14621 ) | ( ~n4697 & n20577 ) | ( n14621 & n20577 ) ;
  assign n30969 = ( ~n1102 & n14187 ) | ( ~n1102 & n30968 ) | ( n14187 & n30968 ) ;
  assign n30970 = ( n7999 & n18915 ) | ( n7999 & ~n21016 ) | ( n18915 & ~n21016 ) ;
  assign n30971 = ( n13035 & ~n25889 ) | ( n13035 & n30970 ) | ( ~n25889 & n30970 ) ;
  assign n30972 = n30815 ^ n8222 ^ 1'b0 ;
  assign n30973 = n25354 ^ n24325 ^ n4905 ;
  assign n30974 = n30973 ^ n28635 ^ n25222 ;
  assign n30975 = n30974 ^ n20626 ^ n13637 ;
  assign n30976 = n23679 | n30975 ;
  assign n30977 = n3413 | n6836 ;
  assign n30979 = n2696 & n15635 ;
  assign n30980 = n30979 ^ n6904 ^ n4795 ;
  assign n30978 = n21050 ^ n19459 ^ n7709 ;
  assign n30981 = n30980 ^ n30978 ^ n22575 ;
  assign n30982 = n23810 ^ n6559 ^ n3303 ;
  assign n30983 = ( ~n9473 & n10483 ) | ( ~n9473 & n14359 ) | ( n10483 & n14359 ) ;
  assign n30984 = n17448 ^ n17203 ^ n1228 ;
  assign n30985 = ( n23485 & n30983 ) | ( n23485 & n30984 ) | ( n30983 & n30984 ) ;
  assign n30986 = ( n3965 & ~n18074 ) | ( n3965 & n30985 ) | ( ~n18074 & n30985 ) ;
  assign n30987 = n30986 ^ n19024 ^ 1'b0 ;
  assign n30988 = ( n8827 & n17917 ) | ( n8827 & ~n30987 ) | ( n17917 & ~n30987 ) ;
  assign n30989 = n29228 ^ n22913 ^ n19594 ;
  assign n30990 = ( n26374 & n26749 ) | ( n26374 & ~n30989 ) | ( n26749 & ~n30989 ) ;
  assign n30991 = n30990 ^ n2588 ^ 1'b0 ;
  assign n30992 = n15469 | n20547 ;
  assign n30993 = n21205 ^ n1830 ^ 1'b0 ;
  assign n30994 = n18433 | n30993 ;
  assign n30995 = n30994 ^ n12290 ^ n7876 ;
  assign n30996 = n21711 ^ n13921 ^ n1470 ;
  assign n30997 = n30996 ^ n15474 ^ n11378 ;
  assign n30998 = n30997 ^ n2247 ^ 1'b0 ;
  assign n30999 = n30995 & ~n30998 ;
  assign n31002 = n20718 ^ n7946 ^ n1766 ;
  assign n31003 = ( n8973 & n22732 ) | ( n8973 & n31002 ) | ( n22732 & n31002 ) ;
  assign n31004 = ( n1430 & n24049 ) | ( n1430 & n31003 ) | ( n24049 & n31003 ) ;
  assign n31000 = n29282 ^ n10873 ^ n8201 ;
  assign n31001 = n16800 & ~n31000 ;
  assign n31005 = n31004 ^ n31001 ^ 1'b0 ;
  assign n31006 = ( n1025 & n8045 ) | ( n1025 & ~n13493 ) | ( n8045 & ~n13493 ) ;
  assign n31007 = n31006 ^ x205 ^ 1'b0 ;
  assign n31008 = n24350 ^ n2558 ^ n1282 ;
  assign n31009 = ( n7596 & n16809 ) | ( n7596 & n27015 ) | ( n16809 & n27015 ) ;
  assign n31010 = n8789 & n11229 ;
  assign n31011 = n12904 & ~n14780 ;
  assign n31012 = ( n11995 & n31010 ) | ( n11995 & n31011 ) | ( n31010 & n31011 ) ;
  assign n31013 = n26212 ^ n24526 ^ n12957 ;
  assign n31014 = ( n1814 & ~n24942 ) | ( n1814 & n31013 ) | ( ~n24942 & n31013 ) ;
  assign n31015 = n31014 ^ n21840 ^ 1'b0 ;
  assign n31016 = ( n1182 & n1224 ) | ( n1182 & ~n8140 ) | ( n1224 & ~n8140 ) ;
  assign n31017 = ( n9899 & n25777 ) | ( n9899 & n31016 ) | ( n25777 & n31016 ) ;
  assign n31018 = n397 & n31017 ;
  assign n31019 = n31018 ^ n15391 ^ n7840 ;
  assign n31022 = n25795 ^ n24094 ^ 1'b0 ;
  assign n31023 = n15008 & ~n31022 ;
  assign n31020 = ( n6283 & n25011 ) | ( n6283 & n27159 ) | ( n25011 & n27159 ) ;
  assign n31021 = n31020 ^ n22922 ^ 1'b0 ;
  assign n31024 = n31023 ^ n31021 ^ n29415 ;
  assign n31025 = ~n11438 & n16911 ;
  assign n31026 = ~n6583 & n31025 ;
  assign n31027 = n31026 ^ n1846 ^ 1'b0 ;
  assign n31028 = n30505 ^ n22320 ^ 1'b0 ;
  assign n31029 = n18672 & n31028 ;
  assign n31030 = ( n25263 & ~n29596 ) | ( n25263 & n31029 ) | ( ~n29596 & n31029 ) ;
  assign n31031 = n2933 ^ n2129 ^ x209 ;
  assign n31032 = n13994 ^ n3235 ^ 1'b0 ;
  assign n31033 = n31031 & ~n31032 ;
  assign n31036 = n14007 ^ n7061 ^ n1753 ;
  assign n31034 = ( n2844 & ~n11372 ) | ( n2844 & n19593 ) | ( ~n11372 & n19593 ) ;
  assign n31035 = n17305 & n31034 ;
  assign n31037 = n31036 ^ n31035 ^ 1'b0 ;
  assign n31038 = n15092 & ~n31037 ;
  assign n31039 = ( n3253 & n7522 ) | ( n3253 & ~n31038 ) | ( n7522 & ~n31038 ) ;
  assign n31040 = ( ~n20619 & n26716 ) | ( ~n20619 & n31039 ) | ( n26716 & n31039 ) ;
  assign n31043 = n998 | n1609 ;
  assign n31044 = n31043 ^ n12679 ^ n1025 ;
  assign n31045 = ( n12456 & n26000 ) | ( n12456 & n31044 ) | ( n26000 & n31044 ) ;
  assign n31041 = n14012 ^ n11704 ^ n954 ;
  assign n31042 = n31041 ^ n25541 ^ n11163 ;
  assign n31046 = n31045 ^ n31042 ^ n20053 ;
  assign n31047 = n16280 ^ n11014 ^ n4421 ;
  assign n31048 = ( n12092 & ~n16366 ) | ( n12092 & n31047 ) | ( ~n16366 & n31047 ) ;
  assign n31049 = ( n9730 & n10214 ) | ( n9730 & ~n31048 ) | ( n10214 & ~n31048 ) ;
  assign n31050 = ( ~n8302 & n11999 ) | ( ~n8302 & n12000 ) | ( n11999 & n12000 ) ;
  assign n31051 = n31050 ^ n12367 ^ n6733 ;
  assign n31052 = n27020 ^ n26526 ^ 1'b0 ;
  assign n31053 = ( ~n28151 & n31051 ) | ( ~n28151 & n31052 ) | ( n31051 & n31052 ) ;
  assign n31054 = n27921 ^ n8829 ^ 1'b0 ;
  assign n31055 = ~n14613 & n15191 ;
  assign n31056 = ~n31054 & n31055 ;
  assign n31057 = ( ~n1174 & n9443 ) | ( ~n1174 & n10595 ) | ( n9443 & n10595 ) ;
  assign n31058 = n31057 ^ n3597 ^ 1'b0 ;
  assign n31059 = ( ~n26823 & n31056 ) | ( ~n26823 & n31058 ) | ( n31056 & n31058 ) ;
  assign n31060 = n18754 ^ n8613 ^ 1'b0 ;
  assign n31061 = n1686 & ~n31060 ;
  assign n31062 = ( n3322 & n9639 ) | ( n3322 & n31061 ) | ( n9639 & n31061 ) ;
  assign n31063 = ( n3728 & n26073 ) | ( n3728 & ~n31062 ) | ( n26073 & ~n31062 ) ;
  assign n31064 = n31063 ^ n28448 ^ n16455 ;
  assign n31065 = n12645 | n28724 ;
  assign n31066 = n11988 | n31065 ;
  assign n31067 = ~n14775 & n29925 ;
  assign n31068 = ~n15182 & n18580 ;
  assign n31069 = ~n31067 & n31068 ;
  assign n31070 = n20892 ^ n2812 ^ 1'b0 ;
  assign n31071 = n31070 ^ n7933 ^ 1'b0 ;
  assign n31072 = n31071 ^ n13891 ^ n5278 ;
  assign n31073 = ( n9732 & n22820 ) | ( n9732 & ~n31072 ) | ( n22820 & ~n31072 ) ;
  assign n31074 = n8951 ^ n629 ^ 1'b0 ;
  assign n31075 = ( n10755 & n11794 ) | ( n10755 & n31074 ) | ( n11794 & n31074 ) ;
  assign n31076 = ( n2952 & n6157 ) | ( n2952 & n6710 ) | ( n6157 & n6710 ) ;
  assign n31077 = ( n8336 & n19369 ) | ( n8336 & n31076 ) | ( n19369 & n31076 ) ;
  assign n31078 = n7723 ^ n5433 ^ 1'b0 ;
  assign n31079 = n31077 | n31078 ;
  assign n31080 = ( n15368 & n26013 ) | ( n15368 & n26124 ) | ( n26013 & n26124 ) ;
  assign n31081 = ( n957 & n2447 ) | ( n957 & n31080 ) | ( n2447 & n31080 ) ;
  assign n31082 = ( n31075 & n31079 ) | ( n31075 & ~n31081 ) | ( n31079 & ~n31081 ) ;
  assign n31083 = n27354 ^ n12420 ^ 1'b0 ;
  assign n31084 = n27321 | n31083 ;
  assign n31085 = n31084 ^ n30856 ^ 1'b0 ;
  assign n31086 = n31085 ^ n5910 ^ n1106 ;
  assign n31087 = n4643 & n5277 ;
  assign n31088 = n27243 & n31087 ;
  assign n31095 = ~n1591 & n6189 ;
  assign n31091 = n26907 ^ n9143 ^ 1'b0 ;
  assign n31092 = n10426 & ~n31091 ;
  assign n31093 = ( n16006 & n16533 ) | ( n16006 & ~n23218 ) | ( n16533 & ~n23218 ) ;
  assign n31094 = ( n27528 & n31092 ) | ( n27528 & n31093 ) | ( n31092 & n31093 ) ;
  assign n31096 = n31095 ^ n31094 ^ n14912 ;
  assign n31089 = n27238 ^ n12245 ^ n1851 ;
  assign n31090 = ( n13077 & n23459 ) | ( n13077 & n31089 ) | ( n23459 & n31089 ) ;
  assign n31097 = n31096 ^ n31090 ^ n1361 ;
  assign n31098 = n12232 ^ n8867 ^ 1'b0 ;
  assign n31099 = n31098 ^ n13207 ^ n5673 ;
  assign n31100 = n28830 ^ n27510 ^ n12899 ;
  assign n31101 = ( n24355 & n24969 ) | ( n24355 & ~n25437 ) | ( n24969 & ~n25437 ) ;
  assign n31102 = ~n13496 & n17234 ;
  assign n31103 = ~n31101 & n31102 ;
  assign n31107 = n9153 ^ n3242 ^ n2789 ;
  assign n31108 = n10950 & n31107 ;
  assign n31109 = n31108 ^ n3331 ^ 1'b0 ;
  assign n31104 = n29719 ^ n22576 ^ 1'b0 ;
  assign n31105 = n27123 & ~n31104 ;
  assign n31106 = ( n13841 & n18541 ) | ( n13841 & ~n31105 ) | ( n18541 & ~n31105 ) ;
  assign n31110 = n31109 ^ n31106 ^ n3625 ;
  assign n31111 = ~n1588 & n23119 ;
  assign n31112 = n31111 ^ n9111 ^ n2234 ;
  assign n31113 = n31112 ^ n16256 ^ n14892 ;
  assign n31114 = ( ~n2224 & n7797 ) | ( ~n2224 & n15693 ) | ( n7797 & n15693 ) ;
  assign n31115 = n31114 ^ n30793 ^ n4321 ;
  assign n31116 = n31115 ^ n14267 ^ n4557 ;
  assign n31118 = n4407 & n12685 ;
  assign n31119 = n406 & n31118 ;
  assign n31120 = n31119 ^ n23511 ^ n2440 ;
  assign n31117 = n1246 | n8541 ;
  assign n31121 = n31120 ^ n31117 ^ 1'b0 ;
  assign n31122 = n31121 ^ n9756 ^ 1'b0 ;
  assign n31123 = n14425 | n31122 ;
  assign n31124 = n19781 | n31123 ;
  assign n31125 = ( n2046 & n4328 ) | ( n2046 & n18066 ) | ( n4328 & n18066 ) ;
  assign n31126 = ( n1422 & ~n9725 ) | ( n1422 & n22418 ) | ( ~n9725 & n22418 ) ;
  assign n31127 = n31126 ^ n14761 ^ n8355 ;
  assign n31128 = n31127 ^ n19263 ^ 1'b0 ;
  assign n31129 = n9060 & n31128 ;
  assign n31130 = ( n1914 & n31125 ) | ( n1914 & n31129 ) | ( n31125 & n31129 ) ;
  assign n31131 = n10863 & n25508 ;
  assign n31132 = n25093 ^ n14838 ^ n10927 ;
  assign n31134 = n31050 ^ n14693 ^ n13477 ;
  assign n31133 = n1278 & n11413 ;
  assign n31135 = n31134 ^ n31133 ^ 1'b0 ;
  assign n31139 = n12021 ^ n940 ^ x105 ;
  assign n31136 = ( n3492 & n3700 ) | ( n3492 & n4450 ) | ( n3700 & n4450 ) ;
  assign n31137 = n10657 ^ n1525 ^ n1326 ;
  assign n31138 = ( n22034 & n31136 ) | ( n22034 & ~n31137 ) | ( n31136 & ~n31137 ) ;
  assign n31140 = n31139 ^ n31138 ^ n11579 ;
  assign n31144 = ( n3743 & n12867 ) | ( n3743 & n18493 ) | ( n12867 & n18493 ) ;
  assign n31142 = ~n6390 & n13891 ;
  assign n31143 = n31142 ^ n17756 ^ 1'b0 ;
  assign n31141 = n9966 ^ n6196 ^ n2225 ;
  assign n31145 = n31144 ^ n31143 ^ n31141 ;
  assign n31146 = n30109 ^ n30048 ^ n12413 ;
  assign n31147 = ( n4795 & ~n23415 ) | ( n4795 & n31146 ) | ( ~n23415 & n31146 ) ;
  assign n31148 = n31147 ^ n5421 ^ n3770 ;
  assign n31149 = n794 ^ x131 ^ 1'b0 ;
  assign n31150 = n5267 & ~n31149 ;
  assign n31151 = n9907 | n31150 ;
  assign n31152 = ( n5361 & ~n6397 ) | ( n5361 & n31151 ) | ( ~n6397 & n31151 ) ;
  assign n31153 = n31107 ^ n3493 ^ n600 ;
  assign n31154 = n9701 & n31153 ;
  assign n31155 = n31154 ^ n11586 ^ 1'b0 ;
  assign n31159 = n19611 ^ n928 ^ x205 ;
  assign n31157 = n12931 ^ n11209 ^ n1440 ;
  assign n31156 = n12910 ^ n8656 ^ n6783 ;
  assign n31158 = n31157 ^ n31156 ^ n8632 ;
  assign n31160 = n31159 ^ n31158 ^ 1'b0 ;
  assign n31161 = ( n286 & n2476 ) | ( n286 & ~n29891 ) | ( n2476 & ~n29891 ) ;
  assign n31162 = n6264 ^ n3001 ^ 1'b0 ;
  assign n31163 = ( n12812 & n31161 ) | ( n12812 & ~n31162 ) | ( n31161 & ~n31162 ) ;
  assign n31164 = ( n2937 & ~n8324 ) | ( n2937 & n16681 ) | ( ~n8324 & n16681 ) ;
  assign n31165 = ( n3468 & n4688 ) | ( n3468 & n31164 ) | ( n4688 & n31164 ) ;
  assign n31166 = n31165 ^ n7851 ^ 1'b0 ;
  assign n31167 = n17583 & ~n31166 ;
  assign n31168 = ( n4128 & n7526 ) | ( n4128 & n25772 ) | ( n7526 & n25772 ) ;
  assign n31169 = n31168 ^ n1453 ^ 1'b0 ;
  assign n31170 = ~n13063 & n31169 ;
  assign n31171 = ( n23446 & n31167 ) | ( n23446 & ~n31170 ) | ( n31167 & ~n31170 ) ;
  assign n31172 = n6629 & n12443 ;
  assign n31173 = ~n31136 & n31172 ;
  assign n31174 = n22570 | n31173 ;
  assign n31175 = n31174 ^ n2375 ^ 1'b0 ;
  assign n31176 = ( n22069 & ~n26702 ) | ( n22069 & n31175 ) | ( ~n26702 & n31175 ) ;
  assign n31179 = n13546 ^ n13407 ^ n7001 ;
  assign n31180 = ( ~n4526 & n11262 ) | ( ~n4526 & n31179 ) | ( n11262 & n31179 ) ;
  assign n31181 = n31180 ^ n11292 ^ n5917 ;
  assign n31177 = n19002 | n19851 ;
  assign n31178 = n21992 & n31177 ;
  assign n31182 = n31181 ^ n31178 ^ 1'b0 ;
  assign n31183 = n14093 | n31182 ;
  assign n31184 = n27562 ^ n11654 ^ n7580 ;
  assign n31185 = n31184 ^ n16928 ^ n7052 ;
  assign n31186 = n22140 ^ n18084 ^ 1'b0 ;
  assign n31187 = n21901 ^ n6389 ^ n5379 ;
  assign n31188 = ( ~n8900 & n24993 ) | ( ~n8900 & n31187 ) | ( n24993 & n31187 ) ;
  assign n31189 = n31188 ^ n26578 ^ 1'b0 ;
  assign n31190 = n31071 ^ n28717 ^ 1'b0 ;
  assign n31191 = n31190 ^ n5872 ^ 1'b0 ;
  assign n31192 = ~n31189 & n31191 ;
  assign n31195 = ( ~n4333 & n11857 ) | ( ~n4333 & n20801 ) | ( n11857 & n20801 ) ;
  assign n31196 = ( n14595 & n28652 ) | ( n14595 & ~n31195 ) | ( n28652 & ~n31195 ) ;
  assign n31197 = n31196 ^ n18072 ^ 1'b0 ;
  assign n31193 = n13167 ^ n6349 ^ 1'b0 ;
  assign n31194 = ~n19985 & n31193 ;
  assign n31198 = n31197 ^ n31194 ^ n13214 ;
  assign n31204 = n6581 & ~n7723 ;
  assign n31205 = ~n3876 & n31204 ;
  assign n31206 = n31205 ^ n5540 ^ n3651 ;
  assign n31207 = ( ~n2416 & n22130 ) | ( ~n2416 & n31206 ) | ( n22130 & n31206 ) ;
  assign n31199 = ~n4481 & n7411 ;
  assign n31200 = ~n2606 & n31199 ;
  assign n31201 = ( n7118 & ~n13454 ) | ( n7118 & n31200 ) | ( ~n13454 & n31200 ) ;
  assign n31202 = n16805 ^ n7061 ^ 1'b0 ;
  assign n31203 = ( n8546 & n31201 ) | ( n8546 & ~n31202 ) | ( n31201 & ~n31202 ) ;
  assign n31208 = n31207 ^ n31203 ^ 1'b0 ;
  assign n31209 = n31198 & ~n31208 ;
  assign n31210 = n8710 ^ n2791 ^ n2441 ;
  assign n31211 = n5971 | n19715 ;
  assign n31212 = ( ~n15377 & n31210 ) | ( ~n15377 & n31211 ) | ( n31210 & n31211 ) ;
  assign n31213 = n12159 | n25419 ;
  assign n31214 = ( n8538 & ~n25368 ) | ( n8538 & n28956 ) | ( ~n25368 & n28956 ) ;
  assign n31215 = ( n14908 & ~n31213 ) | ( n14908 & n31214 ) | ( ~n31213 & n31214 ) ;
  assign n31216 = n16868 ^ n10282 ^ n1721 ;
  assign n31217 = n31216 ^ n19983 ^ n306 ;
  assign n31221 = n12034 & n19484 ;
  assign n31222 = n31221 ^ n28771 ^ n6728 ;
  assign n31218 = n6575 & ~n26641 ;
  assign n31219 = ~n328 & n31218 ;
  assign n31220 = ( n18299 & ~n23588 ) | ( n18299 & n31219 ) | ( ~n23588 & n31219 ) ;
  assign n31223 = n31222 ^ n31220 ^ 1'b0 ;
  assign n31224 = ~n22240 & n31223 ;
  assign n31225 = x211 & n10384 ;
  assign n31226 = n31225 ^ n11948 ^ n9452 ;
  assign n31227 = n6994 & ~n31226 ;
  assign n31228 = n31227 ^ n22320 ^ n11152 ;
  assign n31229 = ( ~n15440 & n31224 ) | ( ~n15440 & n31228 ) | ( n31224 & n31228 ) ;
  assign n31230 = ( ~n5287 & n6841 ) | ( ~n5287 & n7456 ) | ( n6841 & n7456 ) ;
  assign n31231 = n31230 ^ n13865 ^ n2243 ;
  assign n31232 = ~n11455 & n16715 ;
  assign n31233 = ( ~n18392 & n22686 ) | ( ~n18392 & n31232 ) | ( n22686 & n31232 ) ;
  assign n31234 = ( n3554 & n5134 ) | ( n3554 & ~n5350 ) | ( n5134 & ~n5350 ) ;
  assign n31235 = ( ~n31231 & n31233 ) | ( ~n31231 & n31234 ) | ( n31233 & n31234 ) ;
  assign n31236 = n31175 ^ n23305 ^ n3216 ;
  assign n31237 = n12677 & ~n21086 ;
  assign n31238 = ~n24888 & n31237 ;
  assign n31239 = n31238 ^ n4150 ^ 1'b0 ;
  assign n31240 = n15796 ^ n10537 ^ n8454 ;
  assign n31241 = n31240 ^ n9720 ^ n4845 ;
  assign n31242 = ( n11343 & ~n25705 ) | ( n11343 & n31241 ) | ( ~n25705 & n31241 ) ;
  assign n31243 = n24653 ^ n21675 ^ n18103 ;
  assign n31244 = n31243 ^ n28573 ^ n19507 ;
  assign n31247 = n23734 ^ n12392 ^ n1436 ;
  assign n31246 = ( n12528 & n14985 ) | ( n12528 & n27748 ) | ( n14985 & n27748 ) ;
  assign n31248 = n31247 ^ n31246 ^ n11246 ;
  assign n31245 = n10904 & ~n15206 ;
  assign n31249 = n31248 ^ n31245 ^ n9799 ;
  assign n31250 = n23065 ^ n5653 ^ 1'b0 ;
  assign n31251 = ~n24459 & n31250 ;
  assign n31252 = x98 & n18185 ;
  assign n31253 = ( n3292 & n17922 ) | ( n3292 & ~n19691 ) | ( n17922 & ~n19691 ) ;
  assign n31254 = n1226 & ~n31253 ;
  assign n31255 = n28274 & n31254 ;
  assign n31256 = n25680 ^ n813 ^ 1'b0 ;
  assign n31257 = ( x251 & n11123 ) | ( x251 & ~n30435 ) | ( n11123 & ~n30435 ) ;
  assign n31258 = n31257 ^ n10855 ^ n9100 ;
  assign n31259 = n26235 ^ n15822 ^ n3468 ;
  assign n31260 = n22691 ^ n16506 ^ n2429 ;
  assign n31261 = n31260 ^ n13582 ^ n11548 ;
  assign n31262 = ( n12900 & n20014 ) | ( n12900 & ~n31261 ) | ( n20014 & ~n31261 ) ;
  assign n31263 = ( n2403 & ~n3019 ) | ( n2403 & n23770 ) | ( ~n3019 & n23770 ) ;
  assign n31264 = ( ~n17573 & n25646 ) | ( ~n17573 & n31263 ) | ( n25646 & n31263 ) ;
  assign n31265 = n10505 ^ n10098 ^ n5077 ;
  assign n31266 = ( ~n7704 & n31264 ) | ( ~n7704 & n31265 ) | ( n31264 & n31265 ) ;
  assign n31267 = ( n12208 & ~n27600 ) | ( n12208 & n31266 ) | ( ~n27600 & n31266 ) ;
  assign n31268 = n21382 ^ n14734 ^ n1939 ;
  assign n31269 = ( n12941 & n26504 ) | ( n12941 & ~n31268 ) | ( n26504 & ~n31268 ) ;
  assign n31270 = n1410 | n26496 ;
  assign n31271 = n31270 ^ n18079 ^ 1'b0 ;
  assign n31272 = ( n5000 & n8563 ) | ( n5000 & ~n10815 ) | ( n8563 & ~n10815 ) ;
  assign n31273 = n31272 ^ n714 ^ 1'b0 ;
  assign n31274 = n18634 & ~n31273 ;
  assign n31275 = n14081 | n24223 ;
  assign n31276 = n8314 | n29827 ;
  assign n31277 = n31275 & ~n31276 ;
  assign n31278 = ( n975 & n21120 ) | ( n975 & ~n31277 ) | ( n21120 & ~n31277 ) ;
  assign n31279 = n12202 ^ n6706 ^ x46 ;
  assign n31280 = n31279 ^ n23778 ^ n6194 ;
  assign n31281 = n12692 ^ n2016 ^ 1'b0 ;
  assign n31282 = n31281 ^ n19788 ^ 1'b0 ;
  assign n31286 = ( n10607 & n19418 ) | ( n10607 & ~n25495 ) | ( n19418 & ~n25495 ) ;
  assign n31283 = ( ~n838 & n1705 ) | ( ~n838 & n21466 ) | ( n1705 & n21466 ) ;
  assign n31284 = n21941 ^ n11811 ^ n8606 ;
  assign n31285 = n31283 | n31284 ;
  assign n31287 = n31286 ^ n31285 ^ 1'b0 ;
  assign n31291 = ( ~n594 & n918 ) | ( ~n594 & n9457 ) | ( n918 & n9457 ) ;
  assign n31289 = n7102 & n7263 ;
  assign n31290 = n7864 & n31289 ;
  assign n31288 = n6953 ^ n1249 ^ 1'b0 ;
  assign n31292 = n31291 ^ n31290 ^ n31288 ;
  assign n31293 = ( n31282 & n31287 ) | ( n31282 & n31292 ) | ( n31287 & n31292 ) ;
  assign n31294 = ( n18031 & n28055 ) | ( n18031 & n31293 ) | ( n28055 & n31293 ) ;
  assign n31298 = n18257 ^ n10210 ^ 1'b0 ;
  assign n31299 = n13600 & n31298 ;
  assign n31295 = n275 | n13596 ;
  assign n31296 = n31295 ^ n5720 ^ 1'b0 ;
  assign n31297 = n31296 ^ n28477 ^ n10796 ;
  assign n31300 = n31299 ^ n31297 ^ n14097 ;
  assign n31301 = n30143 ^ n15460 ^ n6987 ;
  assign n31302 = ( n6670 & n12148 ) | ( n6670 & ~n27246 ) | ( n12148 & ~n27246 ) ;
  assign n31303 = n6752 & n31302 ;
  assign n31304 = n31301 & n31303 ;
  assign n31305 = n25090 & ~n31304 ;
  assign n31306 = ( n1625 & n4822 ) | ( n1625 & ~n5472 ) | ( n4822 & ~n5472 ) ;
  assign n31307 = n327 | n31306 ;
  assign n31308 = n28347 & n31307 ;
  assign n31309 = n31308 ^ n18236 ^ 1'b0 ;
  assign n31310 = n21335 ^ n14772 ^ n8702 ;
  assign n31311 = n26590 ^ n18145 ^ n14267 ;
  assign n31312 = ( n6559 & ~n31310 ) | ( n6559 & n31311 ) | ( ~n31310 & n31311 ) ;
  assign n31315 = n7209 ^ n1474 ^ 1'b0 ;
  assign n31313 = n7836 ^ n7289 ^ n3143 ;
  assign n31314 = n31313 ^ n10981 ^ n7246 ;
  assign n31316 = n31315 ^ n31314 ^ n7972 ;
  assign n31320 = n27089 ^ n19078 ^ n2152 ;
  assign n31317 = n23587 ^ n1612 ^ 1'b0 ;
  assign n31318 = n31317 ^ n16879 ^ n2505 ;
  assign n31319 = n31318 ^ n7111 ^ n2105 ;
  assign n31321 = n31320 ^ n31319 ^ n5641 ;
  assign n31322 = n31321 ^ n26391 ^ 1'b0 ;
  assign n31323 = ~n2743 & n31322 ;
  assign n31324 = n11197 ^ n6933 ^ 1'b0 ;
  assign n31325 = ~n1663 & n31324 ;
  assign n31326 = ( n15250 & ~n18859 ) | ( n15250 & n31325 ) | ( ~n18859 & n31325 ) ;
  assign n31327 = ( ~n2857 & n15074 ) | ( ~n2857 & n31326 ) | ( n15074 & n31326 ) ;
  assign n31328 = n7110 & ~n15717 ;
  assign n31329 = ( n4034 & ~n17112 ) | ( n4034 & n31328 ) | ( ~n17112 & n31328 ) ;
  assign n31330 = ( ~n25961 & n30017 ) | ( ~n25961 & n31329 ) | ( n30017 & n31329 ) ;
  assign n31331 = ~n29354 & n31330 ;
  assign n31332 = n25034 ^ n24832 ^ n8484 ;
  assign n31333 = n21326 ^ n9188 ^ n5479 ;
  assign n31334 = ( n8149 & ~n22891 ) | ( n8149 & n31333 ) | ( ~n22891 & n31333 ) ;
  assign n31335 = ( n13107 & n15140 ) | ( n13107 & ~n16013 ) | ( n15140 & ~n16013 ) ;
  assign n31336 = n30378 ^ n28852 ^ 1'b0 ;
  assign n31337 = n31335 & n31336 ;
  assign n31338 = n20120 ^ n12551 ^ 1'b0 ;
  assign n31339 = n3653 ^ n1896 ^ 1'b0 ;
  assign n31340 = n31339 ^ n2901 ^ 1'b0 ;
  assign n31341 = n31340 ^ n12250 ^ n10084 ;
  assign n31342 = ( n4043 & n19020 ) | ( n4043 & ~n24990 ) | ( n19020 & ~n24990 ) ;
  assign n31343 = n12739 ^ n10636 ^ n1567 ;
  assign n31344 = n4901 & ~n25846 ;
  assign n31345 = n7327 ^ n3006 ^ n1626 ;
  assign n31346 = ( ~n31343 & n31344 ) | ( ~n31343 & n31345 ) | ( n31344 & n31345 ) ;
  assign n31347 = ( n5034 & n7504 ) | ( n5034 & ~n20105 ) | ( n7504 & ~n20105 ) ;
  assign n31348 = n31347 ^ n18371 ^ n362 ;
  assign n31349 = ( n5044 & n12102 ) | ( n5044 & ~n26441 ) | ( n12102 & ~n26441 ) ;
  assign n31350 = n10149 | n26056 ;
  assign n31351 = n31349 & ~n31350 ;
  assign n31352 = n14821 & ~n28115 ;
  assign n31353 = x106 | n9713 ;
  assign n31354 = ~n6854 & n23478 ;
  assign n31355 = n15630 & n31354 ;
  assign n31356 = n31355 ^ n22632 ^ n17923 ;
  assign n31357 = n31353 & ~n31356 ;
  assign n31358 = n13161 & n31357 ;
  assign n31359 = ( n2068 & n22577 ) | ( n2068 & ~n25368 ) | ( n22577 & ~n25368 ) ;
  assign n31360 = n31359 ^ n23166 ^ n19200 ;
  assign n31361 = ( n4677 & n8895 ) | ( n4677 & ~n12417 ) | ( n8895 & ~n12417 ) ;
  assign n31362 = ( n5027 & ~n13345 ) | ( n5027 & n19146 ) | ( ~n13345 & n19146 ) ;
  assign n31363 = ( n3824 & n7299 ) | ( n3824 & ~n13197 ) | ( n7299 & ~n13197 ) ;
  assign n31364 = n31362 & ~n31363 ;
  assign n31365 = ( n5108 & n17810 ) | ( n5108 & n31364 ) | ( n17810 & n31364 ) ;
  assign n31366 = n31365 ^ n7467 ^ 1'b0 ;
  assign n31367 = n20722 ^ n6413 ^ n939 ;
  assign n31368 = n31367 ^ n17932 ^ n8806 ;
  assign n31370 = ( ~n6684 & n12537 ) | ( ~n6684 & n17702 ) | ( n12537 & n17702 ) ;
  assign n31369 = n13319 ^ n11670 ^ 1'b0 ;
  assign n31371 = n31370 ^ n31369 ^ n17344 ;
  assign n31372 = n31371 ^ n24496 ^ n18177 ;
  assign n31373 = n9789 ^ n8042 ^ n2755 ;
  assign n31374 = n15653 ^ n12166 ^ 1'b0 ;
  assign n31375 = n16954 ^ n7371 ^ 1'b0 ;
  assign n31376 = n8134 & ~n19241 ;
  assign n31377 = ~n31375 & n31376 ;
  assign n31378 = ( n10642 & n31374 ) | ( n10642 & ~n31377 ) | ( n31374 & ~n31377 ) ;
  assign n31382 = n440 & n5965 ;
  assign n31383 = n1568 & n31382 ;
  assign n31384 = n15902 & ~n31383 ;
  assign n31385 = n31384 ^ n16940 ^ 1'b0 ;
  assign n31381 = ( n1432 & n3582 ) | ( n1432 & n13579 ) | ( n3582 & n13579 ) ;
  assign n31379 = ( n7235 & n11335 ) | ( n7235 & ~n12890 ) | ( n11335 & ~n12890 ) ;
  assign n31380 = n31379 ^ n31052 ^ n555 ;
  assign n31386 = n31385 ^ n31381 ^ n31380 ;
  assign n31387 = ( n1551 & n3259 ) | ( n1551 & n20288 ) | ( n3259 & n20288 ) ;
  assign n31388 = n31387 ^ n10379 ^ 1'b0 ;
  assign n31389 = n15284 | n31388 ;
  assign n31390 = n19790 ^ n813 ^ 1'b0 ;
  assign n31391 = n31390 ^ n4733 ^ 1'b0 ;
  assign n31392 = ~n9278 & n31391 ;
  assign n31393 = n31392 ^ n12245 ^ n9041 ;
  assign n31394 = n28625 ^ n21302 ^ n10767 ;
  assign n31395 = n29607 | n31394 ;
  assign n31396 = ~n3177 & n12955 ;
  assign n31397 = ~n27292 & n31396 ;
  assign n31398 = ( n4278 & n28730 ) | ( n4278 & ~n31397 ) | ( n28730 & ~n31397 ) ;
  assign n31399 = n17284 ^ n12745 ^ n2078 ;
  assign n31400 = ~n2779 & n7282 ;
  assign n31401 = ~n14161 & n31400 ;
  assign n31402 = n31401 ^ n26986 ^ 1'b0 ;
  assign n31403 = n658 | n12017 ;
  assign n31404 = n31403 ^ n6202 ^ 1'b0 ;
  assign n31405 = n31404 ^ n22761 ^ n17122 ;
  assign n31406 = ( n9433 & n31402 ) | ( n9433 & ~n31405 ) | ( n31402 & ~n31405 ) ;
  assign n31407 = ( ~n546 & n31399 ) | ( ~n546 & n31406 ) | ( n31399 & n31406 ) ;
  assign n31408 = n10169 | n23408 ;
  assign n31409 = n25203 ^ n18961 ^ x131 ;
  assign n31410 = ( n12344 & n31279 ) | ( n12344 & ~n31409 ) | ( n31279 & ~n31409 ) ;
  assign n31412 = n5240 | n18559 ;
  assign n31413 = n31412 ^ n7852 ^ 1'b0 ;
  assign n31411 = n29479 ^ n16247 ^ n10540 ;
  assign n31414 = n31413 ^ n31411 ^ n2776 ;
  assign n31415 = n22542 ^ n4827 ^ n4233 ;
  assign n31416 = n8389 ^ n7166 ^ n2467 ;
  assign n31417 = n31416 ^ n19002 ^ n5613 ;
  assign n31418 = ( n1272 & n4229 ) | ( n1272 & ~n10590 ) | ( n4229 & ~n10590 ) ;
  assign n31419 = ~n2571 & n31418 ;
  assign n31420 = n19021 ^ n14278 ^ n12797 ;
  assign n31421 = n31420 ^ n31210 ^ n5831 ;
  assign n31422 = n3649 ^ n1389 ^ 1'b0 ;
  assign n31423 = n17064 & ~n31422 ;
  assign n31424 = n29071 ^ n17614 ^ 1'b0 ;
  assign n31425 = ( n5902 & n31423 ) | ( n5902 & n31424 ) | ( n31423 & n31424 ) ;
  assign n31426 = ( ~n2151 & n4644 ) | ( ~n2151 & n6494 ) | ( n4644 & n6494 ) ;
  assign n31427 = ( n6810 & n21557 ) | ( n6810 & ~n28780 ) | ( n21557 & ~n28780 ) ;
  assign n31428 = n29305 ^ n6765 ^ 1'b0 ;
  assign n31429 = ~n17489 & n31428 ;
  assign n31430 = n31429 ^ n11464 ^ n3208 ;
  assign n31431 = ( n31426 & n31427 ) | ( n31426 & ~n31430 ) | ( n31427 & ~n31430 ) ;
  assign n31432 = ( n9692 & n14833 ) | ( n9692 & ~n16264 ) | ( n14833 & ~n16264 ) ;
  assign n31433 = ( n5462 & ~n19558 ) | ( n5462 & n22410 ) | ( ~n19558 & n22410 ) ;
  assign n31434 = n19216 ^ n11622 ^ n3694 ;
  assign n31435 = n1355 & ~n12223 ;
  assign n31436 = n14263 & n31435 ;
  assign n31437 = n20079 ^ n15876 ^ 1'b0 ;
  assign n31438 = ( n15836 & n17752 ) | ( n15836 & ~n17809 ) | ( n17752 & ~n17809 ) ;
  assign n31439 = ( n21789 & n31437 ) | ( n21789 & ~n31438 ) | ( n31437 & ~n31438 ) ;
  assign n31440 = ( n21560 & n29349 ) | ( n21560 & ~n31439 ) | ( n29349 & ~n31439 ) ;
  assign n31444 = n2454 | n4147 ;
  assign n31446 = n17134 ^ n8677 ^ n7940 ;
  assign n31445 = n16011 ^ n8458 ^ 1'b0 ;
  assign n31447 = n31446 ^ n31445 ^ n3519 ;
  assign n31448 = ( ~n2110 & n31444 ) | ( ~n2110 & n31447 ) | ( n31444 & n31447 ) ;
  assign n31449 = ( ~n18794 & n20466 ) | ( ~n18794 & n31448 ) | ( n20466 & n31448 ) ;
  assign n31441 = n23180 ^ n9619 ^ n8935 ;
  assign n31442 = n24287 ^ n14088 ^ n11447 ;
  assign n31443 = ( n10030 & n31441 ) | ( n10030 & ~n31442 ) | ( n31441 & ~n31442 ) ;
  assign n31450 = n31449 ^ n31443 ^ 1'b0 ;
  assign n31451 = n7039 ^ n1108 ^ 1'b0 ;
  assign n31452 = n7948 & ~n31451 ;
  assign n31453 = n31452 ^ n30463 ^ n23482 ;
  assign n31455 = ( ~n5986 & n6042 ) | ( ~n5986 & n6780 ) | ( n6042 & n6780 ) ;
  assign n31456 = n31455 ^ n23504 ^ n21233 ;
  assign n31454 = x89 & ~n21023 ;
  assign n31457 = n31456 ^ n31454 ^ 1'b0 ;
  assign n31458 = ( n15336 & n17120 ) | ( n15336 & n19633 ) | ( n17120 & n19633 ) ;
  assign n31459 = n24335 ^ n18381 ^ 1'b0 ;
  assign n31460 = n23591 ^ n14027 ^ n2891 ;
  assign n31461 = n31460 ^ n18576 ^ n9331 ;
  assign n31462 = ( x76 & n3715 ) | ( x76 & ~n6743 ) | ( n3715 & ~n6743 ) ;
  assign n31463 = n1797 & n31462 ;
  assign n31464 = ( n16041 & n29201 ) | ( n16041 & n31463 ) | ( n29201 & n31463 ) ;
  assign n31465 = n7120 & n16034 ;
  assign n31466 = n31465 ^ n22303 ^ 1'b0 ;
  assign n31474 = n11606 ^ n11083 ^ n466 ;
  assign n31475 = n31474 ^ n9068 ^ n6682 ;
  assign n31469 = n16416 ^ n11064 ^ n972 ;
  assign n31467 = n24642 ^ n15821 ^ n9881 ;
  assign n31468 = n17007 & ~n31467 ;
  assign n31470 = n31469 ^ n31468 ^ 1'b0 ;
  assign n31471 = ( n8241 & n15725 ) | ( n8241 & ~n31470 ) | ( n15725 & ~n31470 ) ;
  assign n31472 = n16544 ^ n9591 ^ 1'b0 ;
  assign n31473 = ~n31471 & n31472 ;
  assign n31476 = n31475 ^ n31473 ^ n6886 ;
  assign n31477 = ( ~n16264 & n24740 ) | ( ~n16264 & n31476 ) | ( n24740 & n31476 ) ;
  assign n31478 = n8947 | n12840 ;
  assign n31479 = n12898 ^ n12150 ^ 1'b0 ;
  assign n31487 = ~n9922 & n21511 ;
  assign n31488 = n31487 ^ n14357 ^ 1'b0 ;
  assign n31485 = n16346 ^ n12723 ^ n8434 ;
  assign n31484 = ~n2953 & n25804 ;
  assign n31481 = ( n922 & n7641 ) | ( n922 & n27354 ) | ( n7641 & n27354 ) ;
  assign n31480 = n5359 | n14621 ;
  assign n31482 = n31481 ^ n31480 ^ 1'b0 ;
  assign n31483 = n9491 & ~n31482 ;
  assign n31486 = n31485 ^ n31484 ^ n31483 ;
  assign n31489 = n31488 ^ n31486 ^ 1'b0 ;
  assign n31490 = ( n12219 & ~n22879 ) | ( n12219 & n31489 ) | ( ~n22879 & n31489 ) ;
  assign n31497 = n23638 ^ n15909 ^ n2481 ;
  assign n31498 = ( n1700 & n2655 ) | ( n1700 & n26979 ) | ( n2655 & n26979 ) ;
  assign n31499 = ( n13806 & ~n31497 ) | ( n13806 & n31498 ) | ( ~n31497 & n31498 ) ;
  assign n31491 = n28166 ^ n10758 ^ 1'b0 ;
  assign n31492 = ~n3454 & n7217 ;
  assign n31493 = n8103 & n31492 ;
  assign n31494 = ( n1379 & n6888 ) | ( n1379 & n12045 ) | ( n6888 & n12045 ) ;
  assign n31495 = ( n13005 & ~n31493 ) | ( n13005 & n31494 ) | ( ~n31493 & n31494 ) ;
  assign n31496 = ( ~n19829 & n31491 ) | ( ~n19829 & n31495 ) | ( n31491 & n31495 ) ;
  assign n31500 = n31499 ^ n31496 ^ n7547 ;
  assign n31501 = ( n10988 & ~n28534 ) | ( n10988 & n31500 ) | ( ~n28534 & n31500 ) ;
  assign n31503 = ( n443 & n3145 ) | ( n443 & n5045 ) | ( n3145 & n5045 ) ;
  assign n31502 = ( ~n1221 & n21979 ) | ( ~n1221 & n29355 ) | ( n21979 & n29355 ) ;
  assign n31504 = n31503 ^ n31502 ^ 1'b0 ;
  assign n31505 = ~n27555 & n31504 ;
  assign n31506 = n31505 ^ n14820 ^ n3087 ;
  assign n31507 = ( n7819 & n14368 ) | ( n7819 & ~n19189 ) | ( n14368 & ~n19189 ) ;
  assign n31508 = n21334 ^ n9384 ^ 1'b0 ;
  assign n31509 = ~n1525 & n31508 ;
  assign n31510 = n31509 ^ n10125 ^ n7106 ;
  assign n31511 = n23442 ^ n23098 ^ 1'b0 ;
  assign n31512 = n13370 & n31511 ;
  assign n31513 = n23491 ^ n8909 ^ n8666 ;
  assign n31514 = n31513 ^ n23810 ^ 1'b0 ;
  assign n31515 = n31512 & ~n31514 ;
  assign n31516 = n18943 & n23384 ;
  assign n31517 = n26715 ^ n15079 ^ 1'b0 ;
  assign n31518 = ( n9767 & n19843 ) | ( n9767 & n26879 ) | ( n19843 & n26879 ) ;
  assign n31519 = ( ~n11984 & n31517 ) | ( ~n11984 & n31518 ) | ( n31517 & n31518 ) ;
  assign n31520 = ( x149 & ~n5813 ) | ( x149 & n10487 ) | ( ~n5813 & n10487 ) ;
  assign n31521 = n31520 ^ n2374 ^ 1'b0 ;
  assign n31522 = n8316 & ~n9676 ;
  assign n31523 = ~n21308 & n31522 ;
  assign n31524 = ( n1422 & n7367 ) | ( n1422 & ~n7592 ) | ( n7367 & ~n7592 ) ;
  assign n31525 = n31524 ^ n1980 ^ 1'b0 ;
  assign n31526 = n877 & n31525 ;
  assign n31527 = ( ~n6243 & n29062 ) | ( ~n6243 & n31526 ) | ( n29062 & n31526 ) ;
  assign n31535 = n12274 ^ n5922 ^ 1'b0 ;
  assign n31536 = n6855 & ~n31535 ;
  assign n31528 = ( n924 & n13438 ) | ( n924 & n19564 ) | ( n13438 & n19564 ) ;
  assign n31530 = n9448 ^ n4775 ^ n3138 ;
  assign n31531 = n20244 ^ n14153 ^ n7860 ;
  assign n31532 = ( n6999 & n31530 ) | ( n6999 & ~n31531 ) | ( n31530 & ~n31531 ) ;
  assign n31529 = n15946 ^ n7862 ^ 1'b0 ;
  assign n31533 = n31532 ^ n31529 ^ n22179 ;
  assign n31534 = ( ~n12288 & n31528 ) | ( ~n12288 & n31533 ) | ( n31528 & n31533 ) ;
  assign n31537 = n31536 ^ n31534 ^ n28912 ;
  assign n31539 = n14404 ^ n4642 ^ 1'b0 ;
  assign n31540 = n31539 ^ n11794 ^ 1'b0 ;
  assign n31538 = n10428 ^ x155 ^ 1'b0 ;
  assign n31541 = n31540 ^ n31538 ^ n17756 ;
  assign n31542 = ( n7351 & n14591 ) | ( n7351 & ~n18107 ) | ( n14591 & ~n18107 ) ;
  assign n31544 = n28655 ^ n14989 ^ n12550 ;
  assign n31545 = ( n17063 & n19347 ) | ( n17063 & n31544 ) | ( n19347 & n31544 ) ;
  assign n31543 = n4653 | n23640 ;
  assign n31546 = n31545 ^ n31543 ^ 1'b0 ;
  assign n31547 = n18336 ^ n2350 ^ x60 ;
  assign n31548 = n31547 ^ n27757 ^ n21111 ;
  assign n31549 = ( n7762 & n8768 ) | ( n7762 & ~n31548 ) | ( n8768 & ~n31548 ) ;
  assign n31550 = n17929 ^ n9278 ^ n4301 ;
  assign n31551 = n19243 ^ n11926 ^ n5275 ;
  assign n31552 = n17001 ^ n7210 ^ 1'b0 ;
  assign n31553 = ~n7236 & n31552 ;
  assign n31554 = n28720 ^ n3958 ^ n2889 ;
  assign n31555 = ( n3398 & n11046 ) | ( n3398 & n31554 ) | ( n11046 & n31554 ) ;
  assign n31556 = n31555 ^ n29181 ^ n22132 ;
  assign n31557 = n5467 | n13561 ;
  assign n31558 = n31557 ^ n26176 ^ 1'b0 ;
  assign n31559 = n31558 ^ n16340 ^ n2372 ;
  assign n31560 = ( n1577 & n2712 ) | ( n1577 & ~n8962 ) | ( n2712 & ~n8962 ) ;
  assign n31562 = n1581 & n3373 ;
  assign n31561 = n24202 ^ n11922 ^ n8565 ;
  assign n31563 = n31562 ^ n31561 ^ n23531 ;
  assign n31564 = ~n31560 & n31563 ;
  assign n31565 = ( n11271 & ~n31559 ) | ( n11271 & n31564 ) | ( ~n31559 & n31564 ) ;
  assign n31566 = n25943 ^ n17418 ^ n11626 ;
  assign n31567 = n27714 ^ n13153 ^ 1'b0 ;
  assign n31568 = n11108 ^ n8160 ^ n461 ;
  assign n31569 = n31568 ^ n8497 ^ n3691 ;
  assign n31570 = ( n12902 & ~n15138 ) | ( n12902 & n22615 ) | ( ~n15138 & n22615 ) ;
  assign n31571 = n4841 | n31570 ;
  assign n31572 = n31569 & ~n31571 ;
  assign n31573 = n27087 ^ n22377 ^ n20318 ;
  assign n31574 = ( n1608 & n20759 ) | ( n1608 & n23793 ) | ( n20759 & n23793 ) ;
  assign n31575 = n31574 ^ n19296 ^ n9856 ;
  assign n31576 = ~n9855 & n12385 ;
  assign n31577 = n31575 & n31576 ;
  assign n31578 = n31577 ^ n23147 ^ 1'b0 ;
  assign n31579 = n11259 ^ x173 ^ 1'b0 ;
  assign n31580 = ~n1945 & n31579 ;
  assign n31581 = ( n1235 & n17082 ) | ( n1235 & ~n31580 ) | ( n17082 & ~n31580 ) ;
  assign n31582 = ( ~n5725 & n16936 ) | ( ~n5725 & n21424 ) | ( n16936 & n21424 ) ;
  assign n31583 = n4227 & ~n5078 ;
  assign n31584 = ( n7695 & n12480 ) | ( n7695 & n31583 ) | ( n12480 & n31583 ) ;
  assign n31585 = n31584 ^ n26354 ^ n15279 ;
  assign n31586 = n393 & n868 ;
  assign n31587 = ~n31585 & n31586 ;
  assign n31588 = ( n4612 & n15903 ) | ( n4612 & n22547 ) | ( n15903 & n22547 ) ;
  assign n31589 = n6019 | n31284 ;
  assign n31590 = ( n19173 & n22026 ) | ( n19173 & ~n31589 ) | ( n22026 & ~n31589 ) ;
  assign n31591 = n29066 ^ n17808 ^ 1'b0 ;
  assign n31592 = ( n5400 & n11345 ) | ( n5400 & n26488 ) | ( n11345 & n26488 ) ;
  assign n31593 = n693 & ~n2265 ;
  assign n31594 = n28422 ^ n14618 ^ 1'b0 ;
  assign n31595 = ( n31592 & n31593 ) | ( n31592 & ~n31594 ) | ( n31593 & ~n31594 ) ;
  assign n31596 = n26683 ^ n19871 ^ n5344 ;
  assign n31597 = n31596 ^ n30625 ^ n10179 ;
  assign n31598 = n31092 ^ n15076 ^ n3034 ;
  assign n31599 = n12312 ^ n7692 ^ n3840 ;
  assign n31600 = ( n11624 & n17247 ) | ( n11624 & n25797 ) | ( n17247 & n25797 ) ;
  assign n31601 = n7660 ^ n7448 ^ 1'b0 ;
  assign n31602 = ~n12262 & n31601 ;
  assign n31603 = n22557 ^ n4961 ^ n4092 ;
  assign n31604 = n31602 & ~n31603 ;
  assign n31605 = n23239 & n26162 ;
  assign n31606 = n15524 & n31605 ;
  assign n31612 = n8039 | n24829 ;
  assign n31613 = n31612 ^ n7605 ^ 1'b0 ;
  assign n31614 = ~n3462 & n31613 ;
  assign n31615 = n31614 ^ n25025 ^ 1'b0 ;
  assign n31610 = n27187 ^ n18123 ^ n6118 ;
  assign n31607 = n21876 ^ n20892 ^ n810 ;
  assign n31608 = n31607 ^ n14794 ^ n8338 ;
  assign n31609 = n31608 ^ n2588 ^ n2330 ;
  assign n31611 = n31610 ^ n31609 ^ n31467 ;
  assign n31616 = n31615 ^ n31611 ^ n26212 ;
  assign n31617 = n25435 ^ n13721 ^ 1'b0 ;
  assign n31618 = n31617 ^ n28300 ^ 1'b0 ;
  assign n31625 = ( n5403 & n12664 ) | ( n5403 & ~n23583 ) | ( n12664 & ~n23583 ) ;
  assign n31626 = ( n1326 & n1682 ) | ( n1326 & n31625 ) | ( n1682 & n31625 ) ;
  assign n31624 = ( n3272 & n10901 ) | ( n3272 & n25429 ) | ( n10901 & n25429 ) ;
  assign n31627 = n31626 ^ n31624 ^ 1'b0 ;
  assign n31628 = n19278 & ~n31627 ;
  assign n31619 = ( n3105 & n5858 ) | ( n3105 & ~n6288 ) | ( n5858 & ~n6288 ) ;
  assign n31620 = ( n1595 & ~n5778 ) | ( n1595 & n31619 ) | ( ~n5778 & n31619 ) ;
  assign n31621 = n31620 ^ n12079 ^ n7482 ;
  assign n31622 = n18065 | n31621 ;
  assign n31623 = n31622 ^ n14888 ^ 1'b0 ;
  assign n31629 = n31628 ^ n31623 ^ n1710 ;
  assign n31630 = ( n5567 & n6831 ) | ( n5567 & n10758 ) | ( n6831 & n10758 ) ;
  assign n31631 = ( n5954 & n14183 ) | ( n5954 & ~n31630 ) | ( n14183 & ~n31630 ) ;
  assign n31632 = ( n6052 & n28706 ) | ( n6052 & n31631 ) | ( n28706 & n31631 ) ;
  assign n31638 = n29780 ^ n8699 ^ 1'b0 ;
  assign n31637 = ( n7454 & ~n10507 ) | ( n7454 & n22160 ) | ( ~n10507 & n22160 ) ;
  assign n31633 = ~n5657 & n12718 ;
  assign n31634 = n29706 & n31633 ;
  assign n31635 = ( n20593 & ~n24403 ) | ( n20593 & n31634 ) | ( ~n24403 & n31634 ) ;
  assign n31636 = ( ~n7098 & n16899 ) | ( ~n7098 & n31635 ) | ( n16899 & n31635 ) ;
  assign n31639 = n31638 ^ n31637 ^ n31636 ;
  assign n31640 = ( n604 & ~n7402 ) | ( n604 & n11128 ) | ( ~n7402 & n11128 ) ;
  assign n31641 = n5574 ^ n3316 ^ n1774 ;
  assign n31642 = n31641 ^ n3124 ^ 1'b0 ;
  assign n31643 = n31642 ^ n11399 ^ 1'b0 ;
  assign n31644 = n31643 ^ n27134 ^ n13146 ;
  assign n31645 = ~n4823 & n4911 ;
  assign n31646 = n31645 ^ n10297 ^ 1'b0 ;
  assign n31647 = ( n1847 & n9496 ) | ( n1847 & n31646 ) | ( n9496 & n31646 ) ;
  assign n31648 = n31647 ^ n12491 ^ n2012 ;
  assign n31649 = n29345 ^ n14652 ^ 1'b0 ;
  assign n31650 = n27192 ^ n17869 ^ 1'b0 ;
  assign n31651 = ~n31649 & n31650 ;
  assign n31652 = n21464 ^ n20940 ^ 1'b0 ;
  assign n31653 = ( ~n5761 & n15812 ) | ( ~n5761 & n31652 ) | ( n15812 & n31652 ) ;
  assign n31654 = n16287 & ~n28678 ;
  assign n31655 = ~n31653 & n31654 ;
  assign n31656 = ( ~n3102 & n10374 ) | ( ~n3102 & n11482 ) | ( n10374 & n11482 ) ;
  assign n31657 = ( ~n21692 & n28511 ) | ( ~n21692 & n29493 ) | ( n28511 & n29493 ) ;
  assign n31658 = n29222 ^ n4707 ^ 1'b0 ;
  assign n31659 = n23320 ^ n8172 ^ 1'b0 ;
  assign n31660 = ( n9133 & n14101 ) | ( n9133 & ~n29258 ) | ( n14101 & ~n29258 ) ;
  assign n31661 = ( ~n18505 & n31659 ) | ( ~n18505 & n31660 ) | ( n31659 & n31660 ) ;
  assign n31662 = ( n4915 & ~n18670 ) | ( n4915 & n31661 ) | ( ~n18670 & n31661 ) ;
  assign n31667 = ( n17114 & n17461 ) | ( n17114 & ~n30896 ) | ( n17461 & ~n30896 ) ;
  assign n31668 = n31667 ^ n18271 ^ n17944 ;
  assign n31663 = n7408 & n14063 ;
  assign n31664 = n31663 ^ n814 ^ 1'b0 ;
  assign n31665 = ( n19551 & n25644 ) | ( n19551 & n31664 ) | ( n25644 & n31664 ) ;
  assign n31666 = n4251 & n31665 ;
  assign n31669 = n31668 ^ n31666 ^ 1'b0 ;
  assign n31671 = n14420 ^ n2947 ^ 1'b0 ;
  assign n31670 = n20593 & ~n27003 ;
  assign n31672 = n31671 ^ n31670 ^ 1'b0 ;
  assign n31673 = ( n1194 & n4661 ) | ( n1194 & n16509 ) | ( n4661 & n16509 ) ;
  assign n31674 = ( ~n8472 & n25173 ) | ( ~n8472 & n31673 ) | ( n25173 & n31673 ) ;
  assign n31675 = n2318 & n28097 ;
  assign n31676 = n31675 ^ n11246 ^ 1'b0 ;
  assign n31677 = n31676 ^ n11225 ^ n10682 ;
  assign n31678 = n21318 ^ n14560 ^ n12985 ;
  assign n31679 = ( n6770 & n14285 ) | ( n6770 & n31678 ) | ( n14285 & n31678 ) ;
  assign n31680 = n31679 ^ n8281 ^ 1'b0 ;
  assign n31681 = n8254 & ~n31680 ;
  assign n31682 = n17704 ^ n1630 ^ 1'b0 ;
  assign n31683 = n4688 & n31682 ;
  assign n31685 = ( n3554 & n4213 ) | ( n3554 & ~n7494 ) | ( n4213 & ~n7494 ) ;
  assign n31684 = n23481 ^ n6071 ^ 1'b0 ;
  assign n31686 = n31685 ^ n31684 ^ n15121 ;
  assign n31687 = n31686 ^ n14420 ^ 1'b0 ;
  assign n31688 = n24822 | n31687 ;
  assign n31689 = n16605 ^ n7212 ^ n6941 ;
  assign n31690 = n31689 ^ n12743 ^ n2427 ;
  assign n31691 = n31690 ^ n28280 ^ n23015 ;
  assign n31692 = ( n11507 & n17191 ) | ( n11507 & n22271 ) | ( n17191 & n22271 ) ;
  assign n31693 = n31692 ^ n15693 ^ n7574 ;
  assign n31694 = n27347 ^ n7834 ^ 1'b0 ;
  assign n31695 = n31694 ^ n7146 ^ n1572 ;
  assign n31698 = n8862 ^ n7215 ^ n5036 ;
  assign n31697 = n3429 & ~n5966 ;
  assign n31699 = n31698 ^ n31697 ^ 1'b0 ;
  assign n31696 = n13713 ^ n8761 ^ n6391 ;
  assign n31700 = n31699 ^ n31696 ^ 1'b0 ;
  assign n31701 = n31695 | n31700 ;
  assign n31702 = n19983 ^ n11320 ^ 1'b0 ;
  assign n31703 = ( ~n12205 & n14638 ) | ( ~n12205 & n20952 ) | ( n14638 & n20952 ) ;
  assign n31704 = ( n3128 & ~n29964 ) | ( n3128 & n31703 ) | ( ~n29964 & n31703 ) ;
  assign n31705 = n31704 ^ n16691 ^ n15749 ;
  assign n31706 = n1337 | n31705 ;
  assign n31707 = n31702 & ~n31706 ;
  assign n31709 = ( n10099 & ~n16437 ) | ( n10099 & n28575 ) | ( ~n16437 & n28575 ) ;
  assign n31708 = ( n3209 & n12831 ) | ( n3209 & ~n14314 ) | ( n12831 & ~n14314 ) ;
  assign n31710 = n31709 ^ n31708 ^ n10467 ;
  assign n31711 = n3755 & ~n15547 ;
  assign n31712 = n31711 ^ n2230 ^ 1'b0 ;
  assign n31713 = n6905 | n31712 ;
  assign n31714 = n31713 ^ n23185 ^ 1'b0 ;
  assign n31715 = ( n7434 & n15072 ) | ( n7434 & n31714 ) | ( n15072 & n31714 ) ;
  assign n31716 = ( n12093 & ~n18641 ) | ( n12093 & n28002 ) | ( ~n18641 & n28002 ) ;
  assign n31717 = n31715 & n31716 ;
  assign n31718 = n19514 & ~n25037 ;
  assign n31719 = ( n10040 & n21268 ) | ( n10040 & n22691 ) | ( n21268 & n22691 ) ;
  assign n31722 = n1396 & ~n2420 ;
  assign n31723 = n31722 ^ n6487 ^ 1'b0 ;
  assign n31724 = n31723 ^ n7446 ^ 1'b0 ;
  assign n31720 = n3357 & ~n3757 ;
  assign n31721 = n31720 ^ n14839 ^ 1'b0 ;
  assign n31725 = n31724 ^ n31721 ^ 1'b0 ;
  assign n31726 = n31719 | n31725 ;
  assign n31727 = x205 & ~n20022 ;
  assign n31728 = n31727 ^ n22651 ^ 1'b0 ;
  assign n31729 = n8436 ^ n4313 ^ n397 ;
  assign n31730 = ( n13331 & ~n19336 ) | ( n13331 & n31729 ) | ( ~n19336 & n31729 ) ;
  assign n31731 = n20410 & n25968 ;
  assign n31732 = ~n9500 & n31731 ;
  assign n31733 = ( ~n8730 & n17999 ) | ( ~n8730 & n31732 ) | ( n17999 & n31732 ) ;
  assign n31734 = ( n20764 & n31730 ) | ( n20764 & n31733 ) | ( n31730 & n31733 ) ;
  assign n31735 = n26805 ^ n18856 ^ n11573 ;
  assign n31736 = n4107 ^ n3108 ^ n2447 ;
  assign n31737 = n18165 ^ n12487 ^ n2074 ;
  assign n31738 = n19218 ^ n12847 ^ n2178 ;
  assign n31739 = ( n31736 & n31737 ) | ( n31736 & ~n31738 ) | ( n31737 & ~n31738 ) ;
  assign n31740 = n16689 ^ n11484 ^ n1347 ;
  assign n31741 = n17957 ^ n9725 ^ n1156 ;
  assign n31742 = n31741 ^ n19120 ^ n14468 ;
  assign n31743 = ( n2633 & ~n31740 ) | ( n2633 & n31742 ) | ( ~n31740 & n31742 ) ;
  assign n31744 = ( n2993 & n31739 ) | ( n2993 & ~n31743 ) | ( n31739 & ~n31743 ) ;
  assign n31746 = n17675 ^ n13228 ^ n4698 ;
  assign n31745 = n13903 ^ n6946 ^ n3328 ;
  assign n31747 = n31746 ^ n31745 ^ n21419 ;
  assign n31748 = n31747 ^ n11802 ^ n9962 ;
  assign n31749 = n22540 & ~n29964 ;
  assign n31750 = n29854 ^ n21573 ^ n18497 ;
  assign n31751 = ( n17162 & n31749 ) | ( n17162 & n31750 ) | ( n31749 & n31750 ) ;
  assign n31752 = ~n5117 & n28507 ;
  assign n31753 = n31752 ^ n27921 ^ 1'b0 ;
  assign n31754 = n17790 | n19068 ;
  assign n31755 = ( n5201 & n5871 ) | ( n5201 & n18658 ) | ( n5871 & n18658 ) ;
  assign n31756 = n15423 ^ n13735 ^ n12673 ;
  assign n31757 = ( n9252 & n31755 ) | ( n9252 & n31756 ) | ( n31755 & n31756 ) ;
  assign n31758 = n26570 ^ n14511 ^ n3568 ;
  assign n31759 = ( n13216 & ~n26483 ) | ( n13216 & n31758 ) | ( ~n26483 & n31758 ) ;
  assign n31760 = ( n5601 & ~n15540 ) | ( n5601 & n28376 ) | ( ~n15540 & n28376 ) ;
  assign n31761 = n11238 ^ n3813 ^ 1'b0 ;
  assign n31762 = ~n23317 & n31761 ;
  assign n31763 = ( ~n963 & n16047 ) | ( ~n963 & n31762 ) | ( n16047 & n31762 ) ;
  assign n31764 = ~n7010 & n31763 ;
  assign n31770 = ~n2237 & n15977 ;
  assign n31768 = n20922 ^ n15303 ^ x231 ;
  assign n31766 = n24667 ^ n21684 ^ n7667 ;
  assign n31765 = n21438 & n27800 ;
  assign n31767 = n31766 ^ n31765 ^ 1'b0 ;
  assign n31769 = n31768 ^ n31767 ^ n8542 ;
  assign n31771 = n31770 ^ n31769 ^ n12053 ;
  assign n31778 = ( ~n1140 & n9299 ) | ( ~n1140 & n16342 ) | ( n9299 & n16342 ) ;
  assign n31772 = n24712 ^ n1499 ^ 1'b0 ;
  assign n31773 = n31772 ^ n9284 ^ 1'b0 ;
  assign n31774 = ( n3739 & n23080 ) | ( n3739 & n31773 ) | ( n23080 & n31773 ) ;
  assign n31775 = n31774 ^ n15524 ^ n1581 ;
  assign n31776 = n8881 | n16088 ;
  assign n31777 = ( n12363 & n31775 ) | ( n12363 & ~n31776 ) | ( n31775 & ~n31776 ) ;
  assign n31779 = n31778 ^ n31777 ^ x231 ;
  assign n31780 = n7095 ^ n4141 ^ 1'b0 ;
  assign n31781 = n31779 | n31780 ;
  assign n31782 = n817 & ~n28996 ;
  assign n31783 = n31782 ^ n23266 ^ n8816 ;
  assign n31784 = ( n13686 & n16817 ) | ( n13686 & ~n31783 ) | ( n16817 & ~n31783 ) ;
  assign n31785 = n31784 ^ n13906 ^ x29 ;
  assign n31786 = n11685 & ~n15133 ;
  assign n31787 = n8835 & ~n9088 ;
  assign n31788 = ~n1095 & n31787 ;
  assign n31789 = n4317 ^ n1845 ^ 1'b0 ;
  assign n31790 = n31723 ^ n19623 ^ 1'b0 ;
  assign n31791 = n11987 | n23908 ;
  assign n31792 = n31791 ^ n10932 ^ 1'b0 ;
  assign n31793 = ( n10932 & n14042 ) | ( n10932 & ~n31792 ) | ( n14042 & ~n31792 ) ;
  assign n31794 = ( n19236 & n31790 ) | ( n19236 & n31793 ) | ( n31790 & n31793 ) ;
  assign n31795 = ( n10191 & ~n21240 ) | ( n10191 & n30321 ) | ( ~n21240 & n30321 ) ;
  assign n31796 = n11280 & ~n31795 ;
  assign n31797 = n11730 & n31796 ;
  assign n31798 = n16334 | n17283 ;
  assign n31799 = n31798 ^ n4145 ^ 1'b0 ;
  assign n31800 = ( n845 & n23253 ) | ( n845 & ~n31799 ) | ( n23253 & ~n31799 ) ;
  assign n31801 = ~n3935 & n23259 ;
  assign n31802 = ~n18777 & n31801 ;
  assign n31803 = ( n6401 & n8938 ) | ( n6401 & n31802 ) | ( n8938 & n31802 ) ;
  assign n31804 = ( n5718 & n7696 ) | ( n5718 & ~n12713 ) | ( n7696 & ~n12713 ) ;
  assign n31805 = n8917 ^ n7693 ^ n7231 ;
  assign n31806 = ( n11242 & n23682 ) | ( n11242 & n31805 ) | ( n23682 & n31805 ) ;
  assign n31807 = n31806 ^ n11126 ^ n5226 ;
  assign n31808 = n31807 ^ n26160 ^ n25441 ;
  assign n31809 = n29884 ^ n24173 ^ n13601 ;
  assign n31810 = n28021 ^ n3873 ^ n2962 ;
  assign n31811 = n21028 ^ n10344 ^ n7058 ;
  assign n31812 = n31811 ^ n25074 ^ 1'b0 ;
  assign n31813 = n25737 | n31812 ;
  assign n31819 = n21183 & ~n21580 ;
  assign n31820 = n31819 ^ n21563 ^ 1'b0 ;
  assign n31821 = n31820 ^ n22411 ^ n16520 ;
  assign n31822 = n31821 ^ n29354 ^ n15390 ;
  assign n31823 = n31822 ^ n2895 ^ 1'b0 ;
  assign n31817 = n16767 ^ n14942 ^ n3243 ;
  assign n31814 = n25412 ^ n2883 ^ n1689 ;
  assign n31815 = n12109 | n31814 ;
  assign n31816 = n31815 ^ n10843 ^ 1'b0 ;
  assign n31818 = n31817 ^ n31816 ^ n10508 ;
  assign n31824 = n31823 ^ n31818 ^ n6267 ;
  assign n31825 = n9042 & ~n22589 ;
  assign n31826 = ~n10604 & n31825 ;
  assign n31827 = n1602 | n31826 ;
  assign n31828 = n6011 & ~n19901 ;
  assign n31829 = ( ~n2679 & n28934 ) | ( ~n2679 & n31828 ) | ( n28934 & n31828 ) ;
  assign n31830 = n31827 & ~n31829 ;
  assign n31831 = n22534 & n31830 ;
  assign n31832 = n29934 ^ n7869 ^ n3105 ;
  assign n31833 = ( n11900 & ~n18609 ) | ( n11900 & n31832 ) | ( ~n18609 & n31832 ) ;
  assign n31834 = x23 & ~n31833 ;
  assign n31835 = ~n31768 & n31834 ;
  assign n31836 = n8963 & ~n23126 ;
  assign n31837 = n31156 & n31836 ;
  assign n31838 = n25108 ^ n18782 ^ n12282 ;
  assign n31839 = ( ~n15423 & n29888 ) | ( ~n15423 & n31621 ) | ( n29888 & n31621 ) ;
  assign n31842 = ( n4794 & n14965 ) | ( n4794 & n19941 ) | ( n14965 & n19941 ) ;
  assign n31840 = ~n13766 & n24379 ;
  assign n31841 = ~n31768 & n31840 ;
  assign n31843 = n31842 ^ n31841 ^ n1963 ;
  assign n31844 = ( n9066 & n12876 ) | ( n9066 & ~n15057 ) | ( n12876 & ~n15057 ) ;
  assign n31845 = n31844 ^ n18865 ^ 1'b0 ;
  assign n31846 = ( n4717 & n12039 ) | ( n4717 & n13146 ) | ( n12039 & n13146 ) ;
  assign n31847 = ( n15912 & n19593 ) | ( n15912 & n31846 ) | ( n19593 & n31846 ) ;
  assign n31848 = n30869 & n31847 ;
  assign n31849 = ( n9766 & n31497 ) | ( n9766 & ~n31848 ) | ( n31497 & ~n31848 ) ;
  assign n31850 = ( n635 & n6672 ) | ( n635 & n12082 ) | ( n6672 & n12082 ) ;
  assign n31851 = n28308 ^ n27390 ^ n5859 ;
  assign n31852 = n30681 ^ n25750 ^ n22935 ;
  assign n31853 = ( n1343 & n4335 ) | ( n1343 & n15106 ) | ( n4335 & n15106 ) ;
  assign n31854 = n31853 ^ n18990 ^ n15070 ;
  assign n31855 = n21447 ^ n7716 ^ 1'b0 ;
  assign n31856 = ( n16465 & ~n28973 ) | ( n16465 & n31855 ) | ( ~n28973 & n31855 ) ;
  assign n31857 = n31856 ^ n25762 ^ 1'b0 ;
  assign n31858 = ( n8222 & ~n12356 ) | ( n8222 & n31857 ) | ( ~n12356 & n31857 ) ;
  assign n31859 = n31858 ^ n16169 ^ n16023 ;
  assign n31860 = n9231 ^ n1684 ^ 1'b0 ;
  assign n31861 = ( ~n912 & n4798 ) | ( ~n912 & n31860 ) | ( n4798 & n31860 ) ;
  assign n31862 = ( ~n6817 & n27310 ) | ( ~n6817 & n31861 ) | ( n27310 & n31861 ) ;
  assign n31864 = n22602 ^ n13977 ^ n9821 ;
  assign n31865 = n31864 ^ n20687 ^ n6340 ;
  assign n31863 = n10690 & ~n30024 ;
  assign n31866 = n31865 ^ n31863 ^ n7907 ;
  assign n31867 = ( n15548 & n19285 ) | ( n15548 & n31866 ) | ( n19285 & n31866 ) ;
  assign n31870 = ~n8220 & n8492 ;
  assign n31871 = ~n8207 & n31870 ;
  assign n31872 = ( n3964 & ~n7023 ) | ( n3964 & n31871 ) | ( ~n7023 & n31871 ) ;
  assign n31868 = n8728 | n10490 ;
  assign n31869 = n31868 ^ n7774 ^ 1'b0 ;
  assign n31873 = n31872 ^ n31869 ^ n7496 ;
  assign n31874 = n2481 & ~n3937 ;
  assign n31875 = n10251 ^ n4608 ^ 1'b0 ;
  assign n31876 = n1204 & ~n31875 ;
  assign n31877 = n31876 ^ n12686 ^ 1'b0 ;
  assign n31878 = n20201 & ~n31877 ;
  assign n31879 = n12724 ^ n4893 ^ n1585 ;
  assign n31880 = ( n1040 & n13145 ) | ( n1040 & n18330 ) | ( n13145 & n18330 ) ;
  assign n31881 = ( n10048 & n11145 ) | ( n10048 & ~n31880 ) | ( n11145 & ~n31880 ) ;
  assign n31882 = ( n21824 & n25875 ) | ( n21824 & n31881 ) | ( n25875 & n31881 ) ;
  assign n31883 = n17278 & ~n17606 ;
  assign n31884 = n31882 & n31883 ;
  assign n31885 = n31884 ^ n7856 ^ n3410 ;
  assign n31886 = ( n1216 & n31879 ) | ( n1216 & ~n31885 ) | ( n31879 & ~n31885 ) ;
  assign n31887 = n6114 ^ n5027 ^ n3006 ;
  assign n31888 = ( n15113 & n19939 ) | ( n15113 & n26157 ) | ( n19939 & n26157 ) ;
  assign n31889 = n8336 & n31888 ;
  assign n31890 = n31887 & n31889 ;
  assign n31891 = ( n10702 & n23873 ) | ( n10702 & ~n31890 ) | ( n23873 & ~n31890 ) ;
  assign n31892 = n23543 ^ n20726 ^ n16152 ;
  assign n31894 = n11163 ^ n3530 ^ n2564 ;
  assign n31893 = n16518 ^ n13336 ^ 1'b0 ;
  assign n31895 = n31894 ^ n31893 ^ n9067 ;
  assign n31896 = ( ~n29797 & n30169 ) | ( ~n29797 & n31895 ) | ( n30169 & n31895 ) ;
  assign n31898 = ( n1535 & n7217 ) | ( n1535 & n19024 ) | ( n7217 & n19024 ) ;
  assign n31897 = n18980 ^ n514 ^ 1'b0 ;
  assign n31899 = n31898 ^ n31897 ^ n18924 ;
  assign n31900 = n19340 ^ n1689 ^ 1'b0 ;
  assign n31901 = ~n4496 & n31900 ;
  assign n31902 = n23686 ^ n18438 ^ n10928 ;
  assign n31903 = x221 & n31902 ;
  assign n31904 = n31903 ^ n6473 ^ 1'b0 ;
  assign n31905 = ( ~n26976 & n31901 ) | ( ~n26976 & n31904 ) | ( n31901 & n31904 ) ;
  assign n31907 = n11412 ^ n8324 ^ n7294 ;
  assign n31906 = n26544 ^ n16831 ^ n774 ;
  assign n31908 = n31907 ^ n31906 ^ n962 ;
  assign n31916 = ( n7828 & n26593 ) | ( n7828 & n29309 ) | ( n26593 & n29309 ) ;
  assign n31912 = n3582 | n7710 ;
  assign n31913 = n15666 ^ n10372 ^ n8040 ;
  assign n31914 = n31913 ^ n10383 ^ n9683 ;
  assign n31915 = n31912 & n31914 ;
  assign n31917 = n31916 ^ n31915 ^ 1'b0 ;
  assign n31918 = ~n13792 & n31917 ;
  assign n31919 = n31918 ^ n28729 ^ 1'b0 ;
  assign n31909 = n13688 & n18314 ;
  assign n31910 = n31909 ^ n3876 ^ 1'b0 ;
  assign n31911 = n14895 & ~n31910 ;
  assign n31920 = n31919 ^ n31911 ^ n18299 ;
  assign n31921 = ( n426 & ~n9229 ) | ( n426 & n23517 ) | ( ~n9229 & n23517 ) ;
  assign n31922 = ( n519 & n1416 ) | ( n519 & ~n2147 ) | ( n1416 & ~n2147 ) ;
  assign n31923 = n16262 & n31922 ;
  assign n31924 = ( n3963 & n16324 ) | ( n3963 & n31923 ) | ( n16324 & n31923 ) ;
  assign n31925 = ( n5453 & ~n31921 ) | ( n5453 & n31924 ) | ( ~n31921 & n31924 ) ;
  assign n31926 = x128 & ~n2930 ;
  assign n31927 = n31926 ^ n23241 ^ n19726 ;
  assign n31928 = ( ~n6969 & n18233 ) | ( ~n6969 & n28996 ) | ( n18233 & n28996 ) ;
  assign n31929 = ~n4864 & n11166 ;
  assign n31930 = n31929 ^ n9945 ^ n6259 ;
  assign n31931 = n31930 ^ n740 ^ x164 ;
  assign n31932 = n5828 & n31931 ;
  assign n31933 = n31932 ^ n26943 ^ 1'b0 ;
  assign n31934 = n6319 | n11622 ;
  assign n31935 = n6171 ^ x68 ^ 1'b0 ;
  assign n31936 = x224 & n31935 ;
  assign n31937 = n12002 ^ n9012 ^ 1'b0 ;
  assign n31938 = n20501 ^ n14038 ^ n2117 ;
  assign n31939 = ( ~n1399 & n31937 ) | ( ~n1399 & n31938 ) | ( n31937 & n31938 ) ;
  assign n31940 = n31936 & ~n31939 ;
  assign n31941 = n28372 ^ n23557 ^ n6626 ;
  assign n31942 = ( n4386 & n22983 ) | ( n4386 & ~n31941 ) | ( n22983 & ~n31941 ) ;
  assign n31943 = n31942 ^ n12890 ^ 1'b0 ;
  assign n31944 = ( n749 & n23302 ) | ( n749 & ~n31943 ) | ( n23302 & ~n31943 ) ;
  assign n31945 = n8219 | n16641 ;
  assign n31947 = n11204 & ~n14569 ;
  assign n31946 = n8633 & n9081 ;
  assign n31948 = n31947 ^ n31946 ^ 1'b0 ;
  assign n31949 = ( n5529 & n11300 ) | ( n5529 & n31948 ) | ( n11300 & n31948 ) ;
  assign n31950 = ( ~n3523 & n27928 ) | ( ~n3523 & n31949 ) | ( n27928 & n31949 ) ;
  assign n31951 = n18921 & n21118 ;
  assign n31952 = ~n8992 & n31951 ;
  assign n31953 = n10126 ^ n2511 ^ 1'b0 ;
  assign n31954 = n11757 & n31953 ;
  assign n31955 = ( ~n17804 & n18060 ) | ( ~n17804 & n31954 ) | ( n18060 & n31954 ) ;
  assign n31956 = n31955 ^ n9906 ^ n2855 ;
  assign n31957 = ( n2687 & ~n27086 ) | ( n2687 & n27881 ) | ( ~n27086 & n27881 ) ;
  assign n31958 = n31806 ^ n28938 ^ n14524 ;
  assign n31959 = n17844 ^ n990 ^ n556 ;
  assign n31960 = ( ~n7137 & n21507 ) | ( ~n7137 & n31959 ) | ( n21507 & n31959 ) ;
  assign n31961 = n10186 ^ n1632 ^ 1'b0 ;
  assign n31962 = ~n4816 & n31961 ;
  assign n31964 = ( n1871 & ~n5963 ) | ( n1871 & n11821 ) | ( ~n5963 & n11821 ) ;
  assign n31965 = n22347 | n31964 ;
  assign n31963 = ( ~n7193 & n21446 ) | ( ~n7193 & n29963 ) | ( n21446 & n29963 ) ;
  assign n31966 = n31965 ^ n31963 ^ n4554 ;
  assign n31967 = n2077 & ~n8694 ;
  assign n31968 = n31967 ^ n7295 ^ 1'b0 ;
  assign n31969 = ( n19021 & ~n19869 ) | ( n19021 & n31968 ) | ( ~n19869 & n31968 ) ;
  assign n31970 = n10289 | n11324 ;
  assign n31971 = n31970 ^ n28562 ^ 1'b0 ;
  assign n31972 = ( n12779 & n29572 ) | ( n12779 & n31971 ) | ( n29572 & n31971 ) ;
  assign n31973 = n26306 ^ n16972 ^ 1'b0 ;
  assign n31974 = n26525 | n31973 ;
  assign n31975 = n28585 ^ n16760 ^ n11804 ;
  assign n31976 = ( n23774 & n24901 ) | ( n23774 & ~n31975 ) | ( n24901 & ~n31975 ) ;
  assign n31977 = ( n4763 & ~n10405 ) | ( n4763 & n23299 ) | ( ~n10405 & n23299 ) ;
  assign n31978 = n31977 ^ n11375 ^ n5118 ;
  assign n31979 = n26173 ^ n3100 ^ n1581 ;
  assign n31980 = n28735 ^ n6507 ^ n1854 ;
  assign n31981 = ( n17242 & n31979 ) | ( n17242 & ~n31980 ) | ( n31979 & ~n31980 ) ;
  assign n31982 = ( ~n17186 & n23463 ) | ( ~n17186 & n31981 ) | ( n23463 & n31981 ) ;
  assign n31983 = n28194 ^ n24753 ^ n2814 ;
  assign n31984 = n10610 & ~n31983 ;
  assign n31985 = n29583 & n31984 ;
  assign n31986 = ( x244 & ~n31982 ) | ( x244 & n31985 ) | ( ~n31982 & n31985 ) ;
  assign n31987 = n18137 & n18444 ;
  assign n31988 = n3491 & n31987 ;
  assign n31989 = n18302 ^ n14334 ^ n5512 ;
  assign n31990 = ( n1390 & n31529 ) | ( n1390 & ~n31989 ) | ( n31529 & ~n31989 ) ;
  assign n31991 = n10301 ^ n2794 ^ 1'b0 ;
  assign n31992 = n11811 | n31991 ;
  assign n31993 = ( n3096 & ~n8885 ) | ( n3096 & n31992 ) | ( ~n8885 & n31992 ) ;
  assign n31994 = n31993 ^ n22058 ^ n11458 ;
  assign n31995 = n17301 & ~n22833 ;
  assign n31996 = ( n13930 & n24819 ) | ( n13930 & ~n31995 ) | ( n24819 & ~n31995 ) ;
  assign n31997 = ( ~n13875 & n17957 ) | ( ~n13875 & n26881 ) | ( n17957 & n26881 ) ;
  assign n31998 = n28489 ^ n9037 ^ n5212 ;
  assign n31999 = ( ~n6071 & n31997 ) | ( ~n6071 & n31998 ) | ( n31997 & n31998 ) ;
  assign n32000 = ( ~n2301 & n16390 ) | ( ~n2301 & n21562 ) | ( n16390 & n21562 ) ;
  assign n32001 = ( n23807 & n31999 ) | ( n23807 & n32000 ) | ( n31999 & n32000 ) ;
  assign n32010 = n11858 & ~n13660 ;
  assign n32002 = n3585 | n6584 ;
  assign n32003 = n13317 | n32002 ;
  assign n32004 = n32003 ^ n8933 ^ n7253 ;
  assign n32005 = n32004 ^ n21911 ^ n2834 ;
  assign n32006 = n32005 ^ n20430 ^ n11540 ;
  assign n32007 = n7468 & ~n32006 ;
  assign n32008 = n32007 ^ n2083 ^ 1'b0 ;
  assign n32009 = ~n1742 & n32008 ;
  assign n32011 = n32010 ^ n32009 ^ n28585 ;
  assign n32013 = n4506 & ~n5689 ;
  assign n32014 = ~n1647 & n32013 ;
  assign n32015 = ( n2626 & n11493 ) | ( n2626 & ~n32014 ) | ( n11493 & ~n32014 ) ;
  assign n32016 = n20783 & ~n32015 ;
  assign n32017 = n11722 & n32016 ;
  assign n32012 = n7622 & n7891 ;
  assign n32018 = n32017 ^ n32012 ^ 1'b0 ;
  assign n32019 = n25419 ^ n13823 ^ n11243 ;
  assign n32020 = n32019 ^ n19233 ^ 1'b0 ;
  assign n32021 = n16300 ^ n12477 ^ n1976 ;
  assign n32022 = n32021 ^ n9350 ^ n6131 ;
  assign n32023 = n32022 ^ n22505 ^ n3250 ;
  assign n32024 = n32023 ^ n31955 ^ n16269 ;
  assign n32025 = n30539 ^ n14839 ^ n9969 ;
  assign n32026 = ( n4708 & n7120 ) | ( n4708 & ~n7780 ) | ( n7120 & ~n7780 ) ;
  assign n32027 = n32026 ^ n18278 ^ n6897 ;
  assign n32028 = ( n6080 & n32025 ) | ( n6080 & n32027 ) | ( n32025 & n32027 ) ;
  assign n32029 = ~n12738 & n18237 ;
  assign n32030 = n4246 | n6257 ;
  assign n32031 = n32030 ^ n3807 ^ 1'b0 ;
  assign n32032 = ~n3110 & n23785 ;
  assign n32033 = n32031 & n32032 ;
  assign n32034 = ( n3231 & n14818 ) | ( n3231 & ~n32033 ) | ( n14818 & ~n32033 ) ;
  assign n32038 = ~n5532 & n17079 ;
  assign n32036 = n12775 ^ n12205 ^ n7698 ;
  assign n32035 = n11403 ^ n11129 ^ n7891 ;
  assign n32037 = n32036 ^ n32035 ^ n19400 ;
  assign n32039 = n32038 ^ n32037 ^ 1'b0 ;
  assign n32040 = n7733 & n8303 ;
  assign n32041 = n25069 & n32040 ;
  assign n32042 = n32041 ^ n6549 ^ 1'b0 ;
  assign n32043 = ~n31493 & n32042 ;
  assign n32044 = n1110 & ~n15475 ;
  assign n32045 = n32044 ^ n20629 ^ 1'b0 ;
  assign n32046 = n2263 & n32045 ;
  assign n32047 = ( n12218 & n32015 ) | ( n12218 & n32046 ) | ( n32015 & n32046 ) ;
  assign n32048 = n13954 | n32047 ;
  assign n32049 = n8555 & ~n32048 ;
  assign n32050 = n10045 ^ n7417 ^ n4211 ;
  assign n32051 = n32050 ^ n23311 ^ n21921 ;
  assign n32052 = ( ~n6467 & n27327 ) | ( ~n6467 & n32051 ) | ( n27327 & n32051 ) ;
  assign n32053 = n14545 ^ n3358 ^ n2130 ;
  assign n32054 = ~n8694 & n26008 ;
  assign n32055 = ( ~n7551 & n8209 ) | ( ~n7551 & n32054 ) | ( n8209 & n32054 ) ;
  assign n32056 = ( n18766 & n21997 ) | ( n18766 & n32055 ) | ( n21997 & n32055 ) ;
  assign n32057 = n14120 & ~n32056 ;
  assign n32058 = ~n19332 & n32057 ;
  assign n32059 = n20312 ^ n5134 ^ 1'b0 ;
  assign n32060 = n28827 & n32059 ;
  assign n32061 = n32060 ^ n30016 ^ 1'b0 ;
  assign n32067 = n7762 | n8983 ;
  assign n32068 = n5805 & ~n32067 ;
  assign n32064 = n6917 | n16060 ;
  assign n32062 = ( n1117 & n18802 ) | ( n1117 & ~n23412 ) | ( n18802 & ~n23412 ) ;
  assign n32063 = ~n29832 & n32062 ;
  assign n32065 = n32064 ^ n32063 ^ 1'b0 ;
  assign n32066 = ~n18626 & n32065 ;
  assign n32069 = n32068 ^ n32066 ^ 1'b0 ;
  assign n32070 = ( n10211 & n17504 ) | ( n10211 & n18495 ) | ( n17504 & n18495 ) ;
  assign n32071 = ( ~n13346 & n22024 ) | ( ~n13346 & n28427 ) | ( n22024 & n28427 ) ;
  assign n32072 = ( n4773 & n6502 ) | ( n4773 & n8422 ) | ( n6502 & n8422 ) ;
  assign n32073 = n6288 & n7067 ;
  assign n32074 = ( n25745 & n32072 ) | ( n25745 & ~n32073 ) | ( n32072 & ~n32073 ) ;
  assign n32075 = ( n27120 & ~n32071 ) | ( n27120 & n32074 ) | ( ~n32071 & n32074 ) ;
  assign n32076 = ( n1774 & ~n15244 ) | ( n1774 & n16629 ) | ( ~n15244 & n16629 ) ;
  assign n32077 = n32076 ^ n31481 ^ n24581 ;
  assign n32078 = ( ~n7523 & n11331 ) | ( ~n7523 & n29831 ) | ( n11331 & n29831 ) ;
  assign n32079 = ( n13273 & n23953 ) | ( n13273 & n28107 ) | ( n23953 & n28107 ) ;
  assign n32080 = ( n17843 & n32078 ) | ( n17843 & ~n32079 ) | ( n32078 & ~n32079 ) ;
  assign n32081 = ( n32075 & n32077 ) | ( n32075 & ~n32080 ) | ( n32077 & ~n32080 ) ;
  assign n32082 = n5429 ^ n986 ^ 1'b0 ;
  assign n32083 = n23928 & ~n32082 ;
  assign n32084 = n10270 ^ n2570 ^ 1'b0 ;
  assign n32085 = n32083 | n32084 ;
  assign n32086 = n8462 ^ n7252 ^ n3305 ;
  assign n32087 = n32086 ^ n18739 ^ n3383 ;
  assign n32088 = n31481 ^ n28830 ^ n8700 ;
  assign n32089 = ( n11634 & ~n32087 ) | ( n11634 & n32088 ) | ( ~n32087 & n32088 ) ;
  assign n32090 = ~n20955 & n32089 ;
  assign n32091 = n32090 ^ n29295 ^ 1'b0 ;
  assign n32092 = n10219 & ~n32091 ;
  assign n32093 = n2317 | n16118 ;
  assign n32094 = n2300 | n31939 ;
  assign n32095 = n27180 & ~n32094 ;
  assign n32096 = n32095 ^ n5189 ^ 1'b0 ;
  assign n32097 = n32096 ^ n19813 ^ n3706 ;
  assign n32098 = n10608 ^ n7045 ^ n3834 ;
  assign n32099 = n18993 | n32098 ;
  assign n32100 = n24299 ^ n8768 ^ n8156 ;
  assign n32101 = ( n707 & n3977 ) | ( n707 & n22576 ) | ( n3977 & n22576 ) ;
  assign n32102 = n26814 ^ n4697 ^ n2562 ;
  assign n32103 = x57 & n32102 ;
  assign n32104 = n32103 ^ n19882 ^ 1'b0 ;
  assign n32105 = n27521 ^ n21002 ^ n7842 ;
  assign n32106 = n26053 ^ n10276 ^ n7394 ;
  assign n32107 = ( n8910 & n32105 ) | ( n8910 & ~n32106 ) | ( n32105 & ~n32106 ) ;
  assign n32108 = ~n23475 & n32107 ;
  assign n32109 = n32108 ^ n4569 ^ 1'b0 ;
  assign n32115 = n10881 ^ n4573 ^ n3696 ;
  assign n32114 = n26370 ^ n18596 ^ 1'b0 ;
  assign n32110 = n19612 ^ n15373 ^ n9748 ;
  assign n32111 = n5689 | n31846 ;
  assign n32112 = n32110 | n32111 ;
  assign n32113 = n32112 ^ n20251 ^ n588 ;
  assign n32116 = n32115 ^ n32114 ^ n32113 ;
  assign n32117 = n32116 ^ n7450 ^ n5414 ;
  assign n32118 = n22462 ^ n15478 ^ n15232 ;
  assign n32119 = n32118 ^ n8849 ^ n6709 ;
  assign n32123 = n17878 ^ n13011 ^ n5483 ;
  assign n32120 = n1203 & ~n16956 ;
  assign n32121 = n3849 & n32120 ;
  assign n32122 = n32121 ^ n23432 ^ n12337 ;
  assign n32124 = n32123 ^ n32122 ^ n5190 ;
  assign n32125 = ~n13694 & n19628 ;
  assign n32126 = ( n13319 & n32124 ) | ( n13319 & ~n32125 ) | ( n32124 & ~n32125 ) ;
  assign n32127 = ( n3094 & n9676 ) | ( n3094 & ~n21193 ) | ( n9676 & ~n21193 ) ;
  assign n32128 = ( n5538 & ~n8219 ) | ( n5538 & n9222 ) | ( ~n8219 & n9222 ) ;
  assign n32129 = n32128 ^ n5419 ^ n4987 ;
  assign n32130 = n32129 ^ n13503 ^ n6102 ;
  assign n32131 = n13586 ^ n12111 ^ n6376 ;
  assign n32132 = n32131 ^ n11410 ^ n11361 ;
  assign n32133 = ~n4208 & n20953 ;
  assign n32134 = n4187 & n32133 ;
  assign n32135 = n16378 | n28442 ;
  assign n32136 = n32134 & ~n32135 ;
  assign n32137 = n14181 ^ n1092 ^ n965 ;
  assign n32138 = n32137 ^ n11940 ^ n868 ;
  assign n32139 = n32138 ^ n16377 ^ 1'b0 ;
  assign n32140 = n20540 | n32139 ;
  assign n32141 = n32140 ^ n29117 ^ n2919 ;
  assign n32142 = n22382 ^ n18177 ^ n3487 ;
  assign n32143 = n26058 ^ n13528 ^ n2647 ;
  assign n32144 = ( n10114 & ~n20902 ) | ( n10114 & n32143 ) | ( ~n20902 & n32143 ) ;
  assign n32147 = n24664 ^ n15397 ^ n4947 ;
  assign n32145 = n10504 & ~n11895 ;
  assign n32146 = n22611 & ~n32145 ;
  assign n32148 = n32147 ^ n32146 ^ 1'b0 ;
  assign n32149 = ( n6669 & ~n12551 ) | ( n6669 & n13073 ) | ( ~n12551 & n13073 ) ;
  assign n32150 = n32149 ^ n15232 ^ n10643 ;
  assign n32151 = n5480 | n8684 ;
  assign n32152 = n32151 ^ n8193 ^ 1'b0 ;
  assign n32153 = n32152 ^ n12986 ^ 1'b0 ;
  assign n32154 = n32150 & ~n32153 ;
  assign n32155 = ~n9821 & n18672 ;
  assign n32156 = n20776 ^ n4614 ^ 1'b0 ;
  assign n32157 = ( n6948 & ~n32155 ) | ( n6948 & n32156 ) | ( ~n32155 & n32156 ) ;
  assign n32163 = n9857 & n28487 ;
  assign n32164 = n32163 ^ n16696 ^ 1'b0 ;
  assign n32158 = ( n5297 & n8642 ) | ( n5297 & ~n26539 ) | ( n8642 & ~n26539 ) ;
  assign n32159 = n32158 ^ n14843 ^ 1'b0 ;
  assign n32160 = ~n5091 & n32159 ;
  assign n32161 = n32160 ^ n7775 ^ 1'b0 ;
  assign n32162 = ( n6597 & n14799 ) | ( n6597 & ~n32161 ) | ( n14799 & ~n32161 ) ;
  assign n32165 = n32164 ^ n32162 ^ 1'b0 ;
  assign n32166 = ( ~n1703 & n12202 ) | ( ~n1703 & n32165 ) | ( n12202 & n32165 ) ;
  assign n32167 = n20750 ^ n6805 ^ n4754 ;
  assign n32168 = n9441 ^ n8753 ^ 1'b0 ;
  assign n32169 = n10302 | n32168 ;
  assign n32170 = n22347 & ~n32169 ;
  assign n32171 = n24352 ^ n15773 ^ n5134 ;
  assign n32172 = n20308 | n25263 ;
  assign n32173 = n19771 & ~n32172 ;
  assign n32174 = n32171 | n32173 ;
  assign n32175 = n32174 ^ n1334 ^ 1'b0 ;
  assign n32176 = n20814 ^ x105 ^ 1'b0 ;
  assign n32177 = n7382 ^ n2820 ^ n296 ;
  assign n32178 = n32177 ^ n19779 ^ 1'b0 ;
  assign n32179 = ~n8958 & n32178 ;
  assign n32180 = n32179 ^ n19557 ^ n11350 ;
  assign n32181 = n32180 ^ n5315 ^ 1'b0 ;
  assign n32182 = ~n6971 & n32181 ;
  assign n32183 = n32182 ^ n26700 ^ n5496 ;
  assign n32184 = n1760 | n9683 ;
  assign n32185 = n32184 ^ n728 ^ 1'b0 ;
  assign n32186 = ( n6858 & n21236 ) | ( n6858 & n32185 ) | ( n21236 & n32185 ) ;
  assign n32187 = n32186 ^ n6256 ^ n4061 ;
  assign n32188 = ( n3783 & n27232 ) | ( n3783 & n32187 ) | ( n27232 & n32187 ) ;
  assign n32189 = ( ~x213 & n768 ) | ( ~x213 & n21713 ) | ( n768 & n21713 ) ;
  assign n32190 = n14751 & n20227 ;
  assign n32191 = ( ~n9631 & n32189 ) | ( ~n9631 & n32190 ) | ( n32189 & n32190 ) ;
  assign n32192 = n23402 ^ n16857 ^ n6994 ;
  assign n32193 = n32192 ^ n31817 ^ 1'b0 ;
  assign n32195 = ( n5504 & ~n16676 ) | ( n5504 & n27292 ) | ( ~n16676 & n27292 ) ;
  assign n32196 = n32195 ^ n17368 ^ n15203 ;
  assign n32194 = n1977 & ~n20660 ;
  assign n32197 = n32196 ^ n32194 ^ 1'b0 ;
  assign n32198 = ( n14048 & ~n18318 ) | ( n14048 & n32197 ) | ( ~n18318 & n32197 ) ;
  assign n32199 = n32198 ^ n19509 ^ n9737 ;
  assign n32200 = ( n8054 & ~n28761 ) | ( n8054 & n28872 ) | ( ~n28761 & n28872 ) ;
  assign n32201 = n32102 ^ n4180 ^ 1'b0 ;
  assign n32202 = n31390 & ~n32201 ;
  assign n32203 = ( n5208 & n14955 ) | ( n5208 & n25910 ) | ( n14955 & n25910 ) ;
  assign n32204 = n22870 & ~n32203 ;
  assign n32205 = n15355 & n32204 ;
  assign n32206 = n7930 ^ n6302 ^ n4403 ;
  assign n32207 = n32206 ^ n27404 ^ n2746 ;
  assign n32208 = n31841 ^ n26387 ^ n25991 ;
  assign n32213 = n12295 ^ n8172 ^ x190 ;
  assign n32214 = n32213 ^ n20843 ^ n10970 ;
  assign n32209 = n14621 ^ n14352 ^ 1'b0 ;
  assign n32210 = ( n18283 & ~n22323 ) | ( n18283 & n26958 ) | ( ~n22323 & n26958 ) ;
  assign n32211 = n32210 ^ n11094 ^ n8182 ;
  assign n32212 = ( n14882 & n32209 ) | ( n14882 & ~n32211 ) | ( n32209 & ~n32211 ) ;
  assign n32215 = n32214 ^ n32212 ^ n29977 ;
  assign n32218 = n1499 | n8742 ;
  assign n32216 = n10112 & ~n16053 ;
  assign n32217 = ( n21488 & ~n23838 ) | ( n21488 & n32216 ) | ( ~n23838 & n32216 ) ;
  assign n32219 = n32218 ^ n32217 ^ n24834 ;
  assign n32220 = ( n8885 & n10028 ) | ( n8885 & ~n27619 ) | ( n10028 & ~n27619 ) ;
  assign n32221 = n32220 ^ n27272 ^ n10045 ;
  assign n32222 = n9353 & ~n17693 ;
  assign n32223 = ~n12005 & n32222 ;
  assign n32224 = n32223 ^ n13631 ^ n11035 ;
  assign n32225 = ( ~n11687 & n26251 ) | ( ~n11687 & n32224 ) | ( n26251 & n32224 ) ;
  assign n32226 = n21053 & n21916 ;
  assign n32227 = n21648 | n32226 ;
  assign n32228 = n32225 & ~n32227 ;
  assign n32229 = n17555 ^ n10957 ^ n5964 ;
  assign n32230 = n32229 ^ n14417 ^ 1'b0 ;
  assign n32231 = n24540 ^ n10828 ^ n4956 ;
  assign n32233 = n26167 ^ n11551 ^ n6621 ;
  assign n32232 = n12801 & ~n16562 ;
  assign n32234 = n32233 ^ n32232 ^ 1'b0 ;
  assign n32235 = n16561 ^ n5575 ^ n328 ;
  assign n32236 = n32235 ^ n14567 ^ n12361 ;
  assign n32237 = n32236 ^ n12804 ^ n1737 ;
  assign n32238 = n19985 ^ n16103 ^ 1'b0 ;
  assign n32239 = ( n337 & n6691 ) | ( n337 & n22249 ) | ( n6691 & n22249 ) ;
  assign n32240 = n24521 ^ n19008 ^ n2102 ;
  assign n32246 = ( n6468 & n8203 ) | ( n6468 & n12562 ) | ( n8203 & n12562 ) ;
  assign n32243 = ( n8701 & ~n11822 ) | ( n8701 & n30078 ) | ( ~n11822 & n30078 ) ;
  assign n32244 = ( n7850 & n30324 ) | ( n7850 & n32243 ) | ( n30324 & n32243 ) ;
  assign n32245 = ( n6622 & n18825 ) | ( n6622 & ~n32244 ) | ( n18825 & ~n32244 ) ;
  assign n32241 = n22266 ^ n8532 ^ n1325 ;
  assign n32242 = ( ~n3057 & n18346 ) | ( ~n3057 & n32241 ) | ( n18346 & n32241 ) ;
  assign n32247 = n32246 ^ n32245 ^ n32242 ;
  assign n32248 = ( n1335 & ~n4853 ) | ( n1335 & n14893 ) | ( ~n4853 & n14893 ) ;
  assign n32249 = n32248 ^ n14543 ^ 1'b0 ;
  assign n32250 = ( n2275 & n21557 ) | ( n2275 & n32249 ) | ( n21557 & n32249 ) ;
  assign n32251 = n25868 ^ n3721 ^ 1'b0 ;
  assign n32252 = ( n451 & n9760 ) | ( n451 & ~n19062 ) | ( n9760 & ~n19062 ) ;
  assign n32253 = ( n4237 & n30634 ) | ( n4237 & n32252 ) | ( n30634 & n32252 ) ;
  assign n32254 = n32253 ^ n16602 ^ n2715 ;
  assign n32255 = n32254 ^ n30925 ^ n6639 ;
  assign n32256 = ( n7390 & n16404 ) | ( n7390 & ~n21428 ) | ( n16404 & ~n21428 ) ;
  assign n32257 = n32256 ^ n6232 ^ n2029 ;
  assign n32258 = n24985 ^ n4374 ^ 1'b0 ;
  assign n32259 = n4360 & n32258 ;
  assign n32260 = n32259 ^ n24604 ^ n19718 ;
  assign n32261 = ( n2257 & n9330 ) | ( n2257 & ~n31111 ) | ( n9330 & ~n31111 ) ;
  assign n32262 = n32261 ^ n19145 ^ 1'b0 ;
  assign n32263 = ~n32260 & n32262 ;
  assign n32264 = n12690 ^ n4150 ^ n792 ;
  assign n32265 = ( n4353 & n12335 ) | ( n4353 & ~n32264 ) | ( n12335 & ~n32264 ) ;
  assign n32266 = ( n6100 & n12716 ) | ( n6100 & n15425 ) | ( n12716 & n15425 ) ;
  assign n32267 = n32266 ^ n13414 ^ n5915 ;
  assign n32268 = ( n766 & n10117 ) | ( n766 & n20316 ) | ( n10117 & n20316 ) ;
  assign n32269 = n32268 ^ n7159 ^ n3823 ;
  assign n32270 = ( n2097 & ~n7862 ) | ( n2097 & n14843 ) | ( ~n7862 & n14843 ) ;
  assign n32271 = ( ~n5297 & n17743 ) | ( ~n5297 & n32270 ) | ( n17743 & n32270 ) ;
  assign n32272 = ( x78 & ~n17139 ) | ( x78 & n31992 ) | ( ~n17139 & n31992 ) ;
  assign n32273 = ( n14970 & ~n23573 ) | ( n14970 & n23801 ) | ( ~n23573 & n23801 ) ;
  assign n32274 = n32273 ^ n24537 ^ 1'b0 ;
  assign n32275 = n11880 ^ n8365 ^ n4210 ;
  assign n32276 = ( ~n9926 & n15113 ) | ( ~n9926 & n32275 ) | ( n15113 & n32275 ) ;
  assign n32277 = ( n9250 & ~n18547 ) | ( n9250 & n31548 ) | ( ~n18547 & n31548 ) ;
  assign n32278 = ( n523 & n1935 ) | ( n523 & ~n27834 ) | ( n1935 & ~n27834 ) ;
  assign n32280 = n5745 ^ n4590 ^ n1793 ;
  assign n32279 = n14985 | n24826 ;
  assign n32281 = n32280 ^ n32279 ^ 1'b0 ;
  assign n32282 = n1595 & n14813 ;
  assign n32283 = ( n892 & n23987 ) | ( n892 & n32282 ) | ( n23987 & n32282 ) ;
  assign n32284 = ( n6408 & n12207 ) | ( n6408 & n31257 ) | ( n12207 & n31257 ) ;
  assign n32285 = n32284 ^ n26200 ^ n25312 ;
  assign n32286 = n5474 ^ n1556 ^ n600 ;
  assign n32287 = n19877 & ~n25603 ;
  assign n32288 = ~n32286 & n32287 ;
  assign n32289 = n7662 | n32288 ;
  assign n32290 = n32289 ^ n31558 ^ n19721 ;
  assign n32291 = n21793 ^ n3130 ^ n1638 ;
  assign n32293 = n15775 ^ n10979 ^ n8121 ;
  assign n32294 = n1344 | n32293 ;
  assign n32295 = n4988 & ~n32294 ;
  assign n32296 = ( ~n1528 & n21439 ) | ( ~n1528 & n32295 ) | ( n21439 & n32295 ) ;
  assign n32292 = n25231 ^ n6572 ^ 1'b0 ;
  assign n32297 = n32296 ^ n32292 ^ n23016 ;
  assign n32298 = ( n1866 & n23774 ) | ( n1866 & ~n32297 ) | ( n23774 & ~n32297 ) ;
  assign n32299 = n16299 ^ n3746 ^ 1'b0 ;
  assign n32300 = n32299 ^ n10196 ^ n1123 ;
  assign n32301 = n32300 ^ n16767 ^ n6497 ;
  assign n32302 = n32301 ^ n3503 ^ n1138 ;
  assign n32303 = n5408 | n12776 ;
  assign n32304 = ( n13048 & n23430 ) | ( n13048 & ~n32303 ) | ( n23430 & ~n32303 ) ;
  assign n32305 = n32304 ^ n4128 ^ 1'b0 ;
  assign n32306 = ( n16642 & ~n32302 ) | ( n16642 & n32305 ) | ( ~n32302 & n32305 ) ;
  assign n32313 = n2992 & n4132 ;
  assign n32307 = n7330 & ~n8665 ;
  assign n32308 = n9787 ^ n2842 ^ 1'b0 ;
  assign n32309 = n2744 & n32308 ;
  assign n32310 = n32309 ^ n6120 ^ n2097 ;
  assign n32311 = ( n18690 & ~n32307 ) | ( n18690 & n32310 ) | ( ~n32307 & n32310 ) ;
  assign n32312 = n32311 ^ n29156 ^ 1'b0 ;
  assign n32314 = n32313 ^ n32312 ^ n2971 ;
  assign n32315 = ~n11634 & n12076 ;
  assign n32316 = ~n1396 & n32315 ;
  assign n32317 = n32316 ^ n25165 ^ n14730 ;
  assign n32318 = n12782 & n30597 ;
  assign n32319 = n11654 & n32318 ;
  assign n32320 = ( n29474 & n31539 ) | ( n29474 & n32319 ) | ( n31539 & n32319 ) ;
  assign n32321 = n23417 ^ n22955 ^ n1560 ;
  assign n32322 = n18956 & ~n32321 ;
  assign n32323 = ~n7681 & n32322 ;
  assign n32324 = n11674 ^ n7613 ^ n7217 ;
  assign n32325 = ( ~n3878 & n24096 ) | ( ~n3878 & n32324 ) | ( n24096 & n32324 ) ;
  assign n32326 = n501 & ~n32325 ;
  assign n32327 = n32326 ^ n16785 ^ 1'b0 ;
  assign n32328 = ( n854 & n14349 ) | ( n854 & ~n17038 ) | ( n14349 & ~n17038 ) ;
  assign n32329 = n32328 ^ n7398 ^ 1'b0 ;
  assign n32330 = n32329 ^ n25388 ^ n19642 ;
  assign n32331 = ( ~n4230 & n29485 ) | ( ~n4230 & n30622 ) | ( n29485 & n30622 ) ;
  assign n32333 = n20223 ^ n4857 ^ 1'b0 ;
  assign n32334 = ~n2831 & n32333 ;
  assign n32332 = ( n8096 & n16145 ) | ( n8096 & n18114 ) | ( n16145 & n18114 ) ;
  assign n32335 = n32334 ^ n32332 ^ n22742 ;
  assign n32336 = n32335 ^ n20159 ^ n11048 ;
  assign n32337 = ( ~n6875 & n9216 ) | ( ~n6875 & n21977 ) | ( n9216 & n21977 ) ;
  assign n32338 = ( n8190 & ~n21420 ) | ( n8190 & n32337 ) | ( ~n21420 & n32337 ) ;
  assign n32339 = n19280 ^ n2169 ^ 1'b0 ;
  assign n32340 = n32339 ^ n12842 ^ 1'b0 ;
  assign n32341 = n32338 & ~n32340 ;
  assign n32342 = n32341 ^ n12419 ^ n5657 ;
  assign n32343 = n18104 ^ n9421 ^ 1'b0 ;
  assign n32344 = n3984 & ~n23726 ;
  assign n32345 = ~n32343 & n32344 ;
  assign n32346 = n21871 ^ n10176 ^ n7572 ;
  assign n32347 = ( ~n2894 & n4753 ) | ( ~n2894 & n32346 ) | ( n4753 & n32346 ) ;
  assign n32348 = n32347 ^ n13226 ^ 1'b0 ;
  assign n32349 = n11215 & ~n18968 ;
  assign n32350 = ~n3790 & n32349 ;
  assign n32351 = n32350 ^ n336 ^ 1'b0 ;
  assign n32352 = x215 & ~n16044 ;
  assign n32353 = ~n24649 & n32352 ;
  assign n32354 = ( ~n4321 & n9773 ) | ( ~n4321 & n32353 ) | ( n9773 & n32353 ) ;
  assign n32355 = n32354 ^ n25720 ^ n2891 ;
  assign n32357 = ~n19031 & n25141 ;
  assign n32358 = n32357 ^ n21183 ^ 1'b0 ;
  assign n32356 = n10275 | n15235 ;
  assign n32359 = n32358 ^ n32356 ^ 1'b0 ;
  assign n32360 = n32359 ^ n18635 ^ 1'b0 ;
  assign n32368 = n27189 ^ n12046 ^ n3673 ;
  assign n32364 = n21543 ^ n9659 ^ n4665 ;
  assign n32365 = ( ~n13194 & n15548 ) | ( ~n13194 & n32364 ) | ( n15548 & n32364 ) ;
  assign n32366 = n32365 ^ n11888 ^ 1'b0 ;
  assign n32367 = ( n6948 & n14400 ) | ( n6948 & ~n32366 ) | ( n14400 & ~n32366 ) ;
  assign n32369 = n32368 ^ n32367 ^ n10830 ;
  assign n32362 = n29257 & n29729 ;
  assign n32361 = n4797 | n6175 ;
  assign n32363 = n32362 ^ n32361 ^ n8887 ;
  assign n32370 = n32369 ^ n32363 ^ n3022 ;
  assign n32371 = n32370 ^ n17985 ^ n1085 ;
  assign n32372 = n25112 ^ n21065 ^ 1'b0 ;
  assign n32373 = n2484 | n32372 ;
  assign n32374 = n32373 ^ n5886 ^ x17 ;
  assign n32381 = n18185 | n20337 ;
  assign n32382 = n5606 | n32381 ;
  assign n32375 = ( x179 & n5814 ) | ( x179 & n13860 ) | ( n5814 & n13860 ) ;
  assign n32376 = ( n2973 & n7856 ) | ( n2973 & ~n32375 ) | ( n7856 & ~n32375 ) ;
  assign n32377 = n32376 ^ n28345 ^ n25314 ;
  assign n32378 = n22282 ^ n21308 ^ n13113 ;
  assign n32379 = n32378 ^ n17969 ^ n5497 ;
  assign n32380 = ( n10864 & ~n32377 ) | ( n10864 & n32379 ) | ( ~n32377 & n32379 ) ;
  assign n32383 = n32382 ^ n32380 ^ n5379 ;
  assign n32384 = n27794 ^ n7145 ^ 1'b0 ;
  assign n32385 = n28438 | n32384 ;
  assign n32386 = n31144 ^ n4667 ^ 1'b0 ;
  assign n32387 = n9309 & ~n32386 ;
  assign n32388 = n32385 | n32387 ;
  assign n32389 = n6900 & ~n23677 ;
  assign n32390 = ~n32388 & n32389 ;
  assign n32391 = n24539 ^ n3339 ^ n1432 ;
  assign n32392 = ~n5632 & n32391 ;
  assign n32393 = n32392 ^ n28388 ^ 1'b0 ;
  assign n32394 = ( ~n8555 & n11820 ) | ( ~n8555 & n15025 ) | ( n11820 & n15025 ) ;
  assign n32395 = n18831 ^ n16334 ^ 1'b0 ;
  assign n32396 = n2932 & n32395 ;
  assign n32397 = ~n32394 & n32396 ;
  assign n32398 = n22180 ^ n19507 ^ n14767 ;
  assign n32399 = ( n2698 & ~n14419 ) | ( n2698 & n32398 ) | ( ~n14419 & n32398 ) ;
  assign n32403 = n17753 ^ n15675 ^ n9001 ;
  assign n32400 = ( ~n2791 & n7227 ) | ( ~n2791 & n12675 ) | ( n7227 & n12675 ) ;
  assign n32401 = n32400 ^ n19724 ^ n3718 ;
  assign n32402 = n16830 & ~n32401 ;
  assign n32404 = n32403 ^ n32402 ^ 1'b0 ;
  assign n32405 = n27119 ^ n21312 ^ n16677 ;
  assign n32406 = n21657 ^ n18193 ^ n7255 ;
  assign n32407 = ( n2105 & n18274 ) | ( n2105 & ~n32406 ) | ( n18274 & ~n32406 ) ;
  assign n32408 = n1983 & n10320 ;
  assign n32409 = n32408 ^ n16979 ^ 1'b0 ;
  assign n32410 = n23710 ^ n17301 ^ n11081 ;
  assign n32411 = n17181 ^ n9218 ^ x20 ;
  assign n32412 = n11455 & ~n13441 ;
  assign n32413 = n9517 & ~n32412 ;
  assign n32414 = n27125 & n32413 ;
  assign n32415 = ~n13351 & n17969 ;
  assign n32416 = ~n19117 & n32415 ;
  assign n32417 = ( n8582 & n8962 ) | ( n8582 & ~n16467 ) | ( n8962 & ~n16467 ) ;
  assign n32418 = n32416 | n32417 ;
  assign n32419 = n32418 ^ n19377 ^ 1'b0 ;
  assign n32420 = ~n32414 & n32419 ;
  assign n32421 = ( ~x173 & n21965 ) | ( ~x173 & n30807 ) | ( n21965 & n30807 ) ;
  assign n32422 = ( n4070 & ~n6778 ) | ( n4070 & n9432 ) | ( ~n6778 & n9432 ) ;
  assign n32423 = n32422 ^ n5658 ^ 1'b0 ;
  assign n32424 = n32421 | n32423 ;
  assign n32425 = ( ~n13783 & n14127 ) | ( ~n13783 & n15175 ) | ( n14127 & n15175 ) ;
  assign n32426 = ( n2691 & n18690 ) | ( n2691 & ~n31749 ) | ( n18690 & ~n31749 ) ;
  assign n32427 = ( n1103 & n7739 ) | ( n1103 & ~n17895 ) | ( n7739 & ~n17895 ) ;
  assign n32428 = n19506 ^ n17617 ^ n11044 ;
  assign n32429 = n2646 | n5333 ;
  assign n32431 = ( n12532 & ~n15213 ) | ( n12532 & n16176 ) | ( ~n15213 & n16176 ) ;
  assign n32432 = ( n17586 & ~n23241 ) | ( n17586 & n32431 ) | ( ~n23241 & n32431 ) ;
  assign n32430 = n4303 & n29452 ;
  assign n32433 = n32432 ^ n32430 ^ 1'b0 ;
  assign n32434 = ( n3757 & n7342 ) | ( n3757 & ~n23964 ) | ( n7342 & ~n23964 ) ;
  assign n32435 = ( n4552 & n10619 ) | ( n4552 & ~n10956 ) | ( n10619 & ~n10956 ) ;
  assign n32436 = ~n8056 & n32435 ;
  assign n32437 = n32436 ^ n6179 ^ 1'b0 ;
  assign n32438 = ( n2232 & n7900 ) | ( n2232 & n11689 ) | ( n7900 & n11689 ) ;
  assign n32439 = ( n32434 & n32437 ) | ( n32434 & n32438 ) | ( n32437 & n32438 ) ;
  assign n32440 = ( ~n1202 & n25882 ) | ( ~n1202 & n32439 ) | ( n25882 & n32439 ) ;
  assign n32441 = ( n6216 & n25378 ) | ( n6216 & n29240 ) | ( n25378 & n29240 ) ;
  assign n32442 = n27772 & ~n32441 ;
  assign n32443 = n21905 ^ n21488 ^ n1791 ;
  assign n32444 = n32443 ^ n30029 ^ n17758 ;
  assign n32445 = n32444 ^ n18219 ^ 1'b0 ;
  assign n32446 = n5178 & n28509 ;
  assign n32448 = ~n1956 & n14307 ;
  assign n32449 = n32448 ^ n9034 ^ 1'b0 ;
  assign n32450 = n32449 ^ n8312 ^ n6577 ;
  assign n32447 = ~n1045 & n4267 ;
  assign n32451 = n32450 ^ n32447 ^ 1'b0 ;
  assign n32452 = ~n4209 & n25211 ;
  assign n32453 = n32452 ^ n26209 ^ 1'b0 ;
  assign n32454 = ( ~n13099 & n30684 ) | ( ~n13099 & n31377 ) | ( n30684 & n31377 ) ;
  assign n32456 = n30383 ^ n15153 ^ n11463 ;
  assign n32455 = n6128 | n29837 ;
  assign n32457 = n32456 ^ n32455 ^ 1'b0 ;
  assign n32458 = n2067 & n32457 ;
  assign n32459 = n32458 ^ n1465 ^ 1'b0 ;
  assign n32460 = n28382 ^ n23995 ^ n4257 ;
  assign n32461 = ( ~n28781 & n32459 ) | ( ~n28781 & n32460 ) | ( n32459 & n32460 ) ;
  assign n32462 = n24358 ^ n12755 ^ n6435 ;
  assign n32463 = n32462 ^ n25079 ^ n18379 ;
  assign n32464 = n27892 ^ n12845 ^ n11445 ;
  assign n32465 = n32464 ^ n15657 ^ n14656 ;
  assign n32466 = n8546 & ~n16228 ;
  assign n32467 = n32466 ^ n20356 ^ 1'b0 ;
  assign n32468 = ( ~n7009 & n15404 ) | ( ~n7009 & n25888 ) | ( n15404 & n25888 ) ;
  assign n32469 = n15329 | n21590 ;
  assign n32470 = n32468 | n32469 ;
  assign n32471 = n9135 ^ n3270 ^ n341 ;
  assign n32472 = ( ~n6325 & n11670 ) | ( ~n6325 & n16995 ) | ( n11670 & n16995 ) ;
  assign n32473 = n13552 ^ n9431 ^ n8393 ;
  assign n32474 = ( n10946 & n11062 ) | ( n10946 & n32473 ) | ( n11062 & n32473 ) ;
  assign n32475 = ( ~n32471 & n32472 ) | ( ~n32471 & n32474 ) | ( n32472 & n32474 ) ;
  assign n32476 = n16842 ^ n12825 ^ n1958 ;
  assign n32477 = ( n14433 & n32026 ) | ( n14433 & ~n32476 ) | ( n32026 & ~n32476 ) ;
  assign n32478 = n32477 ^ n25579 ^ n11889 ;
  assign n32479 = ( n6542 & n13841 ) | ( n6542 & ~n31026 ) | ( n13841 & ~n31026 ) ;
  assign n32480 = n32479 ^ n9499 ^ 1'b0 ;
  assign n32481 = n13280 & ~n32480 ;
  assign n32482 = ~n9954 & n12346 ;
  assign n32483 = ~n32481 & n32482 ;
  assign n32484 = n2037 & n29214 ;
  assign n32485 = n2818 & n32484 ;
  assign n32486 = n18301 | n19180 ;
  assign n32487 = n32486 ^ n10271 ^ 1'b0 ;
  assign n32488 = n32487 ^ n20828 ^ n7942 ;
  assign n32489 = ( ~n3152 & n10688 ) | ( ~n3152 & n23352 ) | ( n10688 & n23352 ) ;
  assign n32490 = n32489 ^ n25012 ^ n24715 ;
  assign n32491 = n5576 ^ n2727 ^ n1007 ;
  assign n32492 = n32491 ^ n4300 ^ 1'b0 ;
  assign n32493 = ( ~n2922 & n7848 ) | ( ~n2922 & n13596 ) | ( n7848 & n13596 ) ;
  assign n32494 = ( n16455 & ~n17381 ) | ( n16455 & n32493 ) | ( ~n17381 & n32493 ) ;
  assign n32495 = n26568 & ~n32494 ;
  assign n32496 = n32495 ^ n22708 ^ 1'b0 ;
  assign n32497 = n2467 & ~n12370 ;
  assign n32498 = n32497 ^ n12693 ^ n860 ;
  assign n32499 = n32498 ^ n26351 ^ n18044 ;
  assign n32500 = n28299 ^ n20832 ^ n11755 ;
  assign n32501 = n30255 ^ n15227 ^ n9277 ;
  assign n32502 = ( n2545 & n32500 ) | ( n2545 & ~n32501 ) | ( n32500 & ~n32501 ) ;
  assign n32503 = ( ~n7825 & n8721 ) | ( ~n7825 & n27060 ) | ( n8721 & n27060 ) ;
  assign n32504 = n742 & n17751 ;
  assign n32505 = n21652 & n32504 ;
  assign n32506 = ( n486 & ~n2717 ) | ( n486 & n5459 ) | ( ~n2717 & n5459 ) ;
  assign n32507 = ~n15934 & n31039 ;
  assign n32508 = ~n32506 & n32507 ;
  assign n32509 = n12169 & ~n32508 ;
  assign n32510 = n16382 ^ n12615 ^ n1443 ;
  assign n32511 = n32510 ^ n28136 ^ n7306 ;
  assign n32512 = n20462 ^ n7636 ^ n800 ;
  assign n32513 = n32512 ^ n27160 ^ n1297 ;
  assign n32514 = n1987 & ~n21009 ;
  assign n32515 = ( n2331 & ~n16836 ) | ( n2331 & n22704 ) | ( ~n16836 & n22704 ) ;
  assign n32516 = n22426 ^ n9540 ^ n8466 ;
  assign n32517 = n16526 ^ n15881 ^ 1'b0 ;
  assign n32518 = x116 & n32517 ;
  assign n32519 = n32518 ^ n1545 ^ 1'b0 ;
  assign n32520 = n14351 | n32519 ;
  assign n32521 = ( ~n26529 & n30597 ) | ( ~n26529 & n32520 ) | ( n30597 & n32520 ) ;
  assign n32522 = n8026 ^ n3733 ^ n2469 ;
  assign n32523 = n1559 & ~n32522 ;
  assign n32524 = ~n3776 & n3878 ;
  assign n32525 = n32524 ^ n11924 ^ 1'b0 ;
  assign n32526 = n32525 ^ n21701 ^ n11925 ;
  assign n32527 = n32526 ^ n22216 ^ n17986 ;
  assign n32528 = ( n1852 & ~n2829 ) | ( n1852 & n14449 ) | ( ~n2829 & n14449 ) ;
  assign n32529 = ~n5839 & n32528 ;
  assign n32530 = n7145 ^ n5106 ^ 1'b0 ;
  assign n32531 = n20251 & n32530 ;
  assign n32532 = ~n502 & n8454 ;
  assign n32533 = n32532 ^ n2659 ^ 1'b0 ;
  assign n32534 = ( n3484 & ~n3623 ) | ( n3484 & n32533 ) | ( ~n3623 & n32533 ) ;
  assign n32535 = ( n6795 & n11179 ) | ( n6795 & ~n32534 ) | ( n11179 & ~n32534 ) ;
  assign n32536 = n3001 | n30268 ;
  assign n32537 = n3471 | n32536 ;
  assign n32538 = n5374 | n32537 ;
  assign n32539 = ( n3631 & ~n10335 ) | ( n3631 & n22477 ) | ( ~n10335 & n22477 ) ;
  assign n32540 = ( n18475 & ~n21522 ) | ( n18475 & n32539 ) | ( ~n21522 & n32539 ) ;
  assign n32541 = n32540 ^ n26386 ^ 1'b0 ;
  assign n32542 = ~n926 & n4513 ;
  assign n32543 = ~n7089 & n32542 ;
  assign n32544 = n11812 & n13559 ;
  assign n32545 = n32543 & n32544 ;
  assign n32546 = ( ~n1408 & n18781 ) | ( ~n1408 & n32545 ) | ( n18781 & n32545 ) ;
  assign n32547 = n12821 | n21730 ;
  assign n32548 = n32546 & ~n32547 ;
  assign n32549 = ~n31074 & n32548 ;
  assign n32550 = n8075 & n8960 ;
  assign n32551 = n32550 ^ n17976 ^ 1'b0 ;
  assign n32552 = n32015 ^ n14854 ^ n623 ;
  assign n32553 = n32311 ^ n30363 ^ 1'b0 ;
  assign n32554 = n32552 | n32553 ;
  assign n32555 = n10222 & n27257 ;
  assign n32556 = ~n17427 & n32555 ;
  assign n32557 = n30278 ^ n25425 ^ n10950 ;
  assign n32558 = n10990 ^ n4030 ^ 1'b0 ;
  assign n32559 = ( n32556 & ~n32557 ) | ( n32556 & n32558 ) | ( ~n32557 & n32558 ) ;
  assign n32560 = n16733 ^ n5661 ^ 1'b0 ;
  assign n32561 = n25650 ^ n19845 ^ n13110 ;
  assign n32562 = n18144 ^ n2967 ^ 1'b0 ;
  assign n32563 = ( n8503 & n17340 ) | ( n8503 & ~n18147 ) | ( n17340 & ~n18147 ) ;
  assign n32564 = n32563 ^ n9352 ^ n4763 ;
  assign n32565 = n5115 ^ n4359 ^ n721 ;
  assign n32566 = n26449 ^ n19403 ^ 1'b0 ;
  assign n32567 = n28345 | n32566 ;
  assign n32568 = n32567 ^ n13947 ^ 1'b0 ;
  assign n32569 = ~n32565 & n32568 ;
  assign n32570 = n22844 ^ n13011 ^ 1'b0 ;
  assign n32571 = ( ~n32564 & n32569 ) | ( ~n32564 & n32570 ) | ( n32569 & n32570 ) ;
  assign n32572 = n32571 ^ n9890 ^ n4031 ;
  assign n32573 = n11763 ^ n3500 ^ 1'b0 ;
  assign n32574 = n32573 ^ n26828 ^ n19412 ;
  assign n32575 = n8177 ^ n4512 ^ x239 ;
  assign n32577 = n30936 ^ n10786 ^ n4088 ;
  assign n32576 = ( ~x79 & n13020 ) | ( ~x79 & n17895 ) | ( n13020 & n17895 ) ;
  assign n32578 = n32577 ^ n32576 ^ 1'b0 ;
  assign n32579 = ~n5379 & n32578 ;
  assign n32580 = ~n18564 & n32579 ;
  assign n32581 = n10441 & ~n14008 ;
  assign n32582 = n16800 ^ n13785 ^ n3843 ;
  assign n32583 = ~n17256 & n24030 ;
  assign n32584 = ( n18211 & n29103 ) | ( n18211 & ~n32583 ) | ( n29103 & ~n32583 ) ;
  assign n32585 = ( n32581 & n32582 ) | ( n32581 & ~n32584 ) | ( n32582 & ~n32584 ) ;
  assign n32586 = n26315 ^ n16582 ^ 1'b0 ;
  assign n32588 = ( n6804 & ~n7236 ) | ( n6804 & n8980 ) | ( ~n7236 & n8980 ) ;
  assign n32589 = n32588 ^ n5452 ^ n767 ;
  assign n32587 = ( n506 & ~n6864 ) | ( n506 & n27528 ) | ( ~n6864 & n27528 ) ;
  assign n32590 = n32589 ^ n32587 ^ 1'b0 ;
  assign n32591 = n5014 & n32590 ;
  assign n32592 = ( n5065 & n5709 ) | ( n5065 & n32591 ) | ( n5709 & n32591 ) ;
  assign n32593 = ( n1698 & n32586 ) | ( n1698 & n32592 ) | ( n32586 & n32592 ) ;
  assign n32594 = n12163 ^ n1017 ^ n342 ;
  assign n32596 = ( ~n1918 & n23344 ) | ( ~n1918 & n28047 ) | ( n23344 & n28047 ) ;
  assign n32595 = ( n2605 & n21165 ) | ( n2605 & n28285 ) | ( n21165 & n28285 ) ;
  assign n32597 = n32596 ^ n32595 ^ 1'b0 ;
  assign n32599 = n3435 & n16061 ;
  assign n32600 = n32599 ^ n16588 ^ 1'b0 ;
  assign n32598 = ( n6138 & n9694 ) | ( n6138 & n23119 ) | ( n9694 & n23119 ) ;
  assign n32601 = n32600 ^ n32598 ^ n4034 ;
  assign n32602 = ( n3301 & n10317 ) | ( n3301 & n13759 ) | ( n10317 & n13759 ) ;
  assign n32603 = n15312 ^ n10787 ^ 1'b0 ;
  assign n32604 = n32603 ^ n26829 ^ 1'b0 ;
  assign n32606 = ( n3413 & n14707 ) | ( n3413 & ~n16708 ) | ( n14707 & ~n16708 ) ;
  assign n32605 = n16109 & n25135 ;
  assign n32607 = n32606 ^ n32605 ^ 1'b0 ;
  assign n32608 = n11674 ^ n2054 ^ n541 ;
  assign n32609 = n18210 ^ n6468 ^ 1'b0 ;
  assign n32610 = ( n29529 & n32608 ) | ( n29529 & ~n32609 ) | ( n32608 & ~n32609 ) ;
  assign n32611 = ( ~n4663 & n11966 ) | ( ~n4663 & n13755 ) | ( n11966 & n13755 ) ;
  assign n32612 = ~n12345 & n12456 ;
  assign n32613 = ( ~n19559 & n32611 ) | ( ~n19559 & n32612 ) | ( n32611 & n32612 ) ;
  assign n32614 = ( ~n16642 & n18724 ) | ( ~n16642 & n20383 ) | ( n18724 & n20383 ) ;
  assign n32615 = n1708 | n25115 ;
  assign n32616 = n32615 ^ n21930 ^ 1'b0 ;
  assign n32617 = n16810 ^ n1395 ^ 1'b0 ;
  assign n32618 = n12643 & n32617 ;
  assign n32619 = n19047 ^ n13918 ^ n10547 ;
  assign n32620 = ~n17559 & n20346 ;
  assign n32621 = n32619 & n32620 ;
  assign n32622 = n9307 ^ n3926 ^ 1'b0 ;
  assign n32623 = n6770 | n32622 ;
  assign n32624 = ( n3707 & ~n13853 ) | ( n3707 & n32623 ) | ( ~n13853 & n32623 ) ;
  assign n32625 = ~n32621 & n32624 ;
  assign n32626 = n32625 ^ n8368 ^ 1'b0 ;
  assign n32627 = n32626 ^ n17203 ^ n14315 ;
  assign n32628 = n19078 ^ n11930 ^ n9482 ;
  assign n32629 = ( ~n9662 & n21213 ) | ( ~n9662 & n32628 ) | ( n21213 & n32628 ) ;
  assign n32630 = n6994 ^ n3983 ^ n523 ;
  assign n32631 = n32630 ^ n23013 ^ 1'b0 ;
  assign n32632 = n5398 & ~n32631 ;
  assign n32633 = n23517 ^ n14782 ^ 1'b0 ;
  assign n32634 = ~n10238 & n32633 ;
  assign n32635 = n32634 ^ n10038 ^ 1'b0 ;
  assign n32636 = ~n15830 & n21469 ;
  assign n32637 = ( n15055 & n30308 ) | ( n15055 & n32636 ) | ( n30308 & n32636 ) ;
  assign n32638 = n26472 ^ n19395 ^ n9353 ;
  assign n32639 = ( n2451 & ~n2930 ) | ( n2451 & n15678 ) | ( ~n2930 & n15678 ) ;
  assign n32640 = ~n24794 & n30822 ;
  assign n32641 = n12711 ^ n7768 ^ n1012 ;
  assign n32642 = n10532 ^ n2287 ^ 1'b0 ;
  assign n32643 = n32641 | n32642 ;
  assign n32644 = n11664 | n32643 ;
  assign n32645 = n14860 & ~n32644 ;
  assign n32647 = ( n9686 & n11845 ) | ( n9686 & n14181 ) | ( n11845 & n14181 ) ;
  assign n32648 = ( ~n14568 & n14697 ) | ( ~n14568 & n32647 ) | ( n14697 & n32647 ) ;
  assign n32649 = n17229 ^ n12730 ^ n10138 ;
  assign n32650 = n8738 & n32649 ;
  assign n32651 = n32648 & n32650 ;
  assign n32646 = ( n14045 & n18361 ) | ( n14045 & n27187 ) | ( n18361 & n27187 ) ;
  assign n32652 = n32651 ^ n32646 ^ n18723 ;
  assign n32654 = n20831 ^ n14858 ^ n2162 ;
  assign n32653 = n4372 ^ n1356 ^ 1'b0 ;
  assign n32655 = n32654 ^ n32653 ^ n9711 ;
  assign n32656 = ( n6398 & n15963 ) | ( n6398 & n31532 ) | ( n15963 & n31532 ) ;
  assign n32657 = n628 & n10863 ;
  assign n32658 = ( n26279 & ~n32656 ) | ( n26279 & n32657 ) | ( ~n32656 & n32657 ) ;
  assign n32659 = n7162 & n10950 ;
  assign n32660 = n32659 ^ n7671 ^ 1'b0 ;
  assign n32661 = ( n8148 & ~n24922 ) | ( n8148 & n32660 ) | ( ~n24922 & n32660 ) ;
  assign n32662 = n32661 ^ n27791 ^ n6996 ;
  assign n32663 = ( n3069 & ~n8980 ) | ( n3069 & n23927 ) | ( ~n8980 & n23927 ) ;
  assign n32665 = n2541 & n17207 ;
  assign n32664 = n31555 ^ n26252 ^ n4885 ;
  assign n32666 = n32665 ^ n32664 ^ 1'b0 ;
  assign n32667 = n32663 & n32666 ;
  assign n32668 = n17515 ^ n10763 ^ n2078 ;
  assign n32669 = ~n22240 & n32668 ;
  assign n32670 = ( ~n19381 & n21259 ) | ( ~n19381 & n32669 ) | ( n21259 & n32669 ) ;
  assign n32671 = n14826 ^ n8702 ^ 1'b0 ;
  assign n32672 = n828 | n32671 ;
  assign n32673 = ( ~n18947 & n25616 ) | ( ~n18947 & n32672 ) | ( n25616 & n32672 ) ;
  assign n32674 = n5119 ^ n3663 ^ 1'b0 ;
  assign n32675 = n20010 ^ n7839 ^ 1'b0 ;
  assign n32676 = n16515 ^ n1581 ^ 1'b0 ;
  assign n32677 = n24768 & ~n32676 ;
  assign n32678 = ( ~n32674 & n32675 ) | ( ~n32674 & n32677 ) | ( n32675 & n32677 ) ;
  assign n32679 = n30615 ^ n28595 ^ 1'b0 ;
  assign n32680 = n32678 & ~n32679 ;
  assign n32681 = n27365 ^ n26492 ^ n8147 ;
  assign n32682 = ( n5748 & n7884 ) | ( n5748 & n26074 ) | ( n7884 & n26074 ) ;
  assign n32683 = ( n21521 & ~n23086 ) | ( n21521 & n32682 ) | ( ~n23086 & n32682 ) ;
  assign n32690 = ~x200 & n9991 ;
  assign n32689 = ( n5466 & n8885 ) | ( n5466 & ~n21422 ) | ( n8885 & ~n21422 ) ;
  assign n32691 = n32690 ^ n32689 ^ 1'b0 ;
  assign n32684 = ( n809 & ~n2895 ) | ( n809 & n3763 ) | ( ~n2895 & n3763 ) ;
  assign n32685 = n32684 ^ n21733 ^ n20574 ;
  assign n32686 = n11550 ^ n9712 ^ 1'b0 ;
  assign n32687 = n32686 ^ n14160 ^ n7503 ;
  assign n32688 = ( n15445 & ~n32685 ) | ( n15445 & n32687 ) | ( ~n32685 & n32687 ) ;
  assign n32692 = n32691 ^ n32688 ^ n8903 ;
  assign n32693 = n19591 ^ n6051 ^ 1'b0 ;
  assign n32694 = n8661 & ~n19592 ;
  assign n32695 = n32694 ^ n16733 ^ 1'b0 ;
  assign n32696 = n15929 ^ n14895 ^ 1'b0 ;
  assign n32697 = ~n22271 & n32696 ;
  assign n32698 = ( ~n16142 & n29167 ) | ( ~n16142 & n32697 ) | ( n29167 & n32697 ) ;
  assign n32699 = ~n11304 & n11443 ;
  assign n32704 = n2681 | n19045 ;
  assign n32705 = n32704 ^ n10858 ^ 1'b0 ;
  assign n32700 = n17564 ^ n17087 ^ n5340 ;
  assign n32701 = n32700 ^ n12288 ^ n403 ;
  assign n32702 = ( n4141 & ~n28702 ) | ( n4141 & n32701 ) | ( ~n28702 & n32701 ) ;
  assign n32703 = ( ~n9072 & n21386 ) | ( ~n9072 & n32702 ) | ( n21386 & n32702 ) ;
  assign n32706 = n32705 ^ n32703 ^ n27365 ;
  assign n32707 = n4515 & ~n23848 ;
  assign n32708 = n24945 ^ n1582 ^ n390 ;
  assign n32709 = n32708 ^ n31596 ^ n25529 ;
  assign n32710 = n14422 ^ n13434 ^ 1'b0 ;
  assign n32711 = n32709 & ~n32710 ;
  assign n32712 = n7295 ^ n5246 ^ n1960 ;
  assign n32713 = ( n13632 & n22428 ) | ( n13632 & ~n32712 ) | ( n22428 & ~n32712 ) ;
  assign n32714 = ( n3082 & ~n9723 ) | ( n3082 & n32713 ) | ( ~n9723 & n32713 ) ;
  assign n32715 = n22107 ^ n10067 ^ n1061 ;
  assign n32716 = ( n516 & n10262 ) | ( n516 & ~n17243 ) | ( n10262 & ~n17243 ) ;
  assign n32717 = n10718 ^ n2404 ^ n2349 ;
  assign n32718 = ( x192 & ~n5331 ) | ( x192 & n32717 ) | ( ~n5331 & n32717 ) ;
  assign n32719 = n32716 | n32718 ;
  assign n32720 = n9535 & ~n32719 ;
  assign n32721 = ( n4603 & n32715 ) | ( n4603 & n32720 ) | ( n32715 & n32720 ) ;
  assign n32722 = ( ~n17878 & n23867 ) | ( ~n17878 & n24940 ) | ( n23867 & n24940 ) ;
  assign n32723 = n32721 & ~n32722 ;
  assign n32724 = ( n9229 & ~n14273 ) | ( n9229 & n23117 ) | ( ~n14273 & n23117 ) ;
  assign n32725 = ( ~n6398 & n22281 ) | ( ~n6398 & n32724 ) | ( n22281 & n32724 ) ;
  assign n32726 = ~n10104 & n16003 ;
  assign n32727 = n23880 & ~n32726 ;
  assign n32728 = ( ~n13696 & n20915 ) | ( ~n13696 & n32373 ) | ( n20915 & n32373 ) ;
  assign n32729 = ( n7819 & ~n17932 ) | ( n7819 & n29045 ) | ( ~n17932 & n29045 ) ;
  assign n32730 = ( n3805 & n6087 ) | ( n3805 & n32729 ) | ( n6087 & n32729 ) ;
  assign n32731 = n2765 & ~n4005 ;
  assign n32732 = n32730 & n32731 ;
  assign n32733 = n32732 ^ n25919 ^ n13763 ;
  assign n32734 = n428 & ~n32733 ;
  assign n32735 = n32734 ^ n11378 ^ 1'b0 ;
  assign n32736 = n2031 & ~n24625 ;
  assign n32737 = ( n4249 & ~n4430 ) | ( n4249 & n5384 ) | ( ~n4430 & n5384 ) ;
  assign n32738 = ( n11867 & n26759 ) | ( n11867 & n32737 ) | ( n26759 & n32737 ) ;
  assign n32742 = n12897 & ~n22764 ;
  assign n32743 = ~n28865 & n32742 ;
  assign n32744 = n3296 & n32743 ;
  assign n32745 = n32744 ^ n5551 ^ n4031 ;
  assign n32739 = n6854 & ~n7111 ;
  assign n32740 = n32739 ^ n8360 ^ n4049 ;
  assign n32741 = n32740 ^ n8618 ^ n1443 ;
  assign n32746 = n32745 ^ n32741 ^ n23272 ;
  assign n32747 = n7116 | n16913 ;
  assign n32748 = n31779 & ~n32747 ;
  assign n32749 = n32748 ^ n4642 ^ 1'b0 ;
  assign n32750 = n9728 | n17064 ;
  assign n32751 = n32750 ^ n15771 ^ 1'b0 ;
  assign n32752 = ( n20731 & n21146 ) | ( n20731 & ~n32751 ) | ( n21146 & ~n32751 ) ;
  assign n32753 = n32752 ^ n18100 ^ n13639 ;
  assign n32754 = n29033 ^ n26244 ^ n13320 ;
  assign n32755 = ( n16834 & ~n17731 ) | ( n16834 & n21006 ) | ( ~n17731 & n21006 ) ;
  assign n32756 = n32755 ^ n14430 ^ n12926 ;
  assign n32757 = n22784 ^ n18974 ^ n5164 ;
  assign n32765 = n25078 ^ n9128 ^ n1844 ;
  assign n32762 = n4150 & n18001 ;
  assign n32763 = n32762 ^ n439 ^ 1'b0 ;
  assign n32764 = n32763 ^ n29956 ^ n25004 ;
  assign n32758 = n28249 ^ n11425 ^ 1'b0 ;
  assign n32759 = n24070 & ~n32758 ;
  assign n32760 = n22206 & n32759 ;
  assign n32761 = ( n27218 & ~n29763 ) | ( n27218 & n32760 ) | ( ~n29763 & n32760 ) ;
  assign n32766 = n32765 ^ n32764 ^ n32761 ;
  assign n32767 = ( n7236 & n12382 ) | ( n7236 & n16735 ) | ( n12382 & n16735 ) ;
  assign n32768 = ~n4734 & n7892 ;
  assign n32769 = n17699 & n32768 ;
  assign n32770 = ( n17568 & n32767 ) | ( n17568 & n32769 ) | ( n32767 & n32769 ) ;
  assign n32771 = ( n8806 & ~n19721 ) | ( n8806 & n31582 ) | ( ~n19721 & n31582 ) ;
  assign n32772 = n25009 ^ n15637 ^ 1'b0 ;
  assign n32773 = ( ~n4695 & n23594 ) | ( ~n4695 & n32772 ) | ( n23594 & n32772 ) ;
  assign n32775 = n9426 ^ n6647 ^ n2568 ;
  assign n32774 = n27706 ^ n22288 ^ n5349 ;
  assign n32776 = n32775 ^ n32774 ^ n8618 ;
  assign n32777 = ~n5135 & n16863 ;
  assign n32778 = n32777 ^ n9776 ^ n6273 ;
  assign n32779 = n26728 & ~n32778 ;
  assign n32780 = n32779 ^ n31613 ^ n5639 ;
  assign n32783 = n15144 ^ n4298 ^ 1'b0 ;
  assign n32781 = ( n3481 & n11828 ) | ( n3481 & ~n13656 ) | ( n11828 & ~n13656 ) ;
  assign n32782 = n32781 ^ n6050 ^ n2992 ;
  assign n32784 = n32783 ^ n32782 ^ n31626 ;
  assign n32785 = n20704 ^ n10435 ^ n5118 ;
  assign n32786 = ~n14362 & n32785 ;
  assign n32787 = ( n1198 & n4995 ) | ( n1198 & ~n6744 ) | ( n4995 & ~n6744 ) ;
  assign n32788 = n32787 ^ n2308 ^ 1'b0 ;
  assign n32789 = n705 & ~n17108 ;
  assign n32790 = n1174 & n5517 ;
  assign n32791 = ( n28956 & n30919 ) | ( n28956 & n32790 ) | ( n30919 & n32790 ) ;
  assign n32792 = n2784 & n8791 ;
  assign n32793 = n32792 ^ n7455 ^ 1'b0 ;
  assign n32794 = ( n3929 & n6936 ) | ( n3929 & ~n18842 ) | ( n6936 & ~n18842 ) ;
  assign n32795 = ( n11465 & n15702 ) | ( n11465 & n32794 ) | ( n15702 & n32794 ) ;
  assign n32796 = n32795 ^ n23974 ^ n21367 ;
  assign n32797 = ( ~n1923 & n25646 ) | ( ~n1923 & n28136 ) | ( n25646 & n28136 ) ;
  assign n32798 = n9641 & ~n32797 ;
  assign n32799 = ~n18935 & n32798 ;
  assign n32800 = ( n12045 & n20527 ) | ( n12045 & n32799 ) | ( n20527 & n32799 ) ;
  assign n32801 = n23199 ^ n13391 ^ n4748 ;
  assign n32802 = n32801 ^ n8172 ^ n6166 ;
  assign n32803 = ( n4242 & ~n13639 ) | ( n4242 & n23253 ) | ( ~n13639 & n23253 ) ;
  assign n32804 = n26853 ^ n7635 ^ 1'b0 ;
  assign n32805 = ( n11046 & n31637 ) | ( n11046 & n32804 ) | ( n31637 & n32804 ) ;
  assign n32806 = ( n7488 & ~n10457 ) | ( n7488 & n28935 ) | ( ~n10457 & n28935 ) ;
  assign n32807 = ( n5857 & n10823 ) | ( n5857 & n24352 ) | ( n10823 & n24352 ) ;
  assign n32808 = n32807 ^ n11135 ^ 1'b0 ;
  assign n32809 = n32808 ^ n14433 ^ n894 ;
  assign n32810 = n2220 | n28888 ;
  assign n32811 = n32810 ^ n1093 ^ 1'b0 ;
  assign n32812 = ( n23238 & n32809 ) | ( n23238 & n32811 ) | ( n32809 & n32811 ) ;
  assign n32813 = n32806 | n32812 ;
  assign n32814 = n26721 ^ n9749 ^ n6149 ;
  assign n32815 = n17901 | n32814 ;
  assign n32816 = ( n4254 & n10082 ) | ( n4254 & ~n17969 ) | ( n10082 & ~n17969 ) ;
  assign n32817 = ( n8260 & ~n27116 ) | ( n8260 & n32816 ) | ( ~n27116 & n32816 ) ;
  assign n32818 = ~n6277 & n9312 ;
  assign n32819 = n32818 ^ n2148 ^ 1'b0 ;
  assign n32820 = ( n5668 & n11922 ) | ( n5668 & n30000 ) | ( n11922 & n30000 ) ;
  assign n32821 = ( n27294 & ~n32819 ) | ( n27294 & n32820 ) | ( ~n32819 & n32820 ) ;
  assign n32822 = n32817 & n32821 ;
  assign n32823 = ( ~n5887 & n7128 ) | ( ~n5887 & n18178 ) | ( n7128 & n18178 ) ;
  assign n32824 = ( ~n1877 & n6975 ) | ( ~n1877 & n20154 ) | ( n6975 & n20154 ) ;
  assign n32825 = n32824 ^ n32624 ^ 1'b0 ;
  assign n32826 = n29452 & ~n32825 ;
  assign n32830 = ( n8050 & ~n8511 ) | ( n8050 & n30444 ) | ( ~n8511 & n30444 ) ;
  assign n32827 = n11140 ^ n451 ^ 1'b0 ;
  assign n32828 = n32827 ^ n10914 ^ 1'b0 ;
  assign n32829 = n32828 ^ n19910 ^ n16682 ;
  assign n32831 = n32830 ^ n32829 ^ n26251 ;
  assign n32832 = n5286 ^ n5082 ^ n4089 ;
  assign n32833 = x115 & ~n4160 ;
  assign n32834 = n12899 & n32833 ;
  assign n32835 = n32834 ^ n22843 ^ n3998 ;
  assign n32836 = ( n15420 & n25781 ) | ( n15420 & n32835 ) | ( n25781 & n32835 ) ;
  assign n32837 = ( n1868 & n32832 ) | ( n1868 & n32836 ) | ( n32832 & n32836 ) ;
  assign n32838 = ( n5196 & ~n27311 ) | ( n5196 & n27885 ) | ( ~n27311 & n27885 ) ;
  assign n32842 = n23848 ^ n21087 ^ n4476 ;
  assign n32841 = ( n867 & n8887 ) | ( n867 & ~n31121 ) | ( n8887 & ~n31121 ) ;
  assign n32843 = n32842 ^ n32841 ^ n3364 ;
  assign n32839 = ( n1739 & n4376 ) | ( n1739 & ~n12580 ) | ( n4376 & ~n12580 ) ;
  assign n32840 = n32839 ^ n17651 ^ n5470 ;
  assign n32844 = n32843 ^ n32840 ^ n16780 ;
  assign n32845 = ( n3732 & n6720 ) | ( n3732 & ~n8711 ) | ( n6720 & ~n8711 ) ;
  assign n32846 = n32845 ^ n31098 ^ 1'b0 ;
  assign n32847 = n21048 & n32846 ;
  assign n32848 = ( n1017 & ~n9387 ) | ( n1017 & n11740 ) | ( ~n9387 & n11740 ) ;
  assign n32849 = n19428 ^ n9976 ^ n9530 ;
  assign n32850 = n32849 ^ n29719 ^ 1'b0 ;
  assign n32851 = ( x222 & ~n3054 ) | ( x222 & n14739 ) | ( ~n3054 & n14739 ) ;
  assign n32852 = ( n969 & n990 ) | ( n969 & n5354 ) | ( n990 & n5354 ) ;
  assign n32853 = ~n24747 & n32852 ;
  assign n32855 = ( n1216 & ~n7693 ) | ( n1216 & n21441 ) | ( ~n7693 & n21441 ) ;
  assign n32856 = n32855 ^ n25646 ^ n5016 ;
  assign n32854 = n800 & ~n4318 ;
  assign n32857 = n32856 ^ n32854 ^ n28059 ;
  assign n32858 = n5190 & ~n25038 ;
  assign n32859 = n32858 ^ n15705 ^ 1'b0 ;
  assign n32862 = n14395 ^ n7716 ^ n1865 ;
  assign n32863 = ( n7473 & n12354 ) | ( n7473 & n32862 ) | ( n12354 & n32862 ) ;
  assign n32864 = n32863 ^ n29992 ^ n8703 ;
  assign n32860 = n30797 ^ n10471 ^ 1'b0 ;
  assign n32861 = n14656 & ~n32860 ;
  assign n32865 = n32864 ^ n32861 ^ n17808 ;
  assign n32866 = n12467 & ~n21120 ;
  assign n32867 = n17215 & ~n32866 ;
  assign n32868 = n32865 & n32867 ;
  assign n32869 = n3743 | n10846 ;
  assign n32870 = n32869 ^ n22622 ^ 1'b0 ;
  assign n32871 = n15511 ^ n7862 ^ n7476 ;
  assign n32872 = ( ~n5587 & n11373 ) | ( ~n5587 & n15010 ) | ( n11373 & n15010 ) ;
  assign n32873 = ~n32871 & n32872 ;
  assign n32874 = n32873 ^ n23051 ^ 1'b0 ;
  assign n32875 = n32874 ^ n15106 ^ 1'b0 ;
  assign n32876 = n32054 ^ n4908 ^ 1'b0 ;
  assign n32877 = ( n26391 & n31190 ) | ( n26391 & ~n32876 ) | ( n31190 & ~n32876 ) ;
  assign n32878 = n9460 ^ n3784 ^ n596 ;
  assign n32879 = ( n8771 & n9912 ) | ( n8771 & ~n17595 ) | ( n9912 & ~n17595 ) ;
  assign n32880 = ( n31016 & ~n32878 ) | ( n31016 & n32879 ) | ( ~n32878 & n32879 ) ;
  assign n32881 = ~n540 & n17678 ;
  assign n32882 = n31709 ^ n31708 ^ n31287 ;
  assign n32883 = ( n6293 & n13833 ) | ( n6293 & ~n15948 ) | ( n13833 & ~n15948 ) ;
  assign n32884 = ( ~n5328 & n13775 ) | ( ~n5328 & n20149 ) | ( n13775 & n20149 ) ;
  assign n32885 = ~n32883 & n32884 ;
  assign n32886 = n21435 ^ n4655 ^ n3623 ;
  assign n32887 = ( n18712 & n31181 ) | ( n18712 & n32886 ) | ( n31181 & n32886 ) ;
  assign n32888 = ( n2276 & ~n19469 ) | ( n2276 & n32887 ) | ( ~n19469 & n32887 ) ;
  assign n32889 = ( n12472 & ~n13733 ) | ( n12472 & n32888 ) | ( ~n13733 & n32888 ) ;
  assign n32890 = n22741 ^ n17742 ^ n5532 ;
  assign n32891 = n32890 ^ n12352 ^ n5371 ;
  assign n32892 = n13995 & n26936 ;
  assign n32893 = n2700 & ~n6508 ;
  assign n32894 = ~n32892 & n32893 ;
  assign n32895 = n9437 ^ n4181 ^ x7 ;
  assign n32896 = n30252 ^ n7419 ^ 1'b0 ;
  assign n32897 = ~n10357 & n32896 ;
  assign n32898 = ( n1276 & n27933 ) | ( n1276 & ~n32897 ) | ( n27933 & ~n32897 ) ;
  assign n32899 = ( n29743 & n32895 ) | ( n29743 & ~n32898 ) | ( n32895 & ~n32898 ) ;
  assign n32900 = n482 & n2020 ;
  assign n32901 = n13496 ^ n8227 ^ 1'b0 ;
  assign n32902 = ( n8798 & ~n32900 ) | ( n8798 & n32901 ) | ( ~n32900 & n32901 ) ;
  assign n32903 = ( ~n12218 & n15778 ) | ( ~n12218 & n32902 ) | ( n15778 & n32902 ) ;
  assign n32904 = n24125 ^ n1576 ^ 1'b0 ;
  assign n32905 = n32904 ^ n19625 ^ 1'b0 ;
  assign n32906 = ~n4829 & n32905 ;
  assign n32907 = ( ~n22139 & n26685 ) | ( ~n22139 & n29603 ) | ( n26685 & n29603 ) ;
  assign n32908 = n15070 & n21375 ;
  assign n32909 = n32908 ^ n20989 ^ n14901 ;
  assign n32910 = n26653 ^ n1197 ^ 1'b0 ;
  assign n32911 = n13843 | n32910 ;
  assign n32912 = ( n553 & ~n15469 ) | ( n553 & n32911 ) | ( ~n15469 & n32911 ) ;
  assign n32913 = ( n11597 & n22112 ) | ( n11597 & n28648 ) | ( n22112 & n28648 ) ;
  assign n32914 = n32913 ^ n17537 ^ n9960 ;
  assign n32915 = n32914 ^ n22185 ^ n7124 ;
  assign n32916 = n22556 & ~n29302 ;
  assign n32917 = n32916 ^ n5820 ^ n2878 ;
  assign n32918 = ( n5016 & n6260 ) | ( n5016 & ~n28603 ) | ( n6260 & ~n28603 ) ;
  assign n32919 = ~n12507 & n29243 ;
  assign n32920 = n32919 ^ n4007 ^ 1'b0 ;
  assign n32921 = ( n10376 & ~n15322 ) | ( n10376 & n32920 ) | ( ~n15322 & n32920 ) ;
  assign n32922 = n32921 ^ n20487 ^ n7312 ;
  assign n32923 = n32922 ^ n27167 ^ n5010 ;
  assign n32924 = n5010 & ~n32923 ;
  assign n32925 = n23126 & n32924 ;
  assign n32926 = ( ~n8893 & n14176 ) | ( ~n8893 & n32925 ) | ( n14176 & n32925 ) ;
  assign n32927 = ( n2012 & n23041 ) | ( n2012 & ~n32926 ) | ( n23041 & ~n32926 ) ;
  assign n32929 = n20049 ^ n5080 ^ 1'b0 ;
  assign n32930 = ~n4091 & n32929 ;
  assign n32928 = ( n1163 & n8031 ) | ( n1163 & ~n18720 ) | ( n8031 & ~n18720 ) ;
  assign n32931 = n32930 ^ n32928 ^ n13777 ;
  assign n32936 = ( n12401 & n14322 ) | ( n12401 & ~n19781 ) | ( n14322 & ~n19781 ) ;
  assign n32932 = n2644 & n11570 ;
  assign n32933 = n32932 ^ n14360 ^ 1'b0 ;
  assign n32934 = n32933 ^ n20985 ^ n10997 ;
  assign n32935 = ( x202 & n28968 ) | ( x202 & n32934 ) | ( n28968 & n32934 ) ;
  assign n32937 = n32936 ^ n32935 ^ n17207 ;
  assign n32938 = n10300 & ~n14094 ;
  assign n32939 = n32938 ^ x48 ^ 1'b0 ;
  assign n32940 = n26681 ^ n9448 ^ 1'b0 ;
  assign n32941 = n15425 ^ n3498 ^ 1'b0 ;
  assign n32942 = n32941 ^ n1909 ^ 1'b0 ;
  assign n32943 = ( n10914 & n24185 ) | ( n10914 & n32942 ) | ( n24185 & n32942 ) ;
  assign n32944 = ~n4453 & n13312 ;
  assign n32945 = ~n32943 & n32944 ;
  assign n32946 = n9443 & n18239 ;
  assign n32947 = ( n1019 & n7435 ) | ( n1019 & ~n13001 ) | ( n7435 & ~n13001 ) ;
  assign n32948 = ( n4984 & n32946 ) | ( n4984 & n32947 ) | ( n32946 & n32947 ) ;
  assign n32949 = ( n7348 & n32945 ) | ( n7348 & ~n32948 ) | ( n32945 & ~n32948 ) ;
  assign n32950 = ( n949 & ~n17860 ) | ( n949 & n27130 ) | ( ~n17860 & n27130 ) ;
  assign n32951 = ~n11654 & n25811 ;
  assign n32952 = n32951 ^ n13374 ^ 1'b0 ;
  assign n32953 = n335 & ~n4181 ;
  assign n32954 = n32953 ^ n13392 ^ 1'b0 ;
  assign n32955 = ( n4256 & ~n19142 ) | ( n4256 & n32954 ) | ( ~n19142 & n32954 ) ;
  assign n32956 = n17624 ^ n11302 ^ n8131 ;
  assign n32957 = ( n4981 & ~n8957 ) | ( n4981 & n32956 ) | ( ~n8957 & n32956 ) ;
  assign n32958 = n31563 ^ n22355 ^ n8907 ;
  assign n32959 = ( ~n32955 & n32957 ) | ( ~n32955 & n32958 ) | ( n32957 & n32958 ) ;
  assign n32961 = n22055 ^ n21241 ^ n13673 ;
  assign n32960 = ( n3343 & n11115 ) | ( n3343 & ~n17727 ) | ( n11115 & ~n17727 ) ;
  assign n32962 = n32961 ^ n32960 ^ n29752 ;
  assign n32963 = n22034 ^ n2805 ^ 1'b0 ;
  assign n32964 = n3339 | n5482 ;
  assign n32965 = n5870 & ~n32964 ;
  assign n32968 = ( n2255 & n2858 ) | ( n2255 & n27719 ) | ( n2858 & n27719 ) ;
  assign n32966 = ~n8692 & n24489 ;
  assign n32967 = n11870 & n32966 ;
  assign n32969 = n32968 ^ n32967 ^ n17969 ;
  assign n32970 = ~n16604 & n32969 ;
  assign n32971 = n32965 & n32970 ;
  assign n32972 = ( ~n3230 & n15822 ) | ( ~n3230 & n26713 ) | ( n15822 & n26713 ) ;
  assign n32973 = ( n893 & n3985 ) | ( n893 & n4679 ) | ( n3985 & n4679 ) ;
  assign n32974 = n32068 ^ n3756 ^ 1'b0 ;
  assign n32975 = n16841 ^ n6387 ^ n1953 ;
  assign n32976 = ( ~n16650 & n32974 ) | ( ~n16650 & n32975 ) | ( n32974 & n32975 ) ;
  assign n32977 = ( ~n32972 & n32973 ) | ( ~n32972 & n32976 ) | ( n32973 & n32976 ) ;
  assign n32979 = n2904 | n13175 ;
  assign n32978 = x96 & n23862 ;
  assign n32980 = n32979 ^ n32978 ^ n22646 ;
  assign n32981 = ( n661 & ~n6634 ) | ( n661 & n32980 ) | ( ~n6634 & n32980 ) ;
  assign n32982 = n6743 & n11675 ;
  assign n32983 = n32982 ^ n19828 ^ n15425 ;
  assign n32984 = ( n32612 & n32783 ) | ( n32612 & ~n32983 ) | ( n32783 & ~n32983 ) ;
  assign n32985 = n15649 ^ n7238 ^ n6279 ;
  assign n32986 = ( ~n661 & n7594 ) | ( ~n661 & n32985 ) | ( n7594 & n32985 ) ;
  assign n32987 = n32986 ^ n4863 ^ n2212 ;
  assign n32988 = n32987 ^ n22602 ^ n22226 ;
  assign n32989 = ( n13241 & n24782 ) | ( n13241 & ~n32988 ) | ( n24782 & ~n32988 ) ;
  assign n32992 = n4091 ^ n2165 ^ 1'b0 ;
  assign n32993 = ~n1002 & n32992 ;
  assign n32991 = ( n1724 & n13250 ) | ( n1724 & ~n14861 ) | ( n13250 & ~n14861 ) ;
  assign n32994 = n32993 ^ n32991 ^ n9473 ;
  assign n32995 = n32994 ^ n17124 ^ 1'b0 ;
  assign n32990 = n5211 & ~n6648 ;
  assign n32996 = n32995 ^ n32990 ^ 1'b0 ;
  assign n32997 = n32996 ^ n28715 ^ n7230 ;
  assign n33000 = ( ~n1139 & n10849 ) | ( ~n1139 & n22692 ) | ( n10849 & n22692 ) ;
  assign n33001 = ( ~n1331 & n15290 ) | ( ~n1331 & n33000 ) | ( n15290 & n33000 ) ;
  assign n33007 = ~n4271 & n9459 ;
  assign n33008 = n33007 ^ n26521 ^ 1'b0 ;
  assign n33009 = ( ~n14298 & n25273 ) | ( ~n14298 & n33008 ) | ( n25273 & n33008 ) ;
  assign n33002 = n5983 & ~n10336 ;
  assign n33003 = n33002 ^ n16271 ^ n1116 ;
  assign n33004 = n33003 ^ n17778 ^ n2343 ;
  assign n33005 = n30129 & ~n33004 ;
  assign n33006 = n33005 ^ n23692 ^ 1'b0 ;
  assign n33010 = n33009 ^ n33006 ^ n25877 ;
  assign n33011 = ( n20085 & n33001 ) | ( n20085 & n33010 ) | ( n33001 & n33010 ) ;
  assign n32998 = ( n835 & n21911 ) | ( n835 & n25435 ) | ( n21911 & n25435 ) ;
  assign n32999 = ~n26445 & n32998 ;
  assign n33012 = n33011 ^ n32999 ^ 1'b0 ;
  assign n33017 = n5376 & n25725 ;
  assign n33018 = ~n6119 & n33017 ;
  assign n33016 = n19264 ^ n9624 ^ n9571 ;
  assign n33014 = n23819 ^ n3801 ^ n2922 ;
  assign n33013 = ( ~n12828 & n17621 ) | ( ~n12828 & n24058 ) | ( n17621 & n24058 ) ;
  assign n33015 = n33014 ^ n33013 ^ n25970 ;
  assign n33019 = n33018 ^ n33016 ^ n33015 ;
  assign n33021 = n9575 ^ n8960 ^ n1352 ;
  assign n33020 = ( n2231 & ~n5831 ) | ( n2231 & n25074 ) | ( ~n5831 & n25074 ) ;
  assign n33022 = n33021 ^ n33020 ^ n22542 ;
  assign n33023 = ( ~n1909 & n6172 ) | ( ~n1909 & n14664 ) | ( n6172 & n14664 ) ;
  assign n33024 = n33023 ^ n29606 ^ n20742 ;
  assign n33025 = ( ~n2766 & n30554 ) | ( ~n2766 & n33024 ) | ( n30554 & n33024 ) ;
  assign n33026 = ( ~n1275 & n20146 ) | ( ~n1275 & n31072 ) | ( n20146 & n31072 ) ;
  assign n33027 = ( n2432 & n7351 ) | ( n2432 & ~n9381 ) | ( n7351 & ~n9381 ) ;
  assign n33028 = ( n5641 & ~n14893 ) | ( n5641 & n33027 ) | ( ~n14893 & n33027 ) ;
  assign n33029 = ( n4965 & n11170 ) | ( n4965 & ~n22270 ) | ( n11170 & ~n22270 ) ;
  assign n33030 = n31561 & n33029 ;
  assign n33031 = n33030 ^ n3376 ^ 1'b0 ;
  assign n33033 = ( ~n2557 & n11388 ) | ( ~n2557 & n13969 ) | ( n11388 & n13969 ) ;
  assign n33032 = n17256 | n28300 ;
  assign n33034 = n33033 ^ n33032 ^ n12807 ;
  assign n33038 = ~n7334 & n15813 ;
  assign n33039 = n33038 ^ n979 ^ 1'b0 ;
  assign n33040 = n19828 & ~n33039 ;
  assign n33041 = n33040 ^ n6052 ^ 1'b0 ;
  assign n33035 = n14099 & ~n25472 ;
  assign n33036 = n33035 ^ n19822 ^ n11457 ;
  assign n33037 = ( n15481 & n28949 ) | ( n15481 & ~n33036 ) | ( n28949 & ~n33036 ) ;
  assign n33042 = n33041 ^ n33037 ^ n4573 ;
  assign n33043 = n20942 ^ n13330 ^ n5583 ;
  assign n33044 = ( n15281 & n20004 ) | ( n15281 & n24711 ) | ( n20004 & n24711 ) ;
  assign n33045 = n31288 ^ n19792 ^ n19634 ;
  assign n33046 = n21504 ^ n2211 ^ 1'b0 ;
  assign n33047 = n24093 ^ n1967 ^ 1'b0 ;
  assign n33048 = ( ~n6898 & n12841 ) | ( ~n6898 & n24075 ) | ( n12841 & n24075 ) ;
  assign n33049 = n9752 ^ n9054 ^ n5643 ;
  assign n33050 = n6801 & n13234 ;
  assign n33051 = ( n23778 & n33049 ) | ( n23778 & ~n33050 ) | ( n33049 & ~n33050 ) ;
  assign n33052 = n20493 ^ n488 ^ 1'b0 ;
  assign n33053 = n4531 | n33052 ;
  assign n33054 = ( ~n9904 & n11771 ) | ( ~n9904 & n15206 ) | ( n11771 & n15206 ) ;
  assign n33055 = ( n290 & ~n6362 ) | ( n290 & n11032 ) | ( ~n6362 & n11032 ) ;
  assign n33056 = ~n1812 & n22288 ;
  assign n33057 = n33056 ^ n33055 ^ 1'b0 ;
  assign n33058 = n15640 ^ n4576 ^ n415 ;
  assign n33059 = ~n32154 & n33058 ;
  assign n33060 = n5261 & n6339 ;
  assign n33061 = n13820 | n31488 ;
  assign n33062 = n5216 | n33061 ;
  assign n33063 = ( ~n19305 & n33060 ) | ( ~n19305 & n33062 ) | ( n33060 & n33062 ) ;
  assign n33068 = ( x59 & n14018 ) | ( x59 & n14941 ) | ( n14018 & n14941 ) ;
  assign n33069 = n33068 ^ n22369 ^ n7115 ;
  assign n33066 = n4116 & ~n24403 ;
  assign n33065 = n26137 ^ n12770 ^ n3262 ;
  assign n33067 = n33066 ^ n33065 ^ n12539 ;
  assign n33070 = n33069 ^ n33067 ^ n15575 ;
  assign n33064 = ( n3834 & n9977 ) | ( n3834 & ~n11987 ) | ( n9977 & ~n11987 ) ;
  assign n33071 = n33070 ^ n33064 ^ n30370 ;
  assign n33072 = ( n22393 & ~n33063 ) | ( n22393 & n33071 ) | ( ~n33063 & n33071 ) ;
  assign n33073 = n17304 ^ n16626 ^ n12501 ;
  assign n33074 = n33073 ^ n8048 ^ 1'b0 ;
  assign n33076 = n11310 ^ n7322 ^ n2381 ;
  assign n33077 = n33076 ^ n8061 ^ 1'b0 ;
  assign n33078 = n16344 & n33077 ;
  assign n33075 = ( x73 & n5667 ) | ( x73 & ~n20595 ) | ( n5667 & ~n20595 ) ;
  assign n33079 = n33078 ^ n33075 ^ n26239 ;
  assign n33080 = n9349 ^ n6067 ^ 1'b0 ;
  assign n33081 = n12852 & ~n21396 ;
  assign n33082 = n33081 ^ n22386 ^ n12543 ;
  assign n33083 = n31486 ^ n12856 ^ n10760 ;
  assign n33084 = n33083 ^ n24524 ^ n11612 ;
  assign n33085 = n1339 & ~n27111 ;
  assign n33086 = n33085 ^ n30302 ^ 1'b0 ;
  assign n33087 = n33086 ^ n11753 ^ n1851 ;
  assign n33088 = n25646 ^ n9711 ^ n3987 ;
  assign n33089 = ( ~n4714 & n24532 ) | ( ~n4714 & n33088 ) | ( n24532 & n33088 ) ;
  assign n33091 = ( n4651 & n9027 ) | ( n4651 & n27240 ) | ( n9027 & n27240 ) ;
  assign n33090 = n5905 ^ n4195 ^ n1541 ;
  assign n33092 = n33091 ^ n33090 ^ n8982 ;
  assign n33094 = n21978 ^ n506 ^ n337 ;
  assign n33093 = ( n685 & n10242 ) | ( n685 & n10617 ) | ( n10242 & n10617 ) ;
  assign n33095 = n33094 ^ n33093 ^ n9488 ;
  assign n33096 = ( n267 & n31272 ) | ( n267 & n33095 ) | ( n31272 & n33095 ) ;
  assign n33097 = ( n14791 & n33092 ) | ( n14791 & n33096 ) | ( n33092 & n33096 ) ;
  assign n33101 = n6872 | n16269 ;
  assign n33102 = n7654 & ~n33101 ;
  assign n33103 = n9681 & ~n33102 ;
  assign n33098 = n4978 & ~n6350 ;
  assign n33099 = n33098 ^ n23302 ^ 1'b0 ;
  assign n33100 = ~n23374 & n33099 ;
  assign n33104 = n33103 ^ n33100 ^ 1'b0 ;
  assign n33105 = n9855 ^ n7726 ^ 1'b0 ;
  assign n33106 = x242 & n33105 ;
  assign n33107 = n28923 ^ n18334 ^ n8412 ;
  assign n33108 = n33107 ^ n11353 ^ n6517 ;
  assign n33109 = n33108 ^ n19275 ^ 1'b0 ;
  assign n33110 = ( n33104 & n33106 ) | ( n33104 & ~n33109 ) | ( n33106 & ~n33109 ) ;
  assign n33111 = ~n5976 & n17258 ;
  assign n33112 = ( ~n4717 & n17236 ) | ( ~n4717 & n33111 ) | ( n17236 & n33111 ) ;
  assign n33113 = n24869 ^ n9069 ^ 1'b0 ;
  assign n33114 = ~n33112 & n33113 ;
  assign n33115 = ( n2445 & n14830 ) | ( n2445 & ~n31471 ) | ( n14830 & ~n31471 ) ;
  assign n33116 = n33115 ^ n3875 ^ n3727 ;
  assign n33117 = ( ~n2734 & n6287 ) | ( ~n2734 & n27204 ) | ( n6287 & n27204 ) ;
  assign n33118 = n33117 ^ n12844 ^ 1'b0 ;
  assign n33119 = ( n11770 & n16201 ) | ( n11770 & n33118 ) | ( n16201 & n33118 ) ;
  assign n33120 = n28154 ^ n19730 ^ n16705 ;
  assign n33121 = n26434 ^ n26244 ^ n14706 ;
  assign n33122 = ( n3253 & n18964 ) | ( n3253 & n19043 ) | ( n18964 & n19043 ) ;
  assign n33123 = n33122 ^ n3685 ^ n1729 ;
  assign n33124 = n12802 ^ n6051 ^ n3908 ;
  assign n33125 = n18104 ^ n17535 ^ 1'b0 ;
  assign n33126 = n33124 & n33125 ;
  assign n33127 = n20929 ^ n3208 ^ 1'b0 ;
  assign n33128 = n33126 & n33127 ;
  assign n33129 = n4272 & ~n31569 ;
  assign n33130 = n17954 & n33129 ;
  assign n33131 = ( n1863 & n11095 ) | ( n1863 & ~n15536 ) | ( n11095 & ~n15536 ) ;
  assign n33132 = n33131 ^ n13391 ^ 1'b0 ;
  assign n33133 = ~n33130 & n33132 ;
  assign n33134 = ( n1402 & n7215 ) | ( n1402 & n27330 ) | ( n7215 & n27330 ) ;
  assign n33135 = n33134 ^ n25421 ^ n9006 ;
  assign n33136 = ( n8162 & n14414 ) | ( n8162 & n28113 ) | ( n14414 & n28113 ) ;
  assign n33137 = n2880 & ~n19786 ;
  assign n33138 = n33137 ^ n671 ^ 1'b0 ;
  assign n33139 = ( ~n2212 & n3627 ) | ( ~n2212 & n7192 ) | ( n3627 & n7192 ) ;
  assign n33140 = n1518 | n33139 ;
  assign n33141 = n9779 | n33140 ;
  assign n33142 = n13072 & ~n33141 ;
  assign n33143 = n33142 ^ n4518 ^ 1'b0 ;
  assign n33144 = n22783 ^ n9081 ^ n6993 ;
  assign n33145 = ~n8806 & n28184 ;
  assign n33146 = n33145 ^ n1435 ^ 1'b0 ;
  assign n33147 = ( n9342 & n22007 ) | ( n9342 & n33146 ) | ( n22007 & n33146 ) ;
  assign n33148 = ~n19397 & n22894 ;
  assign n33149 = ( n33144 & n33147 ) | ( n33144 & ~n33148 ) | ( n33147 & ~n33148 ) ;
  assign n33150 = n27580 ^ n16400 ^ 1'b0 ;
  assign n33151 = n33150 ^ n33067 ^ n14137 ;
  assign n33152 = n31423 ^ n15364 ^ 1'b0 ;
  assign n33153 = ( n13636 & n26824 ) | ( n13636 & n33152 ) | ( n26824 & n33152 ) ;
  assign n33154 = n5996 & ~n27131 ;
  assign n33155 = ~n20021 & n33154 ;
  assign n33156 = n562 & ~n14895 ;
  assign n33157 = n21375 ^ n2138 ^ 1'b0 ;
  assign n33158 = ( n14036 & n24352 ) | ( n14036 & n33157 ) | ( n24352 & n33157 ) ;
  assign n33159 = ( n4226 & ~n15765 ) | ( n4226 & n33158 ) | ( ~n15765 & n33158 ) ;
  assign n33160 = ( n4635 & n6679 ) | ( n4635 & n18537 ) | ( n6679 & n18537 ) ;
  assign n33161 = n33159 & ~n33160 ;
  assign n33162 = ~n2768 & n33161 ;
  assign n33163 = n2364 ^ n371 ^ 1'b0 ;
  assign n33164 = n33163 ^ n31589 ^ n13851 ;
  assign n33166 = ~n14449 & n22257 ;
  assign n33167 = n17157 | n33166 ;
  assign n33168 = n16986 | n33167 ;
  assign n33169 = n33168 ^ n4094 ^ n2060 ;
  assign n33165 = ( ~n15580 & n16533 ) | ( ~n15580 & n23324 ) | ( n16533 & n23324 ) ;
  assign n33170 = n33169 ^ n33165 ^ n7067 ;
  assign n33175 = ( n2820 & ~n12647 ) | ( n2820 & n19375 ) | ( ~n12647 & n19375 ) ;
  assign n33173 = ( n4929 & n8923 ) | ( n4929 & n12900 ) | ( n8923 & n12900 ) ;
  assign n33171 = ( n13133 & n15102 ) | ( n13133 & n32400 ) | ( n15102 & n32400 ) ;
  assign n33172 = n33171 ^ n30873 ^ n15631 ;
  assign n33174 = n33173 ^ n33172 ^ n5414 ;
  assign n33176 = n33175 ^ n33174 ^ 1'b0 ;
  assign n33177 = n33176 ^ n31037 ^ 1'b0 ;
  assign n33178 = n29712 ^ n9892 ^ n6520 ;
  assign n33179 = n33178 ^ n3860 ^ n3446 ;
  assign n33180 = n14201 ^ n1226 ^ 1'b0 ;
  assign n33181 = ~n28942 & n33180 ;
  assign n33182 = ( n7105 & n32892 ) | ( n7105 & n33181 ) | ( n32892 & n33181 ) ;
  assign n33183 = n20408 ^ n16395 ^ 1'b0 ;
  assign n33184 = n6275 & n13877 ;
  assign n33185 = n33184 ^ n30775 ^ 1'b0 ;
  assign n33186 = n33185 ^ n12964 ^ n7636 ;
  assign n33187 = n33186 ^ n19232 ^ n3603 ;
  assign n33191 = n4987 & n7259 ;
  assign n33192 = n33191 ^ n8975 ^ 1'b0 ;
  assign n33193 = n33192 ^ n4207 ^ n1412 ;
  assign n33188 = n28762 ^ n14029 ^ n9678 ;
  assign n33189 = n33188 ^ n10324 ^ 1'b0 ;
  assign n33190 = ~n10935 & n33189 ;
  assign n33194 = n33193 ^ n33190 ^ 1'b0 ;
  assign n33195 = n33194 ^ n14257 ^ n1253 ;
  assign n33196 = n20316 ^ n12742 ^ n6964 ;
  assign n33197 = n31125 ^ n2375 ^ 1'b0 ;
  assign n33198 = n11564 & ~n33197 ;
  assign n33199 = n11179 ^ n7944 ^ n6479 ;
  assign n33200 = ( ~n4673 & n6586 ) | ( ~n4673 & n24087 ) | ( n6586 & n24087 ) ;
  assign n33201 = n33200 ^ n12399 ^ n9051 ;
  assign n33202 = ( ~n6817 & n14820 ) | ( ~n6817 & n33201 ) | ( n14820 & n33201 ) ;
  assign n33203 = ( n20586 & n33199 ) | ( n20586 & n33202 ) | ( n33199 & n33202 ) ;
  assign n33204 = ( ~n33196 & n33198 ) | ( ~n33196 & n33203 ) | ( n33198 & n33203 ) ;
  assign n33206 = n29844 ^ n13625 ^ n7360 ;
  assign n33207 = n845 & n18663 ;
  assign n33208 = ( n28265 & n33206 ) | ( n28265 & n33207 ) | ( n33206 & n33207 ) ;
  assign n33205 = n3565 & ~n13461 ;
  assign n33209 = n33208 ^ n33205 ^ 1'b0 ;
  assign n33210 = ( n1208 & n5527 ) | ( n1208 & n23360 ) | ( n5527 & n23360 ) ;
  assign n33211 = ( n2040 & n11118 ) | ( n2040 & n11159 ) | ( n11118 & n11159 ) ;
  assign n33212 = n21829 ^ n3495 ^ 1'b0 ;
  assign n33213 = n1023 & n33212 ;
  assign n33214 = n33213 ^ n6448 ^ n3773 ;
  assign n33215 = n33214 ^ n15354 ^ n1993 ;
  assign n33216 = n16762 | n24990 ;
  assign n33217 = n2316 | n33216 ;
  assign n33218 = n31695 ^ n13706 ^ 1'b0 ;
  assign n33219 = n11749 & n33218 ;
  assign n33220 = ( n4032 & ~n12587 ) | ( n4032 & n22242 ) | ( ~n12587 & n22242 ) ;
  assign n33224 = n28268 ^ n19285 ^ n2815 ;
  assign n33223 = ( n3105 & n17931 ) | ( n3105 & ~n22600 ) | ( n17931 & ~n22600 ) ;
  assign n33221 = n22495 ^ n18721 ^ n16991 ;
  assign n33222 = n33221 ^ n21678 ^ n14800 ;
  assign n33225 = n33224 ^ n33223 ^ n33222 ;
  assign n33226 = ( n5997 & n15163 ) | ( n5997 & ~n15941 ) | ( n15163 & ~n15941 ) ;
  assign n33227 = ( n3174 & ~n20493 ) | ( n3174 & n28517 ) | ( ~n20493 & n28517 ) ;
  assign n33228 = ( n19080 & n33226 ) | ( n19080 & n33227 ) | ( n33226 & n33227 ) ;
  assign n33229 = ( n1361 & ~n12668 ) | ( n1361 & n33228 ) | ( ~n12668 & n33228 ) ;
  assign n33230 = n13889 ^ n8505 ^ n3102 ;
  assign n33231 = n33230 ^ n24555 ^ n12663 ;
  assign n33232 = n19327 ^ n3067 ^ n1299 ;
  assign n33233 = n21253 & ~n33232 ;
  assign n33234 = n33233 ^ n18543 ^ 1'b0 ;
  assign n33235 = n28681 ^ n10296 ^ n464 ;
  assign n33236 = ~n764 & n33235 ;
  assign n33237 = n33236 ^ n9530 ^ 1'b0 ;
  assign n33240 = n25452 ^ n9012 ^ n4907 ;
  assign n33241 = ( ~n7211 & n7376 ) | ( ~n7211 & n33240 ) | ( n7376 & n33240 ) ;
  assign n33242 = ( n4730 & n13352 ) | ( n4730 & n33241 ) | ( n13352 & n33241 ) ;
  assign n33243 = ~n3150 & n33242 ;
  assign n33244 = n23013 & n33243 ;
  assign n33245 = n24711 | n33244 ;
  assign n33246 = n33245 ^ n23007 ^ 1'b0 ;
  assign n33238 = ( ~n8039 & n13912 ) | ( ~n8039 & n31302 ) | ( n13912 & n31302 ) ;
  assign n33239 = n33238 ^ n19343 ^ n1263 ;
  assign n33247 = n33246 ^ n33239 ^ 1'b0 ;
  assign n33248 = n24485 ^ n15066 ^ n343 ;
  assign n33249 = n926 ^ x144 ^ 1'b0 ;
  assign n33250 = ( n11549 & n12079 ) | ( n11549 & n30325 ) | ( n12079 & n30325 ) ;
  assign n33251 = n18496 ^ n8961 ^ 1'b0 ;
  assign n33252 = ( n9384 & ~n13073 ) | ( n9384 & n17135 ) | ( ~n13073 & n17135 ) ;
  assign n33253 = n5251 ^ n1963 ^ n1591 ;
  assign n33254 = n12038 & ~n33253 ;
  assign n33255 = n26691 ^ n6484 ^ 1'b0 ;
  assign n33256 = n23091 & ~n33255 ;
  assign n33257 = ( n3236 & n23922 ) | ( n3236 & n33256 ) | ( n23922 & n33256 ) ;
  assign n33259 = ( n8343 & n24537 ) | ( n8343 & ~n28372 ) | ( n24537 & ~n28372 ) ;
  assign n33258 = ( n19288 & n26004 ) | ( n19288 & n28752 ) | ( n26004 & n28752 ) ;
  assign n33260 = n33259 ^ n33258 ^ 1'b0 ;
  assign n33261 = n5519 & n11786 ;
  assign n33262 = n33261 ^ n19531 ^ n3266 ;
  assign n33263 = n10420 & n23556 ;
  assign n33264 = ~n27892 & n33263 ;
  assign n33265 = n28475 | n33264 ;
  assign n33266 = n5860 ^ n4018 ^ 1'b0 ;
  assign n33267 = x77 & ~n2548 ;
  assign n33268 = ~n20179 & n33267 ;
  assign n33269 = n761 & n11359 ;
  assign n33270 = ( n641 & ~n13098 ) | ( n641 & n33269 ) | ( ~n13098 & n33269 ) ;
  assign n33271 = n33270 ^ n8060 ^ n6680 ;
  assign n33272 = n6125 ^ n1680 ^ n1595 ;
  assign n33273 = n33272 ^ n23730 ^ 1'b0 ;
  assign n33274 = n31926 & ~n33273 ;
  assign n33275 = n33271 & n33274 ;
  assign n33276 = ( n20427 & ~n24610 ) | ( n20427 & n25437 ) | ( ~n24610 & n25437 ) ;
  assign n33277 = n18208 ^ n12617 ^ n12518 ;
  assign n33278 = n28577 ^ n27150 ^ n24167 ;
  assign n33279 = ( n6051 & ~n6626 ) | ( n6051 & n33278 ) | ( ~n6626 & n33278 ) ;
  assign n33280 = ( ~n19170 & n23556 ) | ( ~n19170 & n33279 ) | ( n23556 & n33279 ) ;
  assign n33283 = n9451 ^ n7535 ^ 1'b0 ;
  assign n33284 = n33283 ^ n8579 ^ 1'b0 ;
  assign n33281 = n16899 ^ n3245 ^ n1682 ;
  assign n33282 = n33281 ^ n341 ^ 1'b0 ;
  assign n33285 = n33284 ^ n33282 ^ n12281 ;
  assign n33286 = ( ~n5079 & n6502 ) | ( ~n5079 & n11872 ) | ( n6502 & n11872 ) ;
  assign n33287 = n778 | n6022 ;
  assign n33288 = n7868 | n33287 ;
  assign n33289 = n33288 ^ n18325 ^ n889 ;
  assign n33290 = n9991 ^ n2692 ^ 1'b0 ;
  assign n33291 = ~n33289 & n33290 ;
  assign n33292 = ( n10896 & n15848 ) | ( n10896 & ~n23544 ) | ( n15848 & ~n23544 ) ;
  assign n33293 = ( n33286 & n33291 ) | ( n33286 & n33292 ) | ( n33291 & n33292 ) ;
  assign n33294 = n25393 ^ n8430 ^ 1'b0 ;
  assign n33295 = ( ~n1055 & n23007 ) | ( ~n1055 & n33294 ) | ( n23007 & n33294 ) ;
  assign n33296 = n5510 & n29124 ;
  assign n33297 = n33296 ^ x19 ^ 1'b0 ;
  assign n33298 = n17248 ^ n14629 ^ n5920 ;
  assign n33299 = n19750 ^ n13750 ^ 1'b0 ;
  assign n33300 = ( n1202 & n1529 ) | ( n1202 & ~n33299 ) | ( n1529 & ~n33299 ) ;
  assign n33301 = n15998 ^ n10853 ^ n5250 ;
  assign n33302 = ( n1777 & n11833 ) | ( n1777 & n29400 ) | ( n11833 & n29400 ) ;
  assign n33303 = n21963 ^ n13176 ^ n8317 ;
  assign n33304 = n33303 ^ n8694 ^ 1'b0 ;
  assign n33305 = n10709 & n33304 ;
  assign n33306 = ~n26344 & n33305 ;
  assign n33307 = n33306 ^ n777 ^ 1'b0 ;
  assign n33308 = n14581 | n33307 ;
  assign n33309 = x86 & ~n4191 ;
  assign n33310 = n33309 ^ n14814 ^ 1'b0 ;
  assign n33311 = n33310 ^ n11174 ^ n5691 ;
  assign n33312 = n18791 ^ n11867 ^ n7235 ;
  assign n33313 = n33312 ^ n21146 ^ n4267 ;
  assign n33314 = ( n8006 & n11382 ) | ( n8006 & n26575 ) | ( n11382 & n26575 ) ;
  assign n33316 = ( n5880 & n13975 ) | ( n5880 & ~n14882 ) | ( n13975 & ~n14882 ) ;
  assign n33315 = n15000 ^ n7192 ^ n3007 ;
  assign n33317 = n33316 ^ n33315 ^ n17266 ;
  assign n33318 = ~n14691 & n23655 ;
  assign n33319 = ~n21059 & n33318 ;
  assign n33320 = ( n6170 & n24933 ) | ( n6170 & ~n33319 ) | ( n24933 & ~n33319 ) ;
  assign n33321 = n2084 & ~n7752 ;
  assign n33322 = n32733 ^ n32300 ^ n264 ;
  assign n33323 = n32742 ^ n18579 ^ n1144 ;
  assign n33324 = ( n3556 & ~n14610 ) | ( n3556 & n19625 ) | ( ~n14610 & n19625 ) ;
  assign n33325 = n6726 & n33324 ;
  assign n33326 = n15930 ^ n2728 ^ 1'b0 ;
  assign n33327 = n33325 & n33326 ;
  assign n33328 = ( ~n26377 & n33323 ) | ( ~n26377 & n33327 ) | ( n33323 & n33327 ) ;
  assign n33329 = n8509 ^ n4422 ^ 1'b0 ;
  assign n33330 = ( n6384 & n17120 ) | ( n6384 & n21044 ) | ( n17120 & n21044 ) ;
  assign n33331 = ( ~n4857 & n6698 ) | ( ~n4857 & n33330 ) | ( n6698 & n33330 ) ;
  assign n33332 = ( n13417 & n17693 ) | ( n13417 & ~n28339 ) | ( n17693 & ~n28339 ) ;
  assign n33333 = n9950 | n33332 ;
  assign n33334 = n33331 & ~n33333 ;
  assign n33335 = n17334 ^ n5761 ^ 1'b0 ;
  assign n33336 = n10415 & n33335 ;
  assign n33337 = n2088 | n15318 ;
  assign n33338 = n33337 ^ n1431 ^ 1'b0 ;
  assign n33339 = n33338 ^ n7280 ^ 1'b0 ;
  assign n33340 = n33336 & ~n33339 ;
  assign n33341 = n1960 | n23848 ;
  assign n33342 = n33340 | n33341 ;
  assign n33343 = n18452 ^ n1069 ^ 1'b0 ;
  assign n33344 = n33343 ^ n24186 ^ n11461 ;
  assign n33345 = n30510 ^ n11933 ^ n9144 ;
  assign n33346 = ( n9892 & ~n19688 ) | ( n9892 & n23676 ) | ( ~n19688 & n23676 ) ;
  assign n33347 = ( n5677 & n17479 ) | ( n5677 & n33346 ) | ( n17479 & n33346 ) ;
  assign n33348 = ( n5667 & n20902 ) | ( n5667 & n28452 ) | ( n20902 & n28452 ) ;
  assign n33349 = n2963 | n33348 ;
  assign n33350 = n30337 ^ n14604 ^ n8097 ;
  assign n33351 = ~n22007 & n33094 ;
  assign n33362 = n30435 ^ n20943 ^ n13541 ;
  assign n33358 = n12570 ^ n9405 ^ n7687 ;
  assign n33359 = n33358 ^ n25680 ^ n4359 ;
  assign n33353 = ( n1455 & ~n21629 ) | ( n1455 & n22294 ) | ( ~n21629 & n22294 ) ;
  assign n33354 = n15908 ^ n15260 ^ n11378 ;
  assign n33355 = n16908 & n33354 ;
  assign n33356 = ~n15281 & n33355 ;
  assign n33357 = ( n1523 & n33353 ) | ( n1523 & n33356 ) | ( n33353 & n33356 ) ;
  assign n33360 = n33359 ^ n33357 ^ n10887 ;
  assign n33361 = ( n13792 & ~n30171 ) | ( n13792 & n33360 ) | ( ~n30171 & n33360 ) ;
  assign n33363 = n33362 ^ n33361 ^ n11535 ;
  assign n33352 = n28905 ^ n16443 ^ n658 ;
  assign n33364 = n33363 ^ n33352 ^ n26449 ;
  assign n33365 = ( ~n31319 & n33351 ) | ( ~n31319 & n33364 ) | ( n33351 & n33364 ) ;
  assign n33366 = n22911 ^ n8716 ^ 1'b0 ;
  assign n33367 = n19498 & n24660 ;
  assign n33368 = n1102 & n33367 ;
  assign n33369 = ( n3096 & ~n33366 ) | ( n3096 & n33368 ) | ( ~n33366 & n33368 ) ;
  assign n33370 = n13943 ^ n13857 ^ n4298 ;
  assign n33371 = n3720 & ~n15222 ;
  assign n33372 = ( n8019 & ~n8570 ) | ( n8019 & n15989 ) | ( ~n8570 & n15989 ) ;
  assign n33373 = n33372 ^ n27657 ^ n6776 ;
  assign n33374 = n6344 ^ n4905 ^ n3365 ;
  assign n33375 = ( ~n11672 & n29580 ) | ( ~n11672 & n33374 ) | ( n29580 & n33374 ) ;
  assign n33376 = n11968 ^ n868 ^ 1'b0 ;
  assign n33377 = n33375 & ~n33376 ;
  assign n33379 = ( n2640 & ~n11034 ) | ( n2640 & n31188 ) | ( ~n11034 & n31188 ) ;
  assign n33378 = n13775 & ~n28475 ;
  assign n33380 = n33379 ^ n33378 ^ 1'b0 ;
  assign n33381 = n10988 ^ n8753 ^ n7408 ;
  assign n33382 = ( ~n2643 & n19452 ) | ( ~n2643 & n33381 ) | ( n19452 & n33381 ) ;
  assign n33383 = ( n7012 & n28910 ) | ( n7012 & n32431 ) | ( n28910 & n32431 ) ;
  assign n33384 = n18924 ^ n5582 ^ 1'b0 ;
  assign n33385 = ( ~n6209 & n19014 ) | ( ~n6209 & n28863 ) | ( n19014 & n28863 ) ;
  assign n33386 = ( n24818 & ~n33284 ) | ( n24818 & n33385 ) | ( ~n33284 & n33385 ) ;
  assign n33387 = ( n7470 & ~n33384 ) | ( n7470 & n33386 ) | ( ~n33384 & n33386 ) ;
  assign n33400 = ( ~n6194 & n18208 ) | ( ~n6194 & n28176 ) | ( n18208 & n28176 ) ;
  assign n33396 = ( n13833 & n15960 ) | ( n13833 & ~n23603 ) | ( n15960 & ~n23603 ) ;
  assign n33397 = ( n3329 & n14339 ) | ( n3329 & n33396 ) | ( n14339 & n33396 ) ;
  assign n33398 = n31077 ^ n3632 ^ 1'b0 ;
  assign n33399 = n33397 & ~n33398 ;
  assign n33401 = n33400 ^ n33399 ^ n28577 ;
  assign n33394 = n12489 ^ n8577 ^ n557 ;
  assign n33389 = x122 & ~n25368 ;
  assign n33390 = ~x23 & n33389 ;
  assign n33388 = n7382 & ~n16604 ;
  assign n33391 = n33390 ^ n33388 ^ 1'b0 ;
  assign n33392 = ~n27648 & n33391 ;
  assign n33393 = n33392 ^ n3629 ^ 1'b0 ;
  assign n33395 = n33394 ^ n33393 ^ n8461 ;
  assign n33402 = n33401 ^ n33395 ^ n12555 ;
  assign n33403 = ( n5719 & n6441 ) | ( n5719 & ~n12005 ) | ( n6441 & ~n12005 ) ;
  assign n33404 = n33403 ^ n26772 ^ n2760 ;
  assign n33405 = ( n14364 & n17055 ) | ( n14364 & n33404 ) | ( n17055 & n33404 ) ;
  assign n33406 = ~n6280 & n30350 ;
  assign n33407 = n33406 ^ n10876 ^ 1'b0 ;
  assign n33408 = n33407 ^ n28440 ^ n22351 ;
  assign n33410 = n20615 | n21778 ;
  assign n33409 = n11798 ^ n1691 ^ 1'b0 ;
  assign n33411 = n33410 ^ n33409 ^ n20934 ;
  assign n33412 = ( n6990 & n11055 ) | ( n6990 & ~n18263 ) | ( n11055 & ~n18263 ) ;
  assign n33413 = ( ~n11251 & n32378 ) | ( ~n11251 & n33412 ) | ( n32378 & n33412 ) ;
  assign n33414 = n33413 ^ n2965 ^ 1'b0 ;
  assign n33416 = n11172 ^ n7603 ^ n3578 ;
  assign n33415 = ( n14776 & n21078 ) | ( n14776 & ~n29823 ) | ( n21078 & ~n29823 ) ;
  assign n33417 = n33416 ^ n33415 ^ n3472 ;
  assign n33418 = n25778 ^ n23044 ^ 1'b0 ;
  assign n33419 = n17480 ^ n16595 ^ n10439 ;
  assign n33420 = n33419 ^ n25954 ^ 1'b0 ;
  assign n33422 = ( n4378 & ~n7143 ) | ( n4378 & n26612 ) | ( ~n7143 & n26612 ) ;
  assign n33421 = ( n826 & ~n4108 ) | ( n826 & n14016 ) | ( ~n4108 & n14016 ) ;
  assign n33423 = n33422 ^ n33421 ^ n11621 ;
  assign n33424 = n33423 ^ n16955 ^ n3926 ;
  assign n33425 = n4509 & n20132 ;
  assign n33426 = ( n1320 & n4168 ) | ( n1320 & ~n20190 ) | ( n4168 & ~n20190 ) ;
  assign n33427 = n33426 ^ n20922 ^ n6279 ;
  assign n33428 = n33427 ^ n28273 ^ 1'b0 ;
  assign n33429 = n12377 ^ n5556 ^ n1928 ;
  assign n33430 = n33429 ^ n24353 ^ n12981 ;
  assign n33433 = ( n2465 & ~n11677 ) | ( n2465 & n12404 ) | ( ~n11677 & n12404 ) ;
  assign n33431 = n15474 ^ n14605 ^ 1'b0 ;
  assign n33432 = n5980 | n33431 ;
  assign n33434 = n33433 ^ n33432 ^ n15038 ;
  assign n33435 = ( n2545 & ~n4687 ) | ( n2545 & n19346 ) | ( ~n4687 & n19346 ) ;
  assign n33436 = ( ~n1157 & n20647 ) | ( ~n1157 & n33435 ) | ( n20647 & n33435 ) ;
  assign n33437 = n7892 | n33436 ;
  assign n33438 = ~n3752 & n33437 ;
  assign n33439 = ~n1310 & n33438 ;
  assign n33440 = n11576 ^ n8750 ^ n2645 ;
  assign n33441 = n33440 ^ n28401 ^ 1'b0 ;
  assign n33442 = n26082 ^ n24755 ^ n11025 ;
  assign n33443 = n23893 | n33442 ;
  assign n33444 = n31888 | n33443 ;
  assign n33445 = n33444 ^ n10590 ^ n9081 ;
  assign n33446 = ( n23465 & n33441 ) | ( n23465 & ~n33445 ) | ( n33441 & ~n33445 ) ;
  assign n33447 = ( ~n10185 & n13245 ) | ( ~n10185 & n18534 ) | ( n13245 & n18534 ) ;
  assign n33448 = ( ~n4136 & n5210 ) | ( ~n4136 & n33447 ) | ( n5210 & n33447 ) ;
  assign n33449 = ( n350 & n14490 ) | ( n350 & n26693 ) | ( n14490 & n26693 ) ;
  assign n33450 = ( n12269 & n16268 ) | ( n12269 & ~n33449 ) | ( n16268 & ~n33449 ) ;
  assign n33451 = n33450 ^ n11037 ^ 1'b0 ;
  assign n33452 = ( n11041 & n12658 ) | ( n11041 & n33451 ) | ( n12658 & n33451 ) ;
  assign n33453 = ( n27983 & n33448 ) | ( n27983 & ~n33452 ) | ( n33448 & ~n33452 ) ;
  assign n33454 = n21304 ^ n5770 ^ x26 ;
  assign n33455 = n8184 | n33454 ;
  assign n33456 = n25033 & ~n33455 ;
  assign n33457 = n13146 | n27940 ;
  assign n33458 = n18200 ^ n13072 ^ 1'b0 ;
  assign n33459 = n33458 ^ n12503 ^ x110 ;
  assign n33460 = ( n10764 & n15191 ) | ( n10764 & ~n21637 ) | ( n15191 & ~n21637 ) ;
  assign n33461 = n33460 ^ n15726 ^ n14392 ;
  assign n33462 = n33461 ^ n25714 ^ n318 ;
  assign n33463 = n27186 ^ n24449 ^ n17683 ;
  assign n33464 = ~x152 & n33463 ;
  assign n33465 = n11926 & ~n33464 ;
  assign n33466 = n33465 ^ n25343 ^ 1'b0 ;
  assign n33467 = n25141 ^ n4244 ^ n2245 ;
  assign n33468 = n33467 ^ n5483 ^ n5415 ;
  assign n33469 = n7943 ^ n5496 ^ n5104 ;
  assign n33470 = ~n2254 & n12223 ;
  assign n33471 = n33470 ^ n8230 ^ 1'b0 ;
  assign n33472 = ~n17028 & n33471 ;
  assign n33473 = n33472 ^ n13308 ^ n8369 ;
  assign n33474 = n29403 ^ n27817 ^ n4219 ;
  assign n33475 = n33474 ^ n8263 ^ n7283 ;
  assign n33476 = n16513 ^ n9532 ^ n6027 ;
  assign n33477 = n33476 ^ n30334 ^ 1'b0 ;
  assign n33478 = n17139 ^ n9933 ^ n8773 ;
  assign n33479 = n11185 & ~n33478 ;
  assign n33480 = n11438 & n33479 ;
  assign n33481 = ( ~n8761 & n11127 ) | ( ~n8761 & n33480 ) | ( n11127 & n33480 ) ;
  assign n33482 = n33146 ^ n29522 ^ n14533 ;
  assign n33483 = ( n4671 & n6728 ) | ( n4671 & ~n28804 ) | ( n6728 & ~n28804 ) ;
  assign n33487 = n19149 ^ n11056 ^ n5595 ;
  assign n33488 = ( n2078 & ~n9797 ) | ( n2078 & n33487 ) | ( ~n9797 & n33487 ) ;
  assign n33484 = ~n7481 & n22384 ;
  assign n33485 = n5043 & n33484 ;
  assign n33486 = n33485 ^ n13452 ^ 1'b0 ;
  assign n33489 = n33488 ^ n33486 ^ n13766 ;
  assign n33490 = n20501 & n24783 ;
  assign n33491 = n20955 ^ x166 ^ 1'b0 ;
  assign n33492 = ( ~n983 & n20096 ) | ( ~n983 & n33491 ) | ( n20096 & n33491 ) ;
  assign n33493 = n20529 ^ n4121 ^ n3335 ;
  assign n33494 = n13263 & ~n33493 ;
  assign n33495 = ( n9072 & n18749 ) | ( n9072 & n33494 ) | ( n18749 & n33494 ) ;
  assign n33499 = ~x175 & n7256 ;
  assign n33498 = ( n9195 & ~n14348 ) | ( n9195 & n14572 ) | ( ~n14348 & n14572 ) ;
  assign n33500 = n33499 ^ n33498 ^ n28108 ;
  assign n33501 = n33500 ^ n23953 ^ n22931 ;
  assign n33496 = n32576 ^ n28266 ^ n7377 ;
  assign n33497 = ~n26059 & n33496 ;
  assign n33502 = n33501 ^ n33497 ^ 1'b0 ;
  assign n33503 = n678 | n2000 ;
  assign n33504 = n33503 ^ n10308 ^ 1'b0 ;
  assign n33505 = n21503 ^ n17476 ^ 1'b0 ;
  assign n33506 = n33505 ^ n25226 ^ x219 ;
  assign n33507 = n33506 ^ n24946 ^ n2258 ;
  assign n33508 = n33507 ^ n15509 ^ 1'b0 ;
  assign n33509 = n33504 & n33508 ;
  assign n33510 = ( x103 & n2684 ) | ( x103 & ~n3263 ) | ( n2684 & ~n3263 ) ;
  assign n33511 = n33510 ^ n5034 ^ n752 ;
  assign n33512 = n33511 ^ n15468 ^ 1'b0 ;
  assign n33513 = ( n22376 & ~n22665 ) | ( n22376 & n25924 ) | ( ~n22665 & n25924 ) ;
  assign n33514 = ( n3564 & ~n11035 ) | ( n3564 & n20967 ) | ( ~n11035 & n20967 ) ;
  assign n33515 = n28206 ^ n9977 ^ n7016 ;
  assign n33516 = n720 | n33515 ;
  assign n33517 = n5788 & ~n22236 ;
  assign n33518 = ~n2944 & n33517 ;
  assign n33519 = n32533 ^ n32431 ^ n21913 ;
  assign n33520 = n20557 ^ n8519 ^ n3151 ;
  assign n33521 = ( ~n8070 & n12926 ) | ( ~n8070 & n33520 ) | ( n12926 & n33520 ) ;
  assign n33522 = n10140 & ~n12616 ;
  assign n33523 = n33522 ^ n2132 ^ 1'b0 ;
  assign n33524 = ( n13703 & ~n32459 ) | ( n13703 & n33523 ) | ( ~n32459 & n33523 ) ;
  assign n33525 = n32630 ^ n25933 ^ 1'b0 ;
  assign n33526 = ~n14675 & n33525 ;
  assign n33527 = n8491 | n11069 ;
  assign n33528 = n33527 ^ n5469 ^ 1'b0 ;
  assign n33529 = ~n33526 & n33528 ;
  assign n33530 = ( n4348 & ~n7534 ) | ( n4348 & n11919 ) | ( ~n7534 & n11919 ) ;
  assign n33531 = ( n1185 & ~n26370 ) | ( n1185 & n33530 ) | ( ~n26370 & n33530 ) ;
  assign n33532 = ~n26359 & n33531 ;
  assign n33533 = ( n11036 & n25137 ) | ( n11036 & n33532 ) | ( n25137 & n33532 ) ;
  assign n33534 = n14736 & ~n33533 ;
  assign n33535 = ~n5268 & n33534 ;
  assign n33536 = ( n505 & ~n23115 ) | ( n505 & n27297 ) | ( ~n23115 & n27297 ) ;
  assign n33537 = ( n3098 & n7207 ) | ( n3098 & n33536 ) | ( n7207 & n33536 ) ;
  assign n33538 = n14566 ^ n7819 ^ n5411 ;
  assign n33539 = ( ~n24786 & n33500 ) | ( ~n24786 & n33538 ) | ( n33500 & n33538 ) ;
  assign n33540 = n17550 ^ n12987 ^ n8022 ;
  assign n33541 = ( n7840 & n9246 ) | ( n7840 & ~n29373 ) | ( n9246 & ~n29373 ) ;
  assign n33542 = n5285 & n12135 ;
  assign n33543 = ~n33541 & n33542 ;
  assign n33544 = n33543 ^ n5657 ^ n3990 ;
  assign n33545 = n27638 ^ n10777 ^ n10072 ;
  assign n33546 = n33545 ^ n27851 ^ n9811 ;
  assign n33547 = ( n19129 & n19375 ) | ( n19129 & ~n22157 ) | ( n19375 & ~n22157 ) ;
  assign n33548 = n15897 ^ n11862 ^ 1'b0 ;
  assign n33549 = ( n3992 & n12872 ) | ( n3992 & n33548 ) | ( n12872 & n33548 ) ;
  assign n33552 = n23650 ^ n13348 ^ 1'b0 ;
  assign n33550 = n29874 ^ n6141 ^ n2348 ;
  assign n33551 = n33524 & ~n33550 ;
  assign n33553 = n33552 ^ n33551 ^ 1'b0 ;
  assign n33554 = n23903 ^ n17689 ^ n12880 ;
  assign n33555 = n4918 ^ n1617 ^ n1462 ;
  assign n33556 = ( n13953 & n16954 ) | ( n13953 & n33555 ) | ( n16954 & n33555 ) ;
  assign n33557 = ( n14978 & n32359 ) | ( n14978 & ~n33556 ) | ( n32359 & ~n33556 ) ;
  assign n33558 = ( ~n5344 & n33554 ) | ( ~n5344 & n33557 ) | ( n33554 & n33557 ) ;
  assign n33559 = ~n1739 & n27513 ;
  assign n33560 = n21028 & n33559 ;
  assign n33561 = ( ~n12439 & n16676 ) | ( ~n12439 & n24338 ) | ( n16676 & n24338 ) ;
  assign n33562 = n982 | n3653 ;
  assign n33563 = n33562 ^ n25514 ^ 1'b0 ;
  assign n33564 = n33563 ^ n10386 ^ n9901 ;
  assign n33565 = ( n3683 & n20986 ) | ( n3683 & ~n33564 ) | ( n20986 & ~n33564 ) ;
  assign n33566 = n19420 & ~n25875 ;
  assign n33567 = n33566 ^ n6606 ^ 1'b0 ;
  assign n33568 = n6910 ^ n6324 ^ n4575 ;
  assign n33569 = n33568 ^ n18547 ^ n15743 ;
  assign n33570 = ( n1347 & n2550 ) | ( n1347 & n14634 ) | ( n2550 & n14634 ) ;
  assign n33571 = ( x47 & n12857 ) | ( x47 & ~n33570 ) | ( n12857 & ~n33570 ) ;
  assign n33572 = n33571 ^ n10059 ^ 1'b0 ;
  assign n33573 = n27303 ^ n21363 ^ n11921 ;
  assign n33574 = n33573 ^ n10185 ^ 1'b0 ;
  assign n33575 = n19356 & n33574 ;
  assign n33576 = n9651 ^ n4327 ^ 1'b0 ;
  assign n33577 = n33576 ^ n9851 ^ n3623 ;
  assign n33578 = n33577 ^ n8561 ^ 1'b0 ;
  assign n33579 = n22660 & ~n25069 ;
  assign n33580 = n33579 ^ n1656 ^ 1'b0 ;
  assign n33581 = n33580 ^ n11869 ^ n4929 ;
  assign n33582 = ( n14374 & n21601 ) | ( n14374 & n33581 ) | ( n21601 & n33581 ) ;
  assign n33584 = n13405 ^ n2089 ^ 1'b0 ;
  assign n33585 = ( n3558 & ~n18849 ) | ( n3558 & n33584 ) | ( ~n18849 & n33584 ) ;
  assign n33583 = ( ~n4037 & n6529 ) | ( ~n4037 & n28077 ) | ( n6529 & n28077 ) ;
  assign n33586 = n33585 ^ n33583 ^ 1'b0 ;
  assign n33589 = n3920 & n7542 ;
  assign n33587 = n24788 ^ n20137 ^ n16062 ;
  assign n33588 = n33587 ^ n29087 ^ n13517 ;
  assign n33590 = n33589 ^ n33588 ^ n19083 ;
  assign n33591 = n2483 | n7363 ;
  assign n33597 = ( n9052 & ~n20735 ) | ( n9052 & n27292 ) | ( ~n20735 & n27292 ) ;
  assign n33593 = ( ~n4970 & n5322 ) | ( ~n4970 & n8315 ) | ( n5322 & n8315 ) ;
  assign n33594 = n21746 ^ n3853 ^ 1'b0 ;
  assign n33595 = ( n21084 & ~n33593 ) | ( n21084 & n33594 ) | ( ~n33593 & n33594 ) ;
  assign n33592 = n17564 ^ n11652 ^ n11232 ;
  assign n33596 = n33595 ^ n33592 ^ n6051 ;
  assign n33598 = n33597 ^ n33596 ^ n5352 ;
  assign n33599 = ( n23380 & n33591 ) | ( n23380 & ~n33598 ) | ( n33591 & ~n33598 ) ;
  assign n33600 = n28810 & ~n33599 ;
  assign n33601 = n22565 ^ n5059 ^ 1'b0 ;
  assign n33602 = n24329 | n33601 ;
  assign n33603 = n8250 ^ n5787 ^ n867 ;
  assign n33604 = ( n6124 & n9343 ) | ( n6124 & ~n11820 ) | ( n9343 & ~n11820 ) ;
  assign n33605 = n4699 ^ n2162 ^ 1'b0 ;
  assign n33606 = ( n12219 & n22273 ) | ( n12219 & n33605 ) | ( n22273 & n33605 ) ;
  assign n33607 = n33606 ^ n15139 ^ 1'b0 ;
  assign n33608 = ( n545 & ~n33604 ) | ( n545 & n33607 ) | ( ~n33604 & n33607 ) ;
  assign n33609 = ~n16322 & n25670 ;
  assign n33610 = ( ~n5974 & n33608 ) | ( ~n5974 & n33609 ) | ( n33608 & n33609 ) ;
  assign n33611 = ( n16275 & n33603 ) | ( n16275 & n33610 ) | ( n33603 & n33610 ) ;
  assign n33612 = ( ~n992 & n13496 ) | ( ~n992 & n13906 ) | ( n13496 & n13906 ) ;
  assign n33613 = n2402 | n33612 ;
  assign n33614 = ~n28316 & n28961 ;
  assign n33615 = n1360 | n23074 ;
  assign n33616 = ( n2374 & ~n33614 ) | ( n2374 & n33615 ) | ( ~n33614 & n33615 ) ;
  assign n33617 = n31959 ^ n6480 ^ 1'b0 ;
  assign n33618 = n9817 & ~n33617 ;
  assign n33619 = n20096 ^ n19733 ^ n7335 ;
  assign n33621 = n20527 ^ n1264 ^ n542 ;
  assign n33620 = n27554 ^ n11310 ^ n7504 ;
  assign n33622 = n33621 ^ n33620 ^ n9744 ;
  assign n33623 = n7477 | n9623 ;
  assign n33624 = ( n13545 & n15542 ) | ( n13545 & ~n33623 ) | ( n15542 & ~n33623 ) ;
  assign n33625 = n28372 ^ n8118 ^ n5554 ;
  assign n33626 = ( ~n6620 & n9054 ) | ( ~n6620 & n33625 ) | ( n9054 & n33625 ) ;
  assign n33627 = n25975 & n33626 ;
  assign n33628 = ( n6455 & n15943 ) | ( n6455 & n33627 ) | ( n15943 & n33627 ) ;
  assign n33629 = n2615 & n21464 ;
  assign n33630 = ( n1182 & ~n3514 ) | ( n1182 & n33629 ) | ( ~n3514 & n33629 ) ;
  assign n33631 = ( ~n33624 & n33628 ) | ( ~n33624 & n33630 ) | ( n33628 & n33630 ) ;
  assign n33632 = n32293 ^ n28150 ^ n1246 ;
  assign n33633 = n4968 & n15353 ;
  assign n33634 = n3350 & n33633 ;
  assign n33635 = n33634 ^ n32623 ^ 1'b0 ;
  assign n33636 = ~n33632 & n33635 ;
  assign n33637 = n11929 | n16731 ;
  assign n33638 = n22698 & n23162 ;
  assign n33639 = n33637 & n33638 ;
  assign n33640 = n33636 | n33639 ;
  assign n33641 = n15685 ^ n15047 ^ n2414 ;
  assign n33642 = n17622 & ~n33641 ;
  assign n33643 = n33642 ^ n7312 ^ 1'b0 ;
  assign n33644 = n3162 | n9149 ;
  assign n33645 = n5271 & ~n33644 ;
  assign n33646 = n33645 ^ n17574 ^ n2676 ;
  assign n33647 = ( n9549 & n28768 ) | ( n9549 & n33646 ) | ( n28768 & n33646 ) ;
  assign n33648 = ~n27352 & n33647 ;
  assign n33649 = ( n8758 & ~n19213 ) | ( n8758 & n33648 ) | ( ~n19213 & n33648 ) ;
  assign n33655 = n29891 ^ n23910 ^ n820 ;
  assign n33651 = n1832 | n31076 ;
  assign n33652 = n12856 & ~n33651 ;
  assign n33653 = n26884 & ~n33652 ;
  assign n33654 = n7636 & n33653 ;
  assign n33656 = n33655 ^ n33654 ^ n8828 ;
  assign n33650 = n10977 & n17667 ;
  assign n33657 = n33656 ^ n33650 ^ 1'b0 ;
  assign n33658 = n18865 ^ n3888 ^ n1647 ;
  assign n33659 = ~n17329 & n33658 ;
  assign n33660 = ~n25461 & n33659 ;
  assign n33661 = n6392 ^ n5552 ^ 1'b0 ;
  assign n33662 = n1361 & ~n33661 ;
  assign n33663 = n33662 ^ n8550 ^ n8434 ;
  assign n33664 = ( n2393 & n2520 ) | ( n2393 & ~n20613 ) | ( n2520 & ~n20613 ) ;
  assign n33665 = n3094 & ~n33664 ;
  assign n33666 = ~n30401 & n33665 ;
  assign n33667 = n27827 | n33666 ;
  assign n33668 = n19183 | n33667 ;
  assign n33669 = ( n24517 & n29773 ) | ( n24517 & n33668 ) | ( n29773 & n33668 ) ;
  assign n33674 = ~n12166 & n13605 ;
  assign n33670 = n13393 & n17001 ;
  assign n33671 = n6240 & n22226 ;
  assign n33672 = n33671 ^ n4699 ^ 1'b0 ;
  assign n33673 = ( n17814 & n33670 ) | ( n17814 & ~n33672 ) | ( n33670 & ~n33672 ) ;
  assign n33675 = n33674 ^ n33673 ^ n12272 ;
  assign n33680 = n10728 ^ n2395 ^ 1'b0 ;
  assign n33676 = n18513 ^ n15955 ^ 1'b0 ;
  assign n33677 = n33676 ^ n12680 ^ 1'b0 ;
  assign n33678 = n2283 & n33677 ;
  assign n33679 = n30141 & n33678 ;
  assign n33681 = n33680 ^ n33679 ^ 1'b0 ;
  assign n33682 = n8184 ^ n4618 ^ 1'b0 ;
  assign n33683 = ( ~n4027 & n16496 ) | ( ~n4027 & n33682 ) | ( n16496 & n33682 ) ;
  assign n33684 = ( ~n2107 & n5971 ) | ( ~n2107 & n33683 ) | ( n5971 & n33683 ) ;
  assign n33685 = n27828 ^ n9641 ^ n1170 ;
  assign n33686 = ( n19371 & ~n21869 ) | ( n19371 & n23041 ) | ( ~n21869 & n23041 ) ;
  assign n33687 = ( n2656 & ~n29806 ) | ( n2656 & n31790 ) | ( ~n29806 & n31790 ) ;
  assign n33688 = x95 & n24810 ;
  assign n33689 = n33688 ^ n1019 ^ 1'b0 ;
  assign n33690 = ( n14684 & n24030 ) | ( n14684 & ~n33689 ) | ( n24030 & ~n33689 ) ;
  assign n33691 = n18394 ^ n9591 ^ n7271 ;
  assign n33692 = ( n5557 & n10332 ) | ( n5557 & n21188 ) | ( n10332 & n21188 ) ;
  assign n33693 = n29097 ^ n19526 ^ 1'b0 ;
  assign n33694 = n18628 ^ n11654 ^ 1'b0 ;
  assign n33695 = ( n33692 & ~n33693 ) | ( n33692 & n33694 ) | ( ~n33693 & n33694 ) ;
  assign n33696 = ( n7306 & ~n12913 ) | ( n7306 & n33695 ) | ( ~n12913 & n33695 ) ;
  assign n33697 = n17874 ^ n8872 ^ n6945 ;
  assign n33698 = n3181 | n33697 ;
  assign n33699 = ( ~n6335 & n15832 ) | ( ~n6335 & n33698 ) | ( n15832 & n33698 ) ;
  assign n33705 = ( n5118 & n5719 ) | ( n5118 & ~n9497 ) | ( n5719 & ~n9497 ) ;
  assign n33700 = n14156 | n25197 ;
  assign n33701 = n18806 & ~n33700 ;
  assign n33702 = ( n13880 & n17496 ) | ( n13880 & n19592 ) | ( n17496 & n19592 ) ;
  assign n33703 = ( ~n5184 & n15947 ) | ( ~n5184 & n33702 ) | ( n15947 & n33702 ) ;
  assign n33704 = ( ~n26032 & n33701 ) | ( ~n26032 & n33703 ) | ( n33701 & n33703 ) ;
  assign n33706 = n33705 ^ n33704 ^ n17873 ;
  assign n33707 = n18318 ^ n15695 ^ 1'b0 ;
  assign n33708 = n8301 | n33707 ;
  assign n33709 = n33708 ^ n14533 ^ n4098 ;
  assign n33710 = n3525 & ~n8590 ;
  assign n33715 = n13758 ^ n13253 ^ n12173 ;
  assign n33712 = ( ~n1444 & n9830 ) | ( ~n1444 & n10992 ) | ( n9830 & n10992 ) ;
  assign n33711 = n14641 ^ n13824 ^ n2384 ;
  assign n33713 = n33712 ^ n33711 ^ 1'b0 ;
  assign n33714 = n6407 & n33713 ;
  assign n33716 = n33715 ^ n33714 ^ n26475 ;
  assign n33717 = ( n19988 & n21128 ) | ( n19988 & n25588 ) | ( n21128 & n25588 ) ;
  assign n33718 = n4462 & n10112 ;
  assign n33719 = n33718 ^ x251 ^ 1'b0 ;
  assign n33720 = ~n33379 & n33719 ;
  assign n33721 = n33720 ^ n28648 ^ n950 ;
  assign n33723 = n27105 ^ n26721 ^ n18849 ;
  assign n33724 = n33723 ^ n12770 ^ n7570 ;
  assign n33722 = n29763 ^ n14659 ^ n12493 ;
  assign n33725 = n33724 ^ n33722 ^ n7692 ;
  assign n33726 = ( x152 & n15460 ) | ( x152 & ~n15732 ) | ( n15460 & ~n15732 ) ;
  assign n33727 = n33726 ^ n10439 ^ 1'b0 ;
  assign n33728 = n7584 ^ n1553 ^ n1179 ;
  assign n33729 = ( n7216 & n13158 ) | ( n7216 & ~n33728 ) | ( n13158 & ~n33728 ) ;
  assign n33730 = ( n14941 & n29516 ) | ( n14941 & ~n33729 ) | ( n29516 & ~n33729 ) ;
  assign n33731 = ( ~n2024 & n3507 ) | ( ~n2024 & n14463 ) | ( n3507 & n14463 ) ;
  assign n33732 = ( n5104 & n5573 ) | ( n5104 & ~n27191 ) | ( n5573 & ~n27191 ) ;
  assign n33733 = n33732 ^ n27595 ^ n12934 ;
  assign n33734 = ( ~n5181 & n9156 ) | ( ~n5181 & n29456 ) | ( n9156 & n29456 ) ;
  assign n33737 = n8272 ^ n3224 ^ 1'b0 ;
  assign n33735 = n20677 ^ n16791 ^ 1'b0 ;
  assign n33736 = n33735 ^ n29228 ^ n15778 ;
  assign n33738 = n33737 ^ n33736 ^ n22850 ;
  assign n33739 = ( n395 & n16735 ) | ( n395 & n33738 ) | ( n16735 & n33738 ) ;
  assign n33740 = ( n954 & n1971 ) | ( n954 & n2307 ) | ( n1971 & n2307 ) ;
  assign n33742 = ~n10934 & n13077 ;
  assign n33743 = ~n6930 & n33742 ;
  assign n33741 = n13555 ^ n6464 ^ n4778 ;
  assign n33744 = n33743 ^ n33741 ^ n5694 ;
  assign n33745 = ( ~n19111 & n33740 ) | ( ~n19111 & n33744 ) | ( n33740 & n33744 ) ;
  assign n33746 = ( n7408 & ~n9268 ) | ( n7408 & n23608 ) | ( ~n9268 & n23608 ) ;
  assign n33747 = ( n4565 & ~n6843 ) | ( n4565 & n8771 ) | ( ~n6843 & n8771 ) ;
  assign n33748 = ( n3680 & n8615 ) | ( n3680 & n9280 ) | ( n8615 & n9280 ) ;
  assign n33749 = n33748 ^ n9266 ^ n2476 ;
  assign n33750 = n17478 | n33749 ;
  assign n33751 = n33747 & ~n33750 ;
  assign n33752 = ( n7070 & ~n14988 ) | ( n7070 & n33751 ) | ( ~n14988 & n33751 ) ;
  assign n33753 = n9816 & ~n11527 ;
  assign n33754 = ~n12044 & n33753 ;
  assign n33755 = ( n5625 & ~n25178 ) | ( n5625 & n33754 ) | ( ~n25178 & n33754 ) ;
  assign n33757 = n29811 ^ n29504 ^ n18790 ;
  assign n33758 = n33757 ^ n4879 ^ 1'b0 ;
  assign n33759 = n33758 ^ n13017 ^ n5353 ;
  assign n33756 = n10014 | n29306 ;
  assign n33760 = n33759 ^ n33756 ^ 1'b0 ;
  assign n33761 = n33760 ^ n18860 ^ 1'b0 ;
  assign n33762 = ( n14888 & n15079 ) | ( n14888 & ~n27131 ) | ( n15079 & ~n27131 ) ;
  assign n33763 = n3793 ^ n3378 ^ n1180 ;
  assign n33764 = n2459 & n4581 ;
  assign n33765 = n1382 & n33764 ;
  assign n33766 = ( n16152 & n16863 ) | ( n16152 & n33765 ) | ( n16863 & n33765 ) ;
  assign n33767 = n33766 ^ n2272 ^ 1'b0 ;
  assign n33768 = n33763 | n33767 ;
  assign n33769 = n25840 & ~n33768 ;
  assign n33770 = ~n4045 & n33769 ;
  assign n33772 = ( n22277 & n23741 ) | ( n22277 & ~n25473 ) | ( n23741 & ~n25473 ) ;
  assign n33771 = n9741 ^ n6382 ^ n4214 ;
  assign n33773 = n33772 ^ n33771 ^ n3872 ;
  assign n33774 = n33773 ^ n31884 ^ 1'b0 ;
  assign n33775 = ~n6746 & n8891 ;
  assign n33776 = ( ~n633 & n9655 ) | ( ~n633 & n33775 ) | ( n9655 & n33775 ) ;
  assign n33777 = n27413 ^ n17731 ^ 1'b0 ;
  assign n33778 = ~n33055 & n33777 ;
  assign n33779 = n33778 ^ n14504 ^ n4784 ;
  assign n33780 = n33779 ^ n25786 ^ n1328 ;
  assign n33781 = n361 & n28782 ;
  assign n33782 = n33781 ^ n2032 ^ 1'b0 ;
  assign n33783 = ( ~n7983 & n33780 ) | ( ~n7983 & n33782 ) | ( n33780 & n33782 ) ;
  assign n33785 = n10452 ^ n9725 ^ x13 ;
  assign n33784 = ( ~n4208 & n8358 ) | ( ~n4208 & n28248 ) | ( n8358 & n28248 ) ;
  assign n33786 = n33785 ^ n33784 ^ n29663 ;
  assign n33787 = n31136 ^ n3397 ^ 1'b0 ;
  assign n33788 = n4399 | n10828 ;
  assign n33789 = ( ~n852 & n9951 ) | ( ~n852 & n33788 ) | ( n9951 & n33788 ) ;
  assign n33790 = n16343 | n22880 ;
  assign n33791 = n10217 | n33790 ;
  assign n33792 = ( n7713 & n14985 ) | ( n7713 & n33791 ) | ( n14985 & n33791 ) ;
  assign n33793 = ~n12821 & n33792 ;
  assign n33794 = n33793 ^ n17967 ^ 1'b0 ;
  assign n33795 = n33794 ^ n15371 ^ x245 ;
  assign n33796 = ( n20028 & n24464 ) | ( n20028 & n33795 ) | ( n24464 & n33795 ) ;
  assign n33797 = n17436 ^ n10932 ^ x4 ;
  assign n33798 = n14237 | n33797 ;
  assign n33799 = n13123 | n23005 ;
  assign n33800 = n33798 & ~n33799 ;
  assign n33801 = ( n15294 & n15667 ) | ( n15294 & n18984 ) | ( n15667 & n18984 ) ;
  assign n33802 = n13886 & ~n21200 ;
  assign n33803 = ~n33801 & n33802 ;
  assign n33804 = n13127 ^ n4698 ^ 1'b0 ;
  assign n33805 = n33804 ^ n9871 ^ n1137 ;
  assign n33806 = ( n8755 & n28316 ) | ( n8755 & ~n32663 ) | ( n28316 & ~n32663 ) ;
  assign n33807 = ( n8724 & n12508 ) | ( n8724 & n18087 ) | ( n12508 & n18087 ) ;
  assign n33808 = n8667 | n9846 ;
  assign n33809 = n33808 ^ n5359 ^ 1'b0 ;
  assign n33810 = ( ~n901 & n15058 ) | ( ~n901 & n33809 ) | ( n15058 & n33809 ) ;
  assign n33813 = ~x9 & n14069 ;
  assign n33811 = n29344 ^ n20238 ^ n12247 ;
  assign n33812 = n28951 & ~n33811 ;
  assign n33814 = n33813 ^ n33812 ^ 1'b0 ;
  assign n33815 = ~n10588 & n28871 ;
  assign n33816 = ~n33814 & n33815 ;
  assign n33819 = n1515 | n3519 ;
  assign n33817 = n19404 ^ n10833 ^ 1'b0 ;
  assign n33818 = n5714 | n33817 ;
  assign n33820 = n33819 ^ n33818 ^ 1'b0 ;
  assign n33821 = n27394 ^ n27371 ^ 1'b0 ;
  assign n33822 = n14900 & n33821 ;
  assign n33823 = ( ~n18327 & n25230 ) | ( ~n18327 & n33822 ) | ( n25230 & n33822 ) ;
  assign n33824 = ~n3504 & n7266 ;
  assign n33825 = n33824 ^ n1172 ^ 1'b0 ;
  assign n33826 = n23235 ^ n7971 ^ n4990 ;
  assign n33827 = n33826 ^ n3328 ^ 1'b0 ;
  assign n33828 = n33825 & ~n33827 ;
  assign n33829 = n27020 ^ n26675 ^ n9743 ;
  assign n33830 = ~n1095 & n33829 ;
  assign n33831 = ( n307 & ~n4754 ) | ( n307 & n23130 ) | ( ~n4754 & n23130 ) ;
  assign n33832 = n25279 & ~n33831 ;
  assign n33833 = n33832 ^ n25273 ^ n12188 ;
  assign n33834 = ( n18362 & n23660 ) | ( n18362 & ~n33833 ) | ( n23660 & ~n33833 ) ;
  assign n33836 = ( n1246 & n9561 ) | ( n1246 & ~n32742 ) | ( n9561 & ~n32742 ) ;
  assign n33837 = ~n5130 & n33836 ;
  assign n33835 = ~n6621 & n25209 ;
  assign n33838 = n33837 ^ n33835 ^ 1'b0 ;
  assign n33839 = n33237 ^ n16194 ^ n6502 ;
  assign n33840 = n30498 ^ n26917 ^ n8647 ;
  assign n33841 = n25140 ^ n14634 ^ n4837 ;
  assign n33842 = n16158 | n33841 ;
  assign n33843 = n33842 ^ n12531 ^ 1'b0 ;
  assign n33844 = ( n20558 & n23624 ) | ( n20558 & n33843 ) | ( n23624 & n33843 ) ;
  assign n33845 = n2095 | n15969 ;
  assign n33846 = n33845 ^ n13348 ^ 1'b0 ;
  assign n33847 = ( n11935 & ~n16362 ) | ( n11935 & n17229 ) | ( ~n16362 & n17229 ) ;
  assign n33849 = n3996 & n6979 ;
  assign n33850 = n33849 ^ n33039 ^ n27564 ;
  assign n33848 = n6285 & ~n26996 ;
  assign n33851 = n33850 ^ n33848 ^ 1'b0 ;
  assign n33852 = n21177 ^ n18748 ^ n6170 ;
  assign n33853 = n1900 & ~n33852 ;
  assign n33854 = n2575 & n33853 ;
  assign n33858 = ( n2919 & ~n5004 ) | ( n2919 & n10302 ) | ( ~n5004 & n10302 ) ;
  assign n33855 = n8281 & n23293 ;
  assign n33856 = n33855 ^ n23809 ^ 1'b0 ;
  assign n33857 = n33856 ^ n29829 ^ n27536 ;
  assign n33859 = n33858 ^ n33857 ^ n8782 ;
  assign n33860 = n5287 | n7522 ;
  assign n33861 = n33860 ^ n8486 ^ 1'b0 ;
  assign n33862 = ( n10859 & n16842 ) | ( n10859 & ~n30407 ) | ( n16842 & ~n30407 ) ;
  assign n33863 = ( n10194 & n33861 ) | ( n10194 & ~n33862 ) | ( n33861 & ~n33862 ) ;
  assign n33864 = ( ~n17276 & n22128 ) | ( ~n17276 & n31143 ) | ( n22128 & n31143 ) ;
  assign n33865 = ( n20223 & n22350 ) | ( n20223 & n33864 ) | ( n22350 & n33864 ) ;
  assign n33866 = n8622 & n21493 ;
  assign n33867 = n33866 ^ n26947 ^ 1'b0 ;
  assign n33868 = n33867 ^ n18245 ^ n11458 ;
  assign n33869 = ( n6383 & n17528 ) | ( n6383 & ~n25221 ) | ( n17528 & ~n25221 ) ;
  assign n33870 = ( ~n11362 & n21003 ) | ( ~n11362 & n33869 ) | ( n21003 & n33869 ) ;
  assign n33871 = ( ~n8282 & n18145 ) | ( ~n8282 & n33870 ) | ( n18145 & n33870 ) ;
  assign n33872 = n24294 ^ n10777 ^ n3884 ;
  assign n33873 = n33872 ^ n10467 ^ 1'b0 ;
  assign n33874 = n17708 ^ n11163 ^ 1'b0 ;
  assign n33875 = n2212 | n33874 ;
  assign n33876 = n20913 ^ n11696 ^ n1077 ;
  assign n33877 = ( ~n2617 & n10278 ) | ( ~n2617 & n28436 ) | ( n10278 & n28436 ) ;
  assign n33878 = n33877 ^ n32009 ^ 1'b0 ;
  assign n33879 = ~n33876 & n33878 ;
  assign n33880 = ( n7546 & n10988 ) | ( n7546 & n17611 ) | ( n10988 & n17611 ) ;
  assign n33881 = n626 & n10301 ;
  assign n33882 = ~n4764 & n33881 ;
  assign n33883 = n30820 ^ n18298 ^ n16607 ;
  assign n33884 = ( ~n7300 & n33882 ) | ( ~n7300 & n33883 ) | ( n33882 & n33883 ) ;
  assign n33889 = n18291 ^ n12349 ^ n8765 ;
  assign n33890 = ( n6438 & n7170 ) | ( n6438 & n33889 ) | ( n7170 & n33889 ) ;
  assign n33885 = n15257 ^ n3035 ^ 1'b0 ;
  assign n33886 = n16829 & ~n33885 ;
  assign n33887 = ( n496 & n2362 ) | ( n496 & ~n33886 ) | ( n2362 & ~n33886 ) ;
  assign n33888 = n25412 & ~n33887 ;
  assign n33891 = n33890 ^ n33888 ^ 1'b0 ;
  assign n33892 = ( n21970 & ~n33884 ) | ( n21970 & n33891 ) | ( ~n33884 & n33891 ) ;
  assign n33893 = n33892 ^ n8722 ^ 1'b0 ;
  assign n33894 = n33880 & ~n33893 ;
  assign n33895 = n13356 & ~n25439 ;
  assign n33896 = ( n4152 & n6338 ) | ( n4152 & n7571 ) | ( n6338 & n7571 ) ;
  assign n33897 = n33896 ^ n11594 ^ 1'b0 ;
  assign n33898 = n22004 ^ n7553 ^ 1'b0 ;
  assign n33899 = ( ~x115 & n4627 ) | ( ~x115 & n10392 ) | ( n4627 & n10392 ) ;
  assign n33900 = ( n3096 & n29825 ) | ( n3096 & n33899 ) | ( n29825 & n33899 ) ;
  assign n33901 = ( n33897 & n33898 ) | ( n33897 & ~n33900 ) | ( n33898 & ~n33900 ) ;
  assign n33902 = ( n2233 & n11310 ) | ( n2233 & ~n12047 ) | ( n11310 & ~n12047 ) ;
  assign n33903 = n28655 ^ n15543 ^ n562 ;
  assign n33904 = ( n13116 & ~n23906 ) | ( n13116 & n33903 ) | ( ~n23906 & n33903 ) ;
  assign n33905 = ( n10104 & n31041 ) | ( n10104 & ~n33904 ) | ( n31041 & ~n33904 ) ;
  assign n33906 = n33905 ^ n22481 ^ n16159 ;
  assign n33907 = ( ~n5616 & n10928 ) | ( ~n5616 & n16710 ) | ( n10928 & n16710 ) ;
  assign n33908 = n33907 ^ n27074 ^ n18721 ;
  assign n33909 = ( ~n1199 & n6468 ) | ( ~n1199 & n33908 ) | ( n6468 & n33908 ) ;
  assign n33910 = n25769 ^ n5312 ^ 1'b0 ;
  assign n33911 = n3682 & ~n33910 ;
  assign n33912 = n33911 ^ n7532 ^ n4511 ;
  assign n33913 = n15425 | n21458 ;
  assign n33914 = n33913 ^ n16675 ^ 1'b0 ;
  assign n33915 = ( n25126 & n33912 ) | ( n25126 & ~n33914 ) | ( n33912 & ~n33914 ) ;
  assign n33916 = n8262 & n17544 ;
  assign n33917 = n10189 ^ n9030 ^ n8413 ;
  assign n33918 = ~n2063 & n3302 ;
  assign n33919 = ( n1753 & n33917 ) | ( n1753 & n33918 ) | ( n33917 & n33918 ) ;
  assign n33922 = n32005 ^ n22353 ^ n13160 ;
  assign n33920 = n9563 & ~n12996 ;
  assign n33921 = ( ~n6549 & n15149 ) | ( ~n6549 & n33920 ) | ( n15149 & n33920 ) ;
  assign n33923 = n33922 ^ n33921 ^ n5648 ;
  assign n33924 = ( n1462 & ~n12651 ) | ( n1462 & n23214 ) | ( ~n12651 & n23214 ) ;
  assign n33925 = ( n6406 & n6539 ) | ( n6406 & n33924 ) | ( n6539 & n33924 ) ;
  assign n33926 = n33925 ^ n8925 ^ n2819 ;
  assign n33927 = n21490 ^ n11109 ^ n685 ;
  assign n33928 = n33926 & n33927 ;
  assign n33929 = n33928 ^ n14392 ^ 1'b0 ;
  assign n33930 = n14773 ^ n4265 ^ 1'b0 ;
  assign n33931 = n13415 ^ n11445 ^ n8881 ;
  assign n33932 = n30183 ^ n3096 ^ 1'b0 ;
  assign n33933 = n33932 ^ n24329 ^ 1'b0 ;
  assign n33934 = n4017 & n33933 ;
  assign n33935 = ~n19316 & n33934 ;
  assign n33936 = ( n3781 & n17801 ) | ( n3781 & n25965 ) | ( n17801 & n25965 ) ;
  assign n33937 = ~n7366 & n16911 ;
  assign n33938 = ~n33936 & n33937 ;
  assign n33944 = n8502 ^ n6446 ^ 1'b0 ;
  assign n33941 = n8438 & ~n15784 ;
  assign n33942 = n14704 & n33941 ;
  assign n33939 = n13197 ^ n12042 ^ 1'b0 ;
  assign n33940 = n6472 | n33939 ;
  assign n33943 = n33942 ^ n33940 ^ n28666 ;
  assign n33945 = n33944 ^ n33943 ^ n17048 ;
  assign n33946 = n16547 ^ n6970 ^ n6381 ;
  assign n33947 = ( n4335 & ~n14736 ) | ( n4335 & n21226 ) | ( ~n14736 & n21226 ) ;
  assign n33948 = ( n775 & n15184 ) | ( n775 & ~n33947 ) | ( n15184 & ~n33947 ) ;
  assign n33949 = ( n8773 & n10247 ) | ( n8773 & ~n17214 ) | ( n10247 & ~n17214 ) ;
  assign n33950 = n33949 ^ n3634 ^ 1'b0 ;
  assign n33951 = n2416 & n8874 ;
  assign n33952 = n33951 ^ n18263 ^ 1'b0 ;
  assign n33953 = n33952 ^ n8034 ^ n634 ;
  assign n33954 = ~n7911 & n21578 ;
  assign n33955 = ( n506 & n14003 ) | ( n506 & ~n33954 ) | ( n14003 & ~n33954 ) ;
  assign n33956 = n27953 & ~n33955 ;
  assign n33957 = ~n30293 & n33956 ;
  assign n33958 = n33957 ^ n24536 ^ n8638 ;
  assign n33959 = n10085 | n15934 ;
  assign n33960 = n33959 ^ n13529 ^ 1'b0 ;
  assign n33961 = n9706 ^ x36 ^ 1'b0 ;
  assign n33962 = ~n14182 & n33961 ;
  assign n33964 = ( ~n1873 & n2537 ) | ( ~n1873 & n7792 ) | ( n2537 & n7792 ) ;
  assign n33965 = n2802 & n33964 ;
  assign n33966 = n33965 ^ n11659 ^ 1'b0 ;
  assign n33963 = ( n1796 & n4657 ) | ( n1796 & n8977 ) | ( n4657 & n8977 ) ;
  assign n33967 = n33966 ^ n33963 ^ n23623 ;
  assign n33968 = ( n9437 & ~n33962 ) | ( n9437 & n33967 ) | ( ~n33962 & n33967 ) ;
  assign n33969 = n7415 ^ n4868 ^ n644 ;
  assign n33970 = n33969 ^ n15010 ^ 1'b0 ;
  assign n33971 = n1170 & ~n2099 ;
  assign n33972 = n33971 ^ n6127 ^ 1'b0 ;
  assign n33973 = n33972 ^ n18410 ^ n15915 ;
  assign n33974 = ( n1806 & n15624 ) | ( n1806 & n33973 ) | ( n15624 & n33973 ) ;
  assign n33975 = ( n21448 & n33970 ) | ( n21448 & ~n33974 ) | ( n33970 & ~n33974 ) ;
  assign n33976 = ( n3476 & n6017 ) | ( n3476 & ~n12051 ) | ( n6017 & ~n12051 ) ;
  assign n33977 = ~n1991 & n11358 ;
  assign n33978 = n33977 ^ n1961 ^ 1'b0 ;
  assign n33979 = n33978 ^ n19545 ^ n16453 ;
  assign n33980 = ( ~n17345 & n33976 ) | ( ~n17345 & n33979 ) | ( n33976 & n33979 ) ;
  assign n33981 = ~n7370 & n14167 ;
  assign n33982 = ~n13306 & n19213 ;
  assign n33983 = n33982 ^ n25988 ^ 1'b0 ;
  assign n33984 = ( n13977 & n33981 ) | ( n13977 & ~n33983 ) | ( n33981 & ~n33983 ) ;
  assign n33985 = ( ~n13634 & n27003 ) | ( ~n13634 & n29975 ) | ( n27003 & n29975 ) ;
  assign n33986 = n10783 ^ n10461 ^ n2232 ;
  assign n33987 = n33986 ^ n21455 ^ n5708 ;
  assign n33988 = n33987 ^ n31291 ^ n2363 ;
  assign n33989 = n6593 & ~n33988 ;
  assign n33990 = n33989 ^ n29948 ^ n7195 ;
  assign n33992 = n10999 ^ n3379 ^ x235 ;
  assign n33991 = n23663 ^ n22950 ^ n9427 ;
  assign n33993 = n33992 ^ n33991 ^ n10072 ;
  assign n33994 = ( n4812 & ~n14354 ) | ( n4812 & n33993 ) | ( ~n14354 & n33993 ) ;
  assign n33995 = ( n13342 & n15548 ) | ( n13342 & n31011 ) | ( n15548 & n31011 ) ;
  assign n33996 = n11963 ^ n8780 ^ n986 ;
  assign n33997 = ( n7345 & n25547 ) | ( n7345 & n33996 ) | ( n25547 & n33996 ) ;
  assign n33998 = ~n33995 & n33997 ;
  assign n33999 = n33998 ^ n3509 ^ 1'b0 ;
  assign n34000 = ( n10831 & n17798 ) | ( n10831 & ~n32226 ) | ( n17798 & ~n32226 ) ;
  assign n34001 = n23331 ^ n12341 ^ n6958 ;
  assign n34002 = n34001 ^ n15760 ^ 1'b0 ;
  assign n34003 = n839 | n11882 ;
  assign n34004 = n14496 ^ n7040 ^ 1'b0 ;
  assign n34005 = n34003 & n34004 ;
  assign n34006 = ~n19923 & n34005 ;
  assign n34007 = n19750 ^ n11696 ^ n1427 ;
  assign n34008 = n34007 ^ n6470 ^ n4017 ;
  assign n34009 = n11913 & ~n34008 ;
  assign n34010 = n34006 & n34009 ;
  assign n34011 = n34010 ^ n13335 ^ n7240 ;
  assign n34015 = n17316 ^ n8507 ^ n4084 ;
  assign n34016 = ( ~n8798 & n12181 ) | ( ~n8798 & n34015 ) | ( n12181 & n34015 ) ;
  assign n34017 = ( n3358 & n11157 ) | ( n3358 & ~n13908 ) | ( n11157 & ~n13908 ) ;
  assign n34018 = ( ~n10138 & n34016 ) | ( ~n10138 & n34017 ) | ( n34016 & n34017 ) ;
  assign n34013 = n977 & ~n1708 ;
  assign n34012 = n27240 ^ n14727 ^ x100 ;
  assign n34014 = n34013 ^ n34012 ^ 1'b0 ;
  assign n34019 = n34018 ^ n34014 ^ n9542 ;
  assign n34021 = n8699 ^ n5803 ^ n3146 ;
  assign n34022 = n34021 ^ n27711 ^ n1405 ;
  assign n34020 = n8950 ^ n7611 ^ n4378 ;
  assign n34023 = n34022 ^ n34020 ^ n20995 ;
  assign n34024 = ~n8092 & n34023 ;
  assign n34025 = ( n8586 & n28735 ) | ( n8586 & n34024 ) | ( n28735 & n34024 ) ;
  assign n34026 = n16003 ^ n1863 ^ 1'b0 ;
  assign n34027 = n18406 & ~n29421 ;
  assign n34028 = n11019 ^ n4116 ^ 1'b0 ;
  assign n34029 = n13807 & ~n24109 ;
  assign n34030 = ~n437 & n34029 ;
  assign n34031 = n19222 ^ n18713 ^ n10446 ;
  assign n34032 = n27447 ^ n25527 ^ n11683 ;
  assign n34033 = n34032 ^ n13999 ^ 1'b0 ;
  assign n34034 = n34031 & ~n34033 ;
  assign n34035 = n29558 ^ n27025 ^ 1'b0 ;
  assign n34036 = n15758 | n34035 ;
  assign n34037 = n12768 ^ n4243 ^ x222 ;
  assign n34038 = n31977 ^ n20166 ^ n10274 ;
  assign n34039 = ( ~n2136 & n5238 ) | ( ~n2136 & n32582 ) | ( n5238 & n32582 ) ;
  assign n34040 = n17886 ^ n7360 ^ 1'b0 ;
  assign n34041 = n27766 & ~n34040 ;
  assign n34042 = n28582 ^ n2716 ^ 1'b0 ;
  assign n34043 = n34042 ^ n15263 ^ n6261 ;
  assign n34044 = x214 | n34043 ;
  assign n34048 = n10368 | n13740 ;
  assign n34045 = n18471 ^ n740 ^ 1'b0 ;
  assign n34046 = n4841 | n34045 ;
  assign n34047 = n34046 ^ n28058 ^ n24172 ;
  assign n34049 = n34048 ^ n34047 ^ n6677 ;
  assign n34050 = ~n19725 & n34022 ;
  assign n34051 = ~n1530 & n34050 ;
  assign n34052 = ( x6 & n15803 ) | ( x6 & ~n34051 ) | ( n15803 & ~n34051 ) ;
  assign n34053 = n33592 ^ n28014 ^ n6042 ;
  assign n34054 = n11687 ^ n2154 ^ 1'b0 ;
  assign n34055 = ( n2903 & ~n5716 ) | ( n2903 & n7451 ) | ( ~n5716 & n7451 ) ;
  assign n34056 = ( n10912 & n20942 ) | ( n10912 & ~n34055 ) | ( n20942 & ~n34055 ) ;
  assign n34057 = ~n1200 & n34056 ;
  assign n34058 = n20229 & n34057 ;
  assign n34059 = n18244 ^ n15952 ^ 1'b0 ;
  assign n34060 = n6824 & n27428 ;
  assign n34061 = n34060 ^ n12962 ^ 1'b0 ;
  assign n34062 = n34059 & n34061 ;
  assign n34063 = ( n34054 & n34058 ) | ( n34054 & n34062 ) | ( n34058 & n34062 ) ;
  assign n34064 = ( n7473 & n11188 ) | ( n7473 & ~n34063 ) | ( n11188 & ~n34063 ) ;
  assign n34065 = n24055 ^ n18470 ^ n17717 ;
  assign n34066 = n26372 ^ n25257 ^ 1'b0 ;
  assign n34067 = n17865 & n34066 ;
  assign n34068 = ( n262 & ~n17241 ) | ( n262 & n17516 ) | ( ~n17241 & n17516 ) ;
  assign n34069 = ( n8436 & ~n10943 ) | ( n8436 & n34068 ) | ( ~n10943 & n34068 ) ;
  assign n34070 = n11611 ^ n10193 ^ n6126 ;
  assign n34071 = n33192 ^ n21362 ^ n6187 ;
  assign n34072 = n4752 & n34071 ;
  assign n34073 = n14393 ^ n1146 ^ 1'b0 ;
  assign n34074 = ( n2162 & n17201 ) | ( n2162 & n34073 ) | ( n17201 & n34073 ) ;
  assign n34075 = ( ~n28286 & n34072 ) | ( ~n28286 & n34074 ) | ( n34072 & n34074 ) ;
  assign n34076 = n6774 | n9424 ;
  assign n34077 = n34076 ^ n4828 ^ 1'b0 ;
  assign n34078 = n21864 ^ n7684 ^ n441 ;
  assign n34081 = ( ~n2566 & n4307 ) | ( ~n2566 & n25185 ) | ( n4307 & n25185 ) ;
  assign n34079 = n12708 & n13802 ;
  assign n34080 = n34079 ^ n12491 ^ 1'b0 ;
  assign n34082 = n34081 ^ n34080 ^ n16140 ;
  assign n34083 = n12312 ^ n9060 ^ n4666 ;
  assign n34084 = ( n3029 & n6391 ) | ( n3029 & ~n13133 ) | ( n6391 & ~n13133 ) ;
  assign n34085 = ~n14318 & n21106 ;
  assign n34086 = n34085 ^ n12570 ^ 1'b0 ;
  assign n34087 = n34086 ^ n17880 ^ 1'b0 ;
  assign n34088 = n23304 & ~n34087 ;
  assign n34089 = ~n34084 & n34088 ;
  assign n34090 = n34083 & n34089 ;
  assign n34091 = ( ~n22566 & n28975 ) | ( ~n22566 & n34090 ) | ( n28975 & n34090 ) ;
  assign n34092 = ~n2596 & n19286 ;
  assign n34093 = ~n33403 & n34092 ;
  assign n34094 = n18395 ^ n15512 ^ n3532 ;
  assign n34095 = n34094 ^ n12415 ^ n11523 ;
  assign n34096 = n15503 & n34095 ;
  assign n34097 = ( n20995 & ~n31167 ) | ( n20995 & n33310 ) | ( ~n31167 & n33310 ) ;
  assign n34098 = n34097 ^ n33052 ^ n26512 ;
  assign n34099 = n13963 ^ n11365 ^ n2268 ;
  assign n34100 = ( n879 & ~n26944 ) | ( n879 & n34099 ) | ( ~n26944 & n34099 ) ;
  assign n34101 = ~n6465 & n18744 ;
  assign n34102 = ( n7708 & ~n20818 ) | ( n7708 & n34101 ) | ( ~n20818 & n34101 ) ;
  assign n34103 = ( ~n2088 & n3462 ) | ( ~n2088 & n3930 ) | ( n3462 & n3930 ) ;
  assign n34104 = n34103 ^ n18610 ^ n16542 ;
  assign n34105 = n24949 ^ n14354 ^ n8710 ;
  assign n34106 = n26672 ^ n13596 ^ 1'b0 ;
  assign n34107 = ~n2916 & n34106 ;
  assign n34108 = ( n12905 & n31502 ) | ( n12905 & ~n34107 ) | ( n31502 & ~n34107 ) ;
  assign n34109 = ( n4045 & n10432 ) | ( n4045 & ~n22124 ) | ( n10432 & ~n22124 ) ;
  assign n34113 = n32961 ^ n17883 ^ n13432 ;
  assign n34110 = n7525 ^ n4953 ^ 1'b0 ;
  assign n34111 = n16354 | n34110 ;
  assign n34112 = n34111 ^ n21252 ^ 1'b0 ;
  assign n34114 = n34113 ^ n34112 ^ n14213 ;
  assign n34119 = n13941 ^ n13515 ^ n1789 ;
  assign n34115 = ( ~n6701 & n16034 ) | ( ~n6701 & n25448 ) | ( n16034 & n25448 ) ;
  assign n34116 = n6566 ^ n3005 ^ 1'b0 ;
  assign n34117 = n19394 & ~n34116 ;
  assign n34118 = ~n34115 & n34117 ;
  assign n34120 = n34119 ^ n34118 ^ 1'b0 ;
  assign n34121 = n1007 & n9037 ;
  assign n34122 = ~n34120 & n34121 ;
  assign n34123 = ~n13654 & n22245 ;
  assign n34124 = n22041 & n34123 ;
  assign n34125 = n25189 ^ n799 ^ 1'b0 ;
  assign n34126 = ( n16984 & ~n18576 ) | ( n16984 & n20009 ) | ( ~n18576 & n20009 ) ;
  assign n34127 = n24985 ^ n18088 ^ n6359 ;
  assign n34128 = ( n20787 & n32672 ) | ( n20787 & n34127 ) | ( n32672 & n34127 ) ;
  assign n34129 = n23450 ^ n15253 ^ n1233 ;
  assign n34130 = ( n19236 & n19300 ) | ( n19236 & ~n34129 ) | ( n19300 & ~n34129 ) ;
  assign n34131 = ( ~x72 & n2895 ) | ( ~x72 & n32985 ) | ( n2895 & n32985 ) ;
  assign n34134 = ( n2718 & n13838 ) | ( n2718 & n23890 ) | ( n13838 & n23890 ) ;
  assign n34132 = n14380 ^ n8080 ^ n7211 ;
  assign n34133 = n34132 ^ n10151 ^ n6632 ;
  assign n34135 = n34134 ^ n34133 ^ n12948 ;
  assign n34136 = ( n538 & n34131 ) | ( n538 & ~n34135 ) | ( n34131 & ~n34135 ) ;
  assign n34137 = ~n10546 & n14665 ;
  assign n34138 = n34137 ^ n28142 ^ 1'b0 ;
  assign n34139 = n34138 ^ n12628 ^ 1'b0 ;
  assign n34140 = n3654 & n34139 ;
  assign n34146 = n23745 ^ n5132 ^ x186 ;
  assign n34144 = n31098 ^ n12294 ^ x57 ;
  assign n34141 = n21674 ^ n13666 ^ n6901 ;
  assign n34142 = ( ~x105 & n2892 ) | ( ~x105 & n34141 ) | ( n2892 & n34141 ) ;
  assign n34143 = n15823 & n34142 ;
  assign n34145 = n34144 ^ n34143 ^ 1'b0 ;
  assign n34147 = n34146 ^ n34145 ^ n11262 ;
  assign n34148 = ( n1587 & ~n5761 ) | ( n1587 & n14364 ) | ( ~n5761 & n14364 ) ;
  assign n34149 = n34148 ^ n11821 ^ n11794 ;
  assign n34150 = ( ~n17119 & n20443 ) | ( ~n17119 & n34149 ) | ( n20443 & n34149 ) ;
  assign n34151 = n33488 ^ n8051 ^ n4075 ;
  assign n34152 = n34151 ^ n24836 ^ n11078 ;
  assign n34157 = ( n8904 & n13462 ) | ( n8904 & ~n26684 ) | ( n13462 & ~n26684 ) ;
  assign n34153 = n5745 & ~n18381 ;
  assign n34154 = n34153 ^ n6634 ^ 1'b0 ;
  assign n34155 = n6018 | n34154 ;
  assign n34156 = n34155 ^ n20622 ^ n3010 ;
  assign n34158 = n34157 ^ n34156 ^ n10639 ;
  assign n34159 = n28202 ^ n24350 ^ 1'b0 ;
  assign n34160 = ( x11 & n27419 ) | ( x11 & ~n34159 ) | ( n27419 & ~n34159 ) ;
  assign n34161 = ~n21665 & n34160 ;
  assign n34162 = ~n17361 & n26218 ;
  assign n34163 = n34162 ^ n6851 ^ 1'b0 ;
  assign n34164 = ( n27885 & n32892 ) | ( n27885 & ~n34163 ) | ( n32892 & ~n34163 ) ;
  assign n34165 = n9752 ^ n8433 ^ n3129 ;
  assign n34166 = n28777 ^ n1757 ^ 1'b0 ;
  assign n34167 = ~n31907 & n34166 ;
  assign n34168 = ( ~n6950 & n34165 ) | ( ~n6950 & n34167 ) | ( n34165 & n34167 ) ;
  assign n34169 = ( n7257 & n12620 ) | ( n7257 & n33024 ) | ( n12620 & n33024 ) ;
  assign n34170 = ( n5593 & ~n13203 ) | ( n5593 & n25296 ) | ( ~n13203 & n25296 ) ;
  assign n34171 = ( n3976 & ~n4160 ) | ( n3976 & n34170 ) | ( ~n4160 & n34170 ) ;
  assign n34172 = ( n5602 & n7526 ) | ( n5602 & n15107 ) | ( n7526 & n15107 ) ;
  assign n34173 = n9230 ^ n623 ^ 1'b0 ;
  assign n34174 = ~n1939 & n3524 ;
  assign n34175 = n34174 ^ x115 ^ 1'b0 ;
  assign n34176 = n34175 ^ n13486 ^ 1'b0 ;
  assign n34177 = n34176 ^ n30522 ^ n17128 ;
  assign n34178 = n28036 ^ n13749 ^ 1'b0 ;
  assign n34179 = n2744 & ~n34178 ;
  assign n34180 = n18981 ^ n11699 ^ 1'b0 ;
  assign n34183 = ( n983 & n5907 ) | ( n983 & ~n14237 ) | ( n5907 & ~n14237 ) ;
  assign n34181 = n16702 | n21589 ;
  assign n34182 = n15643 | n34181 ;
  assign n34184 = n34183 ^ n34182 ^ 1'b0 ;
  assign n34185 = n898 & ~n32828 ;
  assign n34186 = ~n6299 & n34185 ;
  assign n34187 = ( n2338 & ~n34184 ) | ( n2338 & n34186 ) | ( ~n34184 & n34186 ) ;
  assign n34188 = ( ~n3578 & n23774 ) | ( ~n3578 & n30322 ) | ( n23774 & n30322 ) ;
  assign n34189 = ( n4859 & ~n13581 ) | ( n4859 & n14484 ) | ( ~n13581 & n14484 ) ;
  assign n34191 = n9153 ^ n6237 ^ n4591 ;
  assign n34190 = n18065 ^ n15836 ^ n15677 ;
  assign n34192 = n34191 ^ n34190 ^ n11740 ;
  assign n34193 = n34192 ^ n2880 ^ 1'b0 ;
  assign n34194 = n34193 ^ n28812 ^ n12615 ;
  assign n34195 = n14380 & n34194 ;
  assign n34196 = n34195 ^ n1323 ^ 1'b0 ;
  assign n34197 = n6946 | n34196 ;
  assign n34198 = n11776 | n12656 ;
  assign n34199 = n24287 & ~n34198 ;
  assign n34200 = ( n310 & n11911 ) | ( n310 & n23732 ) | ( n11911 & n23732 ) ;
  assign n34201 = n32668 ^ n24825 ^ n1802 ;
  assign n34203 = n20916 ^ n9941 ^ n9327 ;
  assign n34202 = ( n7906 & ~n8928 ) | ( n7906 & n28673 ) | ( ~n8928 & n28673 ) ;
  assign n34204 = n34203 ^ n34202 ^ n3523 ;
  assign n34205 = n12253 & ~n18857 ;
  assign n34206 = ~n6209 & n34205 ;
  assign n34207 = n34206 ^ n10072 ^ 1'b0 ;
  assign n34208 = ( ~n8973 & n11627 ) | ( ~n8973 & n34207 ) | ( n11627 & n34207 ) ;
  assign n34209 = n32369 ^ n14292 ^ n6624 ;
  assign n34210 = ~n34208 & n34209 ;
  assign n34211 = n16934 & ~n23984 ;
  assign n34212 = ~n18873 & n26506 ;
  assign n34213 = n18864 ^ n18010 ^ n4191 ;
  assign n34214 = n32941 ^ n16957 ^ n3632 ;
  assign n34215 = n34213 & n34214 ;
  assign n34217 = ( n1714 & n2953 ) | ( n1714 & ~n6450 ) | ( n2953 & ~n6450 ) ;
  assign n34218 = ( n9431 & n22783 ) | ( n9431 & n34217 ) | ( n22783 & n34217 ) ;
  assign n34216 = n26323 ^ n23408 ^ n4960 ;
  assign n34219 = n34218 ^ n34216 ^ n1464 ;
  assign n34220 = ( n1276 & n18958 ) | ( n1276 & ~n30339 ) | ( n18958 & ~n30339 ) ;
  assign n34221 = ~n25232 & n34220 ;
  assign n34222 = ~n25456 & n34221 ;
  assign n34223 = ( n3697 & ~n24203 ) | ( n3697 & n34222 ) | ( ~n24203 & n34222 ) ;
  assign n34224 = n27086 ^ n20108 ^ n1768 ;
  assign n34225 = n3063 & ~n34224 ;
  assign n34226 = n18046 & n34225 ;
  assign n34227 = n15412 ^ n12964 ^ n529 ;
  assign n34228 = n20299 ^ n20094 ^ n11497 ;
  assign n34230 = ( ~n5846 & n13507 ) | ( ~n5846 & n14794 ) | ( n13507 & n14794 ) ;
  assign n34229 = n1619 | n15843 ;
  assign n34231 = n34230 ^ n34229 ^ 1'b0 ;
  assign n34232 = ( n3892 & n14042 ) | ( n3892 & ~n34231 ) | ( n14042 & ~n34231 ) ;
  assign n34233 = n1128 & ~n11925 ;
  assign n34234 = n34233 ^ n8419 ^ 1'b0 ;
  assign n34235 = n34234 ^ n21719 ^ n7351 ;
  assign n34241 = n888 | n14353 ;
  assign n34242 = n2074 & ~n34241 ;
  assign n34239 = ( ~n6787 & n14427 ) | ( ~n6787 & n28890 ) | ( n14427 & n28890 ) ;
  assign n34240 = n34239 ^ n26818 ^ 1'b0 ;
  assign n34243 = n34242 ^ n34240 ^ n14319 ;
  assign n34236 = n24464 ^ n14147 ^ n6781 ;
  assign n34237 = n34236 ^ n32898 ^ n8873 ;
  assign n34238 = n34237 ^ n11369 ^ n10837 ;
  assign n34244 = n34243 ^ n34238 ^ 1'b0 ;
  assign n34245 = ( n34232 & n34235 ) | ( n34232 & ~n34244 ) | ( n34235 & ~n34244 ) ;
  assign n34246 = n13532 ^ n911 ^ 1'b0 ;
  assign n34247 = n16355 & ~n34246 ;
  assign n34248 = ( n1614 & ~n21939 ) | ( n1614 & n34247 ) | ( ~n21939 & n34247 ) ;
  assign n34249 = ~n18433 & n34248 ;
  assign n34250 = n10337 & n34249 ;
  assign n34251 = ( n7998 & ~n11150 ) | ( n7998 & n34250 ) | ( ~n11150 & n34250 ) ;
  assign n34252 = ( ~n299 & n11481 ) | ( ~n299 & n29733 ) | ( n11481 & n29733 ) ;
  assign n34253 = n34252 ^ n16833 ^ n1953 ;
  assign n34254 = ( n6578 & n15197 ) | ( n6578 & n16689 ) | ( n15197 & n16689 ) ;
  assign n34255 = n34254 ^ n16114 ^ n3516 ;
  assign n34262 = ( n634 & ~n1349 ) | ( n634 & n22655 ) | ( ~n1349 & n22655 ) ;
  assign n34261 = ~n8606 & n20674 ;
  assign n34256 = ( n5306 & n8137 ) | ( n5306 & n11203 ) | ( n8137 & n11203 ) ;
  assign n34257 = n6339 & ~n18825 ;
  assign n34258 = n34257 ^ n12537 ^ n4942 ;
  assign n34259 = ( ~n28595 & n34256 ) | ( ~n28595 & n34258 ) | ( n34256 & n34258 ) ;
  assign n34260 = ( n9520 & ~n25775 ) | ( n9520 & n34259 ) | ( ~n25775 & n34259 ) ;
  assign n34263 = n34262 ^ n34261 ^ n34260 ;
  assign n34264 = ( ~n17123 & n34255 ) | ( ~n17123 & n34263 ) | ( n34255 & n34263 ) ;
  assign n34265 = ( n7323 & n10645 ) | ( n7323 & ~n12109 ) | ( n10645 & ~n12109 ) ;
  assign n34266 = n34265 ^ n5805 ^ n5559 ;
  assign n34267 = n34266 ^ n19822 ^ 1'b0 ;
  assign n34268 = n33472 ^ n27448 ^ n1544 ;
  assign n34278 = n32648 ^ n10713 ^ n2190 ;
  assign n34269 = ( n8272 & n29083 ) | ( n8272 & ~n32956 ) | ( n29083 & ~n32956 ) ;
  assign n34270 = ( n565 & n19219 ) | ( n565 & n34269 ) | ( n19219 & n34269 ) ;
  assign n34271 = n18426 ^ n12161 ^ n4779 ;
  assign n34272 = n9642 ^ n4988 ^ 1'b0 ;
  assign n34273 = n34271 | n34272 ;
  assign n34274 = ~n5414 & n27583 ;
  assign n34275 = n34273 & n34274 ;
  assign n34276 = n34275 ^ n4199 ^ 1'b0 ;
  assign n34277 = n34270 & n34276 ;
  assign n34279 = n34278 ^ n34277 ^ n19817 ;
  assign n34284 = ( n4087 & n7125 ) | ( n4087 & ~n15789 ) | ( n7125 & ~n15789 ) ;
  assign n34281 = n3718 ^ n724 ^ 1'b0 ;
  assign n34282 = ( n9805 & ~n24397 ) | ( n9805 & n34281 ) | ( ~n24397 & n34281 ) ;
  assign n34283 = ~n24291 & n34282 ;
  assign n34285 = n34284 ^ n34283 ^ 1'b0 ;
  assign n34286 = n21643 & ~n34285 ;
  assign n34287 = ~n27583 & n34286 ;
  assign n34280 = ~n5464 & n17165 ;
  assign n34288 = n34287 ^ n34280 ^ 1'b0 ;
  assign n34289 = n16518 ^ n10234 ^ 1'b0 ;
  assign n34290 = ( n2459 & n20624 ) | ( n2459 & n23311 ) | ( n20624 & n23311 ) ;
  assign n34291 = ( n3112 & ~n21718 ) | ( n3112 & n22381 ) | ( ~n21718 & n22381 ) ;
  assign n34292 = n34291 ^ n16032 ^ 1'b0 ;
  assign n34295 = ( n6687 & n8368 ) | ( n6687 & n17329 ) | ( n8368 & n17329 ) ;
  assign n34293 = ~n2666 & n10045 ;
  assign n34294 = n34293 ^ n21191 ^ 1'b0 ;
  assign n34296 = n34295 ^ n34294 ^ n6316 ;
  assign n34297 = ( ~n22107 & n29111 ) | ( ~n22107 & n34296 ) | ( n29111 & n34296 ) ;
  assign n34298 = ~n3653 & n18150 ;
  assign n34299 = n34298 ^ n8800 ^ 1'b0 ;
  assign n34300 = n1849 | n34299 ;
  assign n34301 = n6464 & n14736 ;
  assign n34302 = n34301 ^ n25067 ^ 1'b0 ;
  assign n34303 = n2483 & n34302 ;
  assign n34304 = n3955 ^ n2569 ^ 1'b0 ;
  assign n34305 = ( n4340 & ~n19564 ) | ( n4340 & n34304 ) | ( ~n19564 & n34304 ) ;
  assign n34306 = ( ~n12295 & n18107 ) | ( ~n12295 & n26157 ) | ( n18107 & n26157 ) ;
  assign n34307 = n31898 ^ n14701 ^ n13908 ;
  assign n34308 = n34307 ^ n4603 ^ 1'b0 ;
  assign n34309 = n34306 & ~n34308 ;
  assign n34310 = n32270 ^ n30357 ^ 1'b0 ;
  assign n34311 = n32968 & ~n34310 ;
  assign n34312 = n28848 ^ n6169 ^ n4537 ;
  assign n34313 = ( n5191 & ~n21828 ) | ( n5191 & n33637 ) | ( ~n21828 & n33637 ) ;
  assign n34314 = n5645 & n12429 ;
  assign n34315 = n34314 ^ n10140 ^ 1'b0 ;
  assign n34316 = ~n11746 & n34315 ;
  assign n34317 = n17808 ^ n7401 ^ 1'b0 ;
  assign n34318 = n12839 | n34317 ;
  assign n34319 = n28964 ^ n26950 ^ n5419 ;
  assign n34321 = n6829 | n9492 ;
  assign n34322 = n4911 & ~n34321 ;
  assign n34323 = n34322 ^ n8043 ^ 1'b0 ;
  assign n34320 = n5093 | n34206 ;
  assign n34324 = n34323 ^ n34320 ^ 1'b0 ;
  assign n34325 = n10988 ^ n10375 ^ 1'b0 ;
  assign n34326 = n16920 | n22929 ;
  assign n34327 = n34326 ^ n20332 ^ 1'b0 ;
  assign n34328 = n31029 & n34327 ;
  assign n34329 = ( ~n2640 & n19626 ) | ( ~n2640 & n31562 ) | ( n19626 & n31562 ) ;
  assign n34330 = n34329 ^ n32799 ^ 1'b0 ;
  assign n34332 = ( n2548 & n12100 ) | ( n2548 & ~n28702 ) | ( n12100 & ~n28702 ) ;
  assign n34331 = ( n3680 & n11998 ) | ( n3680 & ~n16247 ) | ( n11998 & ~n16247 ) ;
  assign n34333 = n34332 ^ n34331 ^ n12702 ;
  assign n34334 = n1001 | n2208 ;
  assign n34335 = n34334 ^ n21713 ^ 1'b0 ;
  assign n34336 = ( n8100 & n18768 ) | ( n8100 & ~n34335 ) | ( n18768 & ~n34335 ) ;
  assign n34337 = n24950 ^ n24089 ^ n13683 ;
  assign n34338 = n34337 ^ n13708 ^ n5036 ;
  assign n34339 = n2067 & n16317 ;
  assign n34340 = ( n18152 & ~n18669 ) | ( n18152 & n34339 ) | ( ~n18669 & n34339 ) ;
  assign n34341 = n31047 ^ n21030 ^ n11124 ;
  assign n34342 = n34341 ^ n31050 ^ n9827 ;
  assign n34343 = n33856 ^ n13567 ^ n7898 ;
  assign n34344 = n14570 ^ n11195 ^ n7956 ;
  assign n34345 = n20068 & ~n27322 ;
  assign n34346 = n12376 & n34345 ;
  assign n34347 = n10297 | n34346 ;
  assign n34348 = ( n4957 & n12714 ) | ( n4957 & n30866 ) | ( n12714 & n30866 ) ;
  assign n34349 = n34347 | n34348 ;
  assign n34350 = ( n13573 & n17862 ) | ( n13573 & n18350 ) | ( n17862 & n18350 ) ;
  assign n34351 = ( n4049 & n4763 ) | ( n4049 & ~n20558 ) | ( n4763 & ~n20558 ) ;
  assign n34352 = ( ~n11173 & n16855 ) | ( ~n11173 & n29239 ) | ( n16855 & n29239 ) ;
  assign n34353 = ( ~n34350 & n34351 ) | ( ~n34350 & n34352 ) | ( n34351 & n34352 ) ;
  assign n34354 = n34353 ^ n1676 ^ 1'b0 ;
  assign n34355 = ( ~n11370 & n16101 ) | ( ~n11370 & n23895 ) | ( n16101 & n23895 ) ;
  assign n34356 = n34355 ^ n33595 ^ 1'b0 ;
  assign n34357 = ( ~n5405 & n9429 ) | ( ~n5405 & n29687 ) | ( n9429 & n29687 ) ;
  assign n34358 = n27465 ^ n23007 ^ 1'b0 ;
  assign n34359 = n30022 & ~n34358 ;
  assign n34360 = n34359 ^ n8031 ^ n5739 ;
  assign n34361 = n7435 | n19562 ;
  assign n34362 = n32852 | n34361 ;
  assign n34363 = ( n1815 & n26009 ) | ( n1815 & ~n34362 ) | ( n26009 & ~n34362 ) ;
  assign n34364 = n19344 & n27866 ;
  assign n34365 = ( n6933 & n9153 ) | ( n6933 & n9573 ) | ( n9153 & n9573 ) ;
  assign n34366 = ( n1743 & n11187 ) | ( n1743 & ~n34365 ) | ( n11187 & ~n34365 ) ;
  assign n34367 = n21856 ^ n13288 ^ n2418 ;
  assign n34368 = n34367 ^ n15353 ^ n13558 ;
  assign n34369 = n20901 | n27689 ;
  assign n34370 = n34369 ^ n8600 ^ 1'b0 ;
  assign n34371 = ( n7901 & ~n9317 ) | ( n7901 & n23133 ) | ( ~n9317 & n23133 ) ;
  assign n34372 = n20972 ^ n11447 ^ 1'b0 ;
  assign n34373 = ( n7468 & n14765 ) | ( n7468 & ~n34372 ) | ( n14765 & ~n34372 ) ;
  assign n34374 = ( n2170 & n34371 ) | ( n2170 & ~n34373 ) | ( n34371 & ~n34373 ) ;
  assign n34375 = n33407 ^ n32128 ^ n9220 ;
  assign n34376 = n29895 & n34375 ;
  assign n34377 = n14472 ^ n11812 ^ n3610 ;
  assign n34378 = n34377 ^ n26570 ^ n13140 ;
  assign n34379 = ( n9218 & n26504 ) | ( n9218 & ~n34378 ) | ( n26504 & ~n34378 ) ;
  assign n34380 = n26633 ^ n26394 ^ n16299 ;
  assign n34381 = ( n4784 & ~n10938 ) | ( n4784 & n17251 ) | ( ~n10938 & n17251 ) ;
  assign n34382 = ( n10820 & ~n11348 ) | ( n10820 & n34381 ) | ( ~n11348 & n34381 ) ;
  assign n34383 = ( n8517 & n24108 ) | ( n8517 & n34382 ) | ( n24108 & n34382 ) ;
  assign n34384 = ( n7074 & n7964 ) | ( n7074 & n34383 ) | ( n7964 & n34383 ) ;
  assign n34385 = ( n32260 & ~n34380 ) | ( n32260 & n34384 ) | ( ~n34380 & n34384 ) ;
  assign n34386 = ( n7860 & n11012 ) | ( n7860 & n18173 ) | ( n11012 & n18173 ) ;
  assign n34387 = n34386 ^ n30760 ^ n28663 ;
  assign n34389 = ( n320 & ~n3562 ) | ( n320 & n9372 ) | ( ~n3562 & n9372 ) ;
  assign n34388 = ( n1268 & n23676 ) | ( n1268 & ~n24607 ) | ( n23676 & ~n24607 ) ;
  assign n34390 = n34389 ^ n34388 ^ n19397 ;
  assign n34393 = n15624 ^ n8844 ^ n4690 ;
  assign n34391 = ( n4669 & ~n8357 ) | ( n4669 & n18152 ) | ( ~n8357 & n18152 ) ;
  assign n34392 = x82 & n34391 ;
  assign n34394 = n34393 ^ n34392 ^ 1'b0 ;
  assign n34395 = n34394 ^ n27494 ^ 1'b0 ;
  assign n34396 = n34390 & ~n34395 ;
  assign n34401 = n33422 ^ n20953 ^ n6381 ;
  assign n34397 = ( n2117 & n13647 ) | ( n2117 & ~n18961 ) | ( n13647 & ~n18961 ) ;
  assign n34398 = n34397 ^ n8111 ^ n5172 ;
  assign n34399 = n18245 ^ n15401 ^ 1'b0 ;
  assign n34400 = ~n34398 & n34399 ;
  assign n34402 = n34401 ^ n34400 ^ n10626 ;
  assign n34403 = n24195 | n34402 ;
  assign n34404 = n10295 | n14435 ;
  assign n34405 = n34404 ^ n30608 ^ 1'b0 ;
  assign n34406 = n16683 | n34405 ;
  assign n34407 = n12485 ^ n11246 ^ 1'b0 ;
  assign n34408 = ~n8022 & n34407 ;
  assign n34409 = ( n822 & n7053 ) | ( n822 & n9640 ) | ( n7053 & n9640 ) ;
  assign n34410 = n34409 ^ n11946 ^ 1'b0 ;
  assign n34411 = n4759 & n34410 ;
  assign n34412 = n5507 & ~n24206 ;
  assign n34413 = ~n17591 & n34412 ;
  assign n34414 = ( n13430 & n25766 ) | ( n13430 & ~n34413 ) | ( n25766 & ~n34413 ) ;
  assign n34415 = ( ~n749 & n2626 ) | ( ~n749 & n19338 ) | ( n2626 & n19338 ) ;
  assign n34416 = ( ~n1352 & n2655 ) | ( ~n1352 & n34415 ) | ( n2655 & n34415 ) ;
  assign n34417 = ( n7544 & ~n10660 ) | ( n7544 & n25296 ) | ( ~n10660 & n25296 ) ;
  assign n34418 = n34234 ^ n25871 ^ x49 ;
  assign n34419 = ~n7948 & n34418 ;
  assign n34420 = n7919 | n29862 ;
  assign n34421 = n34420 ^ n19113 ^ n3766 ;
  assign n34422 = ( n34417 & ~n34419 ) | ( n34417 & n34421 ) | ( ~n34419 & n34421 ) ;
  assign n34423 = n4421 & ~n12570 ;
  assign n34424 = n34423 ^ n31977 ^ n17967 ;
  assign n34425 = n20385 ^ n19181 ^ n15741 ;
  assign n34426 = ( ~n7727 & n22672 ) | ( ~n7727 & n34425 ) | ( n22672 & n34425 ) ;
  assign n34427 = ~n10766 & n34426 ;
  assign n34428 = ~n30016 & n34427 ;
  assign n34429 = n6183 & n24827 ;
  assign n34430 = ( n3557 & n24796 ) | ( n3557 & ~n27502 ) | ( n24796 & ~n27502 ) ;
  assign n34431 = ( ~n11295 & n16419 ) | ( ~n11295 & n19485 ) | ( n16419 & n19485 ) ;
  assign n34432 = n28848 ^ n11478 ^ n1120 ;
  assign n34433 = n34431 | n34432 ;
  assign n34434 = n28271 & ~n34433 ;
  assign n34435 = ( ~n1276 & n17102 ) | ( ~n1276 & n30079 ) | ( n17102 & n30079 ) ;
  assign n34436 = n22897 ^ n18859 ^ n6868 ;
  assign n34437 = n34436 ^ n26127 ^ n19413 ;
  assign n34438 = n3708 & n32065 ;
  assign n34439 = n6495 ^ n5897 ^ n713 ;
  assign n34440 = ( n22931 & n34438 ) | ( n22931 & n34439 ) | ( n34438 & n34439 ) ;
  assign n34441 = n28372 ^ n12452 ^ 1'b0 ;
  assign n34442 = n34441 ^ n7513 ^ 1'b0 ;
  assign n34443 = n21534 & n34442 ;
  assign n34444 = n34443 ^ n14512 ^ n6965 ;
  assign n34445 = ( ~n10350 & n10957 ) | ( ~n10350 & n34444 ) | ( n10957 & n34444 ) ;
  assign n34446 = n10335 & ~n34445 ;
  assign n34448 = ~n1157 & n21309 ;
  assign n34449 = n11298 | n34448 ;
  assign n34447 = n26321 & n32142 ;
  assign n34450 = n34449 ^ n34447 ^ 1'b0 ;
  assign n34451 = ( n4675 & ~n10064 ) | ( n4675 & n14181 ) | ( ~n10064 & n14181 ) ;
  assign n34452 = n34451 ^ n8915 ^ 1'b0 ;
  assign n34453 = n6868 ^ n4479 ^ 1'b0 ;
  assign n34454 = ~n32987 & n34453 ;
  assign n34455 = n34454 ^ n29409 ^ n23310 ;
  assign n34456 = n23586 | n23728 ;
  assign n34457 = n34456 ^ n34055 ^ n4739 ;
  assign n34458 = n28391 ^ n6256 ^ n1775 ;
  assign n34459 = ( n5237 & n27556 ) | ( n5237 & n34458 ) | ( n27556 & n34458 ) ;
  assign n34460 = n34459 ^ n18661 ^ 1'b0 ;
  assign n34461 = n8669 & ~n9981 ;
  assign n34462 = n11933 ^ n4882 ^ x110 ;
  assign n34463 = n34462 ^ n662 ^ 1'b0 ;
  assign n34464 = n506 | n27199 ;
  assign n34465 = n34463 & ~n34464 ;
  assign n34466 = ~n8034 & n33396 ;
  assign n34467 = ( n17579 & n21318 ) | ( n17579 & n22391 ) | ( n21318 & n22391 ) ;
  assign n34468 = ( n30955 & n31860 ) | ( n30955 & n34467 ) | ( n31860 & n34467 ) ;
  assign n34469 = n24031 ^ n9226 ^ 1'b0 ;
  assign n34470 = n19675 & n34469 ;
  assign n34471 = n29157 ^ n26043 ^ n2378 ;
  assign n34472 = ( n7973 & n34470 ) | ( n7973 & n34471 ) | ( n34470 & n34471 ) ;
  assign n34473 = ( n14505 & n27686 ) | ( n14505 & n34472 ) | ( n27686 & n34472 ) ;
  assign n34474 = n34269 ^ n16018 ^ n12027 ;
  assign n34475 = ( ~n6866 & n9270 ) | ( ~n6866 & n34474 ) | ( n9270 & n34474 ) ;
  assign n34476 = n34475 ^ n18697 ^ n11521 ;
  assign n34477 = n34476 ^ n1139 ^ n442 ;
  assign n34478 = n24793 ^ n18735 ^ n5458 ;
  assign n34479 = n30022 & ~n31995 ;
  assign n34480 = n34479 ^ n14288 ^ 1'b0 ;
  assign n34481 = ( ~n3694 & n8650 ) | ( ~n3694 & n16115 ) | ( n8650 & n16115 ) ;
  assign n34482 = n34481 ^ n23139 ^ 1'b0 ;
  assign n34483 = n33621 | n34482 ;
  assign n34484 = n34483 ^ n21130 ^ 1'b0 ;
  assign n34491 = n26198 ^ n1140 ^ 1'b0 ;
  assign n34492 = ~n13190 & n34491 ;
  assign n34490 = ~n10061 & n25833 ;
  assign n34493 = n34492 ^ n34490 ^ n3705 ;
  assign n34485 = n2195 & n6856 ;
  assign n34486 = n6096 & n34485 ;
  assign n34487 = ( ~n1438 & n14016 ) | ( ~n1438 & n34486 ) | ( n14016 & n34486 ) ;
  assign n34488 = n34487 ^ n13599 ^ 1'b0 ;
  assign n34489 = n9842 | n34488 ;
  assign n34494 = n34493 ^ n34489 ^ n27287 ;
  assign n34495 = ( n1357 & n13688 ) | ( n1357 & ~n33422 ) | ( n13688 & ~n33422 ) ;
  assign n34496 = n32795 & n34495 ;
  assign n34497 = ( n17377 & n24689 ) | ( n17377 & n27574 ) | ( n24689 & n27574 ) ;
  assign n34500 = n34443 ^ n10147 ^ n3477 ;
  assign n34498 = n27841 ^ n25765 ^ n14317 ;
  assign n34499 = ( ~n12754 & n29072 ) | ( ~n12754 & n34498 ) | ( n29072 & n34498 ) ;
  assign n34501 = n34500 ^ n34499 ^ n5677 ;
  assign n34502 = ( n1308 & n6295 ) | ( n1308 & ~n12372 ) | ( n6295 & ~n12372 ) ;
  assign n34503 = n14455 ^ n7176 ^ n5670 ;
  assign n34504 = n15100 ^ n14387 ^ n6673 ;
  assign n34505 = ( n14999 & n34503 ) | ( n14999 & n34504 ) | ( n34503 & n34504 ) ;
  assign n34506 = ( n1515 & n2809 ) | ( n1515 & ~n23838 ) | ( n2809 & ~n23838 ) ;
  assign n34507 = n34506 ^ n19405 ^ n19227 ;
  assign n34508 = ~n12471 & n34507 ;
  assign n34509 = n34508 ^ n19061 ^ 1'b0 ;
  assign n34510 = n13142 & n34509 ;
  assign n34511 = n30143 ^ n23180 ^ n20319 ;
  assign n34512 = ( n8820 & n25652 ) | ( n8820 & ~n34511 ) | ( n25652 & ~n34511 ) ;
  assign n34513 = ( n6242 & n31885 ) | ( n6242 & ~n34512 ) | ( n31885 & ~n34512 ) ;
  assign n34514 = n28663 ^ n9530 ^ n2171 ;
  assign n34515 = n5854 & ~n19225 ;
  assign n34516 = n34515 ^ n20432 ^ n10485 ;
  assign n34517 = n22858 ^ n9752 ^ n9014 ;
  assign n34518 = ( n12960 & ~n27690 ) | ( n12960 & n34517 ) | ( ~n27690 & n34517 ) ;
  assign n34519 = n15692 ^ n9608 ^ 1'b0 ;
  assign n34520 = ~n32033 & n34519 ;
  assign n34521 = n33920 ^ n26283 ^ n15803 ;
  assign n34522 = n34521 ^ n15933 ^ n5385 ;
  assign n34523 = n30454 ^ n18936 ^ 1'b0 ;
  assign n34524 = n34523 ^ n16204 ^ n2179 ;
  assign n34525 = ( n3412 & n27447 ) | ( n3412 & n34524 ) | ( n27447 & n34524 ) ;
  assign n34533 = n4858 | n25407 ;
  assign n34532 = n13133 & n31774 ;
  assign n34526 = n1940 & ~n7391 ;
  assign n34527 = n34526 ^ n4713 ^ 1'b0 ;
  assign n34528 = n34527 ^ n15225 ^ n4236 ;
  assign n34529 = ( ~n1834 & n11799 ) | ( ~n1834 & n12588 ) | ( n11799 & n12588 ) ;
  assign n34530 = n34529 ^ n4687 ^ 1'b0 ;
  assign n34531 = ( n4675 & n34528 ) | ( n4675 & n34530 ) | ( n34528 & n34530 ) ;
  assign n34534 = n34533 ^ n34532 ^ n34531 ;
  assign n34535 = ( n7915 & ~n17586 ) | ( n7915 & n23105 ) | ( ~n17586 & n23105 ) ;
  assign n34536 = n34535 ^ n14199 ^ n11565 ;
  assign n34537 = ( n12105 & ~n21863 ) | ( n12105 & n34381 ) | ( ~n21863 & n34381 ) ;
  assign n34538 = n27679 ^ n13135 ^ n5079 ;
  assign n34539 = ( n13819 & n17941 ) | ( n13819 & n34538 ) | ( n17941 & n34538 ) ;
  assign n34540 = ( n7789 & ~n34537 ) | ( n7789 & n34539 ) | ( ~n34537 & n34539 ) ;
  assign n34541 = n10652 ^ n8026 ^ 1'b0 ;
  assign n34542 = n22394 ^ n18608 ^ n2963 ;
  assign n34543 = n34541 & n34542 ;
  assign n34544 = ~n33964 & n34543 ;
  assign n34545 = ( ~n1020 & n21213 ) | ( ~n1020 & n28932 ) | ( n21213 & n28932 ) ;
  assign n34546 = ( n12116 & ~n12990 ) | ( n12116 & n23299 ) | ( ~n12990 & n23299 ) ;
  assign n34547 = n34546 ^ n13788 ^ n5716 ;
  assign n34548 = n34547 ^ n12266 ^ n11466 ;
  assign n34549 = n34548 ^ n22852 ^ n11674 ;
  assign n34550 = ( n7757 & ~n15803 ) | ( n7757 & n28058 ) | ( ~n15803 & n28058 ) ;
  assign n34551 = ( n4666 & ~n21555 ) | ( n4666 & n22481 ) | ( ~n21555 & n22481 ) ;
  assign n34552 = ( n7368 & n34550 ) | ( n7368 & ~n34551 ) | ( n34550 & ~n34551 ) ;
  assign n34553 = n14117 ^ n13374 ^ n13211 ;
  assign n34554 = ( n7536 & ~n16142 ) | ( n7536 & n22517 ) | ( ~n16142 & n22517 ) ;
  assign n34555 = n31880 ^ n18658 ^ n12563 ;
  assign n34556 = ( n504 & n7235 ) | ( n504 & n24441 ) | ( n7235 & n24441 ) ;
  assign n34557 = n3820 | n17042 ;
  assign n34558 = n17084 & ~n34557 ;
  assign n34559 = ~n24940 & n32594 ;
  assign n34560 = n34558 & n34559 ;
  assign n34561 = ~n1592 & n23506 ;
  assign n34562 = ( n3090 & n10145 ) | ( n3090 & ~n12129 ) | ( n10145 & ~n12129 ) ;
  assign n34563 = n28556 ^ n24993 ^ n7887 ;
  assign n34564 = n5909 ^ n3207 ^ 1'b0 ;
  assign n34565 = n8868 & ~n34564 ;
  assign n34566 = ( n6904 & n17677 ) | ( n6904 & n34565 ) | ( n17677 & n34565 ) ;
  assign n34567 = n34566 ^ n20639 ^ n4407 ;
  assign n34568 = ( n2195 & n34563 ) | ( n2195 & ~n34567 ) | ( n34563 & ~n34567 ) ;
  assign n34569 = n34568 ^ n26131 ^ 1'b0 ;
  assign n34570 = ( n12201 & n16548 ) | ( n12201 & n24365 ) | ( n16548 & n24365 ) ;
  assign n34572 = ( ~n9426 & n18025 ) | ( ~n9426 & n24970 ) | ( n18025 & n24970 ) ;
  assign n34571 = n11777 & n18447 ;
  assign n34573 = n34572 ^ n34571 ^ 1'b0 ;
  assign n34574 = n9405 | n10687 ;
  assign n34575 = n34574 ^ n4128 ^ 1'b0 ;
  assign n34585 = ~n8669 & n34247 ;
  assign n34578 = n11334 & n12671 ;
  assign n34579 = n34578 ^ n24278 ^ 1'b0 ;
  assign n34580 = n12408 & ~n34579 ;
  assign n34581 = n34580 ^ n1211 ^ 1'b0 ;
  assign n34582 = ( ~n16372 & n28188 ) | ( ~n16372 & n34581 ) | ( n28188 & n34581 ) ;
  assign n34576 = n11888 ^ n6847 ^ 1'b0 ;
  assign n34577 = n34576 ^ n5645 ^ x79 ;
  assign n34583 = n34582 ^ n34577 ^ n5706 ;
  assign n34584 = n34583 ^ n27469 ^ n22340 ;
  assign n34586 = n34585 ^ n34584 ^ n7303 ;
  assign n34592 = n2638 & n20317 ;
  assign n34593 = n34592 ^ n26073 ^ 1'b0 ;
  assign n34590 = ~n4576 & n25378 ;
  assign n34591 = n4459 & n34590 ;
  assign n34594 = n34593 ^ n34591 ^ n6700 ;
  assign n34587 = ( n1739 & n5862 ) | ( n1739 & ~n12291 ) | ( n5862 & ~n12291 ) ;
  assign n34588 = ~n21467 & n34587 ;
  assign n34589 = ( n9068 & n20583 ) | ( n9068 & ~n34588 ) | ( n20583 & ~n34588 ) ;
  assign n34595 = n34594 ^ n34589 ^ n27153 ;
  assign n34598 = n17476 ^ n16272 ^ 1'b0 ;
  assign n34596 = n8927 ^ n6765 ^ 1'b0 ;
  assign n34597 = n34596 ^ n12804 ^ x60 ;
  assign n34599 = n34598 ^ n34597 ^ n18878 ;
  assign n34600 = n10618 ^ n2421 ^ 1'b0 ;
  assign n34601 = ( n1952 & ~n17159 ) | ( n1952 & n34191 ) | ( ~n17159 & n34191 ) ;
  assign n34602 = ( ~x124 & n7842 ) | ( ~x124 & n25643 ) | ( n7842 & n25643 ) ;
  assign n34603 = ( ~n7829 & n34601 ) | ( ~n7829 & n34602 ) | ( n34601 & n34602 ) ;
  assign n34604 = ~n8407 & n28681 ;
  assign n34605 = n34604 ^ n20987 ^ n3360 ;
  assign n34606 = n34508 ^ n26791 ^ n1999 ;
  assign n34607 = n17093 ^ n14787 ^ 1'b0 ;
  assign n34608 = n12638 & ~n34607 ;
  assign n34609 = n34608 ^ n12609 ^ n10049 ;
  assign n34610 = n27749 ^ n24983 ^ 1'b0 ;
  assign n34611 = n20234 ^ n19967 ^ n6004 ;
  assign n34612 = n24430 ^ n6966 ^ 1'b0 ;
  assign n34613 = n34611 | n34612 ;
  assign n34614 = n8981 | n34613 ;
  assign n34615 = ( n10390 & ~n34610 ) | ( n10390 & n34614 ) | ( ~n34610 & n34614 ) ;
  assign n34616 = n34615 ^ n30562 ^ n850 ;
  assign n34617 = ( n6505 & ~n15664 ) | ( n6505 & n31120 ) | ( ~n15664 & n31120 ) ;
  assign n34618 = ( n14180 & n19373 ) | ( n14180 & ~n34617 ) | ( n19373 & ~n34617 ) ;
  assign n34619 = n34618 ^ n9764 ^ 1'b0 ;
  assign n34620 = n20767 & ~n31588 ;
  assign n34621 = n34620 ^ n5218 ^ 1'b0 ;
  assign n34622 = n27949 ^ n13818 ^ 1'b0 ;
  assign n34623 = n34622 ^ n24350 ^ n10428 ;
  assign n34624 = n8551 | n10210 ;
  assign n34625 = n34624 ^ n17841 ^ 1'b0 ;
  assign n34626 = n17065 ^ n5787 ^ 1'b0 ;
  assign n34627 = ~n2524 & n34626 ;
  assign n34628 = ( n25071 & n34625 ) | ( n25071 & ~n34627 ) | ( n34625 & ~n34627 ) ;
  assign n34629 = n7884 ^ n4230 ^ n1044 ;
  assign n34630 = n34629 ^ n26620 ^ n4223 ;
  assign n34631 = ( n4272 & n16178 ) | ( n4272 & n34630 ) | ( n16178 & n34630 ) ;
  assign n34632 = n8118 & ~n34631 ;
  assign n34637 = ( n3990 & n20348 ) | ( n3990 & ~n32781 ) | ( n20348 & ~n32781 ) ;
  assign n34635 = n32186 ^ n9266 ^ n4748 ;
  assign n34633 = x185 & n21972 ;
  assign n34634 = ~n4308 & n34633 ;
  assign n34636 = n34635 ^ n34634 ^ n27375 ;
  assign n34638 = n34637 ^ n34636 ^ n28361 ;
  assign n34639 = n6439 ^ x47 ^ 1'b0 ;
  assign n34640 = n9641 ^ n2162 ^ 1'b0 ;
  assign n34641 = n34640 ^ n16822 ^ 1'b0 ;
  assign n34642 = n34639 & n34641 ;
  assign n34643 = ~n25830 & n34642 ;
  assign n34644 = ( n4749 & n6398 ) | ( n4749 & n15355 ) | ( n6398 & n15355 ) ;
  assign n34645 = n34644 ^ x15 ^ 1'b0 ;
  assign n34646 = ~n32665 & n34645 ;
  assign n34647 = ( n3230 & ~n4520 ) | ( n3230 & n14910 ) | ( ~n4520 & n14910 ) ;
  assign n34648 = n34647 ^ n12233 ^ n11585 ;
  assign n34649 = ( ~n518 & n2566 ) | ( ~n518 & n4081 ) | ( n2566 & n4081 ) ;
  assign n34650 = n18724 ^ n6527 ^ n2832 ;
  assign n34651 = n34649 | n34650 ;
  assign n34652 = n34651 ^ n30627 ^ n12930 ;
  assign n34653 = n19864 ^ n6796 ^ n4452 ;
  assign n34654 = n34653 ^ n24330 ^ n12765 ;
  assign n34655 = ( ~n3305 & n22889 ) | ( ~n3305 & n34654 ) | ( n22889 & n34654 ) ;
  assign n34656 = ( n4670 & n7930 ) | ( n4670 & n14288 ) | ( n7930 & n14288 ) ;
  assign n34657 = n28399 | n34656 ;
  assign n34658 = n24537 ^ n1945 ^ 1'b0 ;
  assign n34659 = n21068 | n34658 ;
  assign n34660 = n34659 ^ n18311 ^ n949 ;
  assign n34661 = ( n17995 & n19780 ) | ( n17995 & n28327 ) | ( n19780 & n28327 ) ;
  assign n34662 = n34661 ^ n22447 ^ n1288 ;
  assign n34663 = n2636 | n27701 ;
  assign n34664 = n1704 | n34663 ;
  assign n34665 = n6842 | n33738 ;
  assign n34666 = ( ~n19862 & n22972 ) | ( ~n19862 & n34665 ) | ( n22972 & n34665 ) ;
  assign n34667 = n33470 ^ n9797 ^ n1707 ;
  assign n34668 = ( ~n12786 & n26021 ) | ( ~n12786 & n34667 ) | ( n26021 & n34667 ) ;
  assign n34672 = ( n441 & n5822 ) | ( n441 & n8338 ) | ( n5822 & n8338 ) ;
  assign n34669 = ( n5215 & ~n12667 ) | ( n5215 & n28065 ) | ( ~n12667 & n28065 ) ;
  assign n34670 = n34669 ^ n19750 ^ 1'b0 ;
  assign n34671 = n21045 & ~n34670 ;
  assign n34673 = n34672 ^ n34671 ^ n15976 ;
  assign n34674 = n3504 & n16023 ;
  assign n34675 = n24566 | n28861 ;
  assign n34676 = n34675 ^ n10308 ^ 1'b0 ;
  assign n34677 = ( n17372 & ~n34674 ) | ( n17372 & n34676 ) | ( ~n34674 & n34676 ) ;
  assign n34678 = n5963 & n16879 ;
  assign n34679 = n34678 ^ n26008 ^ n13668 ;
  assign n34680 = ( n34673 & n34677 ) | ( n34673 & ~n34679 ) | ( n34677 & ~n34679 ) ;
  assign n34681 = n31895 ^ n31574 ^ 1'b0 ;
  assign n34682 = n32177 ^ n22008 ^ 1'b0 ;
  assign n34683 = n2623 & n34682 ;
  assign n34686 = n14062 ^ n13077 ^ n12813 ;
  assign n34684 = n11076 ^ n3617 ^ n1355 ;
  assign n34685 = x27 & ~n34684 ;
  assign n34687 = n34686 ^ n34685 ^ 1'b0 ;
  assign n34688 = n30089 ^ n16573 ^ 1'b0 ;
  assign n34689 = n17000 | n34688 ;
  assign n34690 = n30179 ^ n5784 ^ n3406 ;
  assign n34691 = n17088 ^ n7840 ^ n1512 ;
  assign n34692 = n3843 | n34691 ;
  assign n34693 = ( n16957 & n23199 ) | ( n16957 & ~n26820 ) | ( n23199 & ~n26820 ) ;
  assign n34694 = n34693 ^ n4913 ^ 1'b0 ;
  assign n34695 = n21863 & ~n25994 ;
  assign n34696 = ~n34694 & n34695 ;
  assign n34697 = n34696 ^ n14064 ^ n11143 ;
  assign n34698 = n5834 & ~n34697 ;
  assign n34699 = ( ~n10321 & n15339 ) | ( ~n10321 & n16574 ) | ( n15339 & n16574 ) ;
  assign n34700 = ~n13714 & n25797 ;
  assign n34701 = n34700 ^ n29400 ^ 1'b0 ;
  assign n34702 = ( n5363 & n18590 ) | ( n5363 & n34701 ) | ( n18590 & n34701 ) ;
  assign n34706 = n11351 ^ n4090 ^ n1106 ;
  assign n34705 = n23958 ^ n8426 ^ n512 ;
  assign n34703 = n26492 ^ n20735 ^ n19008 ;
  assign n34704 = n34703 ^ n9936 ^ n4575 ;
  assign n34707 = n34706 ^ n34705 ^ n34704 ;
  assign n34708 = n22845 | n24356 ;
  assign n34711 = ( n6900 & n12259 ) | ( n6900 & ~n16807 ) | ( n12259 & ~n16807 ) ;
  assign n34709 = n30563 ^ n6148 ^ n5270 ;
  assign n34710 = n34709 ^ n19394 ^ n1255 ;
  assign n34712 = n34711 ^ n34710 ^ n20812 ;
  assign n34713 = n29799 ^ n23137 ^ n2233 ;
  assign n34714 = ( ~n15488 & n31355 ) | ( ~n15488 & n32347 ) | ( n31355 & n32347 ) ;
  assign n34716 = ( n9367 & ~n19633 ) | ( n9367 & n32581 ) | ( ~n19633 & n32581 ) ;
  assign n34715 = ~n6573 & n20246 ;
  assign n34717 = n34716 ^ n34715 ^ 1'b0 ;
  assign n34718 = n3774 & n17424 ;
  assign n34719 = n8072 ^ n970 ^ 1'b0 ;
  assign n34720 = ~n6765 & n15135 ;
  assign n34721 = n34720 ^ n2973 ^ 1'b0 ;
  assign n34722 = n34721 ^ n10562 ^ n1614 ;
  assign n34723 = ( n4310 & n34719 ) | ( n4310 & n34722 ) | ( n34719 & n34722 ) ;
  assign n34724 = n30524 ^ n25057 ^ n2981 ;
  assign n34727 = n30487 ^ n26712 ^ n26028 ;
  assign n34725 = n26429 ^ n18924 ^ n4642 ;
  assign n34726 = ( ~x119 & n23730 ) | ( ~x119 & n34725 ) | ( n23730 & n34725 ) ;
  assign n34728 = n34727 ^ n34726 ^ 1'b0 ;
  assign n34729 = n8396 & ~n34728 ;
  assign n34730 = n32736 ^ n7258 ^ 1'b0 ;
  assign n34733 = ( ~n7342 & n11391 ) | ( ~n7342 & n14981 ) | ( n11391 & n14981 ) ;
  assign n34731 = n11361 ^ n10891 ^ 1'b0 ;
  assign n34732 = n14221 & n34731 ;
  assign n34734 = n34733 ^ n34732 ^ n9198 ;
  assign n34735 = n32587 ^ n21482 ^ n3823 ;
  assign n34736 = ( ~n2588 & n17251 ) | ( ~n2588 & n33554 ) | ( n17251 & n33554 ) ;
  assign n34737 = ( n14201 & n19774 ) | ( n14201 & n34736 ) | ( n19774 & n34736 ) ;
  assign n34738 = n34737 ^ n18059 ^ n5012 ;
  assign n34739 = ( n15085 & ~n24858 ) | ( n15085 & n27759 ) | ( ~n24858 & n27759 ) ;
  assign n34740 = ( n34735 & n34738 ) | ( n34735 & ~n34739 ) | ( n34738 & ~n34739 ) ;
  assign n34741 = ( n9559 & n26533 ) | ( n9559 & ~n30429 ) | ( n26533 & ~n30429 ) ;
  assign n34742 = ( ~n283 & n6041 ) | ( ~n283 & n29582 ) | ( n6041 & n29582 ) ;
  assign n34743 = ( n10126 & ~n11302 ) | ( n10126 & n17764 ) | ( ~n11302 & n17764 ) ;
  assign n34744 = ( n14068 & ~n18788 ) | ( n14068 & n30207 ) | ( ~n18788 & n30207 ) ;
  assign n34745 = ( n8773 & n17514 ) | ( n8773 & ~n24751 ) | ( n17514 & ~n24751 ) ;
  assign n34746 = n16977 & n34745 ;
  assign n34747 = ~n14756 & n34746 ;
  assign n34748 = n20761 ^ n15874 ^ 1'b0 ;
  assign n34749 = n18476 ^ n5889 ^ 1'b0 ;
  assign n34750 = ( n1274 & n10128 ) | ( n1274 & n20665 ) | ( n10128 & n20665 ) ;
  assign n34751 = n34541 ^ n12405 ^ n8791 ;
  assign n34752 = ( n4002 & n7522 ) | ( n4002 & ~n23524 ) | ( n7522 & ~n23524 ) ;
  assign n34753 = ( ~n14078 & n16553 ) | ( ~n14078 & n20464 ) | ( n16553 & n20464 ) ;
  assign n34754 = ( n6789 & ~n30431 ) | ( n6789 & n34753 ) | ( ~n30431 & n34753 ) ;
  assign n34755 = n34754 ^ n5147 ^ 1'b0 ;
  assign n34756 = ( ~n17289 & n26231 ) | ( ~n17289 & n33202 ) | ( n26231 & n33202 ) ;
  assign n34757 = n34756 ^ n31980 ^ n11398 ;
  assign n34758 = n1072 & ~n19856 ;
  assign n34759 = ( n9981 & n18789 ) | ( n9981 & ~n27221 ) | ( n18789 & ~n27221 ) ;
  assign n34760 = n12172 | n34759 ;
  assign n34761 = n34760 ^ n8461 ^ 1'b0 ;
  assign n34769 = ( n10860 & n11379 ) | ( n10860 & ~n17431 ) | ( n11379 & ~n17431 ) ;
  assign n34766 = ( ~n22131 & n26945 ) | ( ~n22131 & n30625 ) | ( n26945 & n30625 ) ;
  assign n34765 = n5808 & ~n25143 ;
  assign n34767 = n34766 ^ n34765 ^ 1'b0 ;
  assign n34768 = n1646 & n34767 ;
  assign n34762 = n12003 & n16619 ;
  assign n34763 = n34762 ^ n14641 ^ 1'b0 ;
  assign n34764 = ( n2617 & ~n14948 ) | ( n2617 & n34763 ) | ( ~n14948 & n34763 ) ;
  assign n34770 = n34769 ^ n34768 ^ n34764 ;
  assign n34771 = ( n6465 & ~n14287 ) | ( n6465 & n24994 ) | ( ~n14287 & n24994 ) ;
  assign n34775 = n14099 ^ n5736 ^ n2825 ;
  assign n34772 = n33664 ^ n11004 ^ n10537 ;
  assign n34773 = n13620 | n34772 ;
  assign n34774 = n34773 ^ n16145 ^ 1'b0 ;
  assign n34776 = n34775 ^ n34774 ^ n14518 ;
  assign n34777 = ~n16433 & n32102 ;
  assign n34778 = n2839 & n34777 ;
  assign n34779 = ( n28065 & n28743 ) | ( n28065 & n34778 ) | ( n28743 & n34778 ) ;
  assign n34780 = n11841 ^ n5822 ^ 1'b0 ;
  assign n34781 = n28851 | n34780 ;
  assign n34782 = n26189 ^ n12382 ^ 1'b0 ;
  assign n34783 = ~n19806 & n34782 ;
  assign n34784 = n34783 ^ n9474 ^ 1'b0 ;
  assign n34785 = ( n3633 & n5616 ) | ( n3633 & ~n32987 ) | ( n5616 & ~n32987 ) ;
  assign n34786 = n23277 ^ n7738 ^ n1565 ;
  assign n34787 = n30299 ^ n15003 ^ n10168 ;
  assign n34788 = ( x11 & ~n31036 ) | ( x11 & n34787 ) | ( ~n31036 & n34787 ) ;
  assign n34790 = ~n12516 & n18576 ;
  assign n34791 = n19459 & n34790 ;
  assign n34789 = n10868 & ~n27177 ;
  assign n34792 = n34791 ^ n34789 ^ n8430 ;
  assign n34793 = ~n4093 & n15272 ;
  assign n34794 = ~n10173 & n34793 ;
  assign n34795 = ( n3676 & n14008 ) | ( n3676 & n34794 ) | ( n14008 & n34794 ) ;
  assign n34796 = ( n623 & ~n4379 ) | ( n623 & n6637 ) | ( ~n4379 & n6637 ) ;
  assign n34797 = ( ~n34263 & n34795 ) | ( ~n34263 & n34796 ) | ( n34795 & n34796 ) ;
  assign n34798 = n22803 ^ n5691 ^ 1'b0 ;
  assign n34799 = ( n7292 & n14385 ) | ( n7292 & n34798 ) | ( n14385 & n34798 ) ;
  assign n34800 = ( n10516 & ~n11112 ) | ( n10516 & n11113 ) | ( ~n11112 & n11113 ) ;
  assign n34801 = n1890 & ~n10543 ;
  assign n34802 = n34801 ^ n30826 ^ n2074 ;
  assign n34803 = ( n27643 & ~n34800 ) | ( n27643 & n34802 ) | ( ~n34800 & n34802 ) ;
  assign n34804 = ( n8663 & ~n17217 ) | ( n8663 & n32804 ) | ( ~n17217 & n32804 ) ;
  assign n34805 = n33702 ^ n30419 ^ n21037 ;
  assign n34807 = n29339 ^ n2875 ^ n2063 ;
  assign n34806 = ( ~n15448 & n21165 ) | ( ~n15448 & n22411 ) | ( n21165 & n22411 ) ;
  assign n34808 = n34807 ^ n34806 ^ 1'b0 ;
  assign n34809 = n34808 ^ n28836 ^ n874 ;
  assign n34810 = n30613 ^ n26549 ^ n4901 ;
  assign n34811 = n32680 & n34810 ;
  assign n34812 = n31603 ^ n22169 ^ n19959 ;
  assign n34813 = n34812 ^ n11377 ^ 1'b0 ;
  assign n34814 = n28364 ^ n14313 ^ n11897 ;
  assign n34815 = ( n14589 & n16031 ) | ( n14589 & ~n34814 ) | ( n16031 & ~n34814 ) ;
  assign n34816 = n1663 ^ n1310 ^ 1'b0 ;
  assign n34817 = n16168 ^ n8589 ^ 1'b0 ;
  assign n34818 = n22811 & n34817 ;
  assign n34819 = n3365 & n34818 ;
  assign n34820 = n3421 & n13044 ;
  assign n34821 = n15388 & n34820 ;
  assign n34822 = n17210 | n32300 ;
  assign n34823 = n34822 ^ n20748 ^ n11280 ;
  assign n34824 = ( n21633 & n34821 ) | ( n21633 & n34823 ) | ( n34821 & n34823 ) ;
  assign n34825 = n6202 & ~n34824 ;
  assign n34826 = n34825 ^ n3682 ^ 1'b0 ;
  assign n34827 = n13996 ^ n6321 ^ n5870 ;
  assign n34828 = n21090 ^ n16520 ^ n7084 ;
  assign n34829 = n34828 ^ n28976 ^ n4411 ;
  assign n34830 = ( n1547 & ~n9830 ) | ( n1547 & n20639 ) | ( ~n9830 & n20639 ) ;
  assign n34831 = ( n21713 & n34829 ) | ( n21713 & ~n34830 ) | ( n34829 & ~n34830 ) ;
  assign n34832 = n1991 | n13273 ;
  assign n34833 = n34832 ^ n5310 ^ 1'b0 ;
  assign n34834 = n34833 ^ n19912 ^ 1'b0 ;
  assign n34836 = n7110 ^ n6495 ^ n777 ;
  assign n34835 = ( ~n6223 & n8928 ) | ( ~n6223 & n11937 ) | ( n8928 & n11937 ) ;
  assign n34837 = n34836 ^ n34835 ^ n20558 ;
  assign n34838 = ( n7679 & ~n21668 ) | ( n7679 & n21713 ) | ( ~n21668 & n21713 ) ;
  assign n34839 = n27574 | n28835 ;
  assign n34840 = n17398 | n34839 ;
  assign n34841 = n7150 & ~n34840 ;
  assign n34842 = n6874 & n28422 ;
  assign n34843 = n34842 ^ n19901 ^ n10126 ;
  assign n34844 = n21564 ^ n14861 ^ 1'b0 ;
  assign n34845 = ~n24289 & n34844 ;
  assign n34846 = n34845 ^ n24970 ^ n13399 ;
  assign n34847 = ( n8169 & ~n27324 ) | ( n8169 & n34846 ) | ( ~n27324 & n34846 ) ;
  assign n34848 = ( n2024 & n6335 ) | ( n2024 & n12580 ) | ( n6335 & n12580 ) ;
  assign n34849 = n34848 ^ n19381 ^ n4462 ;
  assign n34850 = n15571 ^ n8782 ^ n2776 ;
  assign n34851 = ~n4591 & n6958 ;
  assign n34852 = n26833 ^ n2967 ^ n1370 ;
  assign n34853 = n31814 ^ n28340 ^ n3215 ;
  assign n34854 = n16951 ^ n6946 ^ 1'b0 ;
  assign n34855 = ( n1103 & n3186 ) | ( n1103 & ~n4581 ) | ( n3186 & ~n4581 ) ;
  assign n34856 = n34855 ^ n9634 ^ 1'b0 ;
  assign n34857 = n24294 | n34856 ;
  assign n34858 = ~n3878 & n24172 ;
  assign n34859 = n5940 & n34858 ;
  assign n34860 = n34859 ^ n23402 ^ n4482 ;
  assign n34861 = n34860 ^ n24244 ^ 1'b0 ;
  assign n34863 = ( n4777 & n6937 ) | ( n4777 & ~n20479 ) | ( n6937 & ~n20479 ) ;
  assign n34864 = ( n8423 & n11671 ) | ( n8423 & n34863 ) | ( n11671 & n34863 ) ;
  assign n34865 = n7596 & n34864 ;
  assign n34866 = n34865 ^ n32690 ^ 1'b0 ;
  assign n34862 = n14635 & ~n17861 ;
  assign n34867 = n34866 ^ n34862 ^ n9563 ;
  assign n34868 = n26879 ^ n8494 ^ n8333 ;
  assign n34869 = n29717 ^ n21107 ^ 1'b0 ;
  assign n34870 = ( n21872 & n26760 ) | ( n21872 & ~n34492 ) | ( n26760 & ~n34492 ) ;
  assign n34871 = n34870 ^ n17016 ^ 1'b0 ;
  assign n34872 = n17087 & n33159 ;
  assign n34873 = ~n8632 & n34872 ;
  assign n34874 = ( n15630 & ~n16193 ) | ( n15630 & n28568 ) | ( ~n16193 & n28568 ) ;
  assign n34875 = n34874 ^ n8471 ^ n4217 ;
  assign n34878 = ( n4194 & n9756 ) | ( n4194 & n11385 ) | ( n9756 & n11385 ) ;
  assign n34876 = n7768 & n31299 ;
  assign n34877 = n23089 & n34876 ;
  assign n34879 = n34878 ^ n34877 ^ n13288 ;
  assign n34880 = n15843 ^ n5521 ^ n2909 ;
  assign n34881 = ( n378 & ~n4323 ) | ( n378 & n20479 ) | ( ~n4323 & n20479 ) ;
  assign n34884 = n13940 ^ n3936 ^ n1410 ;
  assign n34882 = n28624 ^ n16599 ^ 1'b0 ;
  assign n34883 = ~n22633 & n34882 ;
  assign n34885 = n34884 ^ n34883 ^ n26212 ;
  assign n34886 = ( n5764 & n29080 ) | ( n5764 & ~n34885 ) | ( n29080 & ~n34885 ) ;
  assign n34887 = ( n24065 & n34881 ) | ( n24065 & ~n34886 ) | ( n34881 & ~n34886 ) ;
  assign n34888 = ( n1671 & n9066 ) | ( n1671 & ~n34887 ) | ( n9066 & ~n34887 ) ;
  assign n34890 = ( ~n1903 & n9485 ) | ( ~n1903 & n10412 ) | ( n9485 & n10412 ) ;
  assign n34889 = n7420 & n16141 ;
  assign n34891 = n34890 ^ n34889 ^ 1'b0 ;
  assign n34892 = n22255 ^ n488 ^ 1'b0 ;
  assign n34893 = ( n26747 & ~n31678 ) | ( n26747 & n34892 ) | ( ~n31678 & n34892 ) ;
  assign n34894 = n34893 ^ n10840 ^ n7546 ;
  assign n34895 = n9013 & n16471 ;
  assign n34896 = n34895 ^ n7109 ^ 1'b0 ;
  assign n34897 = ( n6023 & n34894 ) | ( n6023 & ~n34896 ) | ( n34894 & ~n34896 ) ;
  assign n34898 = n21059 ^ n2904 ^ 1'b0 ;
  assign n34899 = n6430 & ~n34898 ;
  assign n34903 = ( n1509 & n10551 ) | ( n1509 & ~n11702 ) | ( n10551 & ~n11702 ) ;
  assign n34900 = n9780 & ~n21582 ;
  assign n34901 = n34900 ^ n33792 ^ 1'b0 ;
  assign n34902 = n34901 ^ n26859 ^ n1789 ;
  assign n34904 = n34903 ^ n34902 ^ n25113 ;
  assign n34905 = ( n28625 & ~n34899 ) | ( n28625 & n34904 ) | ( ~n34899 & n34904 ) ;
  assign n34906 = n2393 & ~n10039 ;
  assign n34910 = n14683 ^ n9619 ^ n5110 ;
  assign n34908 = n13049 ^ n5211 ^ 1'b0 ;
  assign n34909 = n34908 ^ n11457 ^ n5391 ;
  assign n34907 = ( n1935 & n19146 ) | ( n1935 & n32444 ) | ( n19146 & n32444 ) ;
  assign n34911 = n34910 ^ n34909 ^ n34907 ;
  assign n34912 = ( n1942 & n6071 ) | ( n1942 & ~n34006 ) | ( n6071 & ~n34006 ) ;
  assign n34913 = ( ~n16584 & n23126 ) | ( ~n16584 & n34912 ) | ( n23126 & n34912 ) ;
  assign n34914 = n31688 | n34913 ;
  assign n34917 = ( ~n5224 & n12452 ) | ( ~n5224 & n13138 ) | ( n12452 & n13138 ) ;
  assign n34915 = n7026 & ~n8007 ;
  assign n34916 = n9810 & n34915 ;
  assign n34918 = n34917 ^ n34916 ^ n5727 ;
  assign n34919 = n21341 ^ n20607 ^ n1091 ;
  assign n34920 = n20450 ^ n14008 ^ n3563 ;
  assign n34921 = n1977 | n8453 ;
  assign n34923 = n27125 ^ n2240 ^ n1462 ;
  assign n34922 = n14524 ^ n8962 ^ n3975 ;
  assign n34924 = n34923 ^ n34922 ^ n3246 ;
  assign n34925 = n34924 ^ n31948 ^ x200 ;
  assign n34944 = ( n4562 & n5035 ) | ( n4562 & ~n18634 ) | ( n5035 & ~n18634 ) ;
  assign n34945 = ( n2468 & ~n7505 ) | ( n2468 & n34944 ) | ( ~n7505 & n34944 ) ;
  assign n34935 = n19454 ^ n2937 ^ 1'b0 ;
  assign n34926 = ~n5243 & n10009 ;
  assign n34927 = n7940 & n34926 ;
  assign n34928 = n9790 ^ n7169 ^ x18 ;
  assign n34929 = n34928 ^ n6436 ^ n6124 ;
  assign n34932 = ( ~n901 & n4885 ) | ( ~n901 & n30889 ) | ( n4885 & n30889 ) ;
  assign n34930 = n21373 ^ n15886 ^ 1'b0 ;
  assign n34931 = ( n29472 & n34213 ) | ( n29472 & ~n34930 ) | ( n34213 & ~n34930 ) ;
  assign n34933 = n34932 ^ n34931 ^ n32879 ;
  assign n34934 = ( n34927 & ~n34929 ) | ( n34927 & n34933 ) | ( ~n34929 & n34933 ) ;
  assign n34936 = n34935 ^ n34934 ^ n6744 ;
  assign n34938 = n12994 ^ n11210 ^ n7144 ;
  assign n34937 = ( ~n571 & n8705 ) | ( ~n571 & n26968 ) | ( n8705 & n26968 ) ;
  assign n34939 = n34938 ^ n34937 ^ n34916 ;
  assign n34940 = n34939 ^ n29696 ^ n29436 ;
  assign n34941 = n30420 & n34940 ;
  assign n34942 = n34936 & n34941 ;
  assign n34943 = n4038 | n34942 ;
  assign n34946 = n34945 ^ n34943 ^ 1'b0 ;
  assign n34947 = ( n8359 & n23377 ) | ( n8359 & n26860 ) | ( n23377 & n26860 ) ;
  assign n34951 = ( ~n2052 & n3208 ) | ( ~n2052 & n7378 ) | ( n3208 & n7378 ) ;
  assign n34952 = ( n1443 & ~n5762 ) | ( n1443 & n34951 ) | ( ~n5762 & n34951 ) ;
  assign n34948 = ( ~n1039 & n1978 ) | ( ~n1039 & n8350 ) | ( n1978 & n8350 ) ;
  assign n34949 = ( ~n4254 & n10895 ) | ( ~n4254 & n34948 ) | ( n10895 & n34948 ) ;
  assign n34950 = n26112 & ~n34949 ;
  assign n34953 = n34952 ^ n34950 ^ 1'b0 ;
  assign n34954 = n16436 | n34953 ;
  assign n34955 = n34947 | n34954 ;
  assign n34956 = ( ~n8822 & n16166 ) | ( ~n8822 & n29542 ) | ( n16166 & n29542 ) ;
  assign n34957 = n34956 ^ n29828 ^ n21967 ;
  assign n34958 = n34957 ^ n17817 ^ n16011 ;
  assign n34959 = n7245 | n10475 ;
  assign n34960 = n13673 & n34959 ;
  assign n34961 = ~n6953 & n34960 ;
  assign n34962 = ~n7096 & n34961 ;
  assign n34963 = n34962 ^ n33795 ^ n30848 ;
  assign n34966 = ( n680 & ~n6328 ) | ( n680 & n23503 ) | ( ~n6328 & n23503 ) ;
  assign n34964 = ( n2147 & n22654 ) | ( n2147 & n30818 ) | ( n22654 & n30818 ) ;
  assign n34965 = ( ~n2429 & n9301 ) | ( ~n2429 & n34964 ) | ( n9301 & n34964 ) ;
  assign n34967 = n34966 ^ n34965 ^ n5304 ;
  assign n34968 = n34438 ^ n15413 ^ 1'b0 ;
  assign n34969 = ( n2322 & ~n23500 ) | ( n2322 & n32537 ) | ( ~n23500 & n32537 ) ;
  assign n34970 = ( n9714 & n11621 ) | ( n9714 & ~n13499 ) | ( n11621 & ~n13499 ) ;
  assign n34971 = n34970 ^ n14962 ^ n5965 ;
  assign n34972 = n34937 ^ n32612 ^ n19646 ;
  assign n34973 = n474 & ~n6827 ;
  assign n34974 = n34973 ^ n34420 ^ n985 ;
  assign n34975 = n18849 ^ n4844 ^ n1141 ;
  assign n34976 = n15511 ^ n15248 ^ n5997 ;
  assign n34977 = ( n1958 & n34975 ) | ( n1958 & ~n34976 ) | ( n34975 & ~n34976 ) ;
  assign n34978 = n14261 ^ n5373 ^ 1'b0 ;
  assign n34979 = n17084 | n34978 ;
  assign n34980 = n34979 ^ n30221 ^ n492 ;
  assign n34981 = ~n294 & n29432 ;
  assign n34982 = n34980 & n34981 ;
  assign n34983 = n3932 & ~n4762 ;
  assign n34984 = n11574 & ~n34023 ;
  assign n34985 = ( n10368 & n12693 ) | ( n10368 & n22855 ) | ( n12693 & n22855 ) ;
  assign n34986 = n21259 ^ n10622 ^ n3254 ;
  assign n34987 = n31042 ^ n18780 ^ n9913 ;
  assign n34988 = ( n6636 & n26999 ) | ( n6636 & n34987 ) | ( n26999 & n34987 ) ;
  assign n34989 = n21649 ^ n18163 ^ n9664 ;
  assign n34990 = ( n1008 & n1523 ) | ( n1008 & ~n28556 ) | ( n1523 & ~n28556 ) ;
  assign n34991 = ( n8585 & n13381 ) | ( n8585 & n15819 ) | ( n13381 & n15819 ) ;
  assign n34992 = n34991 ^ n14718 ^ n4192 ;
  assign n34993 = ( n30690 & n34990 ) | ( n30690 & ~n34992 ) | ( n34990 & ~n34992 ) ;
  assign n34994 = n5087 | n34993 ;
  assign n34995 = n932 & ~n34994 ;
  assign n34996 = n34995 ^ n24904 ^ n18107 ;
  assign n34997 = ( n7755 & n16712 ) | ( n7755 & n19648 ) | ( n16712 & n19648 ) ;
  assign n34998 = n31220 ^ n18765 ^ 1'b0 ;
  assign n34999 = n8038 ^ n6754 ^ n4562 ;
  assign n35000 = n8120 | n34999 ;
  assign n35001 = ( n6740 & ~n17458 ) | ( n6740 & n35000 ) | ( ~n17458 & n35000 ) ;
  assign n35002 = ( n23101 & n34998 ) | ( n23101 & n35001 ) | ( n34998 & n35001 ) ;
  assign n35003 = ( n1411 & n25739 ) | ( n1411 & n28098 ) | ( n25739 & n28098 ) ;
  assign n35004 = n35003 ^ n14954 ^ n10113 ;
  assign n35005 = n23567 ^ n14589 ^ n1580 ;
  assign n35006 = ( ~n7484 & n11508 ) | ( ~n7484 & n17884 ) | ( n11508 & n17884 ) ;
  assign n35007 = ~n13471 & n35006 ;
  assign n35008 = n35005 & n35007 ;
  assign n35009 = n12947 ^ n5815 ^ n4632 ;
  assign n35010 = ( n4167 & n18568 ) | ( n4167 & n35009 ) | ( n18568 & n35009 ) ;
  assign n35011 = ( n7429 & ~n35008 ) | ( n7429 & n35010 ) | ( ~n35008 & n35010 ) ;
  assign n35012 = ( ~n1550 & n2940 ) | ( ~n1550 & n35011 ) | ( n2940 & n35011 ) ;
  assign n35014 = ( n4599 & ~n15666 ) | ( n4599 & n18721 ) | ( ~n15666 & n18721 ) ;
  assign n35013 = n18696 & ~n19379 ;
  assign n35015 = n35014 ^ n35013 ^ 1'b0 ;
  assign n35016 = n33992 ^ n20008 ^ 1'b0 ;
  assign n35017 = n35016 ^ n14777 ^ n4401 ;
  assign n35018 = n20725 & n35017 ;
  assign n35019 = n35018 ^ n7936 ^ 1'b0 ;
  assign n35020 = n24110 ^ n18646 ^ n12420 ;
  assign n35021 = ( n2544 & n17415 ) | ( n2544 & n35020 ) | ( n17415 & n35020 ) ;
  assign n35026 = n24603 ^ n19776 ^ 1'b0 ;
  assign n35024 = n7065 ^ n854 ^ 1'b0 ;
  assign n35025 = n23336 | n35024 ;
  assign n35022 = n2428 | n18290 ;
  assign n35023 = n35022 ^ n24198 ^ n17514 ;
  assign n35027 = n35026 ^ n35025 ^ n35023 ;
  assign n35029 = ~n1779 & n10762 ;
  assign n35028 = n6690 ^ n1711 ^ n691 ;
  assign n35030 = n35029 ^ n35028 ^ n9360 ;
  assign n35031 = n35030 ^ n19172 ^ n13053 ;
  assign n35032 = ( n1075 & n11131 ) | ( n1075 & ~n24861 ) | ( n11131 & ~n24861 ) ;
  assign n35033 = n27305 ^ n5539 ^ n2182 ;
  assign n35037 = n25388 ^ n20257 ^ n14777 ;
  assign n35035 = n1564 & n6603 ;
  assign n35036 = ~n9924 & n35035 ;
  assign n35034 = n10630 ^ n10103 ^ 1'b0 ;
  assign n35038 = n35037 ^ n35036 ^ n35034 ;
  assign n35039 = ( n11375 & n35033 ) | ( n11375 & ~n35038 ) | ( n35033 & ~n35038 ) ;
  assign n35040 = n4924 | n6454 ;
  assign n35041 = n2073 | n15888 ;
  assign n35042 = n2344 & ~n35041 ;
  assign n35043 = n35042 ^ n5156 ^ n4636 ;
  assign n35044 = n2157 ^ n994 ^ 1'b0 ;
  assign n35045 = n11188 | n35044 ;
  assign n35046 = n35045 ^ n23880 ^ n14186 ;
  assign n35047 = ( n3173 & n20630 ) | ( n3173 & ~n35046 ) | ( n20630 & ~n35046 ) ;
  assign n35048 = ( ~n3380 & n4963 ) | ( ~n3380 & n31275 ) | ( n4963 & n31275 ) ;
  assign n35049 = ( n14715 & n25565 ) | ( n14715 & n35048 ) | ( n25565 & n35048 ) ;
  assign n35050 = n28820 ^ n14111 ^ n5098 ;
  assign n35051 = ( n1143 & ~n7975 ) | ( n1143 & n34331 ) | ( ~n7975 & n34331 ) ;
  assign n35052 = n35051 ^ n1355 ^ 1'b0 ;
  assign n35053 = x143 & ~n35052 ;
  assign n35055 = n10094 ^ n7651 ^ n4539 ;
  assign n35054 = n26614 | n30455 ;
  assign n35056 = n35055 ^ n35054 ^ 1'b0 ;
  assign n35057 = n4506 & ~n7717 ;
  assign n35058 = ~n8396 & n35057 ;
  assign n35059 = n35058 ^ n7738 ^ n2402 ;
  assign n35060 = n1197 | n4170 ;
  assign n35061 = n35060 ^ n972 ^ 1'b0 ;
  assign n35062 = n35061 ^ n22065 ^ n20591 ;
  assign n35063 = ~n2271 & n7483 ;
  assign n35064 = n20139 & n35063 ;
  assign n35065 = n35064 ^ n635 ^ 1'b0 ;
  assign n35066 = n35065 ^ n19337 ^ 1'b0 ;
  assign n35067 = ( n2672 & ~n6805 ) | ( n2672 & n35066 ) | ( ~n6805 & n35066 ) ;
  assign n35068 = ( n11321 & n12798 ) | ( n11321 & ~n35067 ) | ( n12798 & ~n35067 ) ;
  assign n35069 = n19799 ^ n5630 ^ 1'b0 ;
  assign n35070 = ~n973 & n35069 ;
  assign n35071 = ( n2946 & n11987 ) | ( n2946 & n35070 ) | ( n11987 & n35070 ) ;
  assign n35072 = ( n2942 & n6656 ) | ( n2942 & n26177 ) | ( n6656 & n26177 ) ;
  assign n35073 = n3721 ^ n2238 ^ n954 ;
  assign n35074 = n35073 ^ n7925 ^ n2883 ;
  assign n35075 = ( ~n10386 & n35072 ) | ( ~n10386 & n35074 ) | ( n35072 & n35074 ) ;
  assign n35076 = ( n20940 & ~n30366 ) | ( n20940 & n30574 ) | ( ~n30366 & n30574 ) ;
  assign n35077 = ( ~n7259 & n28042 ) | ( ~n7259 & n35076 ) | ( n28042 & n35076 ) ;
  assign n35078 = n35077 ^ n3840 ^ 1'b0 ;
  assign n35079 = n17743 ^ n12839 ^ 1'b0 ;
  assign n35080 = n23594 | n35079 ;
  assign n35081 = n31381 & ~n35080 ;
  assign n35082 = ( ~n1390 & n9472 ) | ( ~n1390 & n18283 ) | ( n9472 & n18283 ) ;
  assign n35083 = ( n7066 & n20477 ) | ( n7066 & ~n35082 ) | ( n20477 & ~n35082 ) ;
  assign n35084 = n2285 & n9021 ;
  assign n35085 = ( n447 & n8716 ) | ( n447 & ~n16657 ) | ( n8716 & ~n16657 ) ;
  assign n35086 = n35085 ^ n23907 ^ n4432 ;
  assign n35087 = ( n22468 & n23205 ) | ( n22468 & n32794 ) | ( n23205 & n32794 ) ;
  assign n35088 = n21050 ^ n708 ^ 1'b0 ;
  assign n35089 = n35088 ^ n21563 ^ n12261 ;
  assign n35090 = n7034 & ~n10440 ;
  assign n35091 = ~n12815 & n35090 ;
  assign n35092 = n3779 ^ n373 ^ 1'b0 ;
  assign n35093 = ~n17936 & n35092 ;
  assign n35094 = n35093 ^ n14324 ^ 1'b0 ;
  assign n35095 = n5090 & n16359 ;
  assign n35096 = n35095 ^ n14680 ^ 1'b0 ;
  assign n35097 = x89 & n27150 ;
  assign n35098 = ~n18435 & n35097 ;
  assign n35099 = n35098 ^ n19726 ^ 1'b0 ;
  assign n35100 = n32872 ^ n26442 ^ n4189 ;
  assign n35101 = ( n1869 & n11319 ) | ( n1869 & n35100 ) | ( n11319 & n35100 ) ;
  assign n35102 = x93 | n11214 ;
  assign n35103 = ( n18455 & ~n22267 ) | ( n18455 & n35102 ) | ( ~n22267 & n35102 ) ;
  assign n35104 = n28277 ^ n19593 ^ n728 ;
  assign n35106 = ~n1851 & n21084 ;
  assign n35107 = n35106 ^ n9625 ^ 1'b0 ;
  assign n35105 = ~n5367 & n32787 ;
  assign n35108 = n35107 ^ n35105 ^ n7915 ;
  assign n35111 = n19463 ^ n10079 ^ n5324 ;
  assign n35112 = ( x189 & n963 ) | ( x189 & ~n6172 ) | ( n963 & ~n6172 ) ;
  assign n35113 = ( n1242 & ~n14022 ) | ( n1242 & n31047 ) | ( ~n14022 & n31047 ) ;
  assign n35114 = ( n25616 & n35112 ) | ( n25616 & n35113 ) | ( n35112 & n35113 ) ;
  assign n35115 = ( n9936 & ~n35111 ) | ( n9936 & n35114 ) | ( ~n35111 & n35114 ) ;
  assign n35109 = n32224 ^ n14018 ^ n12005 ;
  assign n35110 = n18173 & n35109 ;
  assign n35116 = n35115 ^ n35110 ^ n25727 ;
  assign n35117 = ( n2882 & n20197 ) | ( n2882 & ~n23608 ) | ( n20197 & ~n23608 ) ;
  assign n35118 = ~n6543 & n35117 ;
  assign n35119 = ( n2424 & ~n3142 ) | ( n2424 & n5549 ) | ( ~n3142 & n5549 ) ;
  assign n35120 = ( n12190 & ~n28572 ) | ( n12190 & n35119 ) | ( ~n28572 & n35119 ) ;
  assign n35121 = ( ~n11153 & n35118 ) | ( ~n11153 & n35120 ) | ( n35118 & n35120 ) ;
  assign n35122 = n35121 ^ n25060 ^ n874 ;
  assign n35123 = n24443 ^ n17244 ^ n2192 ;
  assign n35124 = ( n3000 & n12819 ) | ( n3000 & ~n35123 ) | ( n12819 & ~n35123 ) ;
  assign n35125 = ~n9819 & n13301 ;
  assign n35126 = n28058 & n35125 ;
  assign n35127 = ~n1739 & n12594 ;
  assign n35128 = n10379 & n35127 ;
  assign n35129 = ( n3110 & n4749 ) | ( n3110 & ~n35128 ) | ( n4749 & ~n35128 ) ;
  assign n35132 = n4642 ^ n2941 ^ n1518 ;
  assign n35130 = n11864 ^ n1461 ^ 1'b0 ;
  assign n35131 = n26388 & ~n35130 ;
  assign n35133 = n35132 ^ n35131 ^ n16566 ;
  assign n35134 = n35129 & n35133 ;
  assign n35135 = ( n26604 & ~n35126 ) | ( n26604 & n35134 ) | ( ~n35126 & n35134 ) ;
  assign n35136 = ( ~n6897 & n11470 ) | ( ~n6897 & n20989 ) | ( n11470 & n20989 ) ;
  assign n35137 = n15078 ^ n11383 ^ n7401 ;
  assign n35138 = n12780 | n35137 ;
  assign n35139 = n35138 ^ n11014 ^ 1'b0 ;
  assign n35140 = ~n16193 & n35139 ;
  assign n35141 = ~n17980 & n35140 ;
  assign n35142 = n4206 & ~n6862 ;
  assign n35143 = n35142 ^ n17899 ^ n9418 ;
  assign n35144 = ( n766 & ~n5086 ) | ( n766 & n9651 ) | ( ~n5086 & n9651 ) ;
  assign n35145 = n2850 ^ n871 ^ n724 ;
  assign n35146 = ( n8820 & n35144 ) | ( n8820 & n35145 ) | ( n35144 & n35145 ) ;
  assign n35147 = n35146 ^ n24433 ^ n15583 ;
  assign n35149 = n32003 ^ n4924 ^ 1'b0 ;
  assign n35148 = ( n3232 & ~n16380 ) | ( n3232 & n30806 ) | ( ~n16380 & n30806 ) ;
  assign n35150 = n35149 ^ n35148 ^ n4178 ;
  assign n35151 = ( n2451 & n7301 ) | ( n2451 & ~n18152 ) | ( n7301 & ~n18152 ) ;
  assign n35152 = n35151 ^ n21202 ^ 1'b0 ;
  assign n35153 = n1912 | n4148 ;
  assign n35154 = n14936 | n35153 ;
  assign n35159 = n16310 ^ n3966 ^ 1'b0 ;
  assign n35155 = n14637 ^ n10877 ^ n7293 ;
  assign n35156 = ( n588 & ~n8046 ) | ( n588 & n35155 ) | ( ~n8046 & n35155 ) ;
  assign n35157 = ( ~n14645 & n19343 ) | ( ~n14645 & n35156 ) | ( n19343 & n35156 ) ;
  assign n35158 = n35157 ^ n5460 ^ n2345 ;
  assign n35160 = n35159 ^ n35158 ^ n16945 ;
  assign n35161 = n33890 ^ n27167 ^ n24510 ;
  assign n35162 = ~n4128 & n17479 ;
  assign n35163 = n22781 ^ n18046 ^ 1'b0 ;
  assign n35164 = ( n10158 & n27364 ) | ( n10158 & n28184 ) | ( n27364 & n28184 ) ;
  assign n35165 = n35164 ^ n33926 ^ n8694 ;
  assign n35166 = n35165 ^ n24777 ^ n19809 ;
  assign n35167 = ( n34375 & n35163 ) | ( n34375 & ~n35166 ) | ( n35163 & ~n35166 ) ;
  assign n35168 = n27960 ^ n14987 ^ 1'b0 ;
  assign n35169 = n31738 | n35168 ;
  assign n35170 = ( n375 & n3846 ) | ( n375 & n7722 ) | ( n3846 & n7722 ) ;
  assign n35171 = n35170 ^ n5273 ^ 1'b0 ;
  assign n35172 = ~n28498 & n35171 ;
  assign n35173 = n4147 & n9101 ;
  assign n35174 = ~n20711 & n35173 ;
  assign n35175 = n35174 ^ n26880 ^ n18857 ;
  assign n35176 = n13943 ^ n4500 ^ 1'b0 ;
  assign n35177 = n35175 & ~n35176 ;
  assign n35178 = ( n920 & ~n1844 ) | ( n920 & n4797 ) | ( ~n1844 & n4797 ) ;
  assign n35179 = n25037 ^ n19737 ^ n5600 ;
  assign n35180 = ( n30893 & n35178 ) | ( n30893 & ~n35179 ) | ( n35178 & ~n35179 ) ;
  assign n35181 = n9147 ^ n1030 ^ 1'b0 ;
  assign n35182 = n28355 ^ n7658 ^ n1731 ;
  assign n35183 = n35182 ^ n30881 ^ 1'b0 ;
  assign n35184 = n1347 & n35183 ;
  assign n35185 = ( n25422 & ~n35181 ) | ( n25422 & n35184 ) | ( ~n35181 & n35184 ) ;
  assign n35186 = ( n16130 & n35180 ) | ( n16130 & n35185 ) | ( n35180 & n35185 ) ;
  assign n35187 = n34647 ^ n34209 ^ n22471 ;
  assign n35188 = ( n4472 & ~n5153 ) | ( n4472 & n12776 ) | ( ~n5153 & n12776 ) ;
  assign n35189 = n35188 ^ n11040 ^ n3634 ;
  assign n35190 = n20239 ^ n15198 ^ n9624 ;
  assign n35191 = n26971 & ~n35190 ;
  assign n35192 = n35191 ^ n12804 ^ 1'b0 ;
  assign n35193 = n13902 & n35192 ;
  assign n35194 = n2483 ^ n1366 ^ 1'b0 ;
  assign n35195 = n10509 ^ n724 ^ 1'b0 ;
  assign n35196 = n35195 ^ n22331 ^ 1'b0 ;
  assign n35197 = ~n14048 & n35196 ;
  assign n35198 = ( n9829 & n35194 ) | ( n9829 & ~n35197 ) | ( n35194 & ~n35197 ) ;
  assign n35199 = n35198 ^ n27888 ^ 1'b0 ;
  assign n35200 = n28661 ^ n18113 ^ n8096 ;
  assign n35201 = n35200 ^ n13030 ^ n5973 ;
  assign n35202 = n35201 ^ n23906 ^ n9177 ;
  assign n35203 = n35202 ^ n25698 ^ n23431 ;
  assign n35204 = n5808 & ~n25112 ;
  assign n35205 = n33359 ^ n23290 ^ 1'b0 ;
  assign n35206 = n13249 & n35205 ;
  assign n35207 = n940 | n9801 ;
  assign n35208 = n35207 ^ n2125 ^ 1'b0 ;
  assign n35210 = n6106 ^ n2403 ^ 1'b0 ;
  assign n35211 = ~n16701 & n35210 ;
  assign n35209 = ~n6544 & n30392 ;
  assign n35212 = n35211 ^ n35209 ^ 1'b0 ;
  assign n35214 = n18831 | n25879 ;
  assign n35213 = n21939 ^ n15079 ^ n14156 ;
  assign n35215 = n35214 ^ n35213 ^ 1'b0 ;
  assign n35216 = ( n22607 & ~n23204 ) | ( n22607 & n28638 ) | ( ~n23204 & n28638 ) ;
  assign n35217 = n11613 ^ n4857 ^ 1'b0 ;
  assign n35218 = n12288 ^ n6609 ^ 1'b0 ;
  assign n35219 = ~n28982 & n35218 ;
  assign n35220 = n26820 ^ n16911 ^ n443 ;
  assign n35221 = ( ~n2816 & n23367 ) | ( ~n2816 & n34144 ) | ( n23367 & n34144 ) ;
  assign n35222 = n18598 | n32154 ;
  assign n35223 = n17874 ^ n3281 ^ 1'b0 ;
  assign n35224 = ( n12392 & n21548 ) | ( n12392 & n35223 ) | ( n21548 & n35223 ) ;
  assign n35225 = ( n961 & ~n2103 ) | ( n961 & n35224 ) | ( ~n2103 & n35224 ) ;
  assign n35226 = n5244 ^ n4447 ^ n2405 ;
  assign n35227 = ( n13584 & n14295 ) | ( n13584 & n35226 ) | ( n14295 & n35226 ) ;
  assign n35228 = ( n17178 & ~n26032 ) | ( n17178 & n35227 ) | ( ~n26032 & n35227 ) ;
  assign n35229 = ( n12653 & n29616 ) | ( n12653 & n35228 ) | ( n29616 & n35228 ) ;
  assign n35230 = n21768 ^ n6785 ^ 1'b0 ;
  assign n35231 = n10871 ^ n10141 ^ 1'b0 ;
  assign n35232 = n11553 | n35231 ;
  assign n35233 = n35232 ^ n13113 ^ 1'b0 ;
  assign n35234 = n35233 ^ n10929 ^ 1'b0 ;
  assign n35235 = n13851 & ~n35234 ;
  assign n35236 = ( ~n1183 & n35230 ) | ( ~n1183 & n35235 ) | ( n35230 & n35235 ) ;
  assign n35237 = n28434 | n35236 ;
  assign n35238 = n35237 ^ n10895 ^ 1'b0 ;
  assign n35239 = ( n34014 & ~n35229 ) | ( n34014 & n35238 ) | ( ~n35229 & n35238 ) ;
  assign n35240 = ~n4890 & n29161 ;
  assign n35241 = ~n29100 & n35240 ;
  assign n35242 = n21578 ^ n18385 ^ n1376 ;
  assign n35243 = ( n3354 & ~n4042 ) | ( n3354 & n12150 ) | ( ~n4042 & n12150 ) ;
  assign n35244 = ( n1896 & n3956 ) | ( n1896 & n14317 ) | ( n3956 & n14317 ) ;
  assign n35245 = ( n6335 & n35243 ) | ( n6335 & ~n35244 ) | ( n35243 & ~n35244 ) ;
  assign n35246 = n33908 ^ n9835 ^ 1'b0 ;
  assign n35248 = ( ~n1357 & n6540 ) | ( ~n1357 & n13320 ) | ( n6540 & n13320 ) ;
  assign n35247 = n24209 ^ n8391 ^ n2973 ;
  assign n35249 = n35248 ^ n35247 ^ n29319 ;
  assign n35250 = n28456 ^ n8732 ^ n3112 ;
  assign n35251 = ( n5918 & n24391 ) | ( n5918 & n35250 ) | ( n24391 & n35250 ) ;
  assign n35252 = n18109 & ~n32871 ;
  assign n35253 = n6613 ^ n4777 ^ 1'b0 ;
  assign n35254 = n8598 & n35253 ;
  assign n35255 = n26873 & n35254 ;
  assign n35256 = n24768 ^ n19131 ^ n9646 ;
  assign n35257 = n35256 ^ n23654 ^ n19431 ;
  assign n35258 = ( n32608 & ~n33536 ) | ( n32608 & n35257 ) | ( ~n33536 & n35257 ) ;
  assign n35259 = n17338 & n30196 ;
  assign n35260 = n33732 ^ n23586 ^ n2126 ;
  assign n35261 = n16743 ^ n2879 ^ 1'b0 ;
  assign n35262 = n35260 & n35261 ;
  assign n35263 = n35262 ^ n12516 ^ n751 ;
  assign n35264 = ( n17980 & ~n18856 ) | ( n17980 & n29875 ) | ( ~n18856 & n29875 ) ;
  assign n35265 = n25198 | n30651 ;
  assign n35266 = n6890 & ~n12541 ;
  assign n35267 = n35266 ^ n1778 ^ 1'b0 ;
  assign n35268 = n14016 ^ n4202 ^ n794 ;
  assign n35269 = n21899 & ~n29151 ;
  assign n35270 = ~n11419 & n35269 ;
  assign n35271 = ( n1474 & n21627 ) | ( n1474 & n35270 ) | ( n21627 & n35270 ) ;
  assign n35272 = n13428 & n30043 ;
  assign n35273 = n35272 ^ n25777 ^ 1'b0 ;
  assign n35274 = n35273 ^ n31820 ^ 1'b0 ;
  assign n35275 = ( n4732 & n13269 ) | ( n4732 & ~n18891 ) | ( n13269 & ~n18891 ) ;
  assign n35276 = n35275 ^ n25005 ^ n4678 ;
  assign n35277 = n13785 ^ n8087 ^ n6944 ;
  assign n35278 = n2912 ^ n566 ^ 1'b0 ;
  assign n35279 = n27589 | n35278 ;
  assign n35280 = n4205 ^ n2618 ^ n1343 ;
  assign n35281 = n33163 ^ n10705 ^ 1'b0 ;
  assign n35282 = n19453 | n20557 ;
  assign n35283 = n35282 ^ n29493 ^ 1'b0 ;
  assign n35284 = ( n1580 & n12570 ) | ( n1580 & n35283 ) | ( n12570 & n35283 ) ;
  assign n35285 = ( n8830 & n21176 ) | ( n8830 & n30372 ) | ( n21176 & n30372 ) ;
  assign n35286 = ( x20 & n3314 ) | ( x20 & ~n12751 ) | ( n3314 & ~n12751 ) ;
  assign n35287 = ( n4051 & n29985 ) | ( n4051 & ~n35286 ) | ( n29985 & ~n35286 ) ;
  assign n35288 = ( n3828 & ~n11607 ) | ( n3828 & n35287 ) | ( ~n11607 & n35287 ) ;
  assign n35289 = n14596 ^ n3500 ^ 1'b0 ;
  assign n35290 = n30180 & n35289 ;
  assign n35291 = ( n4384 & n7023 ) | ( n4384 & n12372 ) | ( n7023 & n12372 ) ;
  assign n35292 = n35291 ^ n9347 ^ 1'b0 ;
  assign n35293 = n28715 ^ n28125 ^ 1'b0 ;
  assign n35294 = n33142 & n35293 ;
  assign n35295 = ( n9801 & n35292 ) | ( n9801 & n35294 ) | ( n35292 & n35294 ) ;
  assign n35296 = n9459 | n19633 ;
  assign n35297 = n35296 ^ n6632 ^ 1'b0 ;
  assign n35298 = n33464 ^ n17290 ^ 1'b0 ;
  assign n35299 = n28771 ^ n1269 ^ 1'b0 ;
  assign n35300 = n22350 ^ n22033 ^ n6346 ;
  assign n35301 = n35300 ^ n32619 ^ 1'b0 ;
  assign n35302 = ( n34824 & n35299 ) | ( n34824 & ~n35301 ) | ( n35299 & ~n35301 ) ;
  assign n35303 = ~n766 & n13970 ;
  assign n35304 = ~n6429 & n35303 ;
  assign n35305 = ~n2062 & n5638 ;
  assign n35306 = n35305 ^ n604 ^ 1'b0 ;
  assign n35307 = n21028 ^ n8436 ^ 1'b0 ;
  assign n35308 = n31659 & n35307 ;
  assign n35309 = ( n15275 & n30346 ) | ( n15275 & n35308 ) | ( n30346 & n35308 ) ;
  assign n35310 = ( ~n4100 & n30020 ) | ( ~n4100 & n33624 ) | ( n30020 & n33624 ) ;
  assign n35311 = n18823 | n35310 ;
  assign n35312 = n27670 | n35311 ;
  assign n35313 = ( n7171 & n32636 ) | ( n7171 & n35312 ) | ( n32636 & n35312 ) ;
  assign n35314 = ( n5668 & n15947 ) | ( n5668 & n35131 ) | ( n15947 & n35131 ) ;
  assign n35315 = n15871 & ~n35314 ;
  assign n35316 = ( n14704 & ~n16069 ) | ( n14704 & n21176 ) | ( ~n16069 & n21176 ) ;
  assign n35317 = n12836 ^ n7529 ^ 1'b0 ;
  assign n35318 = ~n4697 & n35317 ;
  assign n35319 = ( n33067 & n35316 ) | ( n33067 & ~n35318 ) | ( n35316 & ~n35318 ) ;
  assign n35320 = ( n4341 & ~n9591 ) | ( n4341 & n16461 ) | ( ~n9591 & n16461 ) ;
  assign n35321 = ( n18114 & n28594 ) | ( n18114 & n35320 ) | ( n28594 & n35320 ) ;
  assign n35322 = n11758 & n35321 ;
  assign n35323 = ~n2957 & n35322 ;
  assign n35324 = n26432 ^ n19488 ^ n14827 ;
  assign n35325 = n21195 ^ n10419 ^ x58 ;
  assign n35326 = n18662 ^ n11709 ^ n10496 ;
  assign n35329 = n27118 ^ n15807 ^ n2127 ;
  assign n35328 = n31281 ^ n18873 ^ n2860 ;
  assign n35327 = n12259 & n13271 ;
  assign n35330 = n35329 ^ n35328 ^ n35327 ;
  assign n35331 = n35330 ^ n29514 ^ n412 ;
  assign n35332 = n34021 ^ n12738 ^ x184 ;
  assign n35333 = n35332 ^ n7496 ^ 1'b0 ;
  assign n35334 = n35333 ^ n22153 ^ n11701 ;
  assign n35335 = n25911 & n35334 ;
  assign n35336 = n2111 & n35335 ;
  assign n35337 = n9900 ^ n1592 ^ 1'b0 ;
  assign n35338 = n12641 & n35337 ;
  assign n35339 = ( n3917 & n33420 ) | ( n3917 & ~n35338 ) | ( n33420 & ~n35338 ) ;
  assign n35340 = n21123 ^ n14513 ^ n13295 ;
  assign n35341 = ( n916 & n14307 ) | ( n916 & n29772 ) | ( n14307 & n29772 ) ;
  assign n35342 = n35341 ^ n21147 ^ 1'b0 ;
  assign n35343 = n35342 ^ n17290 ^ n12102 ;
  assign n35344 = ( n2804 & ~n17627 ) | ( n2804 & n26275 ) | ( ~n17627 & n26275 ) ;
  assign n35345 = ~n27751 & n33630 ;
  assign n35346 = n35345 ^ n5091 ^ 1'b0 ;
  assign n35347 = n13769 & n21728 ;
  assign n35348 = n35347 ^ n5893 ^ 1'b0 ;
  assign n35350 = n30005 ^ n12353 ^ n11698 ;
  assign n35349 = n12251 & n26775 ;
  assign n35351 = n35350 ^ n35349 ^ 1'b0 ;
  assign n35352 = n25827 ^ n1196 ^ n391 ;
  assign n35353 = n1654 & n35352 ;
  assign n35354 = n6879 & ~n35353 ;
  assign n35355 = n10169 & n35354 ;
  assign n35356 = n19083 | n32358 ;
  assign n35357 = ( ~n26824 & n35355 ) | ( ~n26824 & n35356 ) | ( n35355 & n35356 ) ;
  assign n35359 = ( n3651 & n4795 ) | ( n3651 & ~n9320 ) | ( n4795 & ~n9320 ) ;
  assign n35358 = ( n14803 & ~n16339 ) | ( n14803 & n19895 ) | ( ~n16339 & n19895 ) ;
  assign n35360 = n35359 ^ n35358 ^ n33082 ;
  assign n35362 = n27516 ^ n11226 ^ n10800 ;
  assign n35361 = ( n4021 & ~n26275 ) | ( n4021 & n28961 ) | ( ~n26275 & n28961 ) ;
  assign n35363 = n35362 ^ n35361 ^ 1'b0 ;
  assign n35364 = ( n2097 & ~n2206 ) | ( n2097 & n5681 ) | ( ~n2206 & n5681 ) ;
  assign n35365 = ( n5243 & n15723 ) | ( n5243 & n19566 ) | ( n15723 & n19566 ) ;
  assign n35366 = ( n3823 & ~n31020 ) | ( n3823 & n35365 ) | ( ~n31020 & n35365 ) ;
  assign n35367 = n17012 ^ n9571 ^ 1'b0 ;
  assign n35368 = ( n13912 & ~n14992 ) | ( n13912 & n16717 ) | ( ~n14992 & n16717 ) ;
  assign n35369 = ( ~n956 & n3358 ) | ( ~n956 & n18724 ) | ( n3358 & n18724 ) ;
  assign n35370 = ( n11617 & n24838 ) | ( n11617 & ~n29683 ) | ( n24838 & ~n29683 ) ;
  assign n35371 = n35370 ^ n17674 ^ 1'b0 ;
  assign n35372 = n35369 & ~n35371 ;
  assign n35373 = n35372 ^ n18789 ^ n8914 ;
  assign n35374 = ( ~n14057 & n35368 ) | ( ~n14057 & n35373 ) | ( n35368 & n35373 ) ;
  assign n35375 = n27606 ^ n14407 ^ n4248 ;
  assign n35376 = n35375 ^ n20602 ^ n7915 ;
  assign n35377 = n35376 ^ n20117 ^ n15706 ;
  assign n35378 = n26339 ^ n9081 ^ 1'b0 ;
  assign n35379 = n22945 & ~n35378 ;
  assign n35380 = n35379 ^ n29668 ^ n20321 ;
  assign n35381 = ( n1064 & ~n10630 ) | ( n1064 & n22137 ) | ( ~n10630 & n22137 ) ;
  assign n35382 = n35381 ^ n2759 ^ 1'b0 ;
  assign n35383 = ( n9759 & ~n35380 ) | ( n9759 & n35382 ) | ( ~n35380 & n35382 ) ;
  assign n35384 = ~n6755 & n7515 ;
  assign n35385 = n7444 & n35384 ;
  assign n35386 = ( n9328 & n20448 ) | ( n9328 & n22664 ) | ( n20448 & n22664 ) ;
  assign n35387 = ( n1493 & n3181 ) | ( n1493 & ~n26315 ) | ( n3181 & ~n26315 ) ;
  assign n35388 = ( n3950 & ~n10599 ) | ( n3950 & n11229 ) | ( ~n10599 & n11229 ) ;
  assign n35389 = n35387 & n35388 ;
  assign n35390 = ~n35386 & n35389 ;
  assign n35391 = n35390 ^ n4633 ^ 1'b0 ;
  assign n35392 = ~n20683 & n35391 ;
  assign n35393 = ( n17437 & n35385 ) | ( n17437 & ~n35392 ) | ( n35385 & ~n35392 ) ;
  assign n35394 = ( n1041 & ~n33940 ) | ( n1041 & n35393 ) | ( ~n33940 & n35393 ) ;
  assign n35395 = n19438 ^ n9295 ^ n1782 ;
  assign n35396 = ( n6776 & n16603 ) | ( n6776 & n35395 ) | ( n16603 & n35395 ) ;
  assign n35397 = ( n18730 & n19280 ) | ( n18730 & ~n23110 ) | ( n19280 & ~n23110 ) ;
  assign n35398 = n35397 ^ n19544 ^ n1407 ;
  assign n35399 = n17122 | n35398 ;
  assign n35400 = n35399 ^ n14254 ^ 1'b0 ;
  assign n35401 = ( n13284 & ~n16445 ) | ( n13284 & n29817 ) | ( ~n16445 & n29817 ) ;
  assign n35402 = ( n3728 & ~n12826 ) | ( n3728 & n19906 ) | ( ~n12826 & n19906 ) ;
  assign n35403 = ~n15878 & n24887 ;
  assign n35404 = n28009 ^ n14949 ^ n13965 ;
  assign n35405 = ( ~n14305 & n20469 ) | ( ~n14305 & n23230 ) | ( n20469 & n23230 ) ;
  assign n35406 = ~n35404 & n35405 ;
  assign n35407 = ( n5842 & n12803 ) | ( n5842 & ~n20002 ) | ( n12803 & ~n20002 ) ;
  assign n35408 = ( n1212 & n1371 ) | ( n1212 & n35407 ) | ( n1371 & n35407 ) ;
  assign n35409 = n20537 ^ n8663 ^ 1'b0 ;
  assign n35410 = n35408 & n35409 ;
  assign n35412 = n16037 ^ n6122 ^ 1'b0 ;
  assign n35413 = ~n13469 & n35412 ;
  assign n35411 = ~n6365 & n26949 ;
  assign n35414 = n35413 ^ n35411 ^ 1'b0 ;
  assign n35415 = n6570 & ~n18389 ;
  assign n35416 = ~n13520 & n35415 ;
  assign n35417 = ~n12640 & n20747 ;
  assign n35418 = ~n22955 & n35417 ;
  assign n35419 = ( n16214 & n29377 ) | ( n16214 & ~n35418 ) | ( n29377 & ~n35418 ) ;
  assign n35420 = ( n4977 & n35416 ) | ( n4977 & ~n35419 ) | ( n35416 & ~n35419 ) ;
  assign n35421 = n4272 & ~n35420 ;
  assign n35422 = ~n23450 & n35421 ;
  assign n35423 = n17853 ^ n4973 ^ 1'b0 ;
  assign n35424 = n28659 ^ n10709 ^ n2473 ;
  assign n35425 = ~n9294 & n35424 ;
  assign n35426 = ( n1083 & ~n17681 ) | ( n1083 & n25734 ) | ( ~n17681 & n25734 ) ;
  assign n35427 = ~n11755 & n35426 ;
  assign n35428 = n35427 ^ n20101 ^ 1'b0 ;
  assign n35429 = n35428 ^ n22438 ^ n12869 ;
  assign n35430 = n17706 ^ n9553 ^ n3808 ;
  assign n35431 = n35430 ^ n26326 ^ n5094 ;
  assign n35432 = n24619 ^ n8033 ^ 1'b0 ;
  assign n35433 = n35432 ^ n22564 ^ n20758 ;
  assign n35434 = n4452 & ~n6890 ;
  assign n35439 = ( n4947 & ~n8795 ) | ( n4947 & n17361 ) | ( ~n8795 & n17361 ) ;
  assign n35438 = ( ~n2484 & n4079 ) | ( ~n2484 & n13301 ) | ( n4079 & n13301 ) ;
  assign n35435 = n12184 & n32839 ;
  assign n35436 = n35435 ^ n18943 ^ 1'b0 ;
  assign n35437 = ( n2023 & n25574 ) | ( n2023 & ~n35436 ) | ( n25574 & ~n35436 ) ;
  assign n35440 = n35439 ^ n35438 ^ n35437 ;
  assign n35441 = ( n9852 & n13783 ) | ( n9852 & ~n14052 ) | ( n13783 & ~n14052 ) ;
  assign n35442 = ( n4865 & n15393 ) | ( n4865 & n23459 ) | ( n15393 & n23459 ) ;
  assign n35443 = ( ~n424 & n8367 ) | ( ~n424 & n21282 ) | ( n8367 & n21282 ) ;
  assign n35444 = n35227 ^ n12919 ^ n304 ;
  assign n35445 = ( n16053 & n32563 ) | ( n16053 & ~n35444 ) | ( n32563 & ~n35444 ) ;
  assign n35446 = ~n4424 & n8832 ;
  assign n35447 = ( n6666 & n25782 ) | ( n6666 & n32884 ) | ( n25782 & n32884 ) ;
  assign n35448 = ~n13956 & n30634 ;
  assign n35449 = ~n26124 & n35448 ;
  assign n35460 = ~n8082 & n9029 ;
  assign n35461 = n35460 ^ n2022 ^ 1'b0 ;
  assign n35450 = n12250 ^ n9900 ^ n3387 ;
  assign n35451 = ( n525 & ~n8428 ) | ( n525 & n27752 ) | ( ~n8428 & n27752 ) ;
  assign n35452 = n35451 ^ n13107 ^ n3668 ;
  assign n35453 = ( n4795 & n8722 ) | ( n4795 & n10984 ) | ( n8722 & n10984 ) ;
  assign n35454 = ( n17740 & ~n34021 ) | ( n17740 & n35453 ) | ( ~n34021 & n35453 ) ;
  assign n35455 = n35452 & n35454 ;
  assign n35456 = ~x152 & n35455 ;
  assign n35457 = n2148 ^ n1441 ^ 1'b0 ;
  assign n35458 = n35456 & n35457 ;
  assign n35459 = n35450 & n35458 ;
  assign n35462 = n35461 ^ n35459 ^ 1'b0 ;
  assign n35463 = n12532 & ~n35462 ;
  assign n35465 = ( ~n7324 & n11150 ) | ( ~n7324 & n28150 ) | ( n11150 & n28150 ) ;
  assign n35464 = ( n9055 & n15255 ) | ( n9055 & ~n19214 ) | ( n15255 & ~n19214 ) ;
  assign n35466 = n35465 ^ n35464 ^ n7672 ;
  assign n35467 = n16198 ^ n11926 ^ n10789 ;
  assign n35468 = ( n1242 & ~n22581 ) | ( n1242 & n34454 ) | ( ~n22581 & n34454 ) ;
  assign n35469 = ( n868 & ~n15941 ) | ( n868 & n24836 ) | ( ~n15941 & n24836 ) ;
  assign n35470 = n26226 ^ n17675 ^ n2248 ;
  assign n35471 = n35470 ^ n3018 ^ 1'b0 ;
  assign n35472 = n9914 | n19162 ;
  assign n35474 = ( ~x89 & n6714 ) | ( ~x89 & n30432 ) | ( n6714 & n30432 ) ;
  assign n35475 = n3932 & ~n35474 ;
  assign n35476 = n35475 ^ n29900 ^ 1'b0 ;
  assign n35473 = ~n867 & n1060 ;
  assign n35477 = n35476 ^ n35473 ^ 1'b0 ;
  assign n35478 = n24018 ^ n16573 ^ n849 ;
  assign n35479 = n15117 ^ n8569 ^ 1'b0 ;
  assign n35480 = n21433 ^ n18924 ^ n6477 ;
  assign n35481 = ( n5901 & ~n7538 ) | ( n5901 & n16084 ) | ( ~n7538 & n16084 ) ;
  assign n35482 = ( n9491 & n12508 ) | ( n9491 & n19408 ) | ( n12508 & n19408 ) ;
  assign n35483 = ( n22957 & ~n35481 ) | ( n22957 & n35482 ) | ( ~n35481 & n35482 ) ;
  assign n35484 = n26826 ^ n4589 ^ n2653 ;
  assign n35485 = ( ~n15070 & n27744 ) | ( ~n15070 & n35484 ) | ( n27744 & n35484 ) ;
  assign n35486 = n22285 ^ n16406 ^ 1'b0 ;
  assign n35487 = ~n35485 & n35486 ;
  assign n35488 = n20741 ^ n9591 ^ n8382 ;
  assign n35489 = n27417 ^ n9708 ^ 1'b0 ;
  assign n35490 = n3010 & n8376 ;
  assign n35491 = n35490 ^ n29605 ^ n4609 ;
  assign n35492 = n7510 | n27875 ;
  assign n35493 = n20422 & ~n35492 ;
  assign n35494 = ~n15413 & n35493 ;
  assign n35495 = n12653 ^ n9191 ^ n3879 ;
  assign n35496 = ( n18847 & n19081 ) | ( n18847 & ~n35495 ) | ( n19081 & ~n35495 ) ;
  assign n35497 = n6331 & ~n35496 ;
  assign n35498 = n35497 ^ n34031 ^ 1'b0 ;
  assign n35499 = ( n4321 & ~n35494 ) | ( n4321 & n35498 ) | ( ~n35494 & n35498 ) ;
  assign n35500 = n35107 ^ n22024 ^ n14743 ;
  assign n35501 = n471 | n11832 ;
  assign n35502 = ( n9290 & ~n9343 ) | ( n9290 & n23218 ) | ( ~n9343 & n23218 ) ;
  assign n35503 = n35502 ^ n16326 ^ n5460 ;
  assign n35504 = n35503 ^ n17451 ^ n16588 ;
  assign n35505 = n35504 ^ n2858 ^ 1'b0 ;
  assign n35506 = n35501 | n35505 ;
  assign n35507 = n10469 | n21868 ;
  assign n35508 = ( n1349 & ~n7259 ) | ( n1349 & n8440 ) | ( ~n7259 & n8440 ) ;
  assign n35509 = n35507 & ~n35508 ;
  assign n35510 = n27350 ^ n15061 ^ n3521 ;
  assign n35511 = n31574 ^ n11766 ^ n9121 ;
  assign n35512 = n35511 ^ n34591 ^ n5403 ;
  assign n35513 = ~n1897 & n5779 ;
  assign n35514 = n35513 ^ n31253 ^ 1'b0 ;
  assign n35515 = n8596 ^ n7158 ^ 1'b0 ;
  assign n35516 = ( ~n7973 & n8629 ) | ( ~n7973 & n15290 ) | ( n8629 & n15290 ) ;
  assign n35517 = n33925 ^ n5286 ^ 1'b0 ;
  assign n35518 = ~n32965 & n35517 ;
  assign n35519 = ( n14373 & n35516 ) | ( n14373 & n35518 ) | ( n35516 & n35518 ) ;
  assign n35520 = n3332 ^ n3265 ^ 1'b0 ;
  assign n35521 = n35519 | n35520 ;
  assign n35522 = ( x220 & n2474 ) | ( x220 & ~n13481 ) | ( n2474 & ~n13481 ) ;
  assign n35523 = n8243 ^ n3921 ^ n3188 ;
  assign n35524 = n24286 ^ n15948 ^ n14000 ;
  assign n35525 = ( n19634 & n35523 ) | ( n19634 & n35524 ) | ( n35523 & n35524 ) ;
  assign n35526 = n23979 ^ n18760 ^ x28 ;
  assign n35527 = ( n8155 & n9811 ) | ( n8155 & ~n30868 ) | ( n9811 & ~n30868 ) ;
  assign n35528 = n35527 ^ n16830 ^ n656 ;
  assign n35529 = n26032 ^ n10039 ^ 1'b0 ;
  assign n35530 = ( ~n13088 & n14470 ) | ( ~n13088 & n26035 ) | ( n14470 & n26035 ) ;
  assign n35531 = n27436 ^ n9192 ^ n3157 ;
  assign n35532 = ( ~n2941 & n7178 ) | ( ~n2941 & n35531 ) | ( n7178 & n35531 ) ;
  assign n35533 = n35532 ^ n14558 ^ 1'b0 ;
  assign n35534 = ~n35530 & n35533 ;
  assign n35535 = n11870 | n35534 ;
  assign n35536 = n35529 | n35535 ;
  assign n35537 = ( n904 & n22538 ) | ( n904 & ~n25225 ) | ( n22538 & ~n25225 ) ;
  assign n35538 = n29536 & ~n35537 ;
  assign n35539 = n29997 & n35538 ;
  assign n35540 = ( n2324 & n5676 ) | ( n2324 & n6226 ) | ( n5676 & n6226 ) ;
  assign n35541 = ( n5848 & ~n14980 ) | ( n5848 & n35540 ) | ( ~n14980 & n35540 ) ;
  assign n35542 = n29532 ^ n22517 ^ 1'b0 ;
  assign n35543 = ( ~n8258 & n11115 ) | ( ~n8258 & n12166 ) | ( n11115 & n12166 ) ;
  assign n35544 = n24150 ^ n21804 ^ 1'b0 ;
  assign n35545 = ( ~n2550 & n35543 ) | ( ~n2550 & n35544 ) | ( n35543 & n35544 ) ;
  assign n35546 = ( n7463 & n15396 ) | ( n7463 & ~n15677 ) | ( n15396 & ~n15677 ) ;
  assign n35547 = ( n23420 & n33415 ) | ( n23420 & n35546 ) | ( n33415 & n35546 ) ;
  assign n35548 = n1703 & ~n6718 ;
  assign n35549 = n33272 ^ n11144 ^ n5875 ;
  assign n35550 = ( n1744 & ~n26633 ) | ( n1744 & n35549 ) | ( ~n26633 & n35549 ) ;
  assign n35551 = n29962 ^ n15362 ^ n6337 ;
  assign n35552 = n35551 ^ n34397 ^ n23770 ;
  assign n35553 = ( n10282 & ~n27824 ) | ( n10282 & n28489 ) | ( ~n27824 & n28489 ) ;
  assign n35554 = ( n3755 & n29398 ) | ( n3755 & n34377 ) | ( n29398 & n34377 ) ;
  assign n35555 = ( n4286 & n14466 ) | ( n4286 & n16300 ) | ( n14466 & n16300 ) ;
  assign n35556 = n27585 ^ n18384 ^ n16185 ;
  assign n35557 = ( n22572 & ~n35555 ) | ( n22572 & n35556 ) | ( ~n35555 & n35556 ) ;
  assign n35558 = n20983 ^ n11012 ^ 1'b0 ;
  assign n35559 = n9636 | n12324 ;
  assign n35560 = ( n11662 & ~n19311 ) | ( n11662 & n35559 ) | ( ~n19311 & n35559 ) ;
  assign n35561 = n16073 ^ n13290 ^ n10086 ;
  assign n35562 = n32010 ^ n29889 ^ n7150 ;
  assign n35563 = n24491 ^ n4552 ^ 1'b0 ;
  assign n35564 = n35562 & ~n35563 ;
  assign n35565 = n3516 ^ n3111 ^ 1'b0 ;
  assign n35566 = n3115 | n35565 ;
  assign n35567 = ( ~n4145 & n10731 ) | ( ~n4145 & n35566 ) | ( n10731 & n35566 ) ;
  assign n35568 = n35567 ^ n4484 ^ n3279 ;
  assign n35569 = n14707 & ~n21177 ;
  assign n35570 = ~n28983 & n35569 ;
  assign n35571 = n19914 & n35570 ;
  assign n35572 = n35571 ^ n18271 ^ n2505 ;
  assign n35573 = ( n30631 & ~n35568 ) | ( n30631 & n35572 ) | ( ~n35568 & n35572 ) ;
  assign n35574 = n19011 ^ n16925 ^ 1'b0 ;
  assign n35575 = ( ~n3035 & n4704 ) | ( ~n3035 & n35574 ) | ( n4704 & n35574 ) ;
  assign n35576 = ( n6775 & n9469 ) | ( n6775 & ~n35575 ) | ( n9469 & ~n35575 ) ;
  assign n35577 = n33593 ^ n1218 ^ 1'b0 ;
  assign n35578 = n19220 ^ n5943 ^ n4760 ;
  assign n35579 = ( n32820 & n35577 ) | ( n32820 & n35578 ) | ( n35577 & n35578 ) ;
  assign n35580 = n22293 ^ n4042 ^ n471 ;
  assign n35581 = ( n8646 & n14822 ) | ( n8646 & ~n20236 ) | ( n14822 & ~n20236 ) ;
  assign n35582 = ( x54 & n1367 ) | ( x54 & n2647 ) | ( n1367 & n2647 ) ;
  assign n35583 = n35582 ^ n27347 ^ n20533 ;
  assign n35584 = ( ~n1040 & n21764 ) | ( ~n1040 & n35583 ) | ( n21764 & n35583 ) ;
  assign n35585 = n12669 ^ n4843 ^ n2156 ;
  assign n35586 = n35585 ^ n23551 ^ n11615 ;
  assign n35587 = ( ~n6740 & n7253 ) | ( ~n6740 & n26460 ) | ( n7253 & n26460 ) ;
  assign n35589 = ( ~n21158 & n23545 ) | ( ~n21158 & n28744 ) | ( n23545 & n28744 ) ;
  assign n35588 = n18160 ^ n17951 ^ n1733 ;
  assign n35590 = n35589 ^ n35588 ^ n3301 ;
  assign n35591 = ( n10920 & n35587 ) | ( n10920 & ~n35590 ) | ( n35587 & ~n35590 ) ;
  assign n35592 = ( n7463 & n7540 ) | ( n7463 & n15635 ) | ( n7540 & n15635 ) ;
  assign n35593 = n35592 ^ n7166 ^ n1071 ;
  assign n35594 = ( n7473 & n23489 ) | ( n7473 & n35593 ) | ( n23489 & n35593 ) ;
  assign n35595 = n35594 ^ n13173 ^ n3358 ;
  assign n35596 = n11273 ^ n8949 ^ n3143 ;
  assign n35597 = n35596 ^ n31340 ^ n13173 ;
  assign n35598 = n16455 | n22522 ;
  assign n35599 = n35598 ^ n15259 ^ 1'b0 ;
  assign n35600 = n11094 & ~n19383 ;
  assign n35601 = n35600 ^ n32787 ^ 1'b0 ;
  assign n35602 = ( n15135 & n18896 ) | ( n15135 & n35601 ) | ( n18896 & n35601 ) ;
  assign n35603 = ( n16015 & n35599 ) | ( n16015 & n35602 ) | ( n35599 & n35602 ) ;
  assign n35604 = n11698 | n14772 ;
  assign n35605 = n3006 | n35604 ;
  assign n35606 = n35605 ^ n12644 ^ n812 ;
  assign n35607 = ( n35597 & n35603 ) | ( n35597 & ~n35606 ) | ( n35603 & ~n35606 ) ;
  assign n35608 = n5267 & n7030 ;
  assign n35609 = n1364 & n35608 ;
  assign n35610 = n29410 ^ n13361 ^ 1'b0 ;
  assign n35611 = n20032 & ~n35610 ;
  assign n35612 = ( ~n3241 & n15559 ) | ( ~n3241 & n32604 ) | ( n15559 & n32604 ) ;
  assign n35613 = n18391 ^ n14496 ^ n3094 ;
  assign n35614 = ( ~n4362 & n9076 ) | ( ~n4362 & n35613 ) | ( n9076 & n35613 ) ;
  assign n35615 = n35614 ^ n33444 ^ n7490 ;
  assign n35616 = ( ~n14130 & n34413 ) | ( ~n14130 & n35615 ) | ( n34413 & n35615 ) ;
  assign n35617 = n35083 ^ n31688 ^ n27157 ;
  assign n35619 = n6109 ^ n2734 ^ 1'b0 ;
  assign n35620 = n17041 | n35619 ;
  assign n35618 = ~n12350 & n21117 ;
  assign n35621 = n35620 ^ n35618 ^ n17664 ;
  assign n35622 = n15960 ^ n5151 ^ 1'b0 ;
  assign n35623 = n2524 | n35622 ;
  assign n35624 = ( n7949 & n21932 ) | ( n7949 & ~n29446 ) | ( n21932 & ~n29446 ) ;
  assign n35626 = ( ~n1800 & n5479 ) | ( ~n1800 & n26794 ) | ( n5479 & n26794 ) ;
  assign n35625 = ( n749 & n9447 ) | ( n749 & ~n26784 ) | ( n9447 & ~n26784 ) ;
  assign n35627 = n35626 ^ n35625 ^ n35165 ;
  assign n35628 = ( ~n2954 & n5918 ) | ( ~n2954 & n15414 ) | ( n5918 & n15414 ) ;
  assign n35629 = n35628 ^ n2582 ^ 1'b0 ;
  assign n35630 = ~n1367 & n35629 ;
  assign n35631 = ( n3241 & ~n4517 ) | ( n3241 & n35630 ) | ( ~n4517 & n35630 ) ;
  assign n35633 = n19724 ^ n11449 ^ n5645 ;
  assign n35634 = n35633 ^ n6114 ^ n315 ;
  assign n35632 = n7435 | n14127 ;
  assign n35635 = n35634 ^ n35632 ^ 1'b0 ;
  assign n35636 = ( n1276 & n29408 ) | ( n1276 & n35635 ) | ( n29408 & n35635 ) ;
  assign n35637 = n17087 ^ n11477 ^ 1'b0 ;
  assign n35638 = n15952 | n35637 ;
  assign n35639 = n35638 ^ n17077 ^ x229 ;
  assign n35643 = n17835 & ~n26094 ;
  assign n35644 = n35643 ^ n22979 ^ n2590 ;
  assign n35640 = n27634 ^ n21377 ^ n3277 ;
  assign n35641 = n11063 & ~n35640 ;
  assign n35642 = n18261 & n35641 ;
  assign n35645 = n35644 ^ n35642 ^ n10895 ;
  assign n35646 = n28703 ^ n19259 ^ x253 ;
  assign n35647 = ( n6589 & ~n28140 ) | ( n6589 & n29786 ) | ( ~n28140 & n29786 ) ;
  assign n35649 = ( ~n7277 & n10359 ) | ( ~n7277 & n33303 ) | ( n10359 & n33303 ) ;
  assign n35650 = n35649 ^ n13285 ^ 1'b0 ;
  assign n35651 = n14736 & n35650 ;
  assign n35648 = ( n2365 & ~n10449 ) | ( n2365 & n18922 ) | ( ~n10449 & n18922 ) ;
  assign n35652 = n35651 ^ n35648 ^ n16201 ;
  assign n35653 = n25183 ^ n1938 ^ 1'b0 ;
  assign n35654 = n10649 | n35653 ;
  assign n35655 = n35654 ^ n9503 ^ 1'b0 ;
  assign n35656 = n23595 | n35655 ;
  assign n35657 = n8329 ^ n8101 ^ 1'b0 ;
  assign n35658 = ( n10658 & ~n18859 ) | ( n10658 & n35657 ) | ( ~n18859 & n35657 ) ;
  assign n35659 = ( n23331 & n35656 ) | ( n23331 & ~n35658 ) | ( n35656 & ~n35658 ) ;
  assign n35660 = n1676 | n4842 ;
  assign n35661 = n35660 ^ n32630 ^ 1'b0 ;
  assign n35662 = n8850 ^ n5591 ^ 1'b0 ;
  assign n35663 = ( ~n9330 & n25393 ) | ( ~n9330 & n32954 ) | ( n25393 & n32954 ) ;
  assign n35664 = n35663 ^ n7699 ^ 1'b0 ;
  assign n35665 = n33918 ^ n25327 ^ 1'b0 ;
  assign n35666 = n14794 & ~n35665 ;
  assign n35667 = ( ~n7344 & n8573 ) | ( ~n7344 & n35666 ) | ( n8573 & n35666 ) ;
  assign n35668 = n6891 | n9429 ;
  assign n35669 = n35668 ^ n29313 ^ n28509 ;
  assign n35670 = n2487 & ~n4009 ;
  assign n35671 = ~n1028 & n35670 ;
  assign n35672 = n30757 ^ n3031 ^ x151 ;
  assign n35673 = ~n2869 & n35672 ;
  assign n35674 = n8825 & n34909 ;
  assign n35675 = n20577 ^ n10147 ^ 1'b0 ;
  assign n35676 = n6489 & n35675 ;
  assign n35677 = n35676 ^ n15759 ^ n7994 ;
  assign n35678 = ( n6524 & n29616 ) | ( n6524 & n30728 ) | ( n29616 & n30728 ) ;
  assign n35679 = n35677 & ~n35678 ;
  assign n35680 = ( n7496 & n8218 ) | ( n7496 & ~n8643 ) | ( n8218 & ~n8643 ) ;
  assign n35681 = n35680 ^ n8600 ^ 1'b0 ;
  assign n35682 = ( n10417 & n12480 ) | ( n10417 & n35681 ) | ( n12480 & n35681 ) ;
  assign n35683 = ( n8356 & n34990 ) | ( n8356 & ~n35531 ) | ( n34990 & ~n35531 ) ;
  assign n35684 = n35683 ^ n29324 ^ 1'b0 ;
  assign n35685 = n34088 & ~n35684 ;
  assign n35688 = n1207 ^ n706 ^ 1'b0 ;
  assign n35686 = n9766 ^ n7432 ^ x28 ;
  assign n35687 = n35686 ^ n19332 ^ n18111 ;
  assign n35689 = n35688 ^ n35687 ^ 1'b0 ;
  assign n35690 = n20299 & n35689 ;
  assign n35691 = n24650 ^ n2385 ^ 1'b0 ;
  assign n35692 = n28443 | n35691 ;
  assign n35693 = ~n14313 & n15903 ;
  assign n35694 = n16764 & n35693 ;
  assign n35695 = n13175 ^ n9637 ^ n4180 ;
  assign n35696 = n6288 | n35695 ;
  assign n35697 = n35694 & ~n35696 ;
  assign n35698 = n35697 ^ n12109 ^ n1882 ;
  assign n35699 = ( n11140 & n26192 ) | ( n11140 & ~n35112 ) | ( n26192 & ~n35112 ) ;
  assign n35701 = n26210 ^ n9624 ^ n5331 ;
  assign n35700 = n8175 & n15614 ;
  assign n35702 = n35701 ^ n35700 ^ 1'b0 ;
  assign n35703 = ( n12670 & n32266 ) | ( n12670 & ~n35702 ) | ( n32266 & ~n35702 ) ;
  assign n35705 = n11310 ^ n2088 ^ 1'b0 ;
  assign n35704 = ( ~n3139 & n23283 ) | ( ~n3139 & n30931 ) | ( n23283 & n30931 ) ;
  assign n35706 = n35705 ^ n35704 ^ n27057 ;
  assign n35707 = ( n1558 & n19400 ) | ( n1558 & ~n35706 ) | ( n19400 & ~n35706 ) ;
  assign n35708 = n5629 ^ n4716 ^ 1'b0 ;
  assign n35709 = n6460 | n21124 ;
  assign n35710 = n25944 & ~n35709 ;
  assign n35711 = n35708 & ~n35710 ;
  assign n35712 = n35711 ^ n12718 ^ 1'b0 ;
  assign n35713 = n32775 | n35712 ;
  assign n35714 = n4094 | n7294 ;
  assign n35715 = n35714 ^ n7882 ^ 1'b0 ;
  assign n35716 = n17843 & ~n35715 ;
  assign n35717 = ( n2690 & n27430 ) | ( n2690 & n35716 ) | ( n27430 & n35716 ) ;
  assign n35722 = n22284 ^ n9226 ^ n697 ;
  assign n35718 = ( ~n5236 & n6433 ) | ( ~n5236 & n6842 ) | ( n6433 & n6842 ) ;
  assign n35719 = n35718 ^ n23633 ^ n692 ;
  assign n35720 = n5059 & ~n35719 ;
  assign n35721 = n13825 & n35720 ;
  assign n35723 = n35722 ^ n35721 ^ 1'b0 ;
  assign n35724 = n4256 & n33142 ;
  assign n35725 = n35724 ^ n16283 ^ 1'b0 ;
  assign n35726 = ( n2653 & ~n11306 ) | ( n2653 & n33670 ) | ( ~n11306 & n33670 ) ;
  assign n35727 = ( n11814 & n18624 ) | ( n11814 & ~n29311 ) | ( n18624 & ~n29311 ) ;
  assign n35728 = n35029 ^ n33903 ^ n9182 ;
  assign n35729 = n14772 ^ n10681 ^ n5245 ;
  assign n35730 = ( n26343 & ~n35452 ) | ( n26343 & n35729 ) | ( ~n35452 & n35729 ) ;
  assign n35731 = ( n2591 & n24698 ) | ( n2591 & n27510 ) | ( n24698 & n27510 ) ;
  assign n35732 = n13494 ^ n3834 ^ n1071 ;
  assign n35739 = n31547 ^ n29839 ^ 1'b0 ;
  assign n35740 = n15789 & n35739 ;
  assign n35733 = ( ~n2589 & n7139 ) | ( ~n2589 & n29531 ) | ( n7139 & n29531 ) ;
  assign n35734 = n35733 ^ n11580 ^ n1983 ;
  assign n35735 = n35734 ^ n31676 ^ 1'b0 ;
  assign n35736 = ( n5509 & n6373 ) | ( n5509 & ~n27448 ) | ( n6373 & ~n27448 ) ;
  assign n35737 = ( n1960 & n31582 ) | ( n1960 & ~n35736 ) | ( n31582 & ~n35736 ) ;
  assign n35738 = ( x230 & n35735 ) | ( x230 & n35737 ) | ( n35735 & n35737 ) ;
  assign n35741 = n35740 ^ n35738 ^ 1'b0 ;
  assign n35742 = ( n3476 & n4241 ) | ( n3476 & n11160 ) | ( n4241 & n11160 ) ;
  assign n35743 = n35742 ^ n33375 ^ n22698 ;
  assign n35744 = n33083 ^ n22917 ^ n9025 ;
  assign n35745 = ( n4567 & n5304 ) | ( n4567 & ~n12750 ) | ( n5304 & ~n12750 ) ;
  assign n35746 = n35745 ^ n27167 ^ n9922 ;
  assign n35747 = n13631 & n35746 ;
  assign n35748 = n35747 ^ n13065 ^ 1'b0 ;
  assign n35749 = n6201 ^ n3232 ^ x120 ;
  assign n35750 = ( n15469 & n22616 ) | ( n15469 & n35749 ) | ( n22616 & n35749 ) ;
  assign n35751 = n6498 ^ n5950 ^ 1'b0 ;
  assign n35752 = n21642 | n35751 ;
  assign n35753 = n13683 ^ n10241 ^ n4867 ;
  assign n35754 = ( n14723 & ~n16099 ) | ( n14723 & n27528 ) | ( ~n16099 & n27528 ) ;
  assign n35755 = n35754 ^ n35275 ^ n7857 ;
  assign n35756 = n35755 ^ n26093 ^ n2629 ;
  assign n35757 = ( n3982 & n7221 ) | ( n3982 & n9055 ) | ( n7221 & n9055 ) ;
  assign n35758 = n28389 & ~n35757 ;
  assign n35759 = ~n5060 & n35758 ;
  assign n35762 = n4256 & ~n13730 ;
  assign n35760 = n5203 & ~n29863 ;
  assign n35761 = ~n19817 & n35760 ;
  assign n35763 = n35762 ^ n35761 ^ n10797 ;
  assign n35764 = n5291 | n24473 ;
  assign n35765 = ( ~n18741 & n18856 ) | ( ~n18741 & n33591 ) | ( n18856 & n33591 ) ;
  assign n35766 = ( n27476 & ~n35764 ) | ( n27476 & n35765 ) | ( ~n35764 & n35765 ) ;
  assign n35767 = n35766 ^ n23552 ^ n2629 ;
  assign n35768 = ( ~n11235 & n18842 ) | ( ~n11235 & n20190 ) | ( n18842 & n20190 ) ;
  assign n35769 = n35768 ^ n20620 ^ n7639 ;
  assign n35770 = ( n480 & n17563 ) | ( n480 & ~n35769 ) | ( n17563 & ~n35769 ) ;
  assign n35772 = n3505 & ~n24479 ;
  assign n35773 = ~n2790 & n35772 ;
  assign n35774 = n35773 ^ n35585 ^ n15773 ;
  assign n35771 = n28587 ^ n18894 ^ n4841 ;
  assign n35775 = n35774 ^ n35771 ^ n32021 ;
  assign n35776 = n14807 ^ n6665 ^ 1'b0 ;
  assign n35777 = ~n3742 & n10602 ;
  assign n35778 = n35777 ^ n12311 ^ 1'b0 ;
  assign n35779 = n11340 & n35778 ;
  assign n35780 = n35779 ^ n10429 ^ 1'b0 ;
  assign n35781 = n35780 ^ n29724 ^ n16411 ;
  assign n35782 = n19667 & ~n25133 ;
  assign n35783 = n35782 ^ n28651 ^ 1'b0 ;
  assign n35784 = n34300 ^ n14138 ^ 1'b0 ;
  assign n35785 = n35783 & n35784 ;
  assign n35786 = n23840 ^ n20365 ^ n6991 ;
  assign n35787 = n17743 ^ n6399 ^ n1840 ;
  assign n35788 = n35787 ^ n30263 ^ n5971 ;
  assign n35789 = n31144 ^ n23800 ^ 1'b0 ;
  assign n35790 = n35789 ^ n34113 ^ n2692 ;
  assign n35791 = n12252 & n30752 ;
  assign n35792 = n35791 ^ n7102 ^ 1'b0 ;
  assign n35793 = n35792 ^ n22407 ^ n8112 ;
  assign n35794 = ( ~x125 & n25651 ) | ( ~x125 & n35793 ) | ( n25651 & n35793 ) ;
  assign n35795 = ( n619 & ~n8899 ) | ( n619 & n17086 ) | ( ~n8899 & n17086 ) ;
  assign n35796 = ~n1053 & n35795 ;
  assign n35797 = n19848 | n35796 ;
  assign n35798 = n13317 & n21002 ;
  assign n35799 = n35798 ^ n8882 ^ 1'b0 ;
  assign n35800 = ( ~n5895 & n26919 ) | ( ~n5895 & n35799 ) | ( n26919 & n35799 ) ;
  assign n35801 = n35518 ^ n27228 ^ 1'b0 ;
  assign n35802 = n35800 | n35801 ;
  assign n35803 = n23924 ^ n12249 ^ n9972 ;
  assign n35804 = ( x165 & n16128 ) | ( x165 & n16188 ) | ( n16128 & n16188 ) ;
  assign n35805 = n35804 ^ n31263 ^ n23800 ;
  assign n35806 = n35805 ^ n28780 ^ n8169 ;
  assign n35807 = n21244 ^ n1278 ^ 1'b0 ;
  assign n35808 = ( n16446 & ~n35806 ) | ( n16446 & n35807 ) | ( ~n35806 & n35807 ) ;
  assign n35809 = n3835 ^ n2404 ^ 1'b0 ;
  assign n35810 = n10783 & n35809 ;
  assign n35811 = n35810 ^ n20739 ^ n9696 ;
  assign n35812 = ( n4641 & n33413 ) | ( n4641 & n35811 ) | ( n33413 & n35811 ) ;
  assign n35813 = n35742 ^ n12828 ^ n11371 ;
  assign n35814 = ~n7717 & n35813 ;
  assign n35815 = n31488 ^ n24192 ^ n17246 ;
  assign n35816 = ( n17245 & ~n33624 ) | ( n17245 & n34929 ) | ( ~n33624 & n34929 ) ;
  assign n35817 = ( n4688 & ~n6506 ) | ( n4688 & n35816 ) | ( ~n6506 & n35816 ) ;
  assign n35821 = n12438 ^ n10334 ^ 1'b0 ;
  assign n35822 = n32149 & ~n35821 ;
  assign n35820 = n29392 ^ n26717 ^ n22410 ;
  assign n35818 = n21279 ^ n15637 ^ 1'b0 ;
  assign n35819 = n35818 ^ n35000 ^ n2713 ;
  assign n35823 = n35822 ^ n35820 ^ n35819 ;
  assign n35824 = ( ~n18038 & n21016 ) | ( ~n18038 & n33995 ) | ( n21016 & n33995 ) ;
  assign n35825 = ( n6647 & n16517 ) | ( n6647 & n35824 ) | ( n16517 & n35824 ) ;
  assign n35826 = n7902 ^ n7179 ^ 1'b0 ;
  assign n35827 = ( n21311 & ~n28540 ) | ( n21311 & n35826 ) | ( ~n28540 & n35826 ) ;
  assign n35828 = n35827 ^ n29300 ^ n16076 ;
  assign n35829 = ( n16935 & n17916 ) | ( n16935 & n25071 ) | ( n17916 & n25071 ) ;
  assign n35830 = n23374 ^ n4563 ^ 1'b0 ;
  assign n35831 = n12405 & n35830 ;
  assign n35832 = n35831 ^ n17227 ^ 1'b0 ;
  assign n35833 = n31141 ^ n23795 ^ 1'b0 ;
  assign n35834 = ~n31349 & n35833 ;
  assign n35835 = n35834 ^ n25504 ^ n7445 ;
  assign n35836 = n22616 | n35835 ;
  assign n35837 = ( n22511 & ~n35832 ) | ( n22511 & n35836 ) | ( ~n35832 & n35836 ) ;
  assign n35838 = n5289 & ~n20650 ;
  assign n35839 = n35838 ^ n5814 ^ 1'b0 ;
  assign n35840 = n23959 ^ n8967 ^ 1'b0 ;
  assign n35841 = n2820 & ~n35840 ;
  assign n35842 = ( n6247 & n14674 ) | ( n6247 & n19435 ) | ( n14674 & n19435 ) ;
  assign n35852 = ( n2952 & n9646 ) | ( n2952 & n11633 ) | ( n9646 & n11633 ) ;
  assign n35843 = n29951 ^ n13052 ^ n6945 ;
  assign n35844 = n3560 | n7443 ;
  assign n35845 = n3639 & n10112 ;
  assign n35846 = n13328 ^ n9955 ^ n5929 ;
  assign n35847 = n35846 ^ n4552 ^ 1'b0 ;
  assign n35848 = n35845 | n35847 ;
  assign n35849 = n35848 ^ n16169 ^ 1'b0 ;
  assign n35850 = ( n1445 & ~n35844 ) | ( n1445 & n35849 ) | ( ~n35844 & n35849 ) ;
  assign n35851 = ( n8305 & n35843 ) | ( n8305 & n35850 ) | ( n35843 & n35850 ) ;
  assign n35853 = n35852 ^ n35851 ^ n15250 ;
  assign n35854 = ( n806 & n18886 ) | ( n806 & ~n23115 ) | ( n18886 & ~n23115 ) ;
  assign n35855 = n29108 ^ n24397 ^ 1'b0 ;
  assign n35856 = ( ~n22510 & n32840 ) | ( ~n22510 & n35855 ) | ( n32840 & n35855 ) ;
  assign n35861 = ( ~n6437 & n9072 ) | ( ~n6437 & n19611 ) | ( n9072 & n19611 ) ;
  assign n35857 = n5609 & n14152 ;
  assign n35858 = ~n20876 & n31684 ;
  assign n35859 = n35858 ^ n26137 ^ 1'b0 ;
  assign n35860 = ( n29616 & ~n35857 ) | ( n29616 & n35859 ) | ( ~n35857 & n35859 ) ;
  assign n35862 = n35861 ^ n35860 ^ n21608 ;
  assign n35863 = n30027 | n31079 ;
  assign n35864 = x127 & ~n1376 ;
  assign n35866 = n23015 ^ n10091 ^ n4374 ;
  assign n35865 = n2228 | n15772 ;
  assign n35867 = n35866 ^ n35865 ^ n4061 ;
  assign n35868 = n17833 ^ n15087 ^ n8166 ;
  assign n35869 = ( x31 & n8164 ) | ( x31 & n13178 ) | ( n8164 & n13178 ) ;
  assign n35870 = ( ~n6862 & n35868 ) | ( ~n6862 & n35869 ) | ( n35868 & n35869 ) ;
  assign n35871 = ~n1243 & n15304 ;
  assign n35875 = n8395 ^ n1793 ^ n1008 ;
  assign n35874 = n11484 | n17577 ;
  assign n35876 = n35875 ^ n35874 ^ 1'b0 ;
  assign n35872 = n19223 ^ n14072 ^ 1'b0 ;
  assign n35873 = ~n6988 & n35872 ;
  assign n35877 = n35876 ^ n35873 ^ 1'b0 ;
  assign n35878 = n35871 | n35877 ;
  assign n35879 = n35878 ^ n34242 ^ n27131 ;
  assign n35880 = n23512 ^ n9890 ^ 1'b0 ;
  assign n35881 = ( n10416 & n12005 ) | ( n10416 & n16158 ) | ( n12005 & n16158 ) ;
  assign n35882 = n35881 ^ n21856 ^ n9837 ;
  assign n35883 = n35882 ^ n6953 ^ n2432 ;
  assign n35884 = ( n12428 & n16008 ) | ( n12428 & ~n35883 ) | ( n16008 & ~n35883 ) ;
  assign n35885 = n27608 ^ n8980 ^ 1'b0 ;
  assign n35886 = n11329 ^ n5289 ^ 1'b0 ;
  assign n35887 = n8844 | n35886 ;
  assign n35888 = n32528 ^ n7840 ^ 1'b0 ;
  assign n35889 = n18330 & n35888 ;
  assign n35890 = ( n12905 & ~n25798 ) | ( n12905 & n32065 ) | ( ~n25798 & n32065 ) ;
  assign n35891 = ~n5711 & n35890 ;
  assign n35892 = n6834 & ~n10072 ;
  assign n35893 = n15110 ^ n9530 ^ 1'b0 ;
  assign n35894 = n28666 & ~n35893 ;
  assign n35895 = n5504 & n35894 ;
  assign n35896 = ~n35892 & n35895 ;
  assign n35897 = ( n293 & n30120 ) | ( n293 & n35896 ) | ( n30120 & n35896 ) ;
  assign n35902 = n28076 ^ n10115 ^ n3550 ;
  assign n35898 = ( n2374 & ~n10607 ) | ( n2374 & n13297 ) | ( ~n10607 & n13297 ) ;
  assign n35899 = ( n6042 & ~n24661 ) | ( n6042 & n35898 ) | ( ~n24661 & n35898 ) ;
  assign n35900 = n31296 ^ n10982 ^ 1'b0 ;
  assign n35901 = n35899 & n35900 ;
  assign n35903 = n35902 ^ n35901 ^ n5714 ;
  assign n35904 = n4867 & n6773 ;
  assign n35905 = n9168 | n35904 ;
  assign n35906 = n8744 & ~n35905 ;
  assign n35907 = n35906 ^ n993 ^ 1'b0 ;
  assign n35908 = n28858 & n35907 ;
  assign n35909 = n12205 ^ n10433 ^ x29 ;
  assign n35910 = n9306 | n10011 ;
  assign n35911 = n35910 ^ n19348 ^ 1'b0 ;
  assign n35912 = ( n587 & ~n35909 ) | ( n587 & n35911 ) | ( ~n35909 & n35911 ) ;
  assign n35913 = ( ~n6192 & n15621 ) | ( ~n6192 & n33680 ) | ( n15621 & n33680 ) ;
  assign n35914 = n1129 | n7433 ;
  assign n35915 = ( n17841 & n27365 ) | ( n17841 & n28292 ) | ( n27365 & n28292 ) ;
  assign n35918 = ( n1397 & n21337 ) | ( n1397 & n25680 ) | ( n21337 & n25680 ) ;
  assign n35916 = n21300 ^ n11236 ^ n8013 ;
  assign n35917 = n35916 ^ n19739 ^ n7945 ;
  assign n35919 = n35918 ^ n35917 ^ 1'b0 ;
  assign n35920 = ( ~n26169 & n32991 ) | ( ~n26169 & n35919 ) | ( n32991 & n35919 ) ;
  assign n35922 = n8400 | n16865 ;
  assign n35923 = n26189 ^ n5337 ^ 1'b0 ;
  assign n35924 = ~n35922 & n35923 ;
  assign n35925 = n35924 ^ n6476 ^ 1'b0 ;
  assign n35921 = ( ~n2741 & n27191 ) | ( ~n2741 & n32229 ) | ( n27191 & n32229 ) ;
  assign n35926 = n35925 ^ n35921 ^ n27294 ;
  assign n35927 = ( n4465 & n10892 ) | ( n4465 & ~n11475 ) | ( n10892 & ~n11475 ) ;
  assign n35928 = ( ~n23215 & n28260 ) | ( ~n23215 & n35927 ) | ( n28260 & n35927 ) ;
  assign n35929 = n30366 ^ n6609 ^ 1'b0 ;
  assign n35930 = ( ~n16269 & n18895 ) | ( ~n16269 & n35929 ) | ( n18895 & n35929 ) ;
  assign n35931 = n35930 ^ n33498 ^ n29622 ;
  assign n35932 = ( ~n22075 & n35928 ) | ( ~n22075 & n35931 ) | ( n35928 & n35931 ) ;
  assign n35935 = n29117 ^ n9745 ^ n1812 ;
  assign n35933 = ~n17082 & n30384 ;
  assign n35934 = n35933 ^ n27925 ^ n8238 ;
  assign n35936 = n35935 ^ n35934 ^ 1'b0 ;
  assign n35937 = n35932 | n35936 ;
  assign n35940 = ~n9885 & n23018 ;
  assign n35938 = n13971 & ~n16152 ;
  assign n35939 = n35938 ^ n17099 ^ n849 ;
  assign n35941 = n35940 ^ n35939 ^ n30105 ;
  assign n35942 = n35941 ^ n11548 ^ n5778 ;
  assign n35943 = n20508 ^ n15784 ^ n15320 ;
  assign n35944 = ( n13320 & n24544 ) | ( n13320 & n35943 ) | ( n24544 & n35943 ) ;
  assign n35946 = n5664 | n11311 ;
  assign n35947 = n35946 ^ n5755 ^ 1'b0 ;
  assign n35948 = ( n23277 & n24004 ) | ( n23277 & n35947 ) | ( n24004 & n35947 ) ;
  assign n35945 = ( ~n7745 & n29282 ) | ( ~n7745 & n33396 ) | ( n29282 & n33396 ) ;
  assign n35949 = n35948 ^ n35945 ^ n32884 ;
  assign n35950 = n17387 ^ n7646 ^ n6119 ;
  assign n35953 = ( n781 & n4138 ) | ( n781 & n5343 ) | ( n4138 & n5343 ) ;
  assign n35951 = n6529 ^ n3254 ^ n1185 ;
  assign n35952 = ( ~n1483 & n8876 ) | ( ~n1483 & n35951 ) | ( n8876 & n35951 ) ;
  assign n35954 = n35953 ^ n35952 ^ 1'b0 ;
  assign n35955 = ~n26587 & n35954 ;
  assign n35956 = n21006 ^ n12248 ^ n8764 ;
  assign n35957 = ( n6556 & n11776 ) | ( n6556 & n17340 ) | ( n11776 & n17340 ) ;
  assign n35958 = n7923 & ~n35957 ;
  assign n35959 = n35956 & n35958 ;
  assign n35960 = n25807 & ~n27831 ;
  assign n35961 = n35960 ^ n15052 ^ 1'b0 ;
  assign n35962 = n21894 ^ n13985 ^ n8712 ;
  assign n35963 = n5525 ^ n5511 ^ n412 ;
  assign n35964 = n35599 ^ n11862 ^ n9914 ;
  assign n35965 = ( n12929 & ~n35963 ) | ( n12929 & n35964 ) | ( ~n35963 & n35964 ) ;
  assign n35966 = ( ~n7331 & n20339 ) | ( ~n7331 & n27207 ) | ( n20339 & n27207 ) ;
  assign n35968 = ( n7973 & ~n15774 ) | ( n7973 & n19039 ) | ( ~n15774 & n19039 ) ;
  assign n35969 = ( n15152 & n19151 ) | ( n15152 & ~n35968 ) | ( n19151 & ~n35968 ) ;
  assign n35970 = n35969 ^ n17562 ^ n9748 ;
  assign n35967 = n31763 ^ n27404 ^ n23469 ;
  assign n35971 = n35970 ^ n35967 ^ n4941 ;
  assign n35972 = ~n25498 & n27595 ;
  assign n35974 = ( n2206 & n10366 ) | ( n2206 & ~n16556 ) | ( n10366 & ~n16556 ) ;
  assign n35973 = n2714 & ~n11448 ;
  assign n35975 = n35974 ^ n35973 ^ 1'b0 ;
  assign n35981 = n2712 & n12035 ;
  assign n35982 = n32180 & ~n35981 ;
  assign n35978 = ( n1558 & ~n1829 ) | ( n1558 & n15349 ) | ( ~n1829 & n15349 ) ;
  assign n35977 = ( n1047 & n2082 ) | ( n1047 & ~n29746 ) | ( n2082 & ~n29746 ) ;
  assign n35979 = n35978 ^ n35977 ^ n25764 ;
  assign n35976 = n7917 | n10614 ;
  assign n35980 = n35979 ^ n35976 ^ n22459 ;
  assign n35983 = n35982 ^ n35980 ^ n33932 ;
  assign n35984 = n10931 ^ n6256 ^ n3654 ;
  assign n35985 = ( ~n2452 & n10614 ) | ( ~n2452 & n35984 ) | ( n10614 & n35984 ) ;
  assign n35986 = n12528 & n13848 ;
  assign n35987 = n35986 ^ n22527 ^ 1'b0 ;
  assign n35988 = ( n22122 & ~n35985 ) | ( n22122 & n35987 ) | ( ~n35985 & n35987 ) ;
  assign n35989 = ~n3560 & n10535 ;
  assign n35990 = n35989 ^ n6298 ^ 1'b0 ;
  assign n35991 = n35990 ^ n16362 ^ n2668 ;
  assign n35992 = ( ~n3305 & n8955 ) | ( ~n3305 & n35991 ) | ( n8955 & n35991 ) ;
  assign n35993 = ( ~n9309 & n15611 ) | ( ~n9309 & n17904 ) | ( n15611 & n17904 ) ;
  assign n35994 = n25700 ^ n14978 ^ n9014 ;
  assign n35995 = n15268 ^ n13958 ^ 1'b0 ;
  assign n35996 = ~n35994 & n35995 ;
  assign n35997 = n10313 & n28851 ;
  assign n35998 = ( n4227 & n6498 ) | ( n4227 & n23128 ) | ( n6498 & n23128 ) ;
  assign n35999 = n18389 ^ n17648 ^ n9174 ;
  assign n36000 = ( n2592 & n35998 ) | ( n2592 & n35999 ) | ( n35998 & n35999 ) ;
  assign n36004 = n30973 ^ n25162 ^ n5624 ;
  assign n36003 = n33315 ^ n20450 ^ n17143 ;
  assign n36001 = n27681 ^ n19365 ^ 1'b0 ;
  assign n36002 = n36001 ^ n9369 ^ n8701 ;
  assign n36005 = n36004 ^ n36003 ^ n36002 ;
  assign n36006 = n36005 ^ n13730 ^ n8154 ;
  assign n36007 = n29878 ^ n5382 ^ 1'b0 ;
  assign n36008 = ( n2644 & ~n16614 ) | ( n2644 & n27195 ) | ( ~n16614 & n27195 ) ;
  assign n36009 = n12819 ^ n6356 ^ x142 ;
  assign n36010 = ( ~n15655 & n36008 ) | ( ~n15655 & n36009 ) | ( n36008 & n36009 ) ;
  assign n36011 = ( n1074 & n24172 ) | ( n1074 & n27237 ) | ( n24172 & n27237 ) ;
  assign n36012 = n36011 ^ n30021 ^ n6430 ;
  assign n36013 = ( n5510 & ~n14379 ) | ( n5510 & n36012 ) | ( ~n14379 & n36012 ) ;
  assign n36014 = n35792 ^ n22307 ^ 1'b0 ;
  assign n36015 = ~n13171 & n36014 ;
  assign n36016 = ~n23125 & n36015 ;
  assign n36017 = n36016 ^ n3479 ^ 1'b0 ;
  assign n36018 = n36017 ^ n10318 ^ 1'b0 ;
  assign n36019 = n36013 | n36018 ;
  assign n36020 = n24640 ^ n24038 ^ 1'b0 ;
  assign n36021 = n14088 ^ x178 ^ x162 ;
  assign n36022 = ( n3810 & n27669 ) | ( n3810 & ~n35852 ) | ( n27669 & ~n35852 ) ;
  assign n36023 = n36021 & ~n36022 ;
  assign n36024 = n17684 ^ n11459 ^ n1410 ;
  assign n36025 = n36024 ^ n28668 ^ n17884 ;
  assign n36026 = ( ~n23512 & n23798 ) | ( ~n23512 & n28170 ) | ( n23798 & n28170 ) ;
  assign n36027 = n12306 ^ n7738 ^ n3727 ;
  assign n36028 = n12201 & ~n31688 ;
  assign n36029 = n36028 ^ n29272 ^ 1'b0 ;
  assign n36030 = n18897 ^ n16603 ^ n14411 ;
  assign n36031 = n36030 ^ n5112 ^ 1'b0 ;
  assign n36032 = n36031 ^ n31559 ^ n27502 ;
  assign n36033 = n32697 ^ n8423 ^ n3060 ;
  assign n36034 = n24215 ^ n7137 ^ n544 ;
  assign n36035 = ~n14197 & n36034 ;
  assign n36036 = n31724 & ~n34585 ;
  assign n36037 = n36036 ^ n11686 ^ 1'b0 ;
  assign n36038 = ( n637 & ~n19105 ) | ( n637 & n36037 ) | ( ~n19105 & n36037 ) ;
  assign n36039 = n35327 ^ n30546 ^ n2256 ;
  assign n36047 = n7275 & ~n10764 ;
  assign n36043 = ( n2681 & n3505 ) | ( n2681 & ~n19961 ) | ( n3505 & ~n19961 ) ;
  assign n36040 = ( n4640 & n7092 ) | ( n4640 & ~n30000 ) | ( n7092 & ~n30000 ) ;
  assign n36041 = ( n5718 & n16163 ) | ( n5718 & ~n36040 ) | ( n16163 & ~n36040 ) ;
  assign n36042 = n36041 ^ n24031 ^ n669 ;
  assign n36044 = n36043 ^ n36042 ^ 1'b0 ;
  assign n36045 = n5167 & n36044 ;
  assign n36046 = n36045 ^ n22340 ^ n7760 ;
  assign n36048 = n36047 ^ n36046 ^ n7144 ;
  assign n36049 = n36048 ^ n32921 ^ n10258 ;
  assign n36050 = n29203 ^ n4038 ^ 1'b0 ;
  assign n36051 = n10964 & ~n36050 ;
  assign n36052 = n7389 & n31859 ;
  assign n36053 = n36052 ^ n13312 ^ 1'b0 ;
  assign n36054 = ( n22418 & n26878 ) | ( n22418 & ~n27607 ) | ( n26878 & ~n27607 ) ;
  assign n36055 = n36054 ^ n27462 ^ n22919 ;
  assign n36056 = ( n8634 & n19314 ) | ( n8634 & ~n21671 ) | ( n19314 & ~n21671 ) ;
  assign n36057 = ( ~n1033 & n1157 ) | ( ~n1033 & n4304 ) | ( n1157 & n4304 ) ;
  assign n36058 = n36057 ^ n16947 ^ n15881 ;
  assign n36061 = n16160 ^ n10086 ^ 1'b0 ;
  assign n36062 = n19718 & ~n36061 ;
  assign n36059 = ( ~n6795 & n15109 ) | ( ~n6795 & n24163 ) | ( n15109 & n24163 ) ;
  assign n36060 = n36059 ^ n30873 ^ n9090 ;
  assign n36063 = n36062 ^ n36060 ^ n5845 ;
  assign n36064 = ( n14597 & ~n36058 ) | ( n14597 & n36063 ) | ( ~n36058 & n36063 ) ;
  assign n36065 = ( n36055 & n36056 ) | ( n36055 & ~n36064 ) | ( n36056 & ~n36064 ) ;
  assign n36066 = n29828 ^ n19835 ^ 1'b0 ;
  assign n36067 = n35010 ^ n7527 ^ n3305 ;
  assign n36070 = n1212 & ~n29251 ;
  assign n36071 = n9913 & n36070 ;
  assign n36068 = n29099 ^ n21606 ^ n13305 ;
  assign n36069 = ( n22496 & n35117 ) | ( n22496 & ~n36068 ) | ( n35117 & ~n36068 ) ;
  assign n36072 = n36071 ^ n36069 ^ n17320 ;
  assign n36073 = n13308 ^ n11332 ^ n9403 ;
  assign n36076 = n24786 ^ n18580 ^ 1'b0 ;
  assign n36077 = n6434 & n36076 ;
  assign n36075 = n18141 | n33797 ;
  assign n36078 = n36077 ^ n36075 ^ 1'b0 ;
  assign n36074 = n25597 ^ n24403 ^ n2457 ;
  assign n36079 = n36078 ^ n36074 ^ n14620 ;
  assign n36080 = n7269 & n36079 ;
  assign n36081 = n25229 ^ n17076 ^ 1'b0 ;
  assign n36082 = n3429 & ~n36081 ;
  assign n36083 = n21052 ^ n11980 ^ n6295 ;
  assign n36084 = n28330 ^ n24657 ^ n17814 ;
  assign n36085 = ( ~n6434 & n36083 ) | ( ~n6434 & n36084 ) | ( n36083 & n36084 ) ;
  assign n36090 = ~n615 & n20416 ;
  assign n36091 = ( ~n1520 & n16435 ) | ( ~n1520 & n36090 ) | ( n16435 & n36090 ) ;
  assign n36092 = n36091 ^ n12048 ^ n1695 ;
  assign n36087 = n25729 ^ n24733 ^ n12405 ;
  assign n36088 = n36087 ^ n16366 ^ n6642 ;
  assign n36086 = n12498 & n27390 ;
  assign n36089 = n36088 ^ n36086 ^ 1'b0 ;
  assign n36093 = n36092 ^ n36089 ^ n24340 ;
  assign n36094 = ( n11489 & n17056 ) | ( n11489 & ~n18898 ) | ( n17056 & ~n18898 ) ;
  assign n36095 = ( n1693 & n34003 ) | ( n1693 & n36094 ) | ( n34003 & n36094 ) ;
  assign n36096 = n7107 ^ n3838 ^ 1'b0 ;
  assign n36097 = ( ~n24603 & n36095 ) | ( ~n24603 & n36096 ) | ( n36095 & n36096 ) ;
  assign n36098 = n5890 ^ n4566 ^ 1'b0 ;
  assign n36099 = n15859 ^ n383 ^ 1'b0 ;
  assign n36100 = n26684 & ~n32220 ;
  assign n36101 = ( n13865 & ~n27063 ) | ( n13865 & n36100 ) | ( ~n27063 & n36100 ) ;
  assign n36102 = ~n36099 & n36101 ;
  assign n36103 = n2927 & ~n6376 ;
  assign n36104 = n3162 & n36103 ;
  assign n36105 = n36104 ^ n27805 ^ n4829 ;
  assign n36106 = ( ~n1183 & n8770 ) | ( ~n1183 & n21180 ) | ( n8770 & n21180 ) ;
  assign n36107 = ( n1639 & n2631 ) | ( n1639 & n13599 ) | ( n2631 & n13599 ) ;
  assign n36108 = n2565 & n36107 ;
  assign n36109 = ( n1286 & n12526 ) | ( n1286 & n36108 ) | ( n12526 & n36108 ) ;
  assign n36110 = n11501 | n34842 ;
  assign n36111 = n12625 ^ n7403 ^ 1'b0 ;
  assign n36112 = n5057 & ~n36111 ;
  assign n36113 = n36112 ^ n35902 ^ n8160 ;
  assign n36114 = ( ~n12492 & n17614 ) | ( ~n12492 & n32017 ) | ( n17614 & n32017 ) ;
  assign n36115 = ~n4898 & n11687 ;
  assign n36116 = n12599 & n36115 ;
  assign n36117 = n36116 ^ n28490 ^ 1'b0 ;
  assign n36118 = n17633 & ~n36117 ;
  assign n36119 = ( n10660 & ~n22866 ) | ( n10660 & n36118 ) | ( ~n22866 & n36118 ) ;
  assign n36120 = ~n8348 & n14063 ;
  assign n36121 = ~n11716 & n36120 ;
  assign n36122 = n6779 ^ n1685 ^ n979 ;
  assign n36123 = n11034 & ~n15310 ;
  assign n36124 = ( n15559 & n16187 ) | ( n15559 & ~n36123 ) | ( n16187 & ~n36123 ) ;
  assign n36125 = ( n12805 & n25569 ) | ( n12805 & ~n31795 ) | ( n25569 & ~n31795 ) ;
  assign n36126 = ( n11044 & n26450 ) | ( n11044 & ~n36125 ) | ( n26450 & ~n36125 ) ;
  assign n36129 = n33035 ^ n1829 ^ n1112 ;
  assign n36127 = ~n3594 & n25799 ;
  assign n36128 = n36127 ^ n33470 ^ 1'b0 ;
  assign n36130 = n36129 ^ n36128 ^ n19502 ;
  assign n36131 = ( n3357 & n14398 ) | ( n3357 & n24669 ) | ( n14398 & n24669 ) ;
  assign n36132 = n36131 ^ n32941 ^ n32319 ;
  assign n36134 = ( ~n5237 & n27241 ) | ( ~n5237 & n31041 ) | ( n27241 & n31041 ) ;
  assign n36133 = n29004 ^ n14685 ^ n5822 ;
  assign n36135 = n36134 ^ n36133 ^ n5829 ;
  assign n36136 = n23715 ^ n17777 ^ n1194 ;
  assign n36137 = ( n15472 & n19455 ) | ( n15472 & ~n36136 ) | ( n19455 & ~n36136 ) ;
  assign n36138 = n9029 ^ n4057 ^ 1'b0 ;
  assign n36139 = n36138 ^ n24629 ^ n4618 ;
  assign n36140 = ( ~n24994 & n31094 ) | ( ~n24994 & n36139 ) | ( n31094 & n36139 ) ;
  assign n36145 = n35875 ^ n9034 ^ n6130 ;
  assign n36144 = n17867 ^ n14716 ^ n4460 ;
  assign n36141 = ~n12616 & n23555 ;
  assign n36142 = n14257 & n36141 ;
  assign n36143 = ( n800 & n22781 ) | ( n800 & ~n36142 ) | ( n22781 & ~n36142 ) ;
  assign n36146 = n36145 ^ n36144 ^ n36143 ;
  assign n36147 = n36146 ^ n16219 ^ 1'b0 ;
  assign n36148 = x211 & ~n13393 ;
  assign n36149 = ~n3787 & n36148 ;
  assign n36150 = n36149 ^ n4017 ^ 1'b0 ;
  assign n36151 = n36150 ^ n32332 ^ n20826 ;
  assign n36152 = n36151 ^ n16874 ^ n2739 ;
  assign n36153 = ( n29342 & ~n33590 ) | ( n29342 & n36152 ) | ( ~n33590 & n36152 ) ;
  assign n36154 = ~n6588 & n22267 ;
  assign n36155 = n2221 & n36154 ;
  assign n36156 = n669 & n25725 ;
  assign n36157 = n36155 & n36156 ;
  assign n36158 = n20466 | n36157 ;
  assign n36159 = n5294 & ~n36158 ;
  assign n36160 = ( ~n2795 & n12639 ) | ( ~n2795 & n16334 ) | ( n12639 & n16334 ) ;
  assign n36161 = n6533 | n14266 ;
  assign n36162 = n36161 ^ n16758 ^ 1'b0 ;
  assign n36163 = ~n810 & n36162 ;
  assign n36164 = n36163 ^ n7287 ^ 1'b0 ;
  assign n36165 = n36164 ^ n328 ^ 1'b0 ;
  assign n36166 = ~n36160 & n36165 ;
  assign n36167 = n36166 ^ n3873 ^ 1'b0 ;
  assign n36168 = n36167 ^ n8429 ^ 1'b0 ;
  assign n36169 = n3453 & ~n12283 ;
  assign n36175 = ( n2025 & n6136 ) | ( n2025 & n30278 ) | ( n6136 & n30278 ) ;
  assign n36176 = n36175 ^ n26544 ^ n14043 ;
  assign n36177 = n36176 ^ n18147 ^ n13481 ;
  assign n36170 = ( ~n663 & n8442 ) | ( ~n663 & n10106 ) | ( n8442 & n10106 ) ;
  assign n36171 = n36170 ^ n8709 ^ n5721 ;
  assign n36172 = ( n3104 & ~n11645 ) | ( n3104 & n36171 ) | ( ~n11645 & n36171 ) ;
  assign n36173 = n30618 ^ n22040 ^ n9059 ;
  assign n36174 = ( n2426 & n36172 ) | ( n2426 & n36173 ) | ( n36172 & n36173 ) ;
  assign n36178 = n36177 ^ n36174 ^ n35694 ;
  assign n36179 = ( n895 & n36169 ) | ( n895 & ~n36178 ) | ( n36169 & ~n36178 ) ;
  assign n36181 = n27648 ^ n6752 ^ 1'b0 ;
  assign n36180 = ( n4334 & ~n17794 ) | ( n4334 & n29280 ) | ( ~n17794 & n29280 ) ;
  assign n36182 = n36181 ^ n36180 ^ n8973 ;
  assign n36183 = n21188 ^ n21178 ^ n3679 ;
  assign n36184 = n23668 ^ n20346 ^ n18237 ;
  assign n36185 = ( ~n4947 & n21086 ) | ( ~n4947 & n36184 ) | ( n21086 & n36184 ) ;
  assign n36186 = n36185 ^ n27019 ^ n20965 ;
  assign n36187 = ~n639 & n7317 ;
  assign n36191 = n2446 & ~n5580 ;
  assign n36192 = n9443 & n36191 ;
  assign n36193 = n36192 ^ n11647 ^ n3303 ;
  assign n36188 = ( ~n1392 & n5146 ) | ( ~n1392 & n32781 ) | ( n5146 & n32781 ) ;
  assign n36189 = n18365 ^ n6383 ^ n2744 ;
  assign n36190 = ( n30175 & ~n36188 ) | ( n30175 & n36189 ) | ( ~n36188 & n36189 ) ;
  assign n36194 = n36193 ^ n36190 ^ n34418 ;
  assign n36195 = n8562 & ~n14581 ;
  assign n36196 = ~n29561 & n36195 ;
  assign n36197 = ( n3142 & n23967 ) | ( n3142 & n36196 ) | ( n23967 & n36196 ) ;
  assign n36198 = n11404 ^ n4778 ^ 1'b0 ;
  assign n36199 = n1425 | n7402 ;
  assign n36200 = ~n36198 & n36199 ;
  assign n36201 = ( n9041 & n12748 ) | ( n9041 & n36200 ) | ( n12748 & n36200 ) ;
  assign n36206 = ( n5799 & ~n17426 ) | ( n5799 & n23685 ) | ( ~n17426 & n23685 ) ;
  assign n36202 = n23566 ^ n4239 ^ n2162 ;
  assign n36203 = n13776 ^ n9236 ^ n6670 ;
  assign n36204 = n36203 ^ n18062 ^ n7675 ;
  assign n36205 = ( n24486 & ~n36202 ) | ( n24486 & n36204 ) | ( ~n36202 & n36204 ) ;
  assign n36207 = n36206 ^ n36205 ^ n29513 ;
  assign n36208 = ( n9954 & n13482 ) | ( n9954 & n28879 ) | ( n13482 & n28879 ) ;
  assign n36210 = n22288 ^ n20477 ^ 1'b0 ;
  assign n36211 = ~n27013 & n36210 ;
  assign n36209 = n22380 ^ n13532 ^ n9012 ;
  assign n36212 = n36211 ^ n36209 ^ 1'b0 ;
  assign n36213 = ( ~n24291 & n29893 ) | ( ~n24291 & n36212 ) | ( n29893 & n36212 ) ;
  assign n36214 = n36213 ^ n18586 ^ n554 ;
  assign n36215 = n11243 ^ n8881 ^ 1'b0 ;
  assign n36216 = n1866 & n36215 ;
  assign n36217 = ( n4351 & n11375 ) | ( n4351 & ~n12572 ) | ( n11375 & ~n12572 ) ;
  assign n36218 = n25442 ^ n4320 ^ 1'b0 ;
  assign n36219 = ( n15355 & ~n36217 ) | ( n15355 & n36218 ) | ( ~n36217 & n36218 ) ;
  assign n36220 = n34218 ^ n22594 ^ 1'b0 ;
  assign n36221 = n14290 ^ n6356 ^ 1'b0 ;
  assign n36222 = n25426 & n36221 ;
  assign n36223 = ~n36220 & n36222 ;
  assign n36224 = n35697 ^ n6726 ^ 1'b0 ;
  assign n36225 = n13847 | n36224 ;
  assign n36226 = n23241 ^ n13746 ^ 1'b0 ;
  assign n36231 = n14721 ^ n5911 ^ 1'b0 ;
  assign n36230 = n28149 ^ n22784 ^ n15845 ;
  assign n36228 = n20898 ^ n14886 ^ n8397 ;
  assign n36227 = n1558 & n9642 ;
  assign n36229 = n36228 ^ n36227 ^ n8586 ;
  assign n36232 = n36231 ^ n36230 ^ n36229 ;
  assign n36233 = ( ~n27129 & n35843 ) | ( ~n27129 & n36232 ) | ( n35843 & n36232 ) ;
  assign n36234 = n26421 & n35248 ;
  assign n36235 = n36234 ^ n1303 ^ 1'b0 ;
  assign n36237 = n7766 | n12694 ;
  assign n36238 = n36237 ^ n19697 ^ n10210 ;
  assign n36236 = ~n5406 & n15961 ;
  assign n36239 = n36238 ^ n36236 ^ 1'b0 ;
  assign n36240 = ( n1840 & ~n36235 ) | ( n1840 & n36239 ) | ( ~n36235 & n36239 ) ;
  assign n36241 = ( n10316 & n29671 ) | ( n10316 & ~n30065 ) | ( n29671 & ~n30065 ) ;
  assign n36243 = ( n8634 & n17947 ) | ( n8634 & n19523 ) | ( n17947 & n19523 ) ;
  assign n36242 = ( n5683 & n10291 ) | ( n5683 & ~n14427 ) | ( n10291 & ~n14427 ) ;
  assign n36244 = n36243 ^ n36242 ^ n16301 ;
  assign n36245 = ( n8334 & n16740 ) | ( n8334 & n36244 ) | ( n16740 & n36244 ) ;
  assign n36246 = ~n4938 & n21635 ;
  assign n36247 = n10268 & n19418 ;
  assign n36248 = n36247 ^ n19420 ^ n16339 ;
  assign n36249 = ( ~n27013 & n36246 ) | ( ~n27013 & n36248 ) | ( n36246 & n36248 ) ;
  assign n36250 = n29817 ^ n28270 ^ 1'b0 ;
  assign n36251 = n5953 & ~n36250 ;
  assign n36252 = n5185 & ~n33795 ;
  assign n36253 = n3564 & ~n20603 ;
  assign n36254 = n36253 ^ n19714 ^ n10978 ;
  assign n36255 = n5240 | n36254 ;
  assign n36256 = n11127 | n36255 ;
  assign n36257 = ( x195 & ~n7210 ) | ( x195 & n33705 ) | ( ~n7210 & n33705 ) ;
  assign n36258 = ( n2359 & ~n23128 ) | ( n2359 & n33093 ) | ( ~n23128 & n33093 ) ;
  assign n36259 = n36258 ^ n23049 ^ n2417 ;
  assign n36260 = ( n6463 & n36257 ) | ( n6463 & n36259 ) | ( n36257 & n36259 ) ;
  assign n36261 = n36260 ^ n18335 ^ 1'b0 ;
  assign n36262 = n13077 & n36261 ;
  assign n36263 = ( n1282 & n36256 ) | ( n1282 & ~n36262 ) | ( n36256 & ~n36262 ) ;
  assign n36264 = ( n10237 & ~n19390 ) | ( n10237 & n30649 ) | ( ~n19390 & n30649 ) ;
  assign n36265 = n13566 ^ n3641 ^ 1'b0 ;
  assign n36266 = n7236 | n36265 ;
  assign n36267 = ( ~n8184 & n36264 ) | ( ~n8184 & n36266 ) | ( n36264 & n36266 ) ;
  assign n36268 = n36267 ^ n4744 ^ 1'b0 ;
  assign n36269 = n6010 | n22361 ;
  assign n36270 = n36269 ^ n22191 ^ n19333 ;
  assign n36271 = ( n4719 & ~n18470 ) | ( n4719 & n34651 ) | ( ~n18470 & n34651 ) ;
  assign n36272 = ( n3037 & n6059 ) | ( n3037 & n12959 ) | ( n6059 & n12959 ) ;
  assign n36273 = n16262 | n27300 ;
  assign n36274 = ( n18128 & ~n36272 ) | ( n18128 & n36273 ) | ( ~n36272 & n36273 ) ;
  assign n36275 = ( n856 & ~n16610 ) | ( n856 & n33288 ) | ( ~n16610 & n33288 ) ;
  assign n36276 = n36275 ^ n25441 ^ n7600 ;
  assign n36277 = n11684 ^ n5783 ^ n3609 ;
  assign n36278 = n36277 ^ n15740 ^ x196 ;
  assign n36279 = n7046 | n14312 ;
  assign n36280 = n36279 ^ n10382 ^ 1'b0 ;
  assign n36281 = ( ~n2718 & n17289 ) | ( ~n2718 & n36280 ) | ( n17289 & n36280 ) ;
  assign n36282 = ( n16955 & n36278 ) | ( n16955 & ~n36281 ) | ( n36278 & ~n36281 ) ;
  assign n36283 = n4010 | n13583 ;
  assign n36284 = n36283 ^ n7920 ^ 1'b0 ;
  assign n36285 = ~n32702 & n36284 ;
  assign n36286 = ( n7345 & n12629 ) | ( n7345 & ~n18754 ) | ( n12629 & ~n18754 ) ;
  assign n36287 = n11021 ^ n479 ^ 1'b0 ;
  assign n36288 = n36286 & n36287 ;
  assign n36289 = n36288 ^ n9489 ^ n8642 ;
  assign n36290 = n36289 ^ n31347 ^ 1'b0 ;
  assign n36291 = ( n906 & n4103 ) | ( n906 & ~n14347 ) | ( n4103 & ~n14347 ) ;
  assign n36292 = ( n9046 & n26749 ) | ( n9046 & n34678 ) | ( n26749 & n34678 ) ;
  assign n36293 = ( n18742 & n36291 ) | ( n18742 & n36292 ) | ( n36291 & n36292 ) ;
  assign n36294 = ( n1050 & ~n13657 ) | ( n1050 & n29066 ) | ( ~n13657 & n29066 ) ;
  assign n36295 = ( n32569 & ~n36293 ) | ( n32569 & n36294 ) | ( ~n36293 & n36294 ) ;
  assign n36296 = n9265 | n29185 ;
  assign n36297 = n26719 | n36296 ;
  assign n36298 = n13749 ^ n10704 ^ 1'b0 ;
  assign n36299 = n36298 ^ n16103 ^ 1'b0 ;
  assign n36300 = n23101 ^ n16033 ^ n12103 ;
  assign n36301 = n36300 ^ n26986 ^ n14898 ;
  assign n36302 = ( ~n1587 & n3689 ) | ( ~n1587 & n5142 ) | ( n3689 & n5142 ) ;
  assign n36303 = n36302 ^ n16689 ^ n10477 ;
  assign n36304 = n22390 ^ n9205 ^ n8561 ;
  assign n36305 = n36304 ^ n23941 ^ n401 ;
  assign n36306 = n21668 ^ n7696 ^ 1'b0 ;
  assign n36307 = n11965 ^ n10251 ^ n5502 ;
  assign n36308 = ( n25764 & n32604 ) | ( n25764 & ~n36307 ) | ( n32604 & ~n36307 ) ;
  assign n36309 = ( n10467 & n18316 ) | ( n10467 & ~n31446 ) | ( n18316 & ~n31446 ) ;
  assign n36310 = ~n6907 & n36309 ;
  assign n36312 = n4926 ^ n2445 ^ n623 ;
  assign n36311 = n20296 ^ n10649 ^ n4939 ;
  assign n36313 = n36312 ^ n36311 ^ x199 ;
  assign n36314 = n28649 ^ n17891 ^ n17082 ;
  assign n36315 = n10095 ^ n699 ^ 1'b0 ;
  assign n36316 = ~n25896 & n36315 ;
  assign n36317 = ( x84 & n4345 ) | ( x84 & ~n36316 ) | ( n4345 & ~n36316 ) ;
  assign n36318 = n36317 ^ n1528 ^ 1'b0 ;
  assign n36319 = n9366 | n36318 ;
  assign n36320 = ( n13822 & ~n17537 ) | ( n13822 & n19120 ) | ( ~n17537 & n19120 ) ;
  assign n36321 = n36320 ^ n11358 ^ 1'b0 ;
  assign n36322 = n36001 ^ n28871 ^ 1'b0 ;
  assign n36327 = n26394 ^ n11378 ^ n7806 ;
  assign n36328 = n36327 ^ n32890 ^ n13930 ;
  assign n36323 = n11447 & n21430 ;
  assign n36324 = n36323 ^ n18592 ^ n6122 ;
  assign n36325 = n27293 | n36324 ;
  assign n36326 = n19378 | n36325 ;
  assign n36329 = n36328 ^ n36326 ^ 1'b0 ;
  assign n36330 = ( n8352 & n16455 ) | ( n8352 & n20767 ) | ( n16455 & n20767 ) ;
  assign n36331 = n36330 ^ n6923 ^ 1'b0 ;
  assign n36332 = n23251 & n36331 ;
  assign n36333 = n36332 ^ n15776 ^ 1'b0 ;
  assign n36334 = n36333 ^ n26702 ^ n649 ;
  assign n36335 = n32313 ^ n19109 ^ n2756 ;
  assign n36336 = n36335 ^ n26778 ^ 1'b0 ;
  assign n36337 = n14222 | n20341 ;
  assign n36338 = n18258 & ~n36337 ;
  assign n36339 = ( n7303 & n8657 ) | ( n7303 & ~n10230 ) | ( n8657 & ~n10230 ) ;
  assign n36340 = n21081 | n36339 ;
  assign n36341 = n6833 | n36340 ;
  assign n36342 = ( n2635 & n4920 ) | ( n2635 & ~n22553 ) | ( n4920 & ~n22553 ) ;
  assign n36343 = n36342 ^ n12286 ^ n3509 ;
  assign n36344 = n36341 & n36343 ;
  assign n36345 = n36344 ^ n24078 ^ 1'b0 ;
  assign n36346 = n15503 ^ n7875 ^ n7465 ;
  assign n36347 = n11378 & n36346 ;
  assign n36348 = n14271 & n36347 ;
  assign n36349 = ( ~n12730 & n17594 ) | ( ~n12730 & n22682 ) | ( n17594 & n22682 ) ;
  assign n36350 = n17798 ^ n5306 ^ n3708 ;
  assign n36351 = n36350 ^ n10624 ^ 1'b0 ;
  assign n36352 = n4762 | n36351 ;
  assign n36353 = n21383 ^ n11465 ^ n3749 ;
  assign n36354 = n697 & n23655 ;
  assign n36355 = ( x237 & ~n15716 ) | ( x237 & n36354 ) | ( ~n15716 & n36354 ) ;
  assign n36356 = n2012 & n15521 ;
  assign n36357 = n36356 ^ n2970 ^ 1'b0 ;
  assign n36358 = ( ~n6426 & n11203 ) | ( ~n6426 & n36357 ) | ( n11203 & n36357 ) ;
  assign n36359 = n26785 & ~n36358 ;
  assign n36360 = n36359 ^ n23495 ^ 1'b0 ;
  assign n36361 = n36360 ^ n14567 ^ n4281 ;
  assign n36364 = ( n4932 & ~n6031 ) | ( n4932 & n6450 ) | ( ~n6031 & n6450 ) ;
  assign n36365 = n36364 ^ n568 ^ x107 ;
  assign n36362 = ( n1616 & n8038 ) | ( n1616 & n15853 ) | ( n8038 & n15853 ) ;
  assign n36363 = n36362 ^ n16976 ^ 1'b0 ;
  assign n36366 = n36365 ^ n36363 ^ n3223 ;
  assign n36367 = n10383 ^ n7940 ^ n5080 ;
  assign n36368 = n35256 ^ n3134 ^ 1'b0 ;
  assign n36369 = n36367 & n36368 ;
  assign n36370 = ( ~n2677 & n5710 ) | ( ~n2677 & n28394 ) | ( n5710 & n28394 ) ;
  assign n36371 = n36370 ^ n32834 ^ n9454 ;
  assign n36372 = n5048 & n21060 ;
  assign n36373 = ~n36371 & n36372 ;
  assign n36374 = n26048 ^ n16034 ^ n2204 ;
  assign n36375 = ( ~n2911 & n20284 ) | ( ~n2911 & n36374 ) | ( n20284 & n36374 ) ;
  assign n36376 = n20319 & ~n25912 ;
  assign n36377 = n8463 | n16069 ;
  assign n36378 = n36377 ^ n9983 ^ 1'b0 ;
  assign n36379 = n36171 ^ n8936 ^ 1'b0 ;
  assign n36380 = ~n4310 & n36379 ;
  assign n36381 = ( n7149 & n36378 ) | ( n7149 & n36380 ) | ( n36378 & n36380 ) ;
  assign n36382 = ( n19560 & n22827 ) | ( n19560 & n26719 ) | ( n22827 & n26719 ) ;
  assign n36383 = n36382 ^ n1582 ^ 1'b0 ;
  assign n36384 = n20206 ^ n12641 ^ n7172 ;
  assign n36385 = ( n3866 & n34975 ) | ( n3866 & ~n36384 ) | ( n34975 & ~n36384 ) ;
  assign n36386 = n14213 ^ n10476 ^ 1'b0 ;
  assign n36387 = n27826 ^ n8624 ^ 1'b0 ;
  assign n36388 = n11892 & n36387 ;
  assign n36389 = n36388 ^ n22499 ^ n6544 ;
  assign n36390 = ( n15554 & ~n21375 ) | ( n15554 & n24466 ) | ( ~n21375 & n24466 ) ;
  assign n36391 = n36390 ^ n28588 ^ n12476 ;
  assign n36392 = n31923 ^ n26539 ^ n9280 ;
  assign n36394 = n13683 ^ n13404 ^ n4918 ;
  assign n36393 = n18481 | n29664 ;
  assign n36395 = n36394 ^ n36393 ^ 1'b0 ;
  assign n36396 = n36395 ^ n13205 ^ n4604 ;
  assign n36397 = n35485 ^ n25343 ^ n20204 ;
  assign n36398 = ~n7949 & n20787 ;
  assign n36399 = n36398 ^ n6039 ^ 1'b0 ;
  assign n36406 = n11153 ^ n11058 ^ 1'b0 ;
  assign n36407 = n16785 & ~n36406 ;
  assign n36405 = n18397 ^ n16745 ^ 1'b0 ;
  assign n36408 = n36407 ^ n36405 ^ n20245 ;
  assign n36404 = n12359 & ~n28322 ;
  assign n36409 = n36408 ^ n36404 ^ 1'b0 ;
  assign n36401 = n4500 & n35291 ;
  assign n36402 = n12352 & n36401 ;
  assign n36403 = n36402 ^ n23780 ^ n21664 ;
  assign n36400 = n5132 | n23781 ;
  assign n36410 = n36409 ^ n36403 ^ n36400 ;
  assign n36411 = n36399 | n36410 ;
  assign n36412 = n26173 ^ n3033 ^ 1'b0 ;
  assign n36413 = ~n7353 & n36412 ;
  assign n36414 = n36413 ^ n17548 ^ n6534 ;
  assign n36415 = ( n753 & n5475 ) | ( n753 & ~n6306 ) | ( n5475 & ~n6306 ) ;
  assign n36416 = ( n3242 & n12111 ) | ( n3242 & ~n13320 ) | ( n12111 & ~n13320 ) ;
  assign n36417 = ( ~n25218 & n36415 ) | ( ~n25218 & n36416 ) | ( n36415 & n36416 ) ;
  assign n36418 = ( n32293 & n36414 ) | ( n32293 & ~n36417 ) | ( n36414 & ~n36417 ) ;
  assign n36419 = ( ~n11261 & n12818 ) | ( ~n11261 & n21408 ) | ( n12818 & n21408 ) ;
  assign n36420 = n11260 ^ n855 ^ 1'b0 ;
  assign n36421 = ( ~n8668 & n10902 ) | ( ~n8668 & n36420 ) | ( n10902 & n36420 ) ;
  assign n36422 = n36421 ^ n36219 ^ n11935 ;
  assign n36424 = n851 & n18483 ;
  assign n36425 = ~n15113 & n36424 ;
  assign n36426 = ( ~n5170 & n7300 ) | ( ~n5170 & n36425 ) | ( n7300 & n36425 ) ;
  assign n36423 = n21003 ^ n19902 ^ n15807 ;
  assign n36427 = n36426 ^ n36423 ^ n13603 ;
  assign n36428 = ( n6679 & n19268 ) | ( n6679 & ~n21016 ) | ( n19268 & ~n21016 ) ;
  assign n36429 = n6519 | n36428 ;
  assign n36430 = n9333 & ~n21006 ;
  assign n36431 = ~n26891 & n36430 ;
  assign n36432 = n36431 ^ n10485 ^ 1'b0 ;
  assign n36433 = n8505 & n36432 ;
  assign n36434 = n30697 ^ n9786 ^ n7074 ;
  assign n36435 = ( n6167 & n22667 ) | ( n6167 & n34706 ) | ( n22667 & n34706 ) ;
  assign n36436 = ( n13577 & ~n26977 ) | ( n13577 & n29258 ) | ( ~n26977 & n29258 ) ;
  assign n36437 = ( ~n755 & n3375 ) | ( ~n755 & n36436 ) | ( n3375 & n36436 ) ;
  assign n36438 = n19608 ^ n10091 ^ n5278 ;
  assign n36440 = n301 | n12389 ;
  assign n36441 = n36440 ^ n3569 ^ 1'b0 ;
  assign n36439 = ( n9217 & n13442 ) | ( n9217 & ~n16124 ) | ( n13442 & ~n16124 ) ;
  assign n36442 = n36441 ^ n36439 ^ n17054 ;
  assign n36443 = ( n5614 & n7161 ) | ( n5614 & ~n12467 ) | ( n7161 & ~n12467 ) ;
  assign n36444 = ( n4717 & ~n17820 ) | ( n4717 & n20405 ) | ( ~n17820 & n20405 ) ;
  assign n36445 = n36444 ^ n6586 ^ 1'b0 ;
  assign n36446 = n36443 & n36445 ;
  assign n36448 = n36002 ^ n19131 ^ n13953 ;
  assign n36447 = n7648 | n18952 ;
  assign n36449 = n36448 ^ n36447 ^ n19617 ;
  assign n36450 = n22698 ^ n15451 ^ 1'b0 ;
  assign n36451 = ~n5584 & n36450 ;
  assign n36457 = ( n4299 & n8738 ) | ( n4299 & n14979 ) | ( n8738 & n14979 ) ;
  assign n36456 = ( n5697 & ~n7509 ) | ( n5697 & n32708 ) | ( ~n7509 & n32708 ) ;
  assign n36452 = n22623 ^ n6714 ^ n1847 ;
  assign n36453 = ( n7915 & n20582 ) | ( n7915 & ~n36452 ) | ( n20582 & ~n36452 ) ;
  assign n36454 = n36453 ^ n10415 ^ 1'b0 ;
  assign n36455 = ~n29606 & n36454 ;
  assign n36458 = n36457 ^ n36456 ^ n36455 ;
  assign n36459 = ( n2903 & n11134 ) | ( n2903 & n33400 ) | ( n11134 & n33400 ) ;
  assign n36460 = n305 | n3379 ;
  assign n36461 = n4336 | n36460 ;
  assign n36462 = ( n21384 & n25349 ) | ( n21384 & ~n36461 ) | ( n25349 & ~n36461 ) ;
  assign n36463 = ( n13616 & n17641 ) | ( n13616 & ~n36462 ) | ( n17641 & ~n36462 ) ;
  assign n36464 = n28203 ^ n26066 ^ n19113 ;
  assign n36465 = n8267 | n36464 ;
  assign n36467 = n22622 ^ n19858 ^ 1'b0 ;
  assign n36466 = n5474 & n35387 ;
  assign n36468 = n36467 ^ n36466 ^ 1'b0 ;
  assign n36469 = ( n714 & n14872 ) | ( n714 & n29062 ) | ( n14872 & n29062 ) ;
  assign n36470 = n36469 ^ n25462 ^ n24454 ;
  assign n36471 = ( ~n2753 & n17246 ) | ( ~n2753 & n18673 ) | ( n17246 & n18673 ) ;
  assign n36475 = ( n19591 & n25341 ) | ( n19591 & ~n25591 ) | ( n25341 & ~n25591 ) ;
  assign n36472 = ( ~n19271 & n23587 ) | ( ~n19271 & n27744 ) | ( n23587 & n27744 ) ;
  assign n36473 = n20141 ^ n4391 ^ 1'b0 ;
  assign n36474 = n36472 | n36473 ;
  assign n36476 = n36475 ^ n36474 ^ n8548 ;
  assign n36477 = n9619 ^ n6862 ^ 1'b0 ;
  assign n36478 = ( ~n2070 & n27518 ) | ( ~n2070 & n36477 ) | ( n27518 & n36477 ) ;
  assign n36479 = ( n2296 & n9445 ) | ( n2296 & n19402 ) | ( n9445 & n19402 ) ;
  assign n36480 = n36479 ^ n29558 ^ n18631 ;
  assign n36481 = n31216 ^ n18134 ^ n2258 ;
  assign n36482 = ( n4134 & n36480 ) | ( n4134 & n36481 ) | ( n36480 & n36481 ) ;
  assign n36483 = ( n4175 & n14050 ) | ( n4175 & ~n23375 ) | ( n14050 & ~n23375 ) ;
  assign n36484 = n1738 & ~n26980 ;
  assign n36485 = ( ~n21870 & n21978 ) | ( ~n21870 & n27989 ) | ( n21978 & n27989 ) ;
  assign n36486 = ( n10567 & ~n20251 ) | ( n10567 & n36485 ) | ( ~n20251 & n36485 ) ;
  assign n36487 = n36486 ^ n2120 ^ n1255 ;
  assign n36488 = ( n11821 & ~n14747 ) | ( n11821 & n36487 ) | ( ~n14747 & n36487 ) ;
  assign n36489 = n21425 ^ n8735 ^ n5201 ;
  assign n36490 = n33682 ^ n12102 ^ 1'b0 ;
  assign n36491 = n27755 & n36490 ;
  assign n36492 = n31998 ^ n26999 ^ n21317 ;
  assign n36493 = n10492 & ~n34482 ;
  assign n36494 = n36493 ^ n1928 ^ 1'b0 ;
  assign n36495 = n12660 ^ n11431 ^ 1'b0 ;
  assign n36496 = n7189 & n36495 ;
  assign n36497 = n6579 ^ n3039 ^ n1510 ;
  assign n36498 = n36497 ^ n22034 ^ 1'b0 ;
  assign n36499 = n21976 & ~n24947 ;
  assign n36500 = n15358 ^ n10110 ^ x73 ;
  assign n36501 = ( n30650 & n36499 ) | ( n30650 & ~n36500 ) | ( n36499 & ~n36500 ) ;
  assign n36502 = n20973 | n21997 ;
  assign n36503 = n9619 | n36502 ;
  assign n36504 = ( n2401 & ~n8736 ) | ( n2401 & n36503 ) | ( ~n8736 & n36503 ) ;
  assign n36505 = n36504 ^ n1194 ^ 1'b0 ;
  assign n36506 = n36505 ^ n1428 ^ 1'b0 ;
  assign n36508 = n32972 ^ n4140 ^ 1'b0 ;
  assign n36507 = n29963 ^ n4924 ^ n3616 ;
  assign n36509 = n36508 ^ n36507 ^ n16692 ;
  assign n36516 = ~n2196 & n21806 ;
  assign n36512 = ( ~n11647 & n15457 ) | ( ~n11647 & n33664 ) | ( n15457 & n33664 ) ;
  assign n36513 = ~x62 & n36512 ;
  assign n36514 = n36513 ^ n3718 ^ 1'b0 ;
  assign n36515 = ( n4667 & ~n23083 ) | ( n4667 & n36514 ) | ( ~n23083 & n36514 ) ;
  assign n36510 = ( n13825 & n15496 ) | ( n13825 & n24561 ) | ( n15496 & n24561 ) ;
  assign n36511 = ( ~n338 & n11446 ) | ( ~n338 & n36510 ) | ( n11446 & n36510 ) ;
  assign n36517 = n36516 ^ n36515 ^ n36511 ;
  assign n36518 = n31375 ^ n24341 ^ 1'b0 ;
  assign n36519 = ( n15034 & n16970 ) | ( n15034 & n29729 ) | ( n16970 & n29729 ) ;
  assign n36520 = n26693 ^ n8599 ^ n744 ;
  assign n36521 = ( n6906 & n30919 ) | ( n6906 & n36520 ) | ( n30919 & n36520 ) ;
  assign n36522 = n10752 ^ n8294 ^ n3158 ;
  assign n36523 = n8650 & ~n36522 ;
  assign n36524 = ( n5869 & n36521 ) | ( n5869 & ~n36523 ) | ( n36521 & ~n36523 ) ;
  assign n36525 = n8687 | n16781 ;
  assign n36526 = n36525 ^ n32619 ^ n11343 ;
  assign n36527 = ( n5530 & ~n20272 ) | ( n5530 & n20437 ) | ( ~n20272 & n20437 ) ;
  assign n36529 = ( n4014 & n5843 ) | ( n4014 & n5849 ) | ( n5843 & n5849 ) ;
  assign n36530 = ( ~n1647 & n6794 ) | ( ~n1647 & n36529 ) | ( n6794 & n36529 ) ;
  assign n36528 = n24082 ^ n4802 ^ n1111 ;
  assign n36531 = n36530 ^ n36528 ^ n29908 ;
  assign n36532 = n36531 ^ n33903 ^ n12835 ;
  assign n36533 = n36527 & ~n36532 ;
  assign n36534 = n36533 ^ n13681 ^ 1'b0 ;
  assign n36535 = n3687 & ~n36094 ;
  assign n36537 = n25670 ^ n892 ^ 1'b0 ;
  assign n36536 = n4727 & ~n34631 ;
  assign n36538 = n36537 ^ n36536 ^ n2172 ;
  assign n36539 = ( n7925 & n12320 ) | ( n7925 & ~n17211 ) | ( n12320 & ~n17211 ) ;
  assign n36540 = n20517 ^ n5210 ^ 1'b0 ;
  assign n36541 = n34022 & n36540 ;
  assign n36542 = n5791 & n36541 ;
  assign n36543 = n4742 & ~n12590 ;
  assign n36544 = n28263 ^ n22472 ^ n766 ;
  assign n36545 = n35904 ^ n32726 ^ n14063 ;
  assign n36546 = n36545 ^ n14273 ^ n9051 ;
  assign n36547 = n24027 ^ n21139 ^ n20687 ;
  assign n36548 = ( ~n3202 & n7310 ) | ( ~n3202 & n13313 ) | ( n7310 & n13313 ) ;
  assign n36549 = n26152 & ~n36548 ;
  assign n36550 = n7082 | n11886 ;
  assign n36552 = ( n5116 & n12385 ) | ( n5116 & n26561 ) | ( n12385 & n26561 ) ;
  assign n36553 = n36552 ^ n24110 ^ n952 ;
  assign n36551 = n16149 | n29927 ;
  assign n36554 = n36553 ^ n36551 ^ n8322 ;
  assign n36555 = n23122 ^ n8730 ^ n3397 ;
  assign n36557 = n1374 | n3279 ;
  assign n36558 = n36557 ^ n348 ^ 1'b0 ;
  assign n36559 = n12619 & n36558 ;
  assign n36560 = n36559 ^ n33523 ^ n19000 ;
  assign n36556 = n1187 | n4896 ;
  assign n36561 = n36560 ^ n36556 ^ 1'b0 ;
  assign n36562 = n36561 ^ n29804 ^ n6848 ;
  assign n36563 = n36562 ^ n25115 ^ 1'b0 ;
  assign n36564 = n31630 ^ n9132 ^ n5615 ;
  assign n36565 = n36564 ^ n21025 ^ 1'b0 ;
  assign n36566 = ( n10626 & ~n19162 ) | ( n10626 & n36565 ) | ( ~n19162 & n36565 ) ;
  assign n36568 = n27789 ^ n25599 ^ n4216 ;
  assign n36569 = n36568 ^ n8536 ^ 1'b0 ;
  assign n36567 = n4827 | n5556 ;
  assign n36570 = n36569 ^ n36567 ^ n32180 ;
  assign n36571 = ~n6977 & n28494 ;
  assign n36572 = n36571 ^ n5625 ^ 1'b0 ;
  assign n36573 = n33919 ^ n24918 ^ 1'b0 ;
  assign n36574 = n18326 ^ n781 ^ 1'b0 ;
  assign n36575 = ( n6522 & n6709 ) | ( n6522 & ~n20855 ) | ( n6709 & ~n20855 ) ;
  assign n36576 = n21438 ^ n18771 ^ 1'b0 ;
  assign n36577 = n36576 ^ n14041 ^ n3839 ;
  assign n36578 = n36577 ^ n5577 ^ n1868 ;
  assign n36579 = ( n6873 & n13544 ) | ( n6873 & n32022 ) | ( n13544 & n32022 ) ;
  assign n36580 = n11295 & ~n18348 ;
  assign n36581 = n36580 ^ n11767 ^ 1'b0 ;
  assign n36582 = n12765 ^ n8055 ^ 1'b0 ;
  assign n36583 = n8976 & ~n36582 ;
  assign n36584 = n31126 ^ n21616 ^ n1761 ;
  assign n36585 = n11541 | n36584 ;
  assign n36586 = n36583 | n36585 ;
  assign n36587 = x113 | n32459 ;
  assign n36588 = ( n9033 & ~n13779 ) | ( n9033 & n14505 ) | ( ~n13779 & n14505 ) ;
  assign n36589 = n8442 & ~n10017 ;
  assign n36590 = n36589 ^ n10237 ^ 1'b0 ;
  assign n36591 = n36590 ^ n35316 ^ n24411 ;
  assign n36592 = n36591 ^ n3847 ^ n2645 ;
  assign n36593 = n27556 ^ n16882 ^ n1868 ;
  assign n36594 = ~n2215 & n15404 ;
  assign n36595 = n20171 & n36594 ;
  assign n36596 = ( n7130 & ~n31789 ) | ( n7130 & n36595 ) | ( ~n31789 & n36595 ) ;
  assign n36597 = n36593 & ~n36596 ;
  assign n36598 = ~n23235 & n36597 ;
  assign n36599 = n33226 ^ n8475 ^ n6169 ;
  assign n36600 = n9834 & ~n36599 ;
  assign n36601 = ~n6063 & n36600 ;
  assign n36602 = n36601 ^ n16699 ^ n13938 ;
  assign n36603 = n16158 ^ n13564 ^ n11378 ;
  assign n36604 = n36603 ^ n19539 ^ 1'b0 ;
  assign n36605 = n36604 ^ n23781 ^ n20684 ;
  assign n36606 = n1968 & ~n7667 ;
  assign n36607 = n36606 ^ n19469 ^ 1'b0 ;
  assign n36608 = n36607 ^ n9097 ^ n1862 ;
  assign n36609 = n36608 ^ n31937 ^ n8930 ;
  assign n36610 = ~n8019 & n36609 ;
  assign n36611 = n16456 ^ n15492 ^ n699 ;
  assign n36612 = n36611 ^ n33555 ^ n15559 ;
  assign n36613 = ( n28339 & ~n32897 ) | ( n28339 & n36134 ) | ( ~n32897 & n36134 ) ;
  assign n36614 = n36613 ^ n25052 ^ n8154 ;
  assign n36615 = ( n9350 & n30693 ) | ( n9350 & ~n36614 ) | ( n30693 & ~n36614 ) ;
  assign n36617 = n11887 ^ n8707 ^ n1803 ;
  assign n36616 = n14851 ^ n4029 ^ n378 ;
  assign n36618 = n36617 ^ n36616 ^ n7638 ;
  assign n36619 = n11379 ^ n6995 ^ 1'b0 ;
  assign n36620 = n1465 & ~n36619 ;
  assign n36621 = n36620 ^ n27826 ^ n8684 ;
  assign n36622 = n30833 ^ n23891 ^ n3753 ;
  assign n36623 = n4586 & n36622 ;
  assign n36624 = n8983 ^ n5926 ^ n3871 ;
  assign n36625 = n36624 ^ n26759 ^ n8486 ;
  assign n36626 = ( n31484 & n36623 ) | ( n31484 & n36625 ) | ( n36623 & n36625 ) ;
  assign n36627 = n21944 ^ n14743 ^ 1'b0 ;
  assign n36629 = n29756 ^ n6977 ^ x188 ;
  assign n36630 = ( n11582 & n26595 ) | ( n11582 & ~n36629 ) | ( n26595 & ~n36629 ) ;
  assign n36628 = n35567 ^ n24931 ^ 1'b0 ;
  assign n36631 = n36630 ^ n36628 ^ n12766 ;
  assign n36632 = n7507 ^ n7110 ^ 1'b0 ;
  assign n36633 = ( n22510 & n36426 ) | ( n22510 & n36632 ) | ( n36426 & n36632 ) ;
  assign n36634 = n36633 ^ n13465 ^ n3158 ;
  assign n36635 = n28577 ^ n26511 ^ n4556 ;
  assign n36636 = n36635 ^ n24360 ^ n2135 ;
  assign n36637 = ( ~n7352 & n12857 ) | ( ~n7352 & n36636 ) | ( n12857 & n36636 ) ;
  assign n36638 = n2039 | n17574 ;
  assign n36639 = n36637 | n36638 ;
  assign n36640 = ( ~n3864 & n8036 ) | ( ~n3864 & n22887 ) | ( n8036 & n22887 ) ;
  assign n36641 = ( ~x15 & n12284 ) | ( ~x15 & n36640 ) | ( n12284 & n36640 ) ;
  assign n36642 = n36641 ^ n31362 ^ n9452 ;
  assign n36643 = ( n1268 & n2412 ) | ( n1268 & n8268 ) | ( n2412 & n8268 ) ;
  assign n36644 = n29052 ^ n16418 ^ n9177 ;
  assign n36645 = ( n14634 & n36643 ) | ( n14634 & n36644 ) | ( n36643 & n36644 ) ;
  assign n36650 = ( n11899 & ~n17074 ) | ( n11899 & n19381 ) | ( ~n17074 & n19381 ) ;
  assign n36646 = n8427 ^ n6517 ^ n2854 ;
  assign n36647 = n36646 ^ n3659 ^ n2756 ;
  assign n36648 = n14971 | n36647 ;
  assign n36649 = n10661 & ~n36648 ;
  assign n36651 = n36650 ^ n36649 ^ n34842 ;
  assign n36652 = ( x27 & ~n3948 ) | ( x27 & n30198 ) | ( ~n3948 & n30198 ) ;
  assign n36653 = ( n2492 & ~n16981 ) | ( n2492 & n33680 ) | ( ~n16981 & n33680 ) ;
  assign n36654 = ( ~n18818 & n25842 ) | ( ~n18818 & n36653 ) | ( n25842 & n36653 ) ;
  assign n36658 = n2700 & n18328 ;
  assign n36655 = ( n4084 & ~n6134 ) | ( n4084 & n23602 ) | ( ~n6134 & n23602 ) ;
  assign n36656 = n36655 ^ x200 ^ 1'b0 ;
  assign n36657 = n16165 & ~n36656 ;
  assign n36659 = n36658 ^ n36657 ^ n21232 ;
  assign n36660 = n35518 ^ n24610 ^ x75 ;
  assign n36661 = n32782 ^ n13522 ^ 1'b0 ;
  assign n36662 = n25846 | n36661 ;
  assign n36663 = n36662 ^ n8358 ^ 1'b0 ;
  assign n36664 = n15209 ^ n5301 ^ 1'b0 ;
  assign n36665 = n4466 & ~n36664 ;
  assign n36666 = n36665 ^ n20194 ^ n17750 ;
  assign n36667 = n19430 ^ n18878 ^ 1'b0 ;
  assign n36668 = ( n3636 & ~n16700 ) | ( n3636 & n32295 ) | ( ~n16700 & n32295 ) ;
  assign n36669 = ( n12945 & n20870 ) | ( n12945 & n28223 ) | ( n20870 & n28223 ) ;
  assign n36670 = ( ~n35321 & n36668 ) | ( ~n35321 & n36669 ) | ( n36668 & n36669 ) ;
  assign n36671 = ( n4717 & n8068 ) | ( n4717 & ~n20317 ) | ( n8068 & ~n20317 ) ;
  assign n36672 = n30570 ^ n4726 ^ n4666 ;
  assign n36673 = ( ~n18398 & n36671 ) | ( ~n18398 & n36672 ) | ( n36671 & n36672 ) ;
  assign n36676 = n410 | n7297 ;
  assign n36677 = ( n3693 & ~n4697 ) | ( n3693 & n36676 ) | ( ~n4697 & n36676 ) ;
  assign n36674 = n3420 ^ n3377 ^ 1'b0 ;
  assign n36675 = n36674 ^ n2668 ^ 1'b0 ;
  assign n36678 = n36677 ^ n36675 ^ n11037 ;
  assign n36679 = n15777 ^ n4834 ^ 1'b0 ;
  assign n36680 = n36679 ^ n16607 ^ n11772 ;
  assign n36681 = n34071 ^ n30154 ^ 1'b0 ;
  assign n36682 = ~n26236 & n36681 ;
  assign n36683 = n9099 ^ n1941 ^ n1511 ;
  assign n36684 = n36683 ^ n18667 ^ n2569 ;
  assign n36685 = n8140 ^ n4471 ^ n2723 ;
  assign n36686 = n1534 ^ n1256 ^ 1'b0 ;
  assign n36687 = n36686 ^ n25478 ^ n1743 ;
  assign n36688 = n5748 & n36687 ;
  assign n36689 = ~n6331 & n36688 ;
  assign n36690 = ( n4974 & n9485 ) | ( n4974 & ~n36689 ) | ( n9485 & ~n36689 ) ;
  assign n36691 = ( ~n2499 & n29059 ) | ( ~n2499 & n36690 ) | ( n29059 & n36690 ) ;
  assign n36692 = ( n22883 & ~n35117 ) | ( n22883 & n35232 ) | ( ~n35117 & n35232 ) ;
  assign n36693 = n36692 ^ n32539 ^ n30175 ;
  assign n36698 = ( n4871 & ~n9635 ) | ( n4871 & n17063 ) | ( ~n9635 & n17063 ) ;
  assign n36695 = n28269 ^ n13042 ^ 1'b0 ;
  assign n36694 = n6786 & ~n25929 ;
  assign n36696 = n36695 ^ n36694 ^ 1'b0 ;
  assign n36697 = n4726 | n36696 ;
  assign n36699 = n36698 ^ n36697 ^ 1'b0 ;
  assign n36700 = n31887 ^ n3394 ^ 1'b0 ;
  assign n36701 = ( ~n11732 & n22363 ) | ( ~n11732 & n36700 ) | ( n22363 & n36700 ) ;
  assign n36702 = n27436 ^ n24767 ^ n20042 ;
  assign n36703 = ( n7319 & ~n31189 ) | ( n7319 & n36702 ) | ( ~n31189 & n36702 ) ;
  assign n36704 = n1439 & n36655 ;
  assign n36705 = n2334 ^ n2175 ^ 1'b0 ;
  assign n36706 = n1372 ^ n549 ^ 1'b0 ;
  assign n36707 = ~n6951 & n36706 ;
  assign n36708 = ( n287 & n4846 ) | ( n287 & ~n36707 ) | ( n4846 & ~n36707 ) ;
  assign n36709 = ( n6226 & ~n11839 ) | ( n6226 & n36708 ) | ( ~n11839 & n36708 ) ;
  assign n36710 = ( n14902 & ~n27560 ) | ( n14902 & n36709 ) | ( ~n27560 & n36709 ) ;
  assign n36711 = ( n4166 & n28597 ) | ( n4166 & ~n36710 ) | ( n28597 & ~n36710 ) ;
  assign n36712 = ( ~n21061 & n36705 ) | ( ~n21061 & n36711 ) | ( n36705 & n36711 ) ;
  assign n36713 = n26032 ^ n21161 ^ 1'b0 ;
  assign n36714 = ~n1094 & n36713 ;
  assign n36715 = ( n13769 & ~n29696 ) | ( n13769 & n36714 ) | ( ~n29696 & n36714 ) ;
  assign n36716 = n36715 ^ n26628 ^ 1'b0 ;
  assign n36717 = n36211 ^ n10250 ^ n3237 ;
  assign n36718 = n36717 ^ n11260 ^ 1'b0 ;
  assign n36719 = n36474 ^ n22937 ^ 1'b0 ;
  assign n36720 = n19496 & n36719 ;
  assign n36721 = ( ~n6584 & n13321 ) | ( ~n6584 & n26150 ) | ( n13321 & n26150 ) ;
  assign n36722 = ( n3632 & n6178 ) | ( n3632 & ~n24801 ) | ( n6178 & ~n24801 ) ;
  assign n36723 = n9311 ^ n1366 ^ n877 ;
  assign n36724 = n36723 ^ n35260 ^ n16688 ;
  assign n36725 = ( n9958 & n26194 ) | ( n9958 & n33538 ) | ( n26194 & n33538 ) ;
  assign n36726 = ( n2469 & n2939 ) | ( n2469 & ~n30049 ) | ( n2939 & ~n30049 ) ;
  assign n36728 = n799 & ~n9776 ;
  assign n36727 = n22528 ^ n18610 ^ n14152 ;
  assign n36729 = n36728 ^ n36727 ^ n7592 ;
  assign n36731 = n18122 ^ n7455 ^ n787 ;
  assign n36732 = ( n9874 & ~n14111 ) | ( n9874 & n36731 ) | ( ~n14111 & n36731 ) ;
  assign n36733 = n5301 | n6223 ;
  assign n36734 = n25821 | n36733 ;
  assign n36735 = ( ~n24617 & n36732 ) | ( ~n24617 & n36734 ) | ( n36732 & n36734 ) ;
  assign n36730 = n31631 & n33609 ;
  assign n36736 = n36735 ^ n36730 ^ n32600 ;
  assign n36737 = n22519 ^ n4412 ^ 1'b0 ;
  assign n36738 = n8078 & ~n36737 ;
  assign n36739 = n36738 ^ n26533 ^ n17454 ;
  assign n36740 = ~n12173 & n36739 ;
  assign n36741 = n13779 | n30904 ;
  assign n36742 = n36741 ^ n34441 ^ 1'b0 ;
  assign n36743 = n1483 & n3593 ;
  assign n36744 = ( n5899 & ~n20321 ) | ( n5899 & n36743 ) | ( ~n20321 & n36743 ) ;
  assign n36745 = n16047 ^ n14638 ^ 1'b0 ;
  assign n36746 = n1394 & ~n36745 ;
  assign n36747 = n36746 ^ n16244 ^ 1'b0 ;
  assign n36748 = n15520 ^ n7627 ^ 1'b0 ;
  assign n36749 = n36748 ^ n11539 ^ n944 ;
  assign n36750 = n28946 ^ n8038 ^ 1'b0 ;
  assign n36751 = n6974 & ~n36750 ;
  assign n36752 = n36749 | n36751 ;
  assign n36753 = n32359 ^ n23250 ^ n5156 ;
  assign n36754 = n6586 ^ n5527 ^ n853 ;
  assign n36755 = n36754 ^ n11540 ^ n5352 ;
  assign n36756 = n36755 ^ n21441 ^ n6728 ;
  assign n36757 = n32508 ^ n7876 ^ n6424 ;
  assign n36758 = n36307 ^ n2094 ^ n1198 ;
  assign n36759 = ~n10451 & n15370 ;
  assign n36760 = n36759 ^ n2017 ^ 1'b0 ;
  assign n36761 = ( n21705 & n36758 ) | ( n21705 & n36760 ) | ( n36758 & n36760 ) ;
  assign n36762 = n6958 | n10703 ;
  assign n36763 = n22229 ^ n7408 ^ n6299 ;
  assign n36764 = n17677 ^ n13696 ^ n2735 ;
  assign n36765 = n36764 ^ n16381 ^ 1'b0 ;
  assign n36766 = n36765 ^ n16171 ^ 1'b0 ;
  assign n36767 = n36763 & ~n36766 ;
  assign n36768 = ( ~n15179 & n36762 ) | ( ~n15179 & n36767 ) | ( n36762 & n36767 ) ;
  assign n36769 = n27310 ^ n24640 ^ n4153 ;
  assign n36771 = ( n11377 & ~n17022 ) | ( n11377 & n25226 ) | ( ~n17022 & n25226 ) ;
  assign n36770 = n21299 & ~n36510 ;
  assign n36772 = n36771 ^ n36770 ^ n17611 ;
  assign n36773 = n8755 ^ n949 ^ 1'b0 ;
  assign n36774 = ( n1971 & n20156 ) | ( n1971 & ~n36773 ) | ( n20156 & ~n36773 ) ;
  assign n36775 = n27269 ^ n24078 ^ 1'b0 ;
  assign n36776 = n6803 & ~n36775 ;
  assign n36777 = n28665 ^ n10554 ^ 1'b0 ;
  assign n36778 = n36667 ^ n18444 ^ 1'b0 ;
  assign n36779 = n36777 | n36778 ;
  assign n36780 = n27271 ^ n11106 ^ 1'b0 ;
  assign n36782 = n16538 ^ n10978 ^ n2776 ;
  assign n36781 = n11195 | n12108 ;
  assign n36783 = n36782 ^ n36781 ^ 1'b0 ;
  assign n36784 = n36783 ^ n9614 ^ n2172 ;
  assign n36785 = n6109 & n12465 ;
  assign n36786 = ~n3870 & n36785 ;
  assign n36787 = n27413 ^ n7171 ^ n5701 ;
  assign n36788 = n21537 ^ n20049 ^ n1361 ;
  assign n36789 = n20333 ^ n451 ^ 1'b0 ;
  assign n36790 = n34441 ^ n19790 ^ n9186 ;
  assign n36791 = n36790 ^ n9410 ^ n6997 ;
  assign n36792 = n36791 ^ n9384 ^ 1'b0 ;
  assign n36793 = ( ~n14517 & n36789 ) | ( ~n14517 & n36792 ) | ( n36789 & n36792 ) ;
  assign n36794 = ( n6864 & n10768 ) | ( n6864 & ~n18817 ) | ( n10768 & ~n18817 ) ;
  assign n36796 = n34048 ^ n33797 ^ n12885 ;
  assign n36795 = n12108 ^ n7793 ^ n2026 ;
  assign n36797 = n36796 ^ n36795 ^ n14730 ;
  assign n36798 = ~n5235 & n32558 ;
  assign n36799 = n36798 ^ n14357 ^ 1'b0 ;
  assign n36800 = ( n17476 & ~n21363 ) | ( n17476 & n31268 ) | ( ~n21363 & n31268 ) ;
  assign n36801 = n36800 ^ n22756 ^ n16109 ;
  assign n36802 = x179 & n36801 ;
  assign n36803 = ~n16189 & n17451 ;
  assign n36804 = n36803 ^ n6036 ^ 1'b0 ;
  assign n36805 = ~n8791 & n36804 ;
  assign n36806 = n19071 ^ n5699 ^ 1'b0 ;
  assign n36807 = n15431 ^ n4523 ^ n652 ;
  assign n36808 = ( n2832 & n13301 ) | ( n2832 & n28578 ) | ( n13301 & n28578 ) ;
  assign n36809 = n36808 ^ n21436 ^ n5593 ;
  assign n36810 = ( n19325 & n36807 ) | ( n19325 & ~n36809 ) | ( n36807 & ~n36809 ) ;
  assign n36811 = n5967 & ~n9075 ;
  assign n36812 = n36811 ^ n17969 ^ n3867 ;
  assign n36813 = ( ~n14662 & n31433 ) | ( ~n14662 & n36812 ) | ( n31433 & n36812 ) ;
  assign n36814 = ( n8663 & ~n21671 ) | ( n8663 & n28997 ) | ( ~n21671 & n28997 ) ;
  assign n36815 = n36814 ^ n19665 ^ 1'b0 ;
  assign n36816 = n27596 & n36815 ;
  assign n36817 = n36816 ^ n25749 ^ n4809 ;
  assign n36818 = ( n3915 & n10374 ) | ( n3915 & ~n28000 ) | ( n10374 & ~n28000 ) ;
  assign n36819 = n3244 & ~n23130 ;
  assign n36820 = n36819 ^ n28047 ^ 1'b0 ;
  assign n36821 = n4756 ^ n2844 ^ 1'b0 ;
  assign n36822 = n36820 & n36821 ;
  assign n36823 = n22374 ^ n17827 ^ n17771 ;
  assign n36824 = ( n22537 & n25478 ) | ( n22537 & n36823 ) | ( n25478 & n36823 ) ;
  assign n36825 = n36822 & ~n36824 ;
  assign n36826 = n9605 ^ n9433 ^ 1'b0 ;
  assign n36827 = n17664 & ~n36826 ;
  assign n36828 = ( n6069 & ~n27420 ) | ( n6069 & n35957 ) | ( ~n27420 & n35957 ) ;
  assign n36829 = n5180 | n33666 ;
  assign n36830 = n31475 ^ n16834 ^ n15175 ;
  assign n36831 = ( n7968 & ~n16101 ) | ( n7968 & n36830 ) | ( ~n16101 & n36830 ) ;
  assign n36832 = n36831 ^ n16817 ^ 1'b0 ;
  assign n36833 = n12376 ^ n9615 ^ n4388 ;
  assign n36834 = ( n1360 & n9635 ) | ( n1360 & n16937 ) | ( n9635 & n16937 ) ;
  assign n36835 = n36834 ^ n33819 ^ n27406 ;
  assign n36836 = ( n13015 & n36833 ) | ( n13015 & ~n36835 ) | ( n36833 & ~n36835 ) ;
  assign n36837 = n22391 ^ n10605 ^ 1'b0 ;
  assign n36838 = n21829 & ~n36837 ;
  assign n36839 = ( n19264 & n25603 ) | ( n19264 & n36838 ) | ( n25603 & n36838 ) ;
  assign n36840 = n20429 ^ n12034 ^ 1'b0 ;
  assign n36841 = ( n4146 & n12811 ) | ( n4146 & ~n36840 ) | ( n12811 & ~n36840 ) ;
  assign n36842 = n4382 & n18215 ;
  assign n36843 = n36842 ^ n20753 ^ 1'b0 ;
  assign n36844 = ( n16168 & n18796 ) | ( n16168 & n33751 ) | ( n18796 & n33751 ) ;
  assign n36845 = n25091 ^ n14683 ^ n14114 ;
  assign n36846 = n36845 ^ n22563 ^ n15899 ;
  assign n36847 = ( n7197 & n32988 ) | ( n7197 & n36846 ) | ( n32988 & n36846 ) ;
  assign n36848 = n6955 ^ n4460 ^ n336 ;
  assign n36849 = ( ~n1334 & n22426 ) | ( ~n1334 & n36848 ) | ( n22426 & n36848 ) ;
  assign n36850 = n36849 ^ n32098 ^ n6067 ;
  assign n36852 = n2925 | n4755 ;
  assign n36853 = n25376 ^ n12407 ^ 1'b0 ;
  assign n36854 = n7547 & n8507 ;
  assign n36855 = n36853 | n36854 ;
  assign n36856 = n36852 & ~n36855 ;
  assign n36851 = n23587 ^ n10513 ^ n4002 ;
  assign n36857 = n36856 ^ n36851 ^ n13669 ;
  assign n36858 = ( n18037 & ~n18091 ) | ( n18037 & n22928 ) | ( ~n18091 & n22928 ) ;
  assign n36859 = ( n5237 & n24582 ) | ( n5237 & ~n28589 ) | ( n24582 & ~n28589 ) ;
  assign n36860 = ( n11142 & ~n30648 ) | ( n11142 & n36859 ) | ( ~n30648 & n36859 ) ;
  assign n36861 = ( n11808 & ~n12050 ) | ( n11808 & n29432 ) | ( ~n12050 & n29432 ) ;
  assign n36862 = ~n2320 & n11156 ;
  assign n36863 = ( ~n7143 & n28831 ) | ( ~n7143 & n36862 ) | ( n28831 & n36862 ) ;
  assign n36864 = n36863 ^ n25344 ^ x176 ;
  assign n36865 = n1481 & ~n11654 ;
  assign n36866 = n36865 ^ n23548 ^ n18010 ;
  assign n36867 = ( n6975 & n8002 ) | ( n6975 & n12394 ) | ( n8002 & n12394 ) ;
  assign n36868 = n35871 | n36867 ;
  assign n36869 = n10006 ^ n9353 ^ n6287 ;
  assign n36870 = ( ~n23041 & n27476 ) | ( ~n23041 & n36869 ) | ( n27476 & n36869 ) ;
  assign n36871 = ( n22675 & n36614 ) | ( n22675 & n36870 ) | ( n36614 & n36870 ) ;
  assign n36872 = n9253 ^ n7383 ^ 1'b0 ;
  assign n36873 = ( n646 & ~n23891 ) | ( n646 & n31926 ) | ( ~n23891 & n31926 ) ;
  assign n36874 = n36872 & n36873 ;
  assign n36875 = n36874 ^ n15674 ^ 1'b0 ;
  assign n36876 = ~n16405 & n30984 ;
  assign n36877 = n33073 ^ n15740 ^ n13519 ;
  assign n36878 = n36876 & n36877 ;
  assign n36879 = ~n14308 & n36878 ;
  assign n36880 = n20658 ^ n2271 ^ 1'b0 ;
  assign n36881 = ( n2093 & n2802 ) | ( n2093 & n8454 ) | ( n2802 & n8454 ) ;
  assign n36882 = ( n3879 & n10459 ) | ( n3879 & ~n11311 ) | ( n10459 & ~n11311 ) ;
  assign n36884 = n9710 ^ n5187 ^ 1'b0 ;
  assign n36885 = n11672 & ~n36884 ;
  assign n36894 = n13719 | n17235 ;
  assign n36895 = n36894 ^ n17156 ^ 1'b0 ;
  assign n36892 = n9817 & n12124 ;
  assign n36893 = n36892 ^ n9686 ^ n6501 ;
  assign n36887 = n3977 ^ n3500 ^ 1'b0 ;
  assign n36888 = ( n993 & n12162 ) | ( n993 & n28284 ) | ( n12162 & n28284 ) ;
  assign n36889 = ( ~n28427 & n36887 ) | ( ~n28427 & n36888 ) | ( n36887 & n36888 ) ;
  assign n36886 = n5446 & n7348 ;
  assign n36890 = n36889 ^ n36886 ^ 1'b0 ;
  assign n36891 = ( n4744 & n23901 ) | ( n4744 & ~n36890 ) | ( n23901 & ~n36890 ) ;
  assign n36896 = n36895 ^ n36893 ^ n36891 ;
  assign n36897 = ( n7828 & n36885 ) | ( n7828 & ~n36896 ) | ( n36885 & ~n36896 ) ;
  assign n36883 = ( n10957 & ~n16019 ) | ( n10957 & n30698 ) | ( ~n16019 & n30698 ) ;
  assign n36898 = n36897 ^ n36883 ^ n14331 ;
  assign n36899 = ( n7607 & ~n16800 ) | ( n7607 & n26971 ) | ( ~n16800 & n26971 ) ;
  assign n36900 = n6607 ^ n1864 ^ 1'b0 ;
  assign n36901 = ( n1180 & ~n5813 ) | ( n1180 & n7062 ) | ( ~n5813 & n7062 ) ;
  assign n36902 = n36901 ^ n25193 ^ x109 ;
  assign n36903 = n1606 & n36902 ;
  assign n36904 = ~n36900 & n36903 ;
  assign n36905 = n785 & ~n15265 ;
  assign n36906 = ~n25619 & n36905 ;
  assign n36909 = ( n16737 & n24338 ) | ( n16737 & ~n32364 ) | ( n24338 & ~n32364 ) ;
  assign n36910 = n36909 ^ n28465 ^ n23049 ;
  assign n36907 = ( n5385 & n8438 ) | ( n5385 & ~n12405 ) | ( n8438 & ~n12405 ) ;
  assign n36908 = n36907 ^ n32619 ^ n5273 ;
  assign n36911 = n36910 ^ n36908 ^ n32533 ;
  assign n36912 = ( n464 & n5982 ) | ( n464 & ~n16708 ) | ( n5982 & ~n16708 ) ;
  assign n36913 = ( ~n3947 & n9028 ) | ( ~n3947 & n13953 ) | ( n9028 & n13953 ) ;
  assign n36914 = n33015 ^ n11816 ^ n10725 ;
  assign n36915 = n32522 ^ n30268 ^ 1'b0 ;
  assign n36916 = ( ~n4280 & n8381 ) | ( ~n4280 & n36291 ) | ( n8381 & n36291 ) ;
  assign n36917 = ( ~n9048 & n13912 ) | ( ~n9048 & n36916 ) | ( n13912 & n36916 ) ;
  assign n36918 = n29467 ^ n19381 ^ n9269 ;
  assign n36919 = n670 & ~n36918 ;
  assign n36920 = ~n13951 & n36919 ;
  assign n36921 = n16388 ^ n12109 ^ 1'b0 ;
  assign n36922 = n12082 & n36921 ;
  assign n36923 = n26617 ^ n6852 ^ n6197 ;
  assign n36924 = ~n29491 & n36923 ;
  assign n36925 = n36924 ^ n12357 ^ 1'b0 ;
  assign n36926 = n15151 ^ n7205 ^ n4012 ;
  assign n36927 = ( n2152 & n22490 ) | ( n2152 & ~n25141 ) | ( n22490 & ~n25141 ) ;
  assign n36928 = ( n28295 & ~n36926 ) | ( n28295 & n36927 ) | ( ~n36926 & n36927 ) ;
  assign n36929 = ( ~n10354 & n26751 ) | ( ~n10354 & n31854 ) | ( n26751 & n31854 ) ;
  assign n36930 = n25090 ^ n20432 ^ 1'b0 ;
  assign n36931 = n7304 & n36930 ;
  assign n36932 = n29143 & n36931 ;
  assign n36935 = n14824 ^ n12834 ^ n1103 ;
  assign n36933 = n16049 ^ n9588 ^ 1'b0 ;
  assign n36934 = n3940 & ~n36933 ;
  assign n36936 = n36935 ^ n36934 ^ n32945 ;
  assign n36937 = n7580 ^ n4099 ^ n2852 ;
  assign n36938 = n27554 & ~n31690 ;
  assign n36939 = ~n7487 & n36938 ;
  assign n36940 = ( n10172 & n36937 ) | ( n10172 & n36939 ) | ( n36937 & n36939 ) ;
  assign n36941 = n36940 ^ n30575 ^ n8980 ;
  assign n36942 = n7590 & ~n34944 ;
  assign n36943 = n2602 & n36942 ;
  assign n36944 = ~n2777 & n26240 ;
  assign n36945 = n35005 & n36944 ;
  assign n36946 = n7276 & ~n36945 ;
  assign n36947 = n36943 & n36946 ;
  assign n36948 = n32064 ^ n28295 ^ n13409 ;
  assign n36949 = n36948 ^ n24702 ^ 1'b0 ;
  assign n36950 = ( n15306 & ~n18415 ) | ( n15306 & n27563 ) | ( ~n18415 & n27563 ) ;
  assign n36951 = n36950 ^ n32015 ^ n15358 ;
  assign n36954 = n13918 ^ n8835 ^ n3464 ;
  assign n36953 = n11604 & n18920 ;
  assign n36955 = n36954 ^ n36953 ^ 1'b0 ;
  assign n36952 = ( n4653 & n11747 ) | ( n4653 & ~n22057 ) | ( n11747 & ~n22057 ) ;
  assign n36956 = n36955 ^ n36952 ^ 1'b0 ;
  assign n36957 = n31561 ^ n10682 ^ n6624 ;
  assign n36958 = n30873 ^ n4248 ^ x167 ;
  assign n36959 = n36958 ^ n33463 ^ n24163 ;
  assign n36960 = n34567 ^ n33366 ^ x179 ;
  assign n36961 = ( ~n36957 & n36959 ) | ( ~n36957 & n36960 ) | ( n36959 & n36960 ) ;
  assign n36962 = n9372 | n12278 ;
  assign n36963 = n12417 & ~n36962 ;
  assign n36964 = n21053 | n36963 ;
  assign n36965 = n25472 & ~n36964 ;
  assign n36966 = n15481 ^ n9210 ^ 1'b0 ;
  assign n36967 = n36965 | n36966 ;
  assign n36968 = n6126 & n17201 ;
  assign n36969 = n36968 ^ n3239 ^ 1'b0 ;
  assign n36970 = n21441 ^ n17929 ^ n397 ;
  assign n36971 = n36970 ^ n24483 ^ n3097 ;
  assign n36972 = n36971 ^ n6882 ^ n2721 ;
  assign n36973 = n36969 & ~n36972 ;
  assign n36975 = n17913 ^ n16725 ^ 1'b0 ;
  assign n36976 = n7729 | n36975 ;
  assign n36974 = ( ~n14958 & n19771 ) | ( ~n14958 & n24085 ) | ( n19771 & n24085 ) ;
  assign n36977 = n36976 ^ n36974 ^ 1'b0 ;
  assign n36978 = n16322 & ~n19068 ;
  assign n36979 = n5104 & n36978 ;
  assign n36980 = n36979 ^ n13194 ^ n10345 ;
  assign n36981 = ( n542 & n7058 ) | ( n542 & n12089 ) | ( n7058 & n12089 ) ;
  assign n36982 = ~n10626 & n14922 ;
  assign n36983 = n36982 ^ n25031 ^ 1'b0 ;
  assign n36984 = ( n21997 & n36981 ) | ( n21997 & n36983 ) | ( n36981 & n36983 ) ;
  assign n36985 = n36984 ^ n9214 ^ n1608 ;
  assign n36986 = ( n8414 & ~n36100 ) | ( n8414 & n36734 ) | ( ~n36100 & n36734 ) ;
  assign n36987 = n17144 ^ n10731 ^ n1914 ;
  assign n36988 = ( n23784 & ~n27955 ) | ( n23784 & n36987 ) | ( ~n27955 & n36987 ) ;
  assign n36991 = n8395 ^ n5754 ^ 1'b0 ;
  assign n36992 = n2395 | n36991 ;
  assign n36990 = n10607 & ~n24002 ;
  assign n36989 = n18547 ^ n7918 ^ n4409 ;
  assign n36993 = n36992 ^ n36990 ^ n36989 ;
  assign n36994 = ( x223 & ~n24826 ) | ( x223 & n25547 ) | ( ~n24826 & n25547 ) ;
  assign n36995 = n10642 | n27878 ;
  assign n36996 = n36995 ^ n33201 ^ 1'b0 ;
  assign n36997 = n7241 & ~n36996 ;
  assign n36998 = ~n8536 & n36997 ;
  assign n36999 = n25906 ^ n1839 ^ 1'b0 ;
  assign n37000 = n36998 | n36999 ;
  assign n37001 = n9715 ^ n9034 ^ n3239 ;
  assign n37002 = ( n36994 & ~n37000 ) | ( n36994 & n37001 ) | ( ~n37000 & n37001 ) ;
  assign n37007 = ( ~n1068 & n18614 ) | ( ~n1068 & n32816 ) | ( n18614 & n32816 ) ;
  assign n37005 = n29234 ^ n16762 ^ 1'b0 ;
  assign n37006 = ( n3738 & n22682 ) | ( n3738 & ~n37005 ) | ( n22682 & ~n37005 ) ;
  assign n37003 = n21229 ^ n7012 ^ 1'b0 ;
  assign n37004 = n37003 ^ n15534 ^ x148 ;
  assign n37008 = n37007 ^ n37006 ^ n37004 ;
  assign n37009 = n19933 ^ n10316 ^ n10269 ;
  assign n37010 = ( ~n1896 & n35705 ) | ( ~n1896 & n37009 ) | ( n35705 & n37009 ) ;
  assign n37011 = n35762 ^ n30881 ^ n14750 ;
  assign n37012 = n37011 ^ n21851 ^ n15986 ;
  assign n37013 = n17074 ^ n13815 ^ 1'b0 ;
  assign n37014 = n25608 & n37013 ;
  assign n37015 = ( n3588 & ~n16998 ) | ( n3588 & n25499 ) | ( ~n16998 & n25499 ) ;
  assign n37016 = ( n12104 & n37014 ) | ( n12104 & ~n37015 ) | ( n37014 & ~n37015 ) ;
  assign n37017 = n7340 & n7952 ;
  assign n37018 = ( n13823 & n31247 ) | ( n13823 & ~n37017 ) | ( n31247 & ~n37017 ) ;
  assign n37019 = n5183 & ~n37018 ;
  assign n37020 = n37019 ^ n30735 ^ 1'b0 ;
  assign n37021 = n37020 ^ n11808 ^ n11536 ;
  assign n37022 = ( n13175 & n13301 ) | ( n13175 & ~n24607 ) | ( n13301 & ~n24607 ) ;
  assign n37023 = n37022 ^ n18267 ^ 1'b0 ;
  assign n37024 = n35626 ^ n23943 ^ n2200 ;
  assign n37027 = ( n9387 & n23555 ) | ( n9387 & ~n25262 ) | ( n23555 & ~n25262 ) ;
  assign n37025 = n4701 ^ n1857 ^ n1751 ;
  assign n37026 = ( n28020 & n28295 ) | ( n28020 & ~n37025 ) | ( n28295 & ~n37025 ) ;
  assign n37028 = n37027 ^ n37026 ^ n31574 ;
  assign n37029 = ~n37024 & n37028 ;
  assign n37030 = n37029 ^ n22140 ^ n15918 ;
  assign n37031 = ( n1500 & n4618 ) | ( n1500 & ~n5458 ) | ( n4618 & ~n5458 ) ;
  assign n37032 = n37031 ^ n14894 ^ n8426 ;
  assign n37033 = ~n1958 & n6942 ;
  assign n37034 = n37033 ^ n18208 ^ 1'b0 ;
  assign n37035 = ( n16506 & n35620 ) | ( n16506 & ~n37034 ) | ( n35620 & ~n37034 ) ;
  assign n37036 = n37035 ^ n35181 ^ n9061 ;
  assign n37040 = ~n10211 & n20142 ;
  assign n37041 = n6040 & n8539 ;
  assign n37042 = ~n9116 & n37041 ;
  assign n37043 = n37040 | n37042 ;
  assign n37044 = n37043 ^ n18409 ^ 1'b0 ;
  assign n37038 = n26001 ^ n20462 ^ n7770 ;
  assign n37037 = n21201 ^ n8061 ^ n1827 ;
  assign n37039 = n37038 ^ n37037 ^ x141 ;
  assign n37045 = n37044 ^ n37039 ^ n9057 ;
  assign n37047 = n17080 ^ n10881 ^ 1'b0 ;
  assign n37048 = ( ~n3930 & n18906 ) | ( ~n3930 & n37047 ) | ( n18906 & n37047 ) ;
  assign n37046 = n5661 & n7477 ;
  assign n37049 = n37048 ^ n37046 ^ 1'b0 ;
  assign n37050 = n25478 ^ n7832 ^ n2858 ;
  assign n37051 = n37050 ^ n2383 ^ 1'b0 ;
  assign n37052 = ( ~n14156 & n21685 ) | ( ~n14156 & n37051 ) | ( n21685 & n37051 ) ;
  assign n37053 = n9269 | n37052 ;
  assign n37054 = n37053 ^ n22371 ^ 1'b0 ;
  assign n37055 = n12857 ^ n4189 ^ 1'b0 ;
  assign n37056 = n37055 ^ n12394 ^ n10251 ;
  assign n37057 = ( n3069 & ~n30794 ) | ( n3069 & n37056 ) | ( ~n30794 & n37056 ) ;
  assign n37060 = ( ~n9360 & n12898 ) | ( ~n9360 & n14449 ) | ( n12898 & n14449 ) ;
  assign n37058 = n17855 | n28802 ;
  assign n37059 = n37058 ^ n11292 ^ 1'b0 ;
  assign n37061 = n37060 ^ n37059 ^ n28374 ;
  assign n37062 = n9960 & n34840 ;
  assign n37063 = ( ~n4017 & n6339 ) | ( ~n4017 & n17503 ) | ( n6339 & n17503 ) ;
  assign n37064 = n37063 ^ n37047 ^ n26182 ;
  assign n37065 = n26156 | n29479 ;
  assign n37066 = n23191 ^ n2899 ^ n1830 ;
  assign n37069 = n27201 ^ n13509 ^ 1'b0 ;
  assign n37067 = n25185 ^ n2448 ^ 1'b0 ;
  assign n37068 = n4094 & ~n37067 ;
  assign n37070 = n37069 ^ n37068 ^ n19393 ;
  assign n37071 = n17633 & ~n37070 ;
  assign n37072 = n37066 & n37071 ;
  assign n37073 = n538 & ~n29279 ;
  assign n37074 = n9428 & n37073 ;
  assign n37075 = n9566 & ~n13235 ;
  assign n37076 = n37075 ^ n21482 ^ 1'b0 ;
  assign n37077 = ( n3661 & ~n4431 ) | ( n3661 & n19379 ) | ( ~n4431 & n19379 ) ;
  assign n37078 = ( ~n13405 & n37076 ) | ( ~n13405 & n37077 ) | ( n37076 & n37077 ) ;
  assign n37079 = ( n11749 & ~n17537 ) | ( n11749 & n24603 ) | ( ~n17537 & n24603 ) ;
  assign n37080 = n37079 ^ n22528 ^ n5904 ;
  assign n37081 = ( n1747 & n2313 ) | ( n1747 & n5627 ) | ( n2313 & n5627 ) ;
  assign n37082 = ~n31057 & n37081 ;
  assign n37083 = ( n6641 & n26200 ) | ( n6641 & ~n37082 ) | ( n26200 & ~n37082 ) ;
  assign n37084 = ( x100 & n915 ) | ( x100 & n13347 ) | ( n915 & n13347 ) ;
  assign n37085 = n37084 ^ n24030 ^ n7455 ;
  assign n37086 = n37085 ^ n14352 ^ n7979 ;
  assign n37087 = n37086 ^ n23272 ^ n9266 ;
  assign n37088 = n26449 ^ n5721 ^ n3532 ;
  assign n37089 = ( ~n2394 & n13330 ) | ( ~n2394 & n37088 ) | ( n13330 & n37088 ) ;
  assign n37090 = n33997 & ~n37089 ;
  assign n37091 = ~n26149 & n37090 ;
  assign n37092 = ( ~n4209 & n7898 ) | ( ~n4209 & n15713 ) | ( n7898 & n15713 ) ;
  assign n37093 = ( x89 & n20569 ) | ( x89 & ~n21700 ) | ( n20569 & ~n21700 ) ;
  assign n37094 = ~n15960 & n37093 ;
  assign n37095 = ( ~n8681 & n18198 ) | ( ~n8681 & n21563 ) | ( n18198 & n21563 ) ;
  assign n37096 = ( ~n10731 & n17863 ) | ( ~n10731 & n37095 ) | ( n17863 & n37095 ) ;
  assign n37097 = ( n2765 & n22707 ) | ( n2765 & n33289 ) | ( n22707 & n33289 ) ;
  assign n37098 = n32031 ^ n9807 ^ n6400 ;
  assign n37099 = n37098 ^ n14851 ^ 1'b0 ;
  assign n37103 = n3743 & ~n5234 ;
  assign n37104 = n37103 ^ n2352 ^ 1'b0 ;
  assign n37105 = n6364 ^ n4053 ^ n368 ;
  assign n37106 = ( n23670 & n37104 ) | ( n23670 & n37105 ) | ( n37104 & n37105 ) ;
  assign n37107 = ( n29251 & ~n29268 ) | ( n29251 & n37106 ) | ( ~n29268 & n37106 ) ;
  assign n37101 = n18173 ^ n15371 ^ n3975 ;
  assign n37100 = n26930 ^ n17537 ^ n10443 ;
  assign n37102 = n37101 ^ n37100 ^ n24740 ;
  assign n37108 = n37107 ^ n37102 ^ 1'b0 ;
  assign n37109 = ~n30431 & n37108 ;
  assign n37110 = ( n2146 & ~n7521 ) | ( n2146 & n30915 ) | ( ~n7521 & n30915 ) ;
  assign n37111 = ( n10856 & ~n32916 ) | ( n10856 & n37110 ) | ( ~n32916 & n37110 ) ;
  assign n37112 = n29078 ^ n28329 ^ n12632 ;
  assign n37113 = ( n31821 & ~n36162 ) | ( n31821 & n37112 ) | ( ~n36162 & n37112 ) ;
  assign n37114 = ( ~n849 & n3398 ) | ( ~n849 & n6395 ) | ( n3398 & n6395 ) ;
  assign n37115 = n26190 & n37114 ;
  assign n37116 = ( n1245 & n37113 ) | ( n1245 & n37115 ) | ( n37113 & n37115 ) ;
  assign n37118 = ( n4055 & n13609 ) | ( n4055 & ~n27374 ) | ( n13609 & ~n27374 ) ;
  assign n37117 = n16476 | n19425 ;
  assign n37119 = n37118 ^ n37117 ^ n16153 ;
  assign n37120 = n37119 ^ n6194 ^ 1'b0 ;
  assign n37121 = n33926 ^ n30293 ^ n5422 ;
  assign n37122 = n32031 ^ n18283 ^ 1'b0 ;
  assign n37123 = n19090 & n37122 ;
  assign n37124 = n37123 ^ n36358 ^ x118 ;
  assign n37125 = ( ~n9252 & n25294 ) | ( ~n9252 & n29158 ) | ( n25294 & n29158 ) ;
  assign n37126 = n25091 ^ n9832 ^ n5576 ;
  assign n37127 = ( ~n11760 & n18476 ) | ( ~n11760 & n37126 ) | ( n18476 & n37126 ) ;
  assign n37128 = ( n17099 & n33870 ) | ( n17099 & n35051 ) | ( n33870 & n35051 ) ;
  assign n37129 = n24739 ^ n414 ^ 1'b0 ;
  assign n37130 = n29786 ^ n3673 ^ 1'b0 ;
  assign n37131 = n37130 ^ n4424 ^ 1'b0 ;
  assign n37132 = n37131 ^ n27441 ^ 1'b0 ;
  assign n37133 = n37129 | n37132 ;
  assign n37134 = ( n2403 & ~n9292 ) | ( n2403 & n37133 ) | ( ~n9292 & n37133 ) ;
  assign n37135 = n37134 ^ n25979 ^ 1'b0 ;
  assign n37136 = n31664 & ~n37135 ;
  assign n37137 = n3092 & n17371 ;
  assign n37138 = n16652 ^ n14354 ^ 1'b0 ;
  assign n37139 = n37137 | n37138 ;
  assign n37140 = n24294 ^ n7303 ^ n3293 ;
  assign n37141 = ( n2204 & n6031 ) | ( n2204 & n16097 ) | ( n6031 & n16097 ) ;
  assign n37142 = ( n9718 & n37140 ) | ( n9718 & ~n37141 ) | ( n37140 & ~n37141 ) ;
  assign n37143 = n12575 | n13953 ;
  assign n37144 = n37142 & ~n37143 ;
  assign n37145 = ( n11670 & n17591 ) | ( n11670 & n37144 ) | ( n17591 & n37144 ) ;
  assign n37146 = n1093 | n6321 ;
  assign n37147 = n37145 | n37146 ;
  assign n37148 = n22261 ^ n19783 ^ n8969 ;
  assign n37149 = n18008 ^ n11952 ^ n5637 ;
  assign n37150 = ( n18965 & n37148 ) | ( n18965 & n37149 ) | ( n37148 & n37149 ) ;
  assign n37151 = n4458 | n30304 ;
  assign n37152 = n21652 | n37151 ;
  assign n37153 = n16920 ^ n6594 ^ n4839 ;
  assign n37154 = n37153 ^ n27976 ^ n12013 ;
  assign n37155 = ~n25381 & n37154 ;
  assign n37156 = n37155 ^ n13842 ^ 1'b0 ;
  assign n37157 = n16652 & n37156 ;
  assign n37158 = n37157 ^ n21282 ^ 1'b0 ;
  assign n37159 = n31260 ^ n10809 ^ 1'b0 ;
  assign n37160 = n1098 & ~n37159 ;
  assign n37161 = n37160 ^ n16245 ^ 1'b0 ;
  assign n37162 = n13221 ^ n11265 ^ n2934 ;
  assign n37163 = n24582 | n37162 ;
  assign n37164 = n13629 ^ n8821 ^ 1'b0 ;
  assign n37165 = n30109 | n37164 ;
  assign n37166 = ( ~n26801 & n29121 ) | ( ~n26801 & n37165 ) | ( n29121 & n37165 ) ;
  assign n37167 = n5550 ^ n5282 ^ 1'b0 ;
  assign n37168 = ~n11781 & n37167 ;
  assign n37169 = n37168 ^ n19838 ^ 1'b0 ;
  assign n37170 = n14206 & n37169 ;
  assign n37171 = n26370 ^ n23901 ^ n22160 ;
  assign n37175 = ( ~n4010 & n19758 ) | ( ~n4010 & n20122 ) | ( n19758 & n20122 ) ;
  assign n37176 = ( n1528 & n8330 ) | ( n1528 & ~n37175 ) | ( n8330 & ~n37175 ) ;
  assign n37177 = n15643 & ~n37176 ;
  assign n37178 = ~n10535 & n37177 ;
  assign n37172 = n929 | n5665 ;
  assign n37173 = n37172 ^ n27512 ^ 1'b0 ;
  assign n37174 = n37173 ^ n3786 ^ 1'b0 ;
  assign n37179 = n37178 ^ n37174 ^ n15322 ;
  assign n37180 = ( n33626 & ~n37171 ) | ( n33626 & n37179 ) | ( ~n37171 & n37179 ) ;
  assign n37181 = n23466 ^ n7991 ^ n2312 ;
  assign n37182 = ( n7871 & n31740 ) | ( n7871 & ~n37181 ) | ( n31740 & ~n37181 ) ;
  assign n37183 = ( ~n10039 & n28931 ) | ( ~n10039 & n33004 ) | ( n28931 & n33004 ) ;
  assign n37184 = n21890 ^ n10111 ^ 1'b0 ;
  assign n37185 = n2814 | n37184 ;
  assign n37186 = n1318 | n30442 ;
  assign n37187 = n37185 & ~n37186 ;
  assign n37188 = n8410 | n9003 ;
  assign n37189 = n37188 ^ n8219 ^ 1'b0 ;
  assign n37190 = n37189 ^ n9385 ^ 1'b0 ;
  assign n37191 = n14709 | n37190 ;
  assign n37192 = n12387 ^ n11039 ^ 1'b0 ;
  assign n37193 = n16684 ^ n4027 ^ n1173 ;
  assign n37194 = n26773 ^ n21123 ^ 1'b0 ;
  assign n37195 = n29553 ^ n5776 ^ n1275 ;
  assign n37196 = n24568 & ~n37195 ;
  assign n37197 = n2395 ^ n1263 ^ 1'b0 ;
  assign n37198 = n37197 ^ n33158 ^ n7467 ;
  assign n37199 = ( n15258 & n18857 ) | ( n15258 & ~n27035 ) | ( n18857 & ~n27035 ) ;
  assign n37200 = ( n4289 & n32254 ) | ( n4289 & ~n37199 ) | ( n32254 & ~n37199 ) ;
  assign n37207 = n9077 & ~n28599 ;
  assign n37208 = n37207 ^ n16231 ^ 1'b0 ;
  assign n37201 = n14767 ^ n12558 ^ n1092 ;
  assign n37202 = n37201 ^ n23158 ^ n15325 ;
  assign n37203 = ( n20733 & n26237 ) | ( n20733 & ~n37202 ) | ( n26237 & ~n37202 ) ;
  assign n37204 = n20721 ^ n17863 ^ n14314 ;
  assign n37205 = ( n14488 & n37203 ) | ( n14488 & ~n37204 ) | ( n37203 & ~n37204 ) ;
  assign n37206 = n3919 | n37205 ;
  assign n37209 = n37208 ^ n37206 ^ 1'b0 ;
  assign n37210 = n11210 ^ n8606 ^ 1'b0 ;
  assign n37211 = ( n2087 & n7003 ) | ( n2087 & ~n25426 ) | ( n7003 & ~n25426 ) ;
  assign n37212 = ( n17794 & ~n26448 ) | ( n17794 & n37211 ) | ( ~n26448 & n37211 ) ;
  assign n37213 = ( n4824 & n28679 ) | ( n4824 & n37212 ) | ( n28679 & n37212 ) ;
  assign n37214 = n31062 ^ n28775 ^ n26786 ;
  assign n37215 = n26613 ^ n13167 ^ n4536 ;
  assign n37216 = ( n14523 & n31619 ) | ( n14523 & ~n37215 ) | ( n31619 & ~n37215 ) ;
  assign n37217 = n16729 ^ n3265 ^ 1'b0 ;
  assign n37218 = n37216 | n37217 ;
  assign n37219 = n27215 & ~n37218 ;
  assign n37220 = ~n27750 & n37219 ;
  assign n37221 = ~n14668 & n34635 ;
  assign n37222 = n37221 ^ n29622 ^ 1'b0 ;
  assign n37223 = n37222 ^ n23364 ^ 1'b0 ;
  assign n37224 = ( n7587 & ~n30412 ) | ( n7587 & n37223 ) | ( ~n30412 & n37223 ) ;
  assign n37225 = n15594 ^ n12695 ^ n5076 ;
  assign n37226 = ( n13427 & n30321 ) | ( n13427 & n37225 ) | ( n30321 & n37225 ) ;
  assign n37227 = n37226 ^ n25939 ^ n20610 ;
  assign n37228 = n37227 ^ n7594 ^ 1'b0 ;
  assign n37229 = ( ~n10696 & n22443 ) | ( ~n10696 & n36204 ) | ( n22443 & n36204 ) ;
  assign n37230 = n37229 ^ n36504 ^ n24699 ;
  assign n37231 = ( n17070 & ~n17322 ) | ( n17070 & n19881 ) | ( ~n17322 & n19881 ) ;
  assign n37232 = ( n13681 & ~n15540 ) | ( n13681 & n37231 ) | ( ~n15540 & n37231 ) ;
  assign n37233 = n14951 ^ n14879 ^ n4169 ;
  assign n37234 = n2311 & ~n6153 ;
  assign n37235 = ~n37233 & n37234 ;
  assign n37236 = ( n1063 & n12647 ) | ( n1063 & ~n35424 ) | ( n12647 & ~n35424 ) ;
  assign n37237 = n5649 & ~n37236 ;
  assign n37238 = ~n14843 & n37237 ;
  assign n37240 = n24048 ^ n4673 ^ 1'b0 ;
  assign n37241 = n15036 | n37240 ;
  assign n37239 = n32417 ^ n17980 ^ 1'b0 ;
  assign n37242 = n37241 ^ n37239 ^ n1812 ;
  assign n37243 = ( n27311 & ~n37238 ) | ( n27311 & n37242 ) | ( ~n37238 & n37242 ) ;
  assign n37244 = ( n7797 & n26235 ) | ( n7797 & n30083 ) | ( n26235 & n30083 ) ;
  assign n37245 = n23839 ^ n5108 ^ 1'b0 ;
  assign n37246 = ( n7488 & n9072 ) | ( n7488 & n37245 ) | ( n9072 & n37245 ) ;
  assign n37247 = ( n11950 & n37244 ) | ( n11950 & n37246 ) | ( n37244 & n37246 ) ;
  assign n37248 = ( n37235 & n37243 ) | ( n37235 & n37247 ) | ( n37243 & n37247 ) ;
  assign n37249 = ( ~n16280 & n19180 ) | ( ~n16280 & n29439 ) | ( n19180 & n29439 ) ;
  assign n37250 = n3797 | n37249 ;
  assign n37251 = n6265 & ~n37250 ;
  assign n37252 = ( n21009 & ~n25126 ) | ( n21009 & n31002 ) | ( ~n25126 & n31002 ) ;
  assign n37253 = n12634 & n37252 ;
  assign n37254 = ( n10272 & n21691 ) | ( n10272 & ~n26235 ) | ( n21691 & ~n26235 ) ;
  assign n37255 = ( n37251 & n37253 ) | ( n37251 & ~n37254 ) | ( n37253 & ~n37254 ) ;
  assign n37256 = n34365 ^ n12564 ^ n7542 ;
  assign n37257 = ( n887 & n33286 ) | ( n887 & ~n37256 ) | ( n33286 & ~n37256 ) ;
  assign n37258 = n21663 ^ n20350 ^ n1886 ;
  assign n37259 = ( n10222 & ~n12458 ) | ( n10222 & n33292 ) | ( ~n12458 & n33292 ) ;
  assign n37260 = n31531 ^ n4528 ^ n1134 ;
  assign n37261 = n37260 ^ n27626 ^ n16887 ;
  assign n37262 = n7979 ^ n3029 ^ n1162 ;
  assign n37263 = n32913 & n37262 ;
  assign n37264 = n37263 ^ n24649 ^ 1'b0 ;
  assign n37265 = ( ~n5716 & n11464 ) | ( ~n5716 & n37264 ) | ( n11464 & n37264 ) ;
  assign n37266 = ( n4512 & n14956 ) | ( n4512 & ~n37265 ) | ( n14956 & ~n37265 ) ;
  assign n37268 = n14466 ^ n7711 ^ 1'b0 ;
  assign n37269 = n9037 & ~n21444 ;
  assign n37270 = n37268 & n37269 ;
  assign n37267 = n33198 ^ n14273 ^ n3820 ;
  assign n37271 = n37270 ^ n37267 ^ n2823 ;
  assign n37272 = ~n10703 & n36254 ;
  assign n37273 = n19059 ^ n16842 ^ n5183 ;
  assign n37274 = n11647 ^ n1486 ^ 1'b0 ;
  assign n37275 = n37274 ^ n29255 ^ 1'b0 ;
  assign n37276 = n37273 & n37275 ;
  assign n37277 = ~n17664 & n37276 ;
  assign n37278 = ~n10856 & n26359 ;
  assign n37279 = n31858 ^ n22036 ^ n20865 ;
  assign n37280 = ( n6940 & n10956 ) | ( n6940 & n12730 ) | ( n10956 & n12730 ) ;
  assign n37281 = ( n3342 & n6762 ) | ( n3342 & ~n8834 ) | ( n6762 & ~n8834 ) ;
  assign n37282 = ~n8694 & n37281 ;
  assign n37283 = n37282 ^ n5365 ^ 1'b0 ;
  assign n37284 = ( ~n7354 & n18278 ) | ( ~n7354 & n37283 ) | ( n18278 & n37283 ) ;
  assign n37285 = n26829 ^ n25783 ^ 1'b0 ;
  assign n37286 = n29239 ^ n13539 ^ x212 ;
  assign n37287 = ( n6940 & n8646 ) | ( n6940 & n18445 ) | ( n8646 & n18445 ) ;
  assign n37288 = ~n1448 & n8398 ;
  assign n37289 = n37288 ^ n36300 ^ 1'b0 ;
  assign n37290 = n7590 & ~n14264 ;
  assign n37291 = n25439 & n37290 ;
  assign n37292 = ( ~n3014 & n9492 ) | ( ~n3014 & n16142 ) | ( n9492 & n16142 ) ;
  assign n37293 = n37292 ^ n28330 ^ n3971 ;
  assign n37294 = ~n30650 & n37293 ;
  assign n37295 = ~n3670 & n33474 ;
  assign n37296 = n29147 ^ n1032 ^ 1'b0 ;
  assign n37297 = n5407 | n16694 ;
  assign n37298 = n22061 | n37297 ;
  assign n37299 = n37298 ^ n22504 ^ n6981 ;
  assign n37303 = n35589 ^ n28213 ^ n8547 ;
  assign n37300 = n4531 | n33680 ;
  assign n37301 = ( n12585 & n13477 ) | ( n12585 & ~n37300 ) | ( n13477 & ~n37300 ) ;
  assign n37302 = ~n19564 & n37301 ;
  assign n37304 = n37303 ^ n37302 ^ n17488 ;
  assign n37305 = n869 & n8155 ;
  assign n37306 = n37305 ^ n13330 ^ 1'b0 ;
  assign n37307 = n37306 ^ n24027 ^ n8112 ;
  assign n37308 = n37307 ^ n13132 ^ n2404 ;
  assign n37309 = n10041 & ~n37308 ;
  assign n37310 = n37309 ^ n28805 ^ 1'b0 ;
  assign n37311 = n5291 & n6477 ;
  assign n37312 = n37311 ^ n3780 ^ 1'b0 ;
  assign n37313 = n16519 ^ n14832 ^ n10115 ;
  assign n37314 = ( n11536 & n18525 ) | ( n11536 & ~n32668 ) | ( n18525 & ~n32668 ) ;
  assign n37315 = n652 & n22032 ;
  assign n37316 = ( n9011 & ~n17591 ) | ( n9011 & n37315 ) | ( ~n17591 & n37315 ) ;
  assign n37317 = n5358 & n6630 ;
  assign n37318 = n37317 ^ n19961 ^ n6002 ;
  assign n37319 = n14109 ^ n8209 ^ n7503 ;
  assign n37320 = ( n5220 & n37318 ) | ( n5220 & ~n37319 ) | ( n37318 & ~n37319 ) ;
  assign n37321 = n37320 ^ n21966 ^ n15492 ;
  assign n37322 = n37321 ^ n29354 ^ n19530 ;
  assign n37323 = n576 | n5368 ;
  assign n37324 = ( ~n2475 & n10837 ) | ( ~n2475 & n37323 ) | ( n10837 & n37323 ) ;
  assign n37325 = ( ~n6396 & n10049 ) | ( ~n6396 & n21296 ) | ( n10049 & n21296 ) ;
  assign n37326 = ( n21127 & n37324 ) | ( n21127 & n37325 ) | ( n37324 & n37325 ) ;
  assign n37327 = ( n24705 & n31318 ) | ( n24705 & ~n37326 ) | ( n31318 & ~n37326 ) ;
  assign n37328 = n26521 ^ n20019 ^ 1'b0 ;
  assign n37329 = ~n35424 & n37328 ;
  assign n37330 = ( n25294 & n25851 ) | ( n25294 & n37329 ) | ( n25851 & n37329 ) ;
  assign n37331 = n5165 | n22484 ;
  assign n37332 = n30974 | n37331 ;
  assign n37333 = n4614 ^ n4150 ^ 1'b0 ;
  assign n37334 = n5551 | n12172 ;
  assign n37335 = n37333 | n37334 ;
  assign n37336 = n3322 & ~n22796 ;
  assign n37337 = ~n26007 & n37336 ;
  assign n37338 = n11491 & n37337 ;
  assign n37339 = ( n8042 & n37335 ) | ( n8042 & n37338 ) | ( n37335 & n37338 ) ;
  assign n37340 = ( x123 & n1050 ) | ( x123 & ~n3269 ) | ( n1050 & ~n3269 ) ;
  assign n37341 = ( ~n7161 & n24705 ) | ( ~n7161 & n37340 ) | ( n24705 & n37340 ) ;
  assign n37342 = n37341 ^ n5909 ^ 1'b0 ;
  assign n37343 = n24361 ^ n21857 ^ n10193 ;
  assign n37344 = n37343 ^ n15458 ^ n8900 ;
  assign n37345 = n17779 ^ n14193 ^ 1'b0 ;
  assign n37346 = ( n4640 & n13636 ) | ( n4640 & ~n14873 ) | ( n13636 & ~n14873 ) ;
  assign n37347 = ~n18920 & n37346 ;
  assign n37348 = ( ~n7825 & n9260 ) | ( ~n7825 & n24175 ) | ( n9260 & n24175 ) ;
  assign n37349 = ( n3359 & ~n6647 ) | ( n3359 & n24237 ) | ( ~n6647 & n24237 ) ;
  assign n37350 = n37349 ^ n34537 ^ n14543 ;
  assign n37351 = ( n9411 & n32376 ) | ( n9411 & ~n37350 ) | ( n32376 & ~n37350 ) ;
  assign n37353 = n28210 ^ n11588 ^ n5760 ;
  assign n37352 = n9411 | n23027 ;
  assign n37354 = n37353 ^ n37352 ^ 1'b0 ;
  assign n37355 = n4832 ^ n3971 ^ 1'b0 ;
  assign n37356 = x71 & ~n37355 ;
  assign n37357 = n37356 ^ n33843 ^ n19183 ;
  assign n37358 = ( n6103 & n37354 ) | ( n6103 & ~n37357 ) | ( n37354 & ~n37357 ) ;
  assign n37359 = n37351 & ~n37358 ;
  assign n37361 = n17336 & ~n29780 ;
  assign n37362 = ~n9014 & n37361 ;
  assign n37360 = n19200 ^ n3380 ^ 1'b0 ;
  assign n37363 = n37362 ^ n37360 ^ n29890 ;
  assign n37364 = n27378 ^ x247 ^ 1'b0 ;
  assign n37365 = ~n31211 & n37364 ;
  assign n37366 = n29742 ^ n8509 ^ n1030 ;
  assign n37367 = n20079 & ~n23595 ;
  assign n37368 = n33988 ^ n19564 ^ n10683 ;
  assign n37369 = ( n11610 & n37367 ) | ( n11610 & n37368 ) | ( n37367 & n37368 ) ;
  assign n37370 = n37369 ^ n32328 ^ n6958 ;
  assign n37371 = n23185 ^ n13235 ^ n614 ;
  assign n37372 = ( ~n2780 & n7950 ) | ( ~n2780 & n37371 ) | ( n7950 & n37371 ) ;
  assign n37373 = ( n26878 & n33987 ) | ( n26878 & ~n37372 ) | ( n33987 & ~n37372 ) ;
  assign n37374 = n35455 ^ n32210 ^ n27384 ;
  assign n37375 = ( ~n1423 & n10462 ) | ( ~n1423 & n37374 ) | ( n10462 & n37374 ) ;
  assign n37376 = n37375 ^ n36560 ^ n22963 ;
  assign n37377 = n32347 ^ n8653 ^ n3031 ;
  assign n37378 = n26843 ^ n12228 ^ 1'b0 ;
  assign n37379 = n12081 & n37378 ;
  assign n37380 = n23395 ^ n2269 ^ 1'b0 ;
  assign n37381 = n8179 | n37380 ;
  assign n37382 = n37381 ^ n744 ^ n447 ;
  assign n37383 = n19555 & ~n37382 ;
  assign n37384 = ( n1684 & ~n7995 ) | ( n1684 & n17069 ) | ( ~n7995 & n17069 ) ;
  assign n37385 = ( ~n21261 & n24485 ) | ( ~n21261 & n37384 ) | ( n24485 & n37384 ) ;
  assign n37386 = n6746 ^ n5014 ^ x0 ;
  assign n37387 = ~n5271 & n37386 ;
  assign n37388 = n33435 ^ n25253 ^ n1281 ;
  assign n37389 = n37388 ^ n20224 ^ n15499 ;
  assign n37390 = ( ~n4670 & n20086 ) | ( ~n4670 & n37389 ) | ( n20086 & n37389 ) ;
  assign n37391 = n6674 & n37390 ;
  assign n37392 = ~n13117 & n37391 ;
  assign n37393 = n25689 ^ n770 ^ 1'b0 ;
  assign n37394 = ~n16245 & n37393 ;
  assign n37395 = n29711 | n30063 ;
  assign n37396 = n37395 ^ n14749 ^ 1'b0 ;
  assign n37397 = n12378 & ~n37396 ;
  assign n37398 = ~n14106 & n37397 ;
  assign n37399 = n8454 & ~n14484 ;
  assign n37400 = n3505 ^ n1196 ^ 1'b0 ;
  assign n37401 = n800 & n37400 ;
  assign n37402 = ( n260 & ~n6122 ) | ( n260 & n17335 ) | ( ~n6122 & n17335 ) ;
  assign n37403 = ( ~n14978 & n37401 ) | ( ~n14978 & n37402 ) | ( n37401 & n37402 ) ;
  assign n37404 = n37403 ^ n16238 ^ n465 ;
  assign n37406 = n16073 & ~n24745 ;
  assign n37407 = n37406 ^ n23148 ^ n18391 ;
  assign n37405 = n10616 & ~n24483 ;
  assign n37408 = n37407 ^ n37405 ^ 1'b0 ;
  assign n37409 = ~n29602 & n37408 ;
  assign n37410 = n33858 ^ n17606 ^ n15749 ;
  assign n37411 = n33073 ^ n11767 ^ n6723 ;
  assign n37412 = n37411 ^ n33222 ^ n28528 ;
  assign n37413 = n25833 ^ n11032 ^ n5128 ;
  assign n37414 = n17655 & ~n37413 ;
  assign n37415 = n35009 ^ n5389 ^ n1444 ;
  assign n37416 = n37415 ^ n18691 ^ 1'b0 ;
  assign n37417 = n18091 & ~n37416 ;
  assign n37418 = n18324 ^ n10544 ^ n3696 ;
  assign n37419 = n37418 ^ n6421 ^ 1'b0 ;
  assign n37420 = n30465 | n37419 ;
  assign n37421 = ( n6224 & n26667 ) | ( n6224 & ~n37420 ) | ( n26667 & ~n37420 ) ;
  assign n37422 = ( ~n338 & n8389 ) | ( ~n338 & n37421 ) | ( n8389 & n37421 ) ;
  assign n37423 = ( ~n724 & n9295 ) | ( ~n724 & n37422 ) | ( n9295 & n37422 ) ;
  assign n37424 = ( ~n28629 & n29072 ) | ( ~n28629 & n37423 ) | ( n29072 & n37423 ) ;
  assign n37425 = ( n504 & n1174 ) | ( n504 & n20386 ) | ( n1174 & n20386 ) ;
  assign n37426 = ( n6663 & n35742 ) | ( n6663 & ~n37425 ) | ( n35742 & ~n37425 ) ;
  assign n37428 = ~n3624 & n6595 ;
  assign n37429 = n37428 ^ n7951 ^ 1'b0 ;
  assign n37430 = n9531 & ~n19269 ;
  assign n37431 = n37430 ^ n8190 ^ 1'b0 ;
  assign n37432 = n37429 & n37431 ;
  assign n37427 = n27820 ^ n7917 ^ 1'b0 ;
  assign n37433 = n37432 ^ n37427 ^ n8865 ;
  assign n37434 = ( n9075 & n12087 ) | ( n9075 & n37433 ) | ( n12087 & n37433 ) ;
  assign n37435 = n11410 ^ n7837 ^ n2034 ;
  assign n37436 = n37435 ^ n13081 ^ n4814 ;
  assign n37441 = ( n1067 & n1896 ) | ( n1067 & n25377 ) | ( n1896 & n25377 ) ;
  assign n37442 = ( n3563 & n15127 ) | ( n3563 & n37441 ) | ( n15127 & n37441 ) ;
  assign n37437 = ( n12693 & n13108 ) | ( n12693 & n23686 ) | ( n13108 & n23686 ) ;
  assign n37438 = n466 | n12322 ;
  assign n37439 = n37438 ^ n33433 ^ n17632 ;
  assign n37440 = n37437 | n37439 ;
  assign n37443 = n37442 ^ n37440 ^ 1'b0 ;
  assign n37444 = ( n13632 & n23636 ) | ( n13632 & ~n34622 ) | ( n23636 & ~n34622 ) ;
  assign n37445 = ( n30955 & ~n37443 ) | ( n30955 & n37444 ) | ( ~n37443 & n37444 ) ;
  assign n37446 = ( n4412 & ~n22600 ) | ( n4412 & n28280 ) | ( ~n22600 & n28280 ) ;
  assign n37447 = ( n15287 & n25682 ) | ( n15287 & ~n37446 ) | ( n25682 & ~n37446 ) ;
  assign n37448 = n31857 ^ n21715 ^ 1'b0 ;
  assign n37449 = ( n3395 & n13424 ) | ( n3395 & ~n22426 ) | ( n13424 & ~n22426 ) ;
  assign n37450 = ~n14385 & n37449 ;
  assign n37451 = n37450 ^ n10477 ^ 1'b0 ;
  assign n37452 = ( n2800 & n14594 ) | ( n2800 & n37451 ) | ( n14594 & n37451 ) ;
  assign n37455 = n17775 ^ n3383 ^ 1'b0 ;
  assign n37453 = n7178 | n15979 ;
  assign n37454 = n37453 ^ n19123 ^ 1'b0 ;
  assign n37456 = n37455 ^ n37454 ^ n14830 ;
  assign n37457 = n37456 ^ n33049 ^ n4088 ;
  assign n37458 = n28341 ^ n22281 ^ 1'b0 ;
  assign n37459 = n37458 ^ n16817 ^ n16628 ;
  assign n37460 = ( n7337 & n10736 ) | ( n7337 & n30024 ) | ( n10736 & n30024 ) ;
  assign n37461 = n3365 ^ n3063 ^ n1464 ;
  assign n37462 = ( ~n20953 & n37460 ) | ( ~n20953 & n37461 ) | ( n37460 & n37461 ) ;
  assign n37463 = n6876 & ~n37462 ;
  assign n37464 = ( n30703 & n37459 ) | ( n30703 & n37463 ) | ( n37459 & n37463 ) ;
  assign n37465 = ( n1278 & ~n1620 ) | ( n1278 & n14106 ) | ( ~n1620 & n14106 ) ;
  assign n37466 = ( n6721 & ~n10562 ) | ( n6721 & n37465 ) | ( ~n10562 & n37465 ) ;
  assign n37467 = n29756 ^ n16669 ^ n11981 ;
  assign n37468 = ( n6584 & n18946 ) | ( n6584 & ~n37467 ) | ( n18946 & ~n37467 ) ;
  assign n37469 = ( ~n15583 & n37466 ) | ( ~n15583 & n37468 ) | ( n37466 & n37468 ) ;
  assign n37470 = n15929 ^ n14032 ^ 1'b0 ;
  assign n37471 = n25013 & n37470 ;
  assign n37472 = n19939 ^ n12281 ^ n4034 ;
  assign n37473 = n37472 ^ n25026 ^ n22366 ;
  assign n37474 = n36150 ^ n19640 ^ 1'b0 ;
  assign n37475 = n37473 | n37474 ;
  assign n37476 = n32586 ^ n20985 ^ n11461 ;
  assign n37477 = ( n2109 & n2265 ) | ( n2109 & n17731 ) | ( n2265 & n17731 ) ;
  assign n37478 = n29106 & ~n37477 ;
  assign n37479 = n37478 ^ n11251 ^ 1'b0 ;
  assign n37480 = ~n12635 & n12851 ;
  assign n37481 = ( n22566 & n27364 ) | ( n22566 & ~n37480 ) | ( n27364 & ~n37480 ) ;
  assign n37482 = n1114 | n7141 ;
  assign n37483 = ( n4287 & ~n15315 ) | ( n4287 & n36541 ) | ( ~n15315 & n36541 ) ;
  assign n37484 = n5870 | n26769 ;
  assign n37485 = n37484 ^ n23964 ^ 1'b0 ;
  assign n37486 = ( n35857 & ~n37483 ) | ( n35857 & n37485 ) | ( ~n37483 & n37485 ) ;
  assign n37487 = n10147 & ~n14334 ;
  assign n37488 = n37487 ^ n25289 ^ n2303 ;
  assign n37491 = ( n5265 & n9252 ) | ( n5265 & ~n23779 ) | ( n9252 & ~n23779 ) ;
  assign n37489 = n32985 ^ n27343 ^ 1'b0 ;
  assign n37490 = n21046 | n37489 ;
  assign n37492 = n37491 ^ n37490 ^ 1'b0 ;
  assign n37493 = ~n12951 & n14228 ;
  assign n37494 = n3652 | n37493 ;
  assign n37495 = n32677 | n37494 ;
  assign n37498 = n2937 | n21065 ;
  assign n37499 = n19771 & ~n37498 ;
  assign n37500 = ( ~n25888 & n30587 ) | ( ~n25888 & n37499 ) | ( n30587 & n37499 ) ;
  assign n37496 = n31056 ^ n11993 ^ n2721 ;
  assign n37497 = ( n9184 & n13405 ) | ( n9184 & n37496 ) | ( n13405 & n37496 ) ;
  assign n37501 = n37500 ^ n37497 ^ n12249 ;
  assign n37502 = n18189 ^ n1754 ^ 1'b0 ;
  assign n37503 = ( ~n25307 & n35714 ) | ( ~n25307 & n37502 ) | ( n35714 & n37502 ) ;
  assign n37504 = ( n872 & n19526 ) | ( n872 & n23787 ) | ( n19526 & n23787 ) ;
  assign n37505 = ( ~n20276 & n37503 ) | ( ~n20276 & n37504 ) | ( n37503 & n37504 ) ;
  assign n37506 = n16346 ^ n8735 ^ 1'b0 ;
  assign n37507 = n8186 & ~n37506 ;
  assign n37508 = n11461 | n18317 ;
  assign n37509 = ( ~n20594 & n36893 ) | ( ~n20594 & n37508 ) | ( n36893 & n37508 ) ;
  assign n37510 = ( n7571 & n9981 ) | ( n7571 & n25450 ) | ( n9981 & n25450 ) ;
  assign n37511 = ( ~n13853 & n29622 ) | ( ~n13853 & n31887 ) | ( n29622 & n31887 ) ;
  assign n37512 = n37511 ^ n18396 ^ 1'b0 ;
  assign n37513 = n5003 & n37512 ;
  assign n37514 = n37513 ^ n37293 ^ n10763 ;
  assign n37515 = ( n4257 & ~n5180 ) | ( n4257 & n5288 ) | ( ~n5180 & n5288 ) ;
  assign n37516 = n37515 ^ n36521 ^ n13979 ;
  assign n37517 = n7136 & n31309 ;
  assign n37518 = n14220 ^ n4311 ^ n2349 ;
  assign n37519 = n37518 ^ n27042 ^ 1'b0 ;
  assign n37520 = n7431 | n37519 ;
  assign n37521 = n13066 ^ n3480 ^ n439 ;
  assign n37522 = ( n4307 & n11224 ) | ( n4307 & ~n14174 ) | ( n11224 & ~n14174 ) ;
  assign n37523 = ( n14149 & n37521 ) | ( n14149 & n37522 ) | ( n37521 & n37522 ) ;
  assign n37524 = n37523 ^ n31458 ^ 1'b0 ;
  assign n37525 = ~n37520 & n37524 ;
  assign n37526 = n27814 ^ n26141 ^ n8507 ;
  assign n37527 = ( n773 & n4042 ) | ( n773 & ~n9634 ) | ( n4042 & ~n9634 ) ;
  assign n37528 = n1560 & ~n24510 ;
  assign n37529 = ( n3385 & n37527 ) | ( n3385 & ~n37528 ) | ( n37527 & ~n37528 ) ;
  assign n37530 = n37529 ^ n18957 ^ n8429 ;
  assign n37532 = n10170 ^ n7442 ^ 1'b0 ;
  assign n37531 = n34486 ^ n23543 ^ n18936 ;
  assign n37533 = n37532 ^ n37531 ^ n26889 ;
  assign n37534 = n37533 ^ n13844 ^ 1'b0 ;
  assign n37537 = n12564 ^ n6059 ^ n3833 ;
  assign n37538 = n8959 & ~n37537 ;
  assign n37539 = n37538 ^ n25475 ^ 1'b0 ;
  assign n37536 = ( ~n3015 & n9951 ) | ( ~n3015 & n29093 ) | ( n9951 & n29093 ) ;
  assign n37535 = n11106 & n29594 ;
  assign n37540 = n37539 ^ n37536 ^ n37535 ;
  assign n37541 = n35164 ^ n7182 ^ 1'b0 ;
  assign n37542 = n37541 ^ n5985 ^ n529 ;
  assign n37543 = ( n17792 & n36916 ) | ( n17792 & n37542 ) | ( n36916 & n37542 ) ;
  assign n37544 = ( n3241 & n8683 ) | ( n3241 & n37543 ) | ( n8683 & n37543 ) ;
  assign n37545 = ( n2029 & n3796 ) | ( n2029 & ~n4207 ) | ( n3796 & ~n4207 ) ;
  assign n37548 = ( ~n633 & n2462 ) | ( ~n633 & n4731 ) | ( n2462 & n4731 ) ;
  assign n37546 = n12919 | n25073 ;
  assign n37547 = n28720 | n37546 ;
  assign n37549 = n37548 ^ n37547 ^ n7603 ;
  assign n37550 = ( ~n11359 & n37545 ) | ( ~n11359 & n37549 ) | ( n37545 & n37549 ) ;
  assign n37551 = n37550 ^ n15594 ^ n12881 ;
  assign n37553 = n18534 ^ n5674 ^ 1'b0 ;
  assign n37552 = n15943 & ~n32233 ;
  assign n37554 = n37553 ^ n37552 ^ n9041 ;
  assign n37555 = ~n5058 & n11188 ;
  assign n37556 = n12500 ^ n8930 ^ n5189 ;
  assign n37557 = n27815 & ~n37556 ;
  assign n37558 = ( n16122 & n36472 ) | ( n16122 & n37557 ) | ( n36472 & n37557 ) ;
  assign n37559 = n37555 | n37558 ;
  assign n37560 = n37559 ^ n15179 ^ 1'b0 ;
  assign n37561 = n33712 ^ n3904 ^ 1'b0 ;
  assign n37562 = n14918 ^ n12018 ^ n10175 ;
  assign n37563 = n37561 | n37562 ;
  assign n37564 = n37563 ^ n7529 ^ 1'b0 ;
  assign n37566 = n11233 ^ n4071 ^ n1385 ;
  assign n37567 = n37566 ^ n9702 ^ 1'b0 ;
  assign n37568 = n6431 & ~n37567 ;
  assign n37569 = n37568 ^ n2711 ^ 1'b0 ;
  assign n37565 = n23397 ^ n1185 ^ 1'b0 ;
  assign n37570 = n37569 ^ n37565 ^ n3908 ;
  assign n37571 = ( n2423 & n7615 ) | ( n2423 & ~n37570 ) | ( n7615 & ~n37570 ) ;
  assign n37572 = ~n6123 & n17241 ;
  assign n37573 = n7991 & n29148 ;
  assign n37574 = n30142 ^ n7595 ^ 1'b0 ;
  assign n37575 = ~n37573 & n37574 ;
  assign n37576 = ( n2490 & n10002 ) | ( n2490 & ~n20209 ) | ( n10002 & ~n20209 ) ;
  assign n37577 = n29152 ^ n12143 ^ n3791 ;
  assign n37578 = n37577 ^ n36940 ^ 1'b0 ;
  assign n37579 = ( n37575 & n37576 ) | ( n37575 & n37578 ) | ( n37576 & n37578 ) ;
  assign n37580 = ( ~n6287 & n20516 ) | ( ~n6287 & n28493 ) | ( n20516 & n28493 ) ;
  assign n37581 = n27349 ^ n11030 ^ n6099 ;
  assign n37582 = ( ~n18476 & n37580 ) | ( ~n18476 & n37581 ) | ( n37580 & n37581 ) ;
  assign n37583 = n8054 | n23340 ;
  assign n37584 = ~n6029 & n10904 ;
  assign n37585 = n37584 ^ n385 ^ 1'b0 ;
  assign n37587 = ~n6716 & n28164 ;
  assign n37588 = n37587 ^ n11549 ^ 1'b0 ;
  assign n37586 = ( n636 & ~n2233 ) | ( n636 & n26467 ) | ( ~n2233 & n26467 ) ;
  assign n37589 = n37588 ^ n37586 ^ n8581 ;
  assign n37590 = n37589 ^ n32828 ^ n23015 ;
  assign n37591 = ( n9874 & n12728 ) | ( n9874 & ~n23673 ) | ( n12728 & ~n23673 ) ;
  assign n37592 = n19611 ^ n8230 ^ n7262 ;
  assign n37593 = ( n4334 & ~n25474 ) | ( n4334 & n37592 ) | ( ~n25474 & n37592 ) ;
  assign n37594 = n34335 ^ n14261 ^ n2836 ;
  assign n37595 = ( n3248 & n3965 ) | ( n3248 & n37594 ) | ( n3965 & n37594 ) ;
  assign n37596 = n24482 ^ n4920 ^ n3427 ;
  assign n37597 = n37596 ^ n10558 ^ 1'b0 ;
  assign n37598 = ~n37595 & n37597 ;
  assign n37599 = ( n6723 & n6828 ) | ( n6723 & ~n16399 ) | ( n6828 & ~n16399 ) ;
  assign n37600 = n24319 ^ n7331 ^ 1'b0 ;
  assign n37601 = ~n23959 & n37600 ;
  assign n37602 = n37601 ^ n15579 ^ n5048 ;
  assign n37603 = n2148 & ~n3574 ;
  assign n37604 = ( n777 & n16602 ) | ( n777 & ~n37603 ) | ( n16602 & ~n37603 ) ;
  assign n37605 = n9162 ^ n2937 ^ n1075 ;
  assign n37606 = n16178 & n16986 ;
  assign n37607 = n37606 ^ n37169 ^ n20284 ;
  assign n37608 = n12779 | n14466 ;
  assign n37609 = n37608 ^ n3808 ^ 1'b0 ;
  assign n37610 = n37609 ^ n12927 ^ 1'b0 ;
  assign n37611 = n37610 ^ n8076 ^ n1320 ;
  assign n37612 = n4758 & ~n15671 ;
  assign n37613 = ~n37611 & n37612 ;
  assign n37614 = n9771 & n31329 ;
  assign n37615 = n14961 ^ n1482 ^ x41 ;
  assign n37616 = n37615 ^ n32897 ^ n13039 ;
  assign n37617 = ( n12157 & n36895 ) | ( n12157 & n37616 ) | ( n36895 & n37616 ) ;
  assign n37618 = n37617 ^ n26344 ^ n2633 ;
  assign n37619 = ( n10558 & n11565 ) | ( n10558 & ~n34451 ) | ( n11565 & ~n34451 ) ;
  assign n37620 = n37619 ^ n18320 ^ n5167 ;
  assign n37621 = ~n10681 & n12448 ;
  assign n37622 = n37621 ^ n18630 ^ 1'b0 ;
  assign n37623 = ( ~n12873 & n17135 ) | ( ~n12873 & n37622 ) | ( n17135 & n37622 ) ;
  assign n37628 = ( n14644 & n15952 ) | ( n14644 & ~n17087 ) | ( n15952 & ~n17087 ) ;
  assign n37624 = n33139 ^ n12880 ^ n8832 ;
  assign n37625 = n16672 & n37624 ;
  assign n37626 = n24096 & n37625 ;
  assign n37627 = ( n5688 & n7178 ) | ( n5688 & n37626 ) | ( n7178 & n37626 ) ;
  assign n37629 = n37628 ^ n37627 ^ 1'b0 ;
  assign n37630 = n32886 ^ n12125 ^ n4078 ;
  assign n37631 = ( ~n6223 & n25304 ) | ( ~n6223 & n37630 ) | ( n25304 & n37630 ) ;
  assign n37632 = ( n2238 & n37202 ) | ( n2238 & ~n37631 ) | ( n37202 & ~n37631 ) ;
  assign n37633 = ( n19679 & n31716 ) | ( n19679 & ~n32366 ) | ( n31716 & ~n32366 ) ;
  assign n37634 = n1832 & n4538 ;
  assign n37637 = ( n6258 & ~n10768 ) | ( n6258 & n21418 ) | ( ~n10768 & n21418 ) ;
  assign n37638 = n37637 ^ n13424 ^ n3250 ;
  assign n37635 = ( ~n3955 & n6991 ) | ( ~n3955 & n20316 ) | ( n6991 & n20316 ) ;
  assign n37636 = n37635 ^ n18314 ^ n3337 ;
  assign n37639 = n37638 ^ n37636 ^ 1'b0 ;
  assign n37640 = ~n12586 & n37639 ;
  assign n37641 = ~n5566 & n37640 ;
  assign n37642 = n22853 ^ n4100 ^ 1'b0 ;
  assign n37643 = n28721 | n37642 ;
  assign n37644 = n37643 ^ n34806 ^ 1'b0 ;
  assign n37645 = n34990 ^ n17109 ^ n8862 ;
  assign n37646 = ( n473 & n21191 ) | ( n473 & ~n23511 ) | ( n21191 & ~n23511 ) ;
  assign n37647 = ( n13552 & ~n24136 ) | ( n13552 & n34271 ) | ( ~n24136 & n34271 ) ;
  assign n37648 = n37647 ^ n26174 ^ n10158 ;
  assign n37649 = ( n23962 & n37646 ) | ( n23962 & n37648 ) | ( n37646 & n37648 ) ;
  assign n37650 = n16184 ^ n8934 ^ n2800 ;
  assign n37651 = ( n3284 & n10043 ) | ( n3284 & ~n37262 ) | ( n10043 & ~n37262 ) ;
  assign n37652 = ( ~n2151 & n8930 ) | ( ~n2151 & n25942 ) | ( n8930 & n25942 ) ;
  assign n37653 = ~n617 & n28539 ;
  assign n37654 = n37653 ^ n10135 ^ 1'b0 ;
  assign n37655 = n4778 | n19222 ;
  assign n37656 = n33782 ^ n19215 ^ n2799 ;
  assign n37657 = n4117 | n6756 ;
  assign n37658 = n37657 ^ n9907 ^ 1'b0 ;
  assign n37659 = n37658 ^ n19026 ^ n10092 ;
  assign n37660 = ( n2361 & n19342 ) | ( n2361 & ~n21818 ) | ( n19342 & ~n21818 ) ;
  assign n37661 = ( n6988 & n25604 ) | ( n6988 & ~n37660 ) | ( n25604 & ~n37660 ) ;
  assign n37662 = ( n1029 & ~n27283 ) | ( n1029 & n37661 ) | ( ~n27283 & n37661 ) ;
  assign n37663 = ( n19886 & n37659 ) | ( n19886 & n37662 ) | ( n37659 & n37662 ) ;
  assign n37664 = n19783 ^ n14462 ^ n10859 ;
  assign n37665 = ( ~n2493 & n5170 ) | ( ~n2493 & n15833 ) | ( n5170 & n15833 ) ;
  assign n37666 = n6847 ^ n5510 ^ n2148 ;
  assign n37667 = ( ~n20593 & n37665 ) | ( ~n20593 & n37666 ) | ( n37665 & n37666 ) ;
  assign n37668 = ( n28442 & n35922 ) | ( n28442 & n37667 ) | ( n35922 & n37667 ) ;
  assign n37669 = n31704 & ~n37668 ;
  assign n37670 = ~n3357 & n37669 ;
  assign n37671 = ( n2172 & ~n11041 ) | ( n2172 & n37670 ) | ( ~n11041 & n37670 ) ;
  assign n37672 = ( n1344 & n3359 ) | ( n1344 & ~n27684 ) | ( n3359 & ~n27684 ) ;
  assign n37673 = ( n18170 & n21257 ) | ( n18170 & n37672 ) | ( n21257 & n37672 ) ;
  assign n37674 = n17355 | n22430 ;
  assign n37675 = n37674 ^ n3372 ^ 1'b0 ;
  assign n37676 = n37675 ^ n26256 ^ n22029 ;
  assign n37677 = ( n1397 & n9781 ) | ( n1397 & n14861 ) | ( n9781 & n14861 ) ;
  assign n37678 = n37677 ^ n33886 ^ 1'b0 ;
  assign n37679 = n1889 & ~n37678 ;
  assign n37680 = ( n5894 & n8433 ) | ( n5894 & n37679 ) | ( n8433 & n37679 ) ;
  assign n37681 = ( n1156 & ~n30974 ) | ( n1156 & n34080 ) | ( ~n30974 & n34080 ) ;
  assign n37682 = ( n12972 & n25274 ) | ( n12972 & n37681 ) | ( n25274 & n37681 ) ;
  assign n37683 = n5714 ^ n3469 ^ 1'b0 ;
  assign n37684 = ( n16750 & n34796 ) | ( n16750 & ~n37683 ) | ( n34796 & ~n37683 ) ;
  assign n37685 = n37684 ^ n32019 ^ n28781 ;
  assign n37687 = n21601 ^ n5459 ^ n2956 ;
  assign n37686 = n9018 ^ n1414 ^ 1'b0 ;
  assign n37688 = n37687 ^ n37686 ^ n36845 ;
  assign n37689 = n30131 ^ n20232 ^ x100 ;
  assign n37690 = n15790 ^ n4434 ^ 1'b0 ;
  assign n37691 = n9040 & ~n37690 ;
  assign n37692 = n37691 ^ n1810 ^ 1'b0 ;
  assign n37693 = ~n3052 & n37692 ;
  assign n37694 = ( ~n16366 & n37689 ) | ( ~n16366 & n37693 ) | ( n37689 & n37693 ) ;
  assign n37695 = ( n10672 & n31159 ) | ( n10672 & ~n37694 ) | ( n31159 & ~n37694 ) ;
  assign n37696 = n22074 ^ n14273 ^ n13916 ;
  assign n37697 = ~n17657 & n24456 ;
  assign n37698 = n37697 ^ n27472 ^ 1'b0 ;
  assign n37699 = n37698 ^ n16882 ^ n4984 ;
  assign n37700 = ~n845 & n11676 ;
  assign n37701 = n15068 & n37700 ;
  assign n37702 = n33795 ^ n17363 ^ 1'b0 ;
  assign n37703 = n9055 ^ n8155 ^ n2929 ;
  assign n37704 = ( x251 & n2066 ) | ( x251 & n36758 ) | ( n2066 & n36758 ) ;
  assign n37705 = n37704 ^ n17142 ^ n15253 ;
  assign n37706 = ( n3020 & n12235 ) | ( n3020 & ~n37705 ) | ( n12235 & ~n37705 ) ;
  assign n37707 = n33623 ^ n11984 ^ n2688 ;
  assign n37708 = ( ~n18725 & n29482 ) | ( ~n18725 & n37707 ) | ( n29482 & n37707 ) ;
  assign n37709 = n7262 ^ n4191 ^ n1552 ;
  assign n37710 = ( ~n8707 & n17815 ) | ( ~n8707 & n37709 ) | ( n17815 & n37709 ) ;
  assign n37711 = n37710 ^ n25762 ^ n15900 ;
  assign n37712 = ( ~n4625 & n15070 ) | ( ~n4625 & n16493 ) | ( n15070 & n16493 ) ;
  assign n37718 = ( ~n372 & n13735 ) | ( ~n372 & n19750 ) | ( n13735 & n19750 ) ;
  assign n37716 = ( n23157 & n28536 ) | ( n23157 & ~n29299 ) | ( n28536 & ~n29299 ) ;
  assign n37715 = n25486 ^ n16050 ^ n9714 ;
  assign n37717 = n37716 ^ n37715 ^ n24361 ;
  assign n37713 = n15468 ^ n9387 ^ n9278 ;
  assign n37714 = n37713 ^ n28659 ^ n1946 ;
  assign n37719 = n37718 ^ n37717 ^ n37714 ;
  assign n37722 = ( n5853 & n7295 ) | ( n5853 & ~n32160 ) | ( n7295 & ~n32160 ) ;
  assign n37720 = ( n14664 & ~n22758 ) | ( n14664 & n34979 ) | ( ~n22758 & n34979 ) ;
  assign n37721 = n37720 ^ n15860 ^ n1983 ;
  assign n37723 = n37722 ^ n37721 ^ 1'b0 ;
  assign n37724 = ~n19081 & n37723 ;
  assign n37726 = n17235 ^ n12205 ^ 1'b0 ;
  assign n37727 = ~n12474 & n37726 ;
  assign n37725 = n28734 ^ n10124 ^ x242 ;
  assign n37728 = n37727 ^ n37725 ^ n2023 ;
  assign n37729 = n9516 & ~n21521 ;
  assign n37730 = n37729 ^ n35774 ^ n5689 ;
  assign n37731 = n11078 ^ n7262 ^ n5359 ;
  assign n37732 = n2863 ^ n939 ^ 1'b0 ;
  assign n37733 = n37732 ^ n12019 ^ n5377 ;
  assign n37734 = n21271 ^ n21100 ^ n9267 ;
  assign n37735 = ( n2727 & ~n28805 ) | ( n2727 & n37734 ) | ( ~n28805 & n37734 ) ;
  assign n37736 = n11268 ^ n8967 ^ n5081 ;
  assign n37737 = ( n4702 & ~n6080 ) | ( n4702 & n37736 ) | ( ~n6080 & n37736 ) ;
  assign n37738 = n37737 ^ n33096 ^ n8413 ;
  assign n37739 = n21728 ^ n8375 ^ 1'b0 ;
  assign n37740 = n28107 ^ n20688 ^ 1'b0 ;
  assign n37741 = ( n15480 & n16108 ) | ( n15480 & ~n33429 ) | ( n16108 & ~n33429 ) ;
  assign n37742 = n24844 ^ n24080 ^ n5486 ;
  assign n37743 = ( ~n9975 & n28058 ) | ( ~n9975 & n31333 ) | ( n28058 & n31333 ) ;
  assign n37744 = ( n13905 & n20361 ) | ( n13905 & n27542 ) | ( n20361 & n27542 ) ;
  assign n37745 = ( n21533 & n25771 ) | ( n21533 & ~n37744 ) | ( n25771 & ~n37744 ) ;
  assign n37748 = n12518 ^ n6796 ^ 1'b0 ;
  assign n37749 = n1269 | n37748 ;
  assign n37746 = ( n8607 & n14250 ) | ( n8607 & ~n21942 ) | ( n14250 & ~n21942 ) ;
  assign n37747 = n37746 ^ n22374 ^ n887 ;
  assign n37750 = n37749 ^ n37747 ^ n31582 ;
  assign n37751 = n29349 ^ n15917 ^ 1'b0 ;
  assign n37754 = ( ~n5396 & n19132 ) | ( ~n5396 & n27436 ) | ( n19132 & n27436 ) ;
  assign n37755 = n11754 ^ n4429 ^ n537 ;
  assign n37756 = ( ~n15717 & n37754 ) | ( ~n15717 & n37755 ) | ( n37754 & n37755 ) ;
  assign n37757 = n37756 ^ n12622 ^ n10516 ;
  assign n37752 = n14963 | n27617 ;
  assign n37753 = n36425 & ~n37752 ;
  assign n37758 = n37757 ^ n37753 ^ n18905 ;
  assign n37763 = n24644 & n30300 ;
  assign n37764 = n37763 ^ n2680 ^ 1'b0 ;
  assign n37759 = n17387 ^ n708 ^ 1'b0 ;
  assign n37760 = n16524 | n37759 ;
  assign n37761 = n37760 ^ n34339 ^ n894 ;
  assign n37762 = ( ~n1482 & n9381 ) | ( ~n1482 & n37761 ) | ( n9381 & n37761 ) ;
  assign n37765 = n37764 ^ n37762 ^ n23191 ;
  assign n37769 = x225 | n3630 ;
  assign n37770 = ( ~n9036 & n35562 ) | ( ~n9036 & n37769 ) | ( n35562 & n37769 ) ;
  assign n37766 = n14966 ^ n14240 ^ n12994 ;
  assign n37767 = n22058 ^ n6221 ^ 1'b0 ;
  assign n37768 = ( n14854 & ~n37766 ) | ( n14854 & n37767 ) | ( ~n37766 & n37767 ) ;
  assign n37771 = n37770 ^ n37768 ^ n2403 ;
  assign n37772 = n9070 ^ n7316 ^ n6398 ;
  assign n37773 = ~n4109 & n37772 ;
  assign n37774 = ~n6661 & n37773 ;
  assign n37775 = n37774 ^ n27503 ^ n17845 ;
  assign n37776 = n27462 ^ n22504 ^ n15609 ;
  assign n37777 = ( n3689 & ~n35320 ) | ( n3689 & n37776 ) | ( ~n35320 & n37776 ) ;
  assign n37778 = n14007 ^ n4452 ^ 1'b0 ;
  assign n37779 = n37778 ^ n36292 ^ 1'b0 ;
  assign n37780 = n27219 ^ n8459 ^ n5970 ;
  assign n37781 = n15214 ^ n11285 ^ n5962 ;
  assign n37782 = n37781 ^ n22097 ^ n19024 ;
  assign n37783 = n37782 ^ n13317 ^ 1'b0 ;
  assign n37784 = n17245 & ~n37783 ;
  assign n37785 = ~n37780 & n37784 ;
  assign n37786 = ( n2426 & ~n10132 ) | ( n2426 & n18699 ) | ( ~n10132 & n18699 ) ;
  assign n37787 = n6843 & n17562 ;
  assign n37788 = ~n17073 & n37787 ;
  assign n37789 = n37788 ^ n28529 ^ n10666 ;
  assign n37790 = ( n13088 & n14431 ) | ( n13088 & ~n17944 ) | ( n14431 & ~n17944 ) ;
  assign n37791 = n37790 ^ n13364 ^ 1'b0 ;
  assign n37792 = n7055 | n22988 ;
  assign n37793 = n20349 | n37792 ;
  assign n37795 = n33035 ^ n28414 ^ 1'b0 ;
  assign n37796 = n3641 & n37795 ;
  assign n37797 = ( n18241 & ~n28106 ) | ( n18241 & n37796 ) | ( ~n28106 & n37796 ) ;
  assign n37794 = n16230 & n16947 ;
  assign n37798 = n37797 ^ n37794 ^ 1'b0 ;
  assign n37799 = ( n4019 & n37793 ) | ( n4019 & n37798 ) | ( n37793 & n37798 ) ;
  assign n37800 = ( ~n1655 & n13645 ) | ( ~n1655 & n15031 ) | ( n13645 & n15031 ) ;
  assign n37801 = n30639 ^ n19894 ^ 1'b0 ;
  assign n37802 = ( n36218 & n37800 ) | ( n36218 & ~n37801 ) | ( n37800 & ~n37801 ) ;
  assign n37803 = n37802 ^ n28954 ^ 1'b0 ;
  assign n37804 = n8355 ^ n4295 ^ n3181 ;
  assign n37805 = ( n26308 & ~n35761 ) | ( n26308 & n37804 ) | ( ~n35761 & n37804 ) ;
  assign n37806 = n36413 ^ n26464 ^ 1'b0 ;
  assign n37807 = n1312 | n37806 ;
  assign n37808 = n5741 ^ n4762 ^ n557 ;
  assign n37809 = ( ~n16909 & n34254 ) | ( ~n16909 & n37808 ) | ( n34254 & n37808 ) ;
  assign n37810 = n37809 ^ n20762 ^ n13184 ;
  assign n37811 = n37810 ^ n15167 ^ n14007 ;
  assign n37812 = n18534 ^ n10806 ^ n10381 ;
  assign n37813 = n37812 ^ n27551 ^ 1'b0 ;
  assign n37814 = n16829 ^ n13793 ^ n2155 ;
  assign n37815 = ( n905 & ~n15492 ) | ( n905 & n37814 ) | ( ~n15492 & n37814 ) ;
  assign n37817 = n27320 ^ n6302 ^ 1'b0 ;
  assign n37818 = n4579 & ~n37817 ;
  assign n37816 = ( n2393 & ~n5579 ) | ( n2393 & n13406 ) | ( ~n5579 & n13406 ) ;
  assign n37819 = n37818 ^ n37816 ^ n23136 ;
  assign n37820 = n30757 ^ n24278 ^ 1'b0 ;
  assign n37821 = n15219 ^ n12000 ^ n1655 ;
  assign n37822 = ( n24388 & n37820 ) | ( n24388 & ~n37821 ) | ( n37820 & ~n37821 ) ;
  assign n37823 = ( n1276 & ~n17709 ) | ( n1276 & n19675 ) | ( ~n17709 & n19675 ) ;
  assign n37824 = n27662 & n37823 ;
  assign n37825 = n37824 ^ n25903 ^ n5088 ;
  assign n37826 = n9357 ^ n6788 ^ n1098 ;
  assign n37827 = n16956 ^ n13837 ^ 1'b0 ;
  assign n37828 = n26001 & ~n37827 ;
  assign n37829 = n27101 ^ n13731 ^ n356 ;
  assign n37830 = x67 & ~n37829 ;
  assign n37831 = n10390 & n37830 ;
  assign n37832 = n21343 ^ n7126 ^ 1'b0 ;
  assign n37833 = ( n14063 & n19314 ) | ( n14063 & n22369 ) | ( n19314 & n22369 ) ;
  assign n37834 = ( n33811 & ~n37832 ) | ( n33811 & n37833 ) | ( ~n37832 & n37833 ) ;
  assign n37835 = n16163 ^ n6690 ^ n1890 ;
  assign n37836 = n14969 ^ n11269 ^ n4099 ;
  assign n37837 = n37836 ^ n6672 ^ n749 ;
  assign n37838 = n12118 ^ n9185 ^ n4213 ;
  assign n37839 = ( ~n7866 & n26919 ) | ( ~n7866 & n37838 ) | ( n26919 & n37838 ) ;
  assign n37840 = n9758 ^ n7567 ^ n3341 ;
  assign n37841 = ~n21258 & n37840 ;
  assign n37842 = n34254 ^ n33907 ^ n28954 ;
  assign n37843 = n16788 ^ n14026 ^ n9798 ;
  assign n37844 = ( ~n17154 & n21428 ) | ( ~n17154 & n37843 ) | ( n21428 & n37843 ) ;
  assign n37847 = ( n714 & n4914 ) | ( n714 & n5183 ) | ( n4914 & n5183 ) ;
  assign n37845 = n16438 ^ n15848 ^ n6054 ;
  assign n37846 = n37845 ^ n22080 ^ n8998 ;
  assign n37848 = n37847 ^ n37846 ^ n13968 ;
  assign n37849 = ( ~n3348 & n22279 ) | ( ~n3348 & n37848 ) | ( n22279 & n37848 ) ;
  assign n37850 = ~n7145 & n7466 ;
  assign n37851 = ~n15098 & n37850 ;
  assign n37852 = ( n26152 & n30825 ) | ( n26152 & n37851 ) | ( n30825 & n37851 ) ;
  assign n37853 = n29738 ^ n14682 ^ n13192 ;
  assign n37854 = n6090 & n28344 ;
  assign n37855 = n37854 ^ n15263 ^ n8304 ;
  assign n37856 = n15085 & n37855 ;
  assign n37857 = n37856 ^ n34278 ^ n31476 ;
  assign n37858 = n16762 ^ n15689 ^ n561 ;
  assign n37859 = n37858 ^ n22607 ^ 1'b0 ;
  assign n37860 = ( n3336 & n23087 ) | ( n3336 & n37859 ) | ( n23087 & n37859 ) ;
  assign n37861 = n17885 ^ n12031 ^ 1'b0 ;
  assign n37862 = ( n13481 & n14685 ) | ( n13481 & ~n37861 ) | ( n14685 & ~n37861 ) ;
  assign n37864 = n11261 & ~n19553 ;
  assign n37863 = ( n943 & n11046 ) | ( n943 & n33583 ) | ( n11046 & n33583 ) ;
  assign n37865 = n37864 ^ n37863 ^ 1'b0 ;
  assign n37866 = n37862 & n37865 ;
  assign n37867 = n20654 ^ n6224 ^ n889 ;
  assign n37868 = n34529 & n37867 ;
  assign n37869 = ~n6280 & n16221 ;
  assign n37870 = n37869 ^ n14801 ^ 1'b0 ;
  assign n37871 = n37870 ^ n821 ^ 1'b0 ;
  assign n37872 = n20660 | n37871 ;
  assign n37873 = ( n3187 & n17706 ) | ( n3187 & n21010 ) | ( n17706 & n21010 ) ;
  assign n37874 = ~n37872 & n37873 ;
  assign n37875 = ( ~n7230 & n9912 ) | ( ~n7230 & n14214 ) | ( n9912 & n14214 ) ;
  assign n37876 = n19844 ^ n11044 ^ 1'b0 ;
  assign n37877 = n10605 | n37876 ;
  assign n37878 = n37875 & ~n37877 ;
  assign n37879 = n37878 ^ n12191 ^ n270 ;
  assign n37880 = ( n8492 & n23266 ) | ( n8492 & ~n32343 ) | ( n23266 & ~n32343 ) ;
  assign n37881 = ( n10215 & ~n20909 ) | ( n10215 & n37880 ) | ( ~n20909 & n37880 ) ;
  assign n37882 = n10040 ^ n7948 ^ n5136 ;
  assign n37883 = n37882 ^ n11690 ^ n1454 ;
  assign n37884 = n37883 ^ n37004 ^ n32476 ;
  assign n37885 = n9703 & n30685 ;
  assign n37886 = n37885 ^ n9012 ^ 1'b0 ;
  assign n37887 = n32668 | n37886 ;
  assign n37888 = n11888 ^ n11695 ^ x249 ;
  assign n37889 = n24925 & n37888 ;
  assign n37890 = n37889 ^ n3078 ^ 1'b0 ;
  assign n37891 = n37890 ^ n6721 ^ n1945 ;
  assign n37892 = ( ~n337 & n21935 ) | ( ~n337 & n37891 ) | ( n21935 & n37891 ) ;
  assign n37893 = n37892 ^ n19654 ^ n8827 ;
  assign n37895 = ( ~n5777 & n16211 ) | ( ~n5777 & n37323 ) | ( n16211 & n37323 ) ;
  assign n37894 = n31057 ^ n17638 ^ 1'b0 ;
  assign n37896 = n37895 ^ n37894 ^ n2246 ;
  assign n37897 = ( n24543 & ~n30142 ) | ( n24543 & n33620 ) | ( ~n30142 & n33620 ) ;
  assign n37898 = ~n372 & n1600 ;
  assign n37899 = n37898 ^ n13296 ^ 1'b0 ;
  assign n37900 = n37899 ^ n26794 ^ n6937 ;
  assign n37901 = n21264 & n37900 ;
  assign n37902 = ~n3877 & n37901 ;
  assign n37903 = n8487 ^ n4829 ^ 1'b0 ;
  assign n37904 = n32316 | n37903 ;
  assign n37905 = n6460 | n37904 ;
  assign n37906 = n12686 & ~n37905 ;
  assign n37907 = ( ~n4243 & n17438 ) | ( ~n4243 & n19270 ) | ( n17438 & n19270 ) ;
  assign n37908 = ( n13130 & n24202 ) | ( n13130 & n37907 ) | ( n24202 & n37907 ) ;
  assign n37909 = ( n31321 & n33814 ) | ( n31321 & n37908 ) | ( n33814 & n37908 ) ;
  assign n37910 = n1217 & ~n16194 ;
  assign n37911 = n1592 & n37910 ;
  assign n37912 = n11995 ^ n10926 ^ n1780 ;
  assign n37913 = ~n37911 & n37912 ;
  assign n37914 = ~x209 & n37913 ;
  assign n37915 = n35061 ^ n34048 ^ n2216 ;
  assign n37916 = ( ~n9332 & n37914 ) | ( ~n9332 & n37915 ) | ( n37914 & n37915 ) ;
  assign n37917 = n5095 ^ n1749 ^ 1'b0 ;
  assign n37918 = n37917 ^ n22945 ^ n1050 ;
  assign n37919 = ( x93 & n12665 ) | ( x93 & n37918 ) | ( n12665 & n37918 ) ;
  assign n37920 = n32855 ^ n23422 ^ n13591 ;
  assign n37921 = n37920 ^ n10708 ^ 1'b0 ;
  assign n37924 = n1170 ^ n1085 ^ 1'b0 ;
  assign n37923 = n22288 ^ n19129 ^ n2700 ;
  assign n37925 = n37924 ^ n37923 ^ n4497 ;
  assign n37926 = x139 & n37925 ;
  assign n37922 = ~n17700 & n20031 ;
  assign n37927 = n37926 ^ n37922 ^ 1'b0 ;
  assign n37928 = n1422 & ~n1424 ;
  assign n37929 = ~n12492 & n37928 ;
  assign n37930 = n24276 ^ n24088 ^ n10438 ;
  assign n37931 = ( n4556 & n23809 ) | ( n4556 & ~n34612 ) | ( n23809 & ~n34612 ) ;
  assign n37932 = n37930 | n37931 ;
  assign n37933 = n23286 ^ n10822 ^ 1'b0 ;
  assign n37934 = n6597 | n37933 ;
  assign n37935 = n37934 ^ n7909 ^ n5800 ;
  assign n37940 = ( n1787 & n8341 ) | ( n1787 & n19810 ) | ( n8341 & n19810 ) ;
  assign n37941 = ~n27491 & n37940 ;
  assign n37942 = n37941 ^ n3208 ^ 1'b0 ;
  assign n37936 = ~n1928 & n13458 ;
  assign n37937 = n37936 ^ n2863 ^ 1'b0 ;
  assign n37938 = ( ~n324 & n8046 ) | ( ~n324 & n25040 ) | ( n8046 & n25040 ) ;
  assign n37939 = ( n15713 & n37937 ) | ( n15713 & n37938 ) | ( n37937 & n37938 ) ;
  assign n37943 = n37942 ^ n37939 ^ x186 ;
  assign n37944 = n26825 ^ n15767 ^ n7980 ;
  assign n37945 = n23200 ^ n19670 ^ n1919 ;
  assign n37946 = n36188 ^ n11818 ^ n3770 ;
  assign n37947 = n17576 | n37878 ;
  assign n37948 = n37947 ^ n16493 ^ 1'b0 ;
  assign n37949 = ( n12283 & n25158 ) | ( n12283 & n37948 ) | ( n25158 & n37948 ) ;
  assign n37950 = n5199 | n8973 ;
  assign n37951 = n30026 & ~n37950 ;
  assign n37952 = n37951 ^ n31712 ^ n12267 ;
  assign n37953 = n37952 ^ n22428 ^ 1'b0 ;
  assign n37954 = n37953 ^ n10716 ^ n8573 ;
  assign n37955 = n7975 ^ n7505 ^ n6112 ;
  assign n37956 = ( n8470 & ~n10412 ) | ( n8470 & n33692 ) | ( ~n10412 & n33692 ) ;
  assign n37957 = n37956 ^ n33039 ^ n17668 ;
  assign n37958 = ( n22713 & ~n37955 ) | ( n22713 & n37957 ) | ( ~n37955 & n37957 ) ;
  assign n37959 = ~n9475 & n37958 ;
  assign n37960 = n28044 ^ n15644 ^ 1'b0 ;
  assign n37961 = n7130 | n23806 ;
  assign n37962 = n37961 ^ n10339 ^ 1'b0 ;
  assign n37963 = ( n31107 & n32025 ) | ( n31107 & ~n37962 ) | ( n32025 & ~n37962 ) ;
  assign n37964 = n32993 ^ n22635 ^ n1729 ;
  assign n37965 = n37964 ^ n4962 ^ 1'b0 ;
  assign n37966 = ( ~n8028 & n17235 ) | ( ~n8028 & n37965 ) | ( n17235 & n37965 ) ;
  assign n37967 = ~n6431 & n33791 ;
  assign n37968 = n37967 ^ n32156 ^ n16757 ;
  assign n37969 = ~n3405 & n33159 ;
  assign n37970 = ~n25693 & n37969 ;
  assign n37971 = ( n21113 & n24768 ) | ( n21113 & n37970 ) | ( n24768 & n37970 ) ;
  assign n37972 = n28408 ^ n9199 ^ n1891 ;
  assign n37973 = n37972 ^ n31558 ^ n2328 ;
  assign n37974 = ~n37971 & n37973 ;
  assign n37975 = n11186 | n20166 ;
  assign n37976 = n10444 | n37975 ;
  assign n37977 = n22074 ^ n3401 ^ 1'b0 ;
  assign n37978 = ( x110 & n36481 ) | ( x110 & n37977 ) | ( n36481 & n37977 ) ;
  assign n37979 = ( n28673 & n37976 ) | ( n28673 & ~n37978 ) | ( n37976 & ~n37978 ) ;
  assign n37980 = n37979 ^ n29340 ^ n9723 ;
  assign n37981 = n37890 ^ n15392 ^ n5430 ;
  assign n37983 = ( n1233 & n8895 ) | ( n1233 & ~n27991 ) | ( n8895 & ~n27991 ) ;
  assign n37982 = n23695 ^ n23203 ^ 1'b0 ;
  assign n37984 = n37983 ^ n37982 ^ n23781 ;
  assign n37985 = ( ~n12325 & n22565 ) | ( ~n12325 & n29310 ) | ( n22565 & n29310 ) ;
  assign n37986 = n6303 & n19317 ;
  assign n37987 = n37986 ^ n34048 ^ n369 ;
  assign n37988 = n37985 & ~n37987 ;
  assign n37989 = n36629 & n37988 ;
  assign n37990 = n32456 ^ n31520 ^ n4656 ;
  assign n37991 = ( ~n10703 & n17691 ) | ( ~n10703 & n30639 ) | ( n17691 & n30639 ) ;
  assign n37992 = ( n4593 & n17489 ) | ( n4593 & n37991 ) | ( n17489 & n37991 ) ;
  assign n37993 = ( n2135 & n37990 ) | ( n2135 & ~n37992 ) | ( n37990 & ~n37992 ) ;
  assign n37994 = n37993 ^ n15064 ^ 1'b0 ;
  assign n37995 = ~n16693 & n37994 ;
  assign n37996 = ~n24871 & n33256 ;
  assign n37997 = n13942 | n25566 ;
  assign n37998 = n37997 ^ n20272 ^ 1'b0 ;
  assign n37999 = ( n9425 & n28304 ) | ( n9425 & n37998 ) | ( n28304 & n37998 ) ;
  assign n38000 = n9851 ^ n9809 ^ n2210 ;
  assign n38001 = n38000 ^ n27856 ^ n14182 ;
  assign n38002 = n22752 ^ n15404 ^ n11902 ;
  assign n38003 = ( ~n16194 & n38001 ) | ( ~n16194 & n38002 ) | ( n38001 & n38002 ) ;
  assign n38004 = ( ~n19384 & n37999 ) | ( ~n19384 & n38003 ) | ( n37999 & n38003 ) ;
  assign n38005 = ( n1178 & n7124 ) | ( n1178 & n7455 ) | ( n7124 & n7455 ) ;
  assign n38006 = n38005 ^ n30444 ^ n4476 ;
  assign n38007 = n25786 ^ n12547 ^ n1484 ;
  assign n38008 = n38007 ^ n19999 ^ n6470 ;
  assign n38009 = n38008 ^ n13923 ^ n9131 ;
  assign n38010 = n36576 ^ n13471 ^ 1'b0 ;
  assign n38011 = n2613 & n21070 ;
  assign n38012 = n38011 ^ n23929 ^ 1'b0 ;
  assign n38013 = n11004 ^ n1993 ^ 1'b0 ;
  assign n38014 = ~n25228 & n38013 ;
  assign n38015 = ( ~n1833 & n2724 ) | ( ~n1833 & n38014 ) | ( n2724 & n38014 ) ;
  assign n38016 = n5935 ^ n1760 ^ 1'b0 ;
  assign n38017 = n24733 & n38016 ;
  assign n38018 = n38017 ^ n26510 ^ n25700 ;
  assign n38019 = n36118 ^ n19673 ^ n2482 ;
  assign n38020 = n32106 ^ n19978 ^ x119 ;
  assign n38021 = n38020 ^ n5301 ^ 1'b0 ;
  assign n38022 = ( n2954 & n5170 ) | ( n2954 & n7948 ) | ( n5170 & n7948 ) ;
  assign n38023 = n38022 ^ n9596 ^ n1815 ;
  assign n38024 = n29221 & n34812 ;
  assign n38025 = n38023 & n38024 ;
  assign n38026 = ( n28792 & n33557 ) | ( n28792 & ~n38025 ) | ( n33557 & ~n38025 ) ;
  assign n38027 = ( n5100 & n11136 ) | ( n5100 & n30244 ) | ( n11136 & n30244 ) ;
  assign n38028 = ( x234 & ~n4715 ) | ( x234 & n5387 ) | ( ~n4715 & n5387 ) ;
  assign n38029 = ( ~n3454 & n30996 ) | ( ~n3454 & n38028 ) | ( n30996 & n38028 ) ;
  assign n38030 = ( n1840 & n24598 ) | ( n1840 & n35148 ) | ( n24598 & n35148 ) ;
  assign n38031 = ( ~n8683 & n21700 ) | ( ~n8683 & n37140 ) | ( n21700 & n37140 ) ;
  assign n38032 = ( n5347 & n14186 ) | ( n5347 & n38031 ) | ( n14186 & n38031 ) ;
  assign n38033 = n7474 & n38032 ;
  assign n38034 = n38033 ^ n1889 ^ 1'b0 ;
  assign n38035 = n23833 ^ n19313 ^ 1'b0 ;
  assign n38039 = ( n1123 & n2563 ) | ( n1123 & n3278 ) | ( n2563 & n3278 ) ;
  assign n38036 = ( ~n7630 & n16905 ) | ( ~n7630 & n28577 ) | ( n16905 & n28577 ) ;
  assign n38037 = n26142 ^ n6047 ^ 1'b0 ;
  assign n38038 = ~n38036 & n38037 ;
  assign n38040 = n38039 ^ n38038 ^ n26243 ;
  assign n38041 = n38040 ^ n18067 ^ n10350 ;
  assign n38042 = ( ~n441 & n18158 ) | ( ~n441 & n26351 ) | ( n18158 & n26351 ) ;
  assign n38043 = ( ~x76 & n382 ) | ( ~x76 & n38042 ) | ( n382 & n38042 ) ;
  assign n38044 = ( n6804 & ~n18495 ) | ( n6804 & n26575 ) | ( ~n18495 & n26575 ) ;
  assign n38045 = ( n3581 & ~n6622 ) | ( n3581 & n6650 ) | ( ~n6622 & n6650 ) ;
  assign n38046 = n35600 ^ n19867 ^ 1'b0 ;
  assign n38047 = n38046 ^ n22998 ^ 1'b0 ;
  assign n38048 = n14622 ^ n9897 ^ n2709 ;
  assign n38049 = ( n1605 & n12247 ) | ( n1605 & n38048 ) | ( n12247 & n38048 ) ;
  assign n38050 = ( ~n13645 & n18248 ) | ( ~n13645 & n38049 ) | ( n18248 & n38049 ) ;
  assign n38051 = n23340 & ~n38050 ;
  assign n38055 = n11032 ^ n5766 ^ 1'b0 ;
  assign n38056 = n5050 & n38055 ;
  assign n38052 = n31641 ^ n25750 ^ n16525 ;
  assign n38053 = ~n2212 & n11931 ;
  assign n38054 = ~n38052 & n38053 ;
  assign n38057 = n38056 ^ n38054 ^ n2832 ;
  assign n38058 = n13822 ^ n8270 ^ n7572 ;
  assign n38059 = n38058 ^ n4765 ^ n1197 ;
  assign n38060 = ( n5842 & ~n14576 ) | ( n5842 & n34791 ) | ( ~n14576 & n34791 ) ;
  assign n38061 = n22912 ^ n14373 ^ 1'b0 ;
  assign n38062 = ( n4350 & n24039 ) | ( n4350 & n25376 ) | ( n24039 & n25376 ) ;
  assign n38063 = ~n16044 & n19878 ;
  assign n38064 = n1044 & n38063 ;
  assign n38065 = ( ~n1973 & n30696 ) | ( ~n1973 & n36831 ) | ( n30696 & n36831 ) ;
  assign n38066 = n8878 & n17974 ;
  assign n38067 = n37225 ^ n23761 ^ n4793 ;
  assign n38068 = ( ~n4425 & n7101 ) | ( ~n4425 & n11645 ) | ( n7101 & n11645 ) ;
  assign n38069 = ( n10177 & n38067 ) | ( n10177 & n38068 ) | ( n38067 & n38068 ) ;
  assign n38070 = n25626 ^ n3713 ^ 1'b0 ;
  assign n38071 = n11631 & n38070 ;
  assign n38072 = ( n4954 & n5325 ) | ( n4954 & ~n14076 ) | ( n5325 & ~n14076 ) ;
  assign n38073 = ( n24701 & n38071 ) | ( n24701 & ~n38072 ) | ( n38071 & ~n38072 ) ;
  assign n38074 = n19317 ^ n17869 ^ n4770 ;
  assign n38075 = ( n12743 & n14004 ) | ( n12743 & ~n38074 ) | ( n14004 & ~n38074 ) ;
  assign n38077 = n13271 ^ n10925 ^ n1964 ;
  assign n38078 = n20022 | n38077 ;
  assign n38079 = n8150 & ~n38078 ;
  assign n38076 = n32936 ^ n2147 ^ 1'b0 ;
  assign n38080 = n38079 ^ n38076 ^ 1'b0 ;
  assign n38081 = n33978 ^ n30735 ^ n11814 ;
  assign n38082 = n38081 ^ n17551 ^ n6063 ;
  assign n38083 = n38082 ^ n36095 ^ n1328 ;
  assign n38084 = n17863 & n29775 ;
  assign n38085 = n14951 & n38084 ;
  assign n38086 = ( n4745 & ~n5408 ) | ( n4745 & n6649 ) | ( ~n5408 & n6649 ) ;
  assign n38087 = ( ~n3727 & n31190 ) | ( ~n3727 & n31712 ) | ( n31190 & n31712 ) ;
  assign n38088 = n32767 ^ n20049 ^ n11499 ;
  assign n38089 = n26903 & ~n38088 ;
  assign n38090 = n38089 ^ n21957 ^ 1'b0 ;
  assign n38091 = ( n28077 & n38087 ) | ( n28077 & n38090 ) | ( n38087 & n38090 ) ;
  assign n38093 = ( n4396 & n14203 ) | ( n4396 & n17641 ) | ( n14203 & n17641 ) ;
  assign n38092 = n28528 ^ n24853 ^ n15946 ;
  assign n38094 = n38093 ^ n38092 ^ n15767 ;
  assign n38095 = ( n6673 & n32664 ) | ( n6673 & n36876 ) | ( n32664 & n36876 ) ;
  assign n38096 = ( n5170 & n6177 ) | ( n5170 & ~n31491 ) | ( n6177 & ~n31491 ) ;
  assign n38097 = ~n14412 & n33708 ;
  assign n38098 = ~n18389 & n38097 ;
  assign n38099 = ( n11260 & n18318 ) | ( n11260 & ~n24089 ) | ( n18318 & ~n24089 ) ;
  assign n38100 = n38099 ^ n17801 ^ 1'b0 ;
  assign n38101 = n14439 ^ n9525 ^ n1922 ;
  assign n38102 = ( n7051 & n20692 ) | ( n7051 & ~n38101 ) | ( n20692 & ~n38101 ) ;
  assign n38103 = ( n3587 & ~n4876 ) | ( n3587 & n37273 ) | ( ~n4876 & n37273 ) ;
  assign n38104 = ( n25572 & n30250 ) | ( n25572 & n34563 ) | ( n30250 & n34563 ) ;
  assign n38105 = n7189 ^ n1481 ^ 1'b0 ;
  assign n38106 = ~n7869 & n38105 ;
  assign n38107 = n38106 ^ n33555 ^ 1'b0 ;
  assign n38108 = n38107 ^ n7248 ^ n1233 ;
  assign n38109 = n9200 | n14533 ;
  assign n38110 = n7627 | n38109 ;
  assign n38111 = ( n1143 & n3719 ) | ( n1143 & n15347 ) | ( n3719 & n15347 ) ;
  assign n38112 = n19962 & n38111 ;
  assign n38113 = n38112 ^ n19408 ^ 1'b0 ;
  assign n38114 = n38113 ^ n30517 ^ n17282 ;
  assign n38115 = ( n2755 & n38110 ) | ( n2755 & ~n38114 ) | ( n38110 & ~n38114 ) ;
  assign n38116 = n20958 ^ n17679 ^ 1'b0 ;
  assign n38117 = ~n20559 & n20807 ;
  assign n38118 = n38117 ^ n35906 ^ n19337 ;
  assign n38119 = n4549 ^ n4267 ^ 1'b0 ;
  assign n38120 = n5747 & ~n38119 ;
  assign n38121 = n38120 ^ n16419 ^ n13637 ;
  assign n38122 = n37637 ^ n14921 ^ n10563 ;
  assign n38123 = n15533 | n38122 ;
  assign n38124 = n10072 ^ n4403 ^ 1'b0 ;
  assign n38125 = ~n38123 & n38124 ;
  assign n38126 = ( ~n689 & n11692 ) | ( ~n689 & n38125 ) | ( n11692 & n38125 ) ;
  assign n38127 = n27970 ^ n27258 ^ 1'b0 ;
  assign n38128 = ~n2722 & n38127 ;
  assign n38129 = n5432 | n11048 ;
  assign n38130 = n38129 ^ n1306 ^ 1'b0 ;
  assign n38131 = n23950 ^ n6293 ^ 1'b0 ;
  assign n38132 = n3781 | n38131 ;
  assign n38133 = ( n31641 & n38130 ) | ( n31641 & n38132 ) | ( n38130 & n38132 ) ;
  assign n38134 = n35353 ^ n32096 ^ n30366 ;
  assign n38135 = n38134 ^ n32524 ^ n1484 ;
  assign n38136 = n29246 ^ n7371 ^ n1396 ;
  assign n38137 = n31829 ^ n17214 ^ n8610 ;
  assign n38138 = n4741 & ~n15723 ;
  assign n38139 = n637 & n38138 ;
  assign n38140 = ( n8060 & n10168 ) | ( n8060 & n38139 ) | ( n10168 & n38139 ) ;
  assign n38141 = ( ~n318 & n2593 ) | ( ~n318 & n17108 ) | ( n2593 & n17108 ) ;
  assign n38142 = ( n4946 & n24147 ) | ( n4946 & n38141 ) | ( n24147 & n38141 ) ;
  assign n38143 = n23289 ^ n6542 ^ 1'b0 ;
  assign n38144 = ( n8689 & ~n36870 ) | ( n8689 & n38143 ) | ( ~n36870 & n38143 ) ;
  assign n38145 = ( ~n11647 & n14376 ) | ( ~n11647 & n35630 ) | ( n14376 & n35630 ) ;
  assign n38146 = ( n4229 & n34006 ) | ( n4229 & ~n38145 ) | ( n34006 & ~n38145 ) ;
  assign n38147 = ~n15596 & n19145 ;
  assign n38148 = n38147 ^ n26713 ^ 1'b0 ;
  assign n38149 = ( n34504 & ~n36022 ) | ( n34504 & n38148 ) | ( ~n36022 & n38148 ) ;
  assign n38150 = ( n434 & n20066 ) | ( n434 & ~n21557 ) | ( n20066 & ~n21557 ) ;
  assign n38151 = n20129 & n38150 ;
  assign n38152 = ( n1599 & ~n9984 ) | ( n1599 & n19922 ) | ( ~n9984 & n19922 ) ;
  assign n38153 = ( n9198 & n11802 ) | ( n9198 & ~n38152 ) | ( n11802 & ~n38152 ) ;
  assign n38154 = ( ~n6394 & n18298 ) | ( ~n6394 & n38153 ) | ( n18298 & n38153 ) ;
  assign n38155 = n34801 ^ n9608 ^ n5115 ;
  assign n38156 = n19268 ^ n14968 ^ n2815 ;
  assign n38157 = ( n19656 & ~n24302 ) | ( n19656 & n38156 ) | ( ~n24302 & n38156 ) ;
  assign n38158 = n38157 ^ n7970 ^ n1890 ;
  assign n38159 = n35107 ^ n29690 ^ n3990 ;
  assign n38160 = ( n2222 & n4406 ) | ( n2222 & n6662 ) | ( n4406 & n6662 ) ;
  assign n38161 = n38160 ^ n18741 ^ 1'b0 ;
  assign n38162 = n38161 ^ n20911 ^ n2899 ;
  assign n38163 = ( n37684 & n38159 ) | ( n37684 & n38162 ) | ( n38159 & n38162 ) ;
  assign n38164 = n28775 ^ n4742 ^ n788 ;
  assign n38165 = ( n5271 & n9763 ) | ( n5271 & n38164 ) | ( n9763 & n38164 ) ;
  assign n38166 = ( n10226 & n35148 ) | ( n10226 & n37143 ) | ( n35148 & n37143 ) ;
  assign n38167 = n38166 ^ n6929 ^ 1'b0 ;
  assign n38168 = n26713 ^ n18894 ^ n6616 ;
  assign n38169 = n6208 ^ n3480 ^ n2093 ;
  assign n38170 = ~n7869 & n38169 ;
  assign n38171 = n38170 ^ n29724 ^ n23253 ;
  assign n38172 = n22874 ^ n6923 ^ n6789 ;
  assign n38173 = ( ~n12702 & n15287 ) | ( ~n12702 & n32346 ) | ( n15287 & n32346 ) ;
  assign n38174 = n12503 | n38173 ;
  assign n38175 = n19420 ^ n1859 ^ 1'b0 ;
  assign n38176 = n18933 & n38175 ;
  assign n38177 = n2504 & ~n16750 ;
  assign n38178 = n31980 & n38177 ;
  assign n38179 = ( n7888 & n38176 ) | ( n7888 & n38178 ) | ( n38176 & n38178 ) ;
  assign n38180 = n38179 ^ n13388 ^ 1'b0 ;
  assign n38181 = ( n557 & n922 ) | ( n557 & n11825 ) | ( n922 & n11825 ) ;
  assign n38182 = n14455 ^ n11053 ^ n9301 ;
  assign n38183 = n38182 ^ n20201 ^ n14461 ;
  assign n38184 = n38181 & n38183 ;
  assign n38185 = n33009 ^ n12577 ^ n6961 ;
  assign n38186 = n1902 | n7024 ;
  assign n38187 = n38185 | n38186 ;
  assign n38188 = n36043 ^ n31942 ^ n18618 ;
  assign n38189 = ( n16465 & ~n22031 ) | ( n16465 & n38188 ) | ( ~n22031 & n38188 ) ;
  assign n38190 = ~n736 & n27755 ;
  assign n38191 = ( n7466 & n13084 ) | ( n7466 & ~n19417 ) | ( n13084 & ~n19417 ) ;
  assign n38192 = n38191 ^ n8789 ^ n1900 ;
  assign n38193 = n38192 ^ n889 ^ 1'b0 ;
  assign n38194 = ( n3259 & ~n22855 ) | ( n3259 & n25012 ) | ( ~n22855 & n25012 ) ;
  assign n38195 = n18285 ^ n16229 ^ n375 ;
  assign n38196 = ( n1900 & n4908 ) | ( n1900 & n38195 ) | ( n4908 & n38195 ) ;
  assign n38197 = n6102 & ~n27204 ;
  assign n38198 = n38197 ^ n11328 ^ 1'b0 ;
  assign n38199 = ( n27649 & n28880 ) | ( n27649 & ~n38198 ) | ( n28880 & ~n38198 ) ;
  assign n38200 = n21215 | n38199 ;
  assign n38201 = ( n7989 & ~n8854 ) | ( n7989 & n34693 ) | ( ~n8854 & n34693 ) ;
  assign n38202 = n14364 | n15810 ;
  assign n38203 = n6771 | n14465 ;
  assign n38204 = n24228 ^ n6963 ^ 1'b0 ;
  assign n38205 = ~n17696 & n38204 ;
  assign n38206 = ( n19623 & ~n35501 ) | ( n19623 & n38205 ) | ( ~n35501 & n38205 ) ;
  assign n38207 = ( n15987 & n16044 ) | ( n15987 & n27723 ) | ( n16044 & n27723 ) ;
  assign n38208 = n26442 ^ n22603 ^ 1'b0 ;
  assign n38209 = ( n29099 & n35158 ) | ( n29099 & ~n38208 ) | ( n35158 & ~n38208 ) ;
  assign n38213 = n9564 ^ n5297 ^ n2658 ;
  assign n38212 = ( n9382 & n10964 ) | ( n9382 & ~n23136 ) | ( n10964 & ~n23136 ) ;
  assign n38210 = n19965 ^ n14956 ^ n4571 ;
  assign n38211 = n38210 ^ n27766 ^ 1'b0 ;
  assign n38214 = n38213 ^ n38212 ^ n38211 ;
  assign n38215 = ( n8163 & ~n21038 ) | ( n8163 & n38214 ) | ( ~n21038 & n38214 ) ;
  assign n38216 = n38215 ^ n32793 ^ 1'b0 ;
  assign n38217 = ~n27293 & n38216 ;
  assign n38218 = ( ~n20940 & n30454 ) | ( ~n20940 & n33066 ) | ( n30454 & n33066 ) ;
  assign n38219 = n38218 ^ n26249 ^ n4044 ;
  assign n38220 = ( n10763 & n32121 ) | ( n10763 & n38219 ) | ( n32121 & n38219 ) ;
  assign n38221 = ~n17464 & n30565 ;
  assign n38222 = n32968 ^ n3823 ^ 1'b0 ;
  assign n38223 = n7625 ^ n7549 ^ 1'b0 ;
  assign n38224 = n12538 & ~n38223 ;
  assign n38225 = ( n1017 & n3012 ) | ( n1017 & n19150 ) | ( n3012 & n19150 ) ;
  assign n38226 = ( n10094 & n38224 ) | ( n10094 & n38225 ) | ( n38224 & n38225 ) ;
  assign n38227 = n2598 ^ n781 ^ 1'b0 ;
  assign n38228 = ~n38226 & n38227 ;
  assign n38229 = n5953 ^ n2005 ^ 1'b0 ;
  assign n38230 = n36008 & ~n38229 ;
  assign n38231 = n38230 ^ n26529 ^ n7304 ;
  assign n38232 = ( n1353 & ~n6290 ) | ( n1353 & n38231 ) | ( ~n6290 & n38231 ) ;
  assign n38233 = n20152 ^ n12397 ^ n5940 ;
  assign n38234 = n38233 ^ n36291 ^ 1'b0 ;
  assign n38235 = ( n1928 & n12936 ) | ( n1928 & ~n23389 ) | ( n12936 & ~n23389 ) ;
  assign n38236 = n7304 ^ n4910 ^ n3395 ;
  assign n38237 = ~n34306 & n38236 ;
  assign n38238 = n22635 ^ n2108 ^ 1'b0 ;
  assign n38239 = n8339 & ~n19961 ;
  assign n38240 = ( n1618 & n38238 ) | ( n1618 & n38239 ) | ( n38238 & n38239 ) ;
  assign n38241 = n38237 & ~n38240 ;
  assign n38242 = ( n6648 & ~n31162 ) | ( n6648 & n33340 ) | ( ~n31162 & n33340 ) ;
  assign n38243 = ( ~n16328 & n20597 ) | ( ~n16328 & n38242 ) | ( n20597 & n38242 ) ;
  assign n38244 = n38243 ^ n8903 ^ n2938 ;
  assign n38245 = n16948 ^ n4871 ^ n4320 ;
  assign n38246 = n8800 | n10919 ;
  assign n38247 = n38246 ^ n11172 ^ 1'b0 ;
  assign n38248 = ~n14317 & n38247 ;
  assign n38249 = n38245 & n38248 ;
  assign n38250 = ( n4610 & n11446 ) | ( n4610 & ~n21370 ) | ( n11446 & ~n21370 ) ;
  assign n38251 = n7940 ^ n6341 ^ 1'b0 ;
  assign n38252 = n22937 ^ n15887 ^ 1'b0 ;
  assign n38253 = n18492 & n38252 ;
  assign n38254 = n38253 ^ n31739 ^ n6120 ;
  assign n38255 = n38254 ^ n9307 ^ n1978 ;
  assign n38256 = n3936 & n19666 ;
  assign n38257 = ~n33849 & n38256 ;
  assign n38258 = ( n18389 & ~n20919 ) | ( n18389 & n22097 ) | ( ~n20919 & n22097 ) ;
  assign n38259 = ( n4842 & n21979 ) | ( n4842 & ~n23538 ) | ( n21979 & ~n23538 ) ;
  assign n38260 = n20810 ^ n15288 ^ n11767 ;
  assign n38261 = ( n38258 & n38259 ) | ( n38258 & n38260 ) | ( n38259 & n38260 ) ;
  assign n38262 = n38261 ^ n31585 ^ n22963 ;
  assign n38263 = ( n1183 & ~n18910 ) | ( n1183 & n29390 ) | ( ~n18910 & n29390 ) ;
  assign n38264 = n38263 ^ n29948 ^ n24663 ;
  assign n38265 = n38264 ^ n10885 ^ n6134 ;
  assign n38269 = n6178 ^ n3873 ^ n473 ;
  assign n38266 = ~n3612 & n7047 ;
  assign n38267 = n3199 & n38266 ;
  assign n38268 = ( n19813 & ~n26811 ) | ( n19813 & n38267 ) | ( ~n26811 & n38267 ) ;
  assign n38270 = n38269 ^ n38268 ^ n21578 ;
  assign n38271 = ~n25912 & n38270 ;
  assign n38272 = ( n20074 & ~n20973 ) | ( n20074 & n31010 ) | ( ~n20973 & n31010 ) ;
  assign n38273 = ( n9881 & n11987 ) | ( n9881 & ~n16041 ) | ( n11987 & ~n16041 ) ;
  assign n38274 = n38273 ^ n27862 ^ n10070 ;
  assign n38275 = ( x79 & n13004 ) | ( x79 & ~n38274 ) | ( n13004 & ~n38274 ) ;
  assign n38276 = ( n5673 & ~n10548 ) | ( n5673 & n12686 ) | ( ~n10548 & n12686 ) ;
  assign n38277 = n19776 ^ n3702 ^ n1276 ;
  assign n38278 = n8359 & n21719 ;
  assign n38279 = ~n38277 & n38278 ;
  assign n38280 = n27084 & n38279 ;
  assign n38281 = n38280 ^ n11497 ^ 1'b0 ;
  assign n38282 = n32582 | n38281 ;
  assign n38283 = n34682 ^ n14531 ^ n10560 ;
  assign n38284 = ( n9490 & ~n11100 ) | ( n9490 & n38283 ) | ( ~n11100 & n38283 ) ;
  assign n38285 = n18451 ^ n13824 ^ n706 ;
  assign n38286 = ( n4032 & ~n36782 ) | ( n4032 & n38285 ) | ( ~n36782 & n38285 ) ;
  assign n38287 = n4623 & n19930 ;
  assign n38288 = n38287 ^ n8914 ^ 1'b0 ;
  assign n38289 = n38288 ^ n15155 ^ n4987 ;
  assign n38290 = ( n1259 & ~n1439 ) | ( n1259 & n38289 ) | ( ~n1439 & n38289 ) ;
  assign n38291 = ( x104 & ~n1073 ) | ( x104 & n14746 ) | ( ~n1073 & n14746 ) ;
  assign n38292 = ~n4078 & n10068 ;
  assign n38293 = n38292 ^ n19158 ^ n6805 ;
  assign n38294 = n4221 & n27284 ;
  assign n38295 = n38294 ^ n3284 ^ 1'b0 ;
  assign n38296 = n38295 ^ n23815 ^ 1'b0 ;
  assign n38297 = n2142 & n38296 ;
  assign n38300 = x183 & ~n34985 ;
  assign n38301 = n38300 ^ n8071 ^ 1'b0 ;
  assign n38298 = n22701 ^ n2339 ^ 1'b0 ;
  assign n38299 = n3400 | n38298 ;
  assign n38302 = n38301 ^ n38299 ^ 1'b0 ;
  assign n38303 = ( n694 & ~n15833 ) | ( n694 & n28799 ) | ( ~n15833 & n28799 ) ;
  assign n38304 = n4919 ^ n1896 ^ 1'b0 ;
  assign n38305 = ( ~n7995 & n23950 ) | ( ~n7995 & n32795 ) | ( n23950 & n32795 ) ;
  assign n38306 = ( n2240 & n6579 ) | ( n2240 & ~n7023 ) | ( n6579 & ~n7023 ) ;
  assign n38307 = n38306 ^ n23457 ^ x100 ;
  assign n38308 = n14659 | n38307 ;
  assign n38309 = ( n30300 & n38305 ) | ( n30300 & ~n38308 ) | ( n38305 & ~n38308 ) ;
  assign n38310 = ( ~n15790 & n32302 ) | ( ~n15790 & n38309 ) | ( n32302 & n38309 ) ;
  assign n38311 = n21037 ^ n13616 ^ n4586 ;
  assign n38312 = n16495 ^ n15604 ^ 1'b0 ;
  assign n38313 = n15286 & n19476 ;
  assign n38314 = n38313 ^ n21145 ^ 1'b0 ;
  assign n38315 = ( n38311 & n38312 ) | ( n38311 & n38314 ) | ( n38312 & n38314 ) ;
  assign n38316 = n7242 ^ n5862 ^ n1748 ;
  assign n38317 = n38316 ^ n29102 ^ n5591 ;
  assign n38318 = ( n2027 & n17044 ) | ( n2027 & ~n22691 ) | ( n17044 & ~n22691 ) ;
  assign n38319 = n12604 | n29051 ;
  assign n38320 = n29302 | n38319 ;
  assign n38321 = n38320 ^ n29013 ^ 1'b0 ;
  assign n38322 = n38318 & ~n38321 ;
  assign n38323 = ( n8872 & n9140 ) | ( n8872 & ~n15681 ) | ( n9140 & ~n15681 ) ;
  assign n38324 = n38323 ^ n30105 ^ n10811 ;
  assign n38325 = n38324 ^ n20473 ^ 1'b0 ;
  assign n38326 = n4937 & n29519 ;
  assign n38327 = n7921 ^ n941 ^ 1'b0 ;
  assign n38328 = n38327 ^ n37619 ^ n16302 ;
  assign n38329 = n25903 & ~n36790 ;
  assign n38330 = n27879 | n38329 ;
  assign n38331 = n4356 & n18124 ;
  assign n38332 = n38331 ^ n12233 ^ 1'b0 ;
  assign n38333 = ( n2136 & ~n9503 ) | ( n2136 & n15915 ) | ( ~n9503 & n15915 ) ;
  assign n38334 = n14127 | n38333 ;
  assign n38335 = n38334 ^ n31724 ^ 1'b0 ;
  assign n38336 = n24570 ^ n9792 ^ 1'b0 ;
  assign n38337 = ( n6329 & n20316 ) | ( n6329 & n38336 ) | ( n20316 & n38336 ) ;
  assign n38338 = n8982 ^ n7078 ^ n296 ;
  assign n38339 = n38338 ^ n2506 ^ 1'b0 ;
  assign n38340 = n8967 & ~n24101 ;
  assign n38341 = n18963 | n27354 ;
  assign n38342 = n38341 ^ n14140 ^ n5550 ;
  assign n38343 = n38342 ^ n24582 ^ n18716 ;
  assign n38344 = ( ~n12438 & n18952 ) | ( ~n12438 & n31821 ) | ( n18952 & n31821 ) ;
  assign n38345 = n10298 & ~n38344 ;
  assign n38346 = n1257 & n38345 ;
  assign n38347 = ( n16995 & n38343 ) | ( n16995 & ~n38346 ) | ( n38343 & ~n38346 ) ;
  assign n38348 = n13508 ^ n3519 ^ 1'b0 ;
  assign n38349 = n9915 ^ n8585 ^ n6108 ;
  assign n38350 = n38349 ^ n38258 ^ n3789 ;
  assign n38351 = n12423 ^ n6492 ^ 1'b0 ;
  assign n38352 = n9577 & n38351 ;
  assign n38353 = n38350 & n38352 ;
  assign n38354 = n34319 ^ n11978 ^ n1454 ;
  assign n38355 = n4025 | n34964 ;
  assign n38356 = n1571 & ~n38355 ;
  assign n38357 = ( n19877 & ~n29012 ) | ( n19877 & n38356 ) | ( ~n29012 & n38356 ) ;
  assign n38358 = n22327 ^ n3298 ^ 1'b0 ;
  assign n38359 = ( n7212 & ~n7991 ) | ( n7212 & n38358 ) | ( ~n7991 & n38358 ) ;
  assign n38360 = ( n2100 & n6130 ) | ( n2100 & n10853 ) | ( n6130 & n10853 ) ;
  assign n38361 = ( ~n3966 & n4806 ) | ( ~n3966 & n38360 ) | ( n4806 & n38360 ) ;
  assign n38362 = ( n11176 & n31283 ) | ( n11176 & n38361 ) | ( n31283 & n38361 ) ;
  assign n38363 = n5493 ^ n2112 ^ 1'b0 ;
  assign n38364 = n8820 | n38363 ;
  assign n38365 = n16454 ^ n16374 ^ 1'b0 ;
  assign n38366 = n9841 & ~n38365 ;
  assign n38367 = n27866 & n38366 ;
  assign n38368 = n30691 & n38367 ;
  assign n38369 = n29813 ^ n10537 ^ n8407 ;
  assign n38370 = n38369 ^ n33291 ^ n16813 ;
  assign n38371 = n30125 ^ n5861 ^ n1920 ;
  assign n38372 = n38370 & n38371 ;
  assign n38373 = ~n32968 & n38372 ;
  assign n38374 = n7485 & n14448 ;
  assign n38375 = n38374 ^ n995 ^ 1'b0 ;
  assign n38376 = n38375 ^ n25672 ^ n20274 ;
  assign n38377 = ( x186 & ~n11434 ) | ( x186 & n19771 ) | ( ~n11434 & n19771 ) ;
  assign n38378 = n38377 ^ n25804 ^ n8014 ;
  assign n38379 = ( n17764 & ~n27503 ) | ( n17764 & n38378 ) | ( ~n27503 & n38378 ) ;
  assign n38380 = ( ~n14468 & n22040 ) | ( ~n14468 & n35228 ) | ( n22040 & n35228 ) ;
  assign n38381 = n38380 ^ n12693 ^ 1'b0 ;
  assign n38382 = n707 | n7979 ;
  assign n38383 = n38382 ^ n11230 ^ 1'b0 ;
  assign n38384 = n38383 ^ n17494 ^ n13191 ;
  assign n38385 = ( n784 & n4018 ) | ( n784 & ~n6249 ) | ( n4018 & ~n6249 ) ;
  assign n38386 = ( n8760 & n11462 ) | ( n8760 & ~n38385 ) | ( n11462 & ~n38385 ) ;
  assign n38387 = ( n2267 & n24259 ) | ( n2267 & n38386 ) | ( n24259 & n38386 ) ;
  assign n38388 = n13014 | n38387 ;
  assign n38389 = n36425 ^ n10031 ^ n4202 ;
  assign n38391 = n31620 ^ n9348 ^ n1875 ;
  assign n38390 = n36407 ^ n31880 ^ n7962 ;
  assign n38392 = n38391 ^ n38390 ^ n16204 ;
  assign n38393 = ( n6058 & n9568 ) | ( n6058 & ~n17794 ) | ( n9568 & ~n17794 ) ;
  assign n38394 = n34339 ^ n29080 ^ n17979 ;
  assign n38395 = ( n30645 & n38393 ) | ( n30645 & n38394 ) | ( n38393 & n38394 ) ;
  assign n38396 = n38077 ^ n34611 ^ n7403 ;
  assign n38397 = ( n13349 & ~n25796 ) | ( n13349 & n26243 ) | ( ~n25796 & n26243 ) ;
  assign n38398 = n7842 | n38397 ;
  assign n38399 = n38396 | n38398 ;
  assign n38401 = n15432 ^ n8019 ^ n4298 ;
  assign n38402 = n26008 ^ n12283 ^ n8549 ;
  assign n38403 = n38402 ^ n26265 ^ n13561 ;
  assign n38404 = n38401 & n38403 ;
  assign n38405 = n9221 & n38404 ;
  assign n38400 = ~n6609 & n36555 ;
  assign n38406 = n38405 ^ n38400 ^ 1'b0 ;
  assign n38407 = ( n1476 & n4245 ) | ( n1476 & n17965 ) | ( n4245 & n17965 ) ;
  assign n38408 = n5015 | n38407 ;
  assign n38409 = ( n2651 & ~n9248 ) | ( n2651 & n22974 ) | ( ~n9248 & n22974 ) ;
  assign n38417 = n12247 ^ n8699 ^ n2484 ;
  assign n38416 = n2680 & n13481 ;
  assign n38418 = n38417 ^ n38416 ^ n18026 ;
  assign n38411 = n20658 ^ n7065 ^ n1899 ;
  assign n38410 = ~n1501 & n33936 ;
  assign n38412 = n38411 ^ n38410 ^ 1'b0 ;
  assign n38413 = ~n799 & n38412 ;
  assign n38414 = n33478 | n38413 ;
  assign n38415 = n23234 | n38414 ;
  assign n38419 = n38418 ^ n38415 ^ n1336 ;
  assign n38420 = n32913 ^ n7411 ^ n977 ;
  assign n38421 = ~n37987 & n38420 ;
  assign n38422 = n21711 ^ n5933 ^ n4547 ;
  assign n38423 = n38422 ^ n12794 ^ 1'b0 ;
  assign n38424 = n16686 | n38423 ;
  assign n38425 = ( n18746 & n20443 ) | ( n18746 & ~n38424 ) | ( n20443 & ~n38424 ) ;
  assign n38426 = n7787 ^ n1647 ^ n701 ;
  assign n38427 = ( n8188 & n15840 ) | ( n8188 & n38426 ) | ( n15840 & n38426 ) ;
  assign n38428 = ( n3689 & n17987 ) | ( n3689 & n38427 ) | ( n17987 & n38427 ) ;
  assign n38429 = n10028 ^ n8679 ^ n5527 ;
  assign n38430 = n6447 ^ n1208 ^ 1'b0 ;
  assign n38431 = n11983 | n38430 ;
  assign n38432 = n8821 & ~n38431 ;
  assign n38433 = ~n38429 & n38432 ;
  assign n38434 = n30848 ^ n26229 ^ n23628 ;
  assign n38435 = n38434 ^ n19061 ^ 1'b0 ;
  assign n38438 = ( n23037 & n27796 ) | ( n23037 & ~n31871 ) | ( n27796 & ~n31871 ) ;
  assign n38436 = n2026 & n7230 ;
  assign n38437 = n2838 & ~n38436 ;
  assign n38439 = n38438 ^ n38437 ^ 1'b0 ;
  assign n38440 = n38439 ^ n29467 ^ n17340 ;
  assign n38441 = n2484 & ~n12092 ;
  assign n38442 = n5108 ^ n4034 ^ n346 ;
  assign n38443 = ( n7265 & n20507 ) | ( n7265 & n38442 ) | ( n20507 & n38442 ) ;
  assign n38444 = n24670 ^ n18952 ^ n9454 ;
  assign n38445 = n38444 ^ n14149 ^ n10125 ;
  assign n38446 = ( n38210 & n38443 ) | ( n38210 & n38445 ) | ( n38443 & n38445 ) ;
  assign n38447 = n23365 ^ n9898 ^ n7487 ;
  assign n38448 = n37304 ^ n26501 ^ n22701 ;
  assign n38449 = n31555 ^ n8261 ^ n305 ;
  assign n38450 = n27294 ^ n9848 ^ n941 ;
  assign n38451 = n12565 ^ n10372 ^ n4241 ;
  assign n38452 = ( n16374 & n38450 ) | ( n16374 & n38451 ) | ( n38450 & n38451 ) ;
  assign n38453 = n7039 & n23558 ;
  assign n38454 = n7667 & n38453 ;
  assign n38455 = n14791 ^ n9486 ^ 1'b0 ;
  assign n38456 = n27055 | n38455 ;
  assign n38457 = ( n15242 & n26913 ) | ( n15242 & n33897 ) | ( n26913 & n33897 ) ;
  assign n38458 = n7969 & n32775 ;
  assign n38459 = ~n38457 & n38458 ;
  assign n38460 = ~n9230 & n36620 ;
  assign n38461 = n25448 & n38460 ;
  assign n38462 = ( ~n7366 & n24777 ) | ( ~n7366 & n38461 ) | ( n24777 & n38461 ) ;
  assign n38463 = ( n1800 & n4714 ) | ( n1800 & n38462 ) | ( n4714 & n38462 ) ;
  assign n38464 = ( n22807 & n28320 ) | ( n22807 & n38463 ) | ( n28320 & n38463 ) ;
  assign n38465 = n20186 ^ n18891 ^ n17684 ;
  assign n38466 = n26722 ^ n16693 ^ 1'b0 ;
  assign n38467 = ( ~n19998 & n38465 ) | ( ~n19998 & n38466 ) | ( n38465 & n38466 ) ;
  assign n38469 = n9315 ^ n2472 ^ n783 ;
  assign n38468 = n30639 ^ n16895 ^ n8295 ;
  assign n38470 = n38469 ^ n38468 ^ n15809 ;
  assign n38471 = n3630 | n7244 ;
  assign n38472 = n2165 & ~n38471 ;
  assign n38473 = ( n1331 & n16623 ) | ( n1331 & n38472 ) | ( n16623 & n38472 ) ;
  assign n38474 = n18397 ^ n3614 ^ 1'b0 ;
  assign n38475 = ( n38470 & ~n38473 ) | ( n38470 & n38474 ) | ( ~n38473 & n38474 ) ;
  assign n38476 = ( n12960 & n23964 ) | ( n12960 & ~n37298 ) | ( n23964 & ~n37298 ) ;
  assign n38477 = ~n4598 & n7180 ;
  assign n38478 = n12699 | n38477 ;
  assign n38479 = n29257 ^ n14564 ^ 1'b0 ;
  assign n38480 = ~n25298 & n38479 ;
  assign n38481 = ( n394 & n14038 ) | ( n394 & ~n14221 ) | ( n14038 & ~n14221 ) ;
  assign n38482 = n38481 ^ n11907 ^ 1'b0 ;
  assign n38483 = n14175 ^ n13995 ^ n1787 ;
  assign n38484 = n38483 ^ n9524 ^ n8434 ;
  assign n38485 = n38484 ^ n2757 ^ n1156 ;
  assign n38486 = n31135 ^ n5985 ^ 1'b0 ;
  assign n38487 = ( n8340 & n22819 ) | ( n8340 & n37717 ) | ( n22819 & n37717 ) ;
  assign n38488 = n2533 ^ n992 ^ 1'b0 ;
  assign n38489 = n38488 ^ n37687 ^ n37354 ;
  assign n38490 = ~n2903 & n17410 ;
  assign n38491 = ~n23365 & n38490 ;
  assign n38492 = n28357 ^ n8135 ^ n6388 ;
  assign n38493 = ( x182 & ~n25419 ) | ( x182 & n38492 ) | ( ~n25419 & n38492 ) ;
  assign n38495 = ( n13741 & n20202 ) | ( n13741 & ~n26974 ) | ( n20202 & ~n26974 ) ;
  assign n38494 = ( n10797 & ~n15280 ) | ( n10797 & n29517 ) | ( ~n15280 & n29517 ) ;
  assign n38496 = n38495 ^ n38494 ^ n17448 ;
  assign n38497 = n23538 ^ n9229 ^ 1'b0 ;
  assign n38498 = ( n13663 & n16010 ) | ( n13663 & ~n38497 ) | ( n16010 & ~n38497 ) ;
  assign n38499 = n16003 ^ n3320 ^ n3041 ;
  assign n38500 = ( n19835 & n35677 ) | ( n19835 & ~n38499 ) | ( n35677 & ~n38499 ) ;
  assign n38501 = ~n2046 & n38500 ;
  assign n38502 = ( x152 & n5445 ) | ( x152 & n22654 ) | ( n5445 & n22654 ) ;
  assign n38503 = ~n8918 & n38502 ;
  assign n38504 = n38503 ^ n21806 ^ 1'b0 ;
  assign n38506 = n18837 ^ n13995 ^ n12266 ;
  assign n38505 = n4759 & ~n7683 ;
  assign n38507 = n38506 ^ n38505 ^ n10251 ;
  assign n38508 = n37140 ^ n23102 ^ 1'b0 ;
  assign n38509 = n11666 ^ n4247 ^ 1'b0 ;
  assign n38513 = ~n3992 & n21856 ;
  assign n38514 = ( n5357 & n13677 ) | ( n5357 & ~n38513 ) | ( n13677 & ~n38513 ) ;
  assign n38510 = n25900 ^ n3353 ^ 1'b0 ;
  assign n38511 = ( ~n10981 & n29381 ) | ( ~n10981 & n38510 ) | ( n29381 & n38510 ) ;
  assign n38512 = n38511 ^ n25370 ^ n10221 ;
  assign n38515 = n38514 ^ n38512 ^ n6809 ;
  assign n38516 = ( n13043 & ~n16500 ) | ( n13043 & n33196 ) | ( ~n16500 & n33196 ) ;
  assign n38517 = n19492 & ~n38516 ;
  assign n38518 = n38517 ^ n17810 ^ n9397 ;
  assign n38519 = n32744 ^ n13430 ^ n3071 ;
  assign n38520 = ( n33728 & n38518 ) | ( n33728 & ~n38519 ) | ( n38518 & ~n38519 ) ;
  assign n38521 = n38520 ^ n32244 ^ n27857 ;
  assign n38522 = n30012 ^ n25144 ^ 1'b0 ;
  assign n38523 = n29316 & ~n38522 ;
  assign n38526 = n23241 ^ n11936 ^ n2202 ;
  assign n38527 = n38526 ^ n27928 ^ n12152 ;
  assign n38528 = ~n11453 & n38527 ;
  assign n38524 = ( n3321 & ~n22983 ) | ( n3321 & n30443 ) | ( ~n22983 & n30443 ) ;
  assign n38525 = ~n10430 & n38524 ;
  assign n38529 = n38528 ^ n38525 ^ 1'b0 ;
  assign n38530 = ( n3526 & n7063 ) | ( n3526 & ~n24767 ) | ( n7063 & ~n24767 ) ;
  assign n38531 = ( n6024 & ~n18409 ) | ( n6024 & n36485 ) | ( ~n18409 & n36485 ) ;
  assign n38532 = ( n20006 & n38530 ) | ( n20006 & n38531 ) | ( n38530 & n38531 ) ;
  assign n38535 = ( n5267 & n9286 ) | ( n5267 & n14421 ) | ( n9286 & n14421 ) ;
  assign n38533 = ( n535 & n7073 ) | ( n535 & ~n13226 ) | ( n7073 & ~n13226 ) ;
  assign n38534 = n38533 ^ n18258 ^ n7262 ;
  assign n38536 = n38535 ^ n38534 ^ n1972 ;
  assign n38537 = n8090 & n18453 ;
  assign n38538 = ~n6836 & n38537 ;
  assign n38539 = ( n27595 & ~n32249 ) | ( n27595 & n38538 ) | ( ~n32249 & n38538 ) ;
  assign n38540 = n38539 ^ n12334 ^ n7892 ;
  assign n38546 = n6119 ^ n3609 ^ n409 ;
  assign n38547 = n38546 ^ n12857 ^ n3823 ;
  assign n38543 = ( n340 & ~n1460 ) | ( n340 & n28905 ) | ( ~n1460 & n28905 ) ;
  assign n38544 = n38543 ^ n32385 ^ n24276 ;
  assign n38541 = n22959 ^ n10846 ^ 1'b0 ;
  assign n38542 = n5719 & ~n38541 ;
  assign n38545 = n38544 ^ n38542 ^ n13188 ;
  assign n38548 = n38547 ^ n38545 ^ 1'b0 ;
  assign n38549 = n5877 & ~n23557 ;
  assign n38550 = ~n28229 & n38549 ;
  assign n38551 = n38550 ^ n38244 ^ n20053 ;
  assign n38552 = ~n12516 & n24080 ;
  assign n38553 = ~n13328 & n38552 ;
  assign n38554 = n38553 ^ n21083 ^ 1'b0 ;
  assign n38555 = n4825 ^ n1499 ^ 1'b0 ;
  assign n38556 = n38554 & ~n38555 ;
  assign n38560 = ( n5049 & n12079 ) | ( n5049 & ~n16311 ) | ( n12079 & ~n16311 ) ;
  assign n38558 = n22598 ^ n17276 ^ 1'b0 ;
  assign n38559 = n20491 & ~n38558 ;
  assign n38557 = ( n13979 & ~n34351 ) | ( n13979 & n38288 ) | ( ~n34351 & n38288 ) ;
  assign n38561 = n38560 ^ n38559 ^ n38557 ;
  assign n38562 = n34431 | n38561 ;
  assign n38563 = n20638 | n38562 ;
  assign n38564 = n13823 | n37052 ;
  assign n38565 = n36647 & ~n38564 ;
  assign n38566 = n38563 & n38565 ;
  assign n38567 = n38566 ^ n29712 ^ n3029 ;
  assign n38568 = ( n3095 & ~n5477 ) | ( n3095 & n10829 ) | ( ~n5477 & n10829 ) ;
  assign n38569 = n38568 ^ n35568 ^ n5270 ;
  assign n38570 = ( ~n2519 & n10184 ) | ( ~n2519 & n30471 ) | ( n10184 & n30471 ) ;
  assign n38571 = n25755 ^ n22566 ^ 1'b0 ;
  assign n38572 = n18162 ^ n12027 ^ n10668 ;
  assign n38573 = n38572 ^ n32546 ^ n990 ;
  assign n38574 = ( n16807 & n19205 ) | ( n16807 & ~n34182 ) | ( n19205 & ~n34182 ) ;
  assign n38575 = ( n7029 & n19714 ) | ( n7029 & ~n29607 ) | ( n19714 & ~n29607 ) ;
  assign n38576 = ( n4458 & n13297 ) | ( n4458 & n19344 ) | ( n13297 & n19344 ) ;
  assign n38577 = ( n8479 & n10259 ) | ( n8479 & n27258 ) | ( n10259 & n27258 ) ;
  assign n38579 = ( n3400 & n10049 ) | ( n3400 & n17555 ) | ( n10049 & n17555 ) ;
  assign n38580 = n10502 ^ n5257 ^ 1'b0 ;
  assign n38581 = ~n38579 & n38580 ;
  assign n38578 = ( n6134 & ~n8958 ) | ( n6134 & n9897 ) | ( ~n8958 & n9897 ) ;
  assign n38582 = n38581 ^ n38578 ^ n528 ;
  assign n38583 = ( n7105 & n10036 ) | ( n7105 & n16450 ) | ( n10036 & n16450 ) ;
  assign n38584 = n38583 ^ n20078 ^ n14121 ;
  assign n38585 = ( n17803 & n22642 ) | ( n17803 & ~n38584 ) | ( n22642 & ~n38584 ) ;
  assign n38586 = n31806 ^ n17247 ^ n14988 ;
  assign n38587 = n16187 | n38586 ;
  assign n38590 = ( ~n833 & n2565 ) | ( ~n833 & n4028 ) | ( n2565 & n4028 ) ;
  assign n38591 = ( ~n2396 & n10728 ) | ( ~n2396 & n38590 ) | ( n10728 & n38590 ) ;
  assign n38588 = n12808 ^ n9297 ^ n2782 ;
  assign n38589 = n732 | n38588 ;
  assign n38592 = n38591 ^ n38589 ^ 1'b0 ;
  assign n38593 = n14117 ^ n7055 ^ n4213 ;
  assign n38594 = n38593 ^ n18308 ^ n9557 ;
  assign n38595 = n24311 | n38594 ;
  assign n38596 = n28865 & ~n38595 ;
  assign n38597 = ( n994 & ~n4856 ) | ( n994 & n5964 ) | ( ~n4856 & n5964 ) ;
  assign n38598 = n38597 ^ n9642 ^ n5694 ;
  assign n38599 = n25185 ^ n15742 ^ n7951 ;
  assign n38600 = n16053 ^ n8794 ^ n5203 ;
  assign n38601 = n38600 ^ n9174 ^ n3783 ;
  assign n38602 = ~n11486 & n16706 ;
  assign n38603 = n38602 ^ n424 ^ 1'b0 ;
  assign n38604 = ( ~n38599 & n38601 ) | ( ~n38599 & n38603 ) | ( n38601 & n38603 ) ;
  assign n38605 = n38598 & n38604 ;
  assign n38606 = n37173 ^ n32387 ^ n299 ;
  assign n38607 = n38606 ^ n11761 ^ n5180 ;
  assign n38608 = n32064 ^ n10380 ^ x41 ;
  assign n38609 = n38608 ^ n26394 ^ n17351 ;
  assign n38610 = ( n19598 & ~n29399 ) | ( n19598 & n32604 ) | ( ~n29399 & n32604 ) ;
  assign n38615 = ( n1295 & n9535 ) | ( n1295 & ~n11724 ) | ( n9535 & ~n11724 ) ;
  assign n38616 = ~n34581 & n38615 ;
  assign n38611 = n20929 & ~n28982 ;
  assign n38612 = n38611 ^ n17582 ^ 1'b0 ;
  assign n38613 = n34220 & ~n38612 ;
  assign n38614 = n38613 ^ n3204 ^ 1'b0 ;
  assign n38617 = n38616 ^ n38614 ^ n17391 ;
  assign n38618 = ( ~n14381 & n19226 ) | ( ~n14381 & n19747 ) | ( n19226 & n19747 ) ;
  assign n38619 = ( ~n5613 & n15412 ) | ( ~n5613 & n34794 ) | ( n15412 & n34794 ) ;
  assign n38620 = ( ~n12508 & n25696 ) | ( ~n12508 & n38619 ) | ( n25696 & n38619 ) ;
  assign n38621 = n35424 ^ n5993 ^ 1'b0 ;
  assign n38622 = ( n2645 & ~n4079 ) | ( n2645 & n24242 ) | ( ~n4079 & n24242 ) ;
  assign n38623 = ( ~n5238 & n6149 ) | ( ~n5238 & n38622 ) | ( n6149 & n38622 ) ;
  assign n38624 = n10390 ^ n3107 ^ n2167 ;
  assign n38625 = ~n12290 & n28357 ;
  assign n38626 = n38625 ^ n32533 ^ 1'b0 ;
  assign n38627 = n38626 ^ n12399 ^ n5059 ;
  assign n38628 = ( n12228 & ~n38624 ) | ( n12228 & n38627 ) | ( ~n38624 & n38627 ) ;
  assign n38629 = ( ~n4419 & n26682 ) | ( ~n4419 & n28899 ) | ( n26682 & n28899 ) ;
  assign n38630 = ( n5716 & n8936 ) | ( n5716 & n30539 ) | ( n8936 & n30539 ) ;
  assign n38631 = n10692 ^ n5287 ^ 1'b0 ;
  assign n38632 = ~n4109 & n38631 ;
  assign n38633 = n37548 & n38632 ;
  assign n38634 = n38630 & n38633 ;
  assign n38635 = n38634 ^ n24680 ^ n10549 ;
  assign n38636 = ( n918 & ~n1355 ) | ( n918 & n7029 ) | ( ~n1355 & n7029 ) ;
  assign n38637 = n38636 ^ n19611 ^ n747 ;
  assign n38638 = ( n1518 & n33620 ) | ( n1518 & ~n38637 ) | ( n33620 & ~n38637 ) ;
  assign n38639 = ~n13377 & n23218 ;
  assign n38642 = n21120 | n26725 ;
  assign n38643 = n38642 ^ n22854 ^ 1'b0 ;
  assign n38640 = ( n11998 & ~n12196 ) | ( n11998 & n33021 ) | ( ~n12196 & n33021 ) ;
  assign n38641 = ( n3152 & n17898 ) | ( n3152 & ~n38640 ) | ( n17898 & ~n38640 ) ;
  assign n38644 = n38643 ^ n38641 ^ n17080 ;
  assign n38645 = n15064 | n38644 ;
  assign n38646 = n38639 & ~n38645 ;
  assign n38647 = n13741 ^ n4570 ^ 1'b0 ;
  assign n38648 = n5686 | n38647 ;
  assign n38651 = ( n26327 & n26429 ) | ( n26327 & ~n31221 ) | ( n26429 & ~n31221 ) ;
  assign n38649 = n15145 ^ n7540 ^ n2161 ;
  assign n38650 = n38649 ^ n18525 ^ n17122 ;
  assign n38652 = n38651 ^ n38650 ^ n4667 ;
  assign n38659 = ~n1812 & n37707 ;
  assign n38660 = n38659 ^ x148 ^ 1'b0 ;
  assign n38653 = n18683 ^ n5354 ^ n3626 ;
  assign n38654 = n15242 ^ n12899 ^ n9322 ;
  assign n38655 = n38654 ^ n28154 ^ n21756 ;
  assign n38656 = n10788 | n38655 ;
  assign n38657 = n6542 & ~n38656 ;
  assign n38658 = ( n30546 & ~n38653 ) | ( n30546 & n38657 ) | ( ~n38653 & n38657 ) ;
  assign n38661 = n38660 ^ n38658 ^ n13687 ;
  assign n38662 = n38195 ^ n38145 ^ n7957 ;
  assign n38663 = n5804 & n27354 ;
  assign n38664 = ( n33712 & n34932 ) | ( n33712 & ~n38663 ) | ( n34932 & ~n38663 ) ;
  assign n38665 = ( n5937 & ~n18424 ) | ( n5937 & n25416 ) | ( ~n18424 & n25416 ) ;
  assign n38669 = n4151 & n35388 ;
  assign n38668 = n4016 & ~n18023 ;
  assign n38670 = n38669 ^ n38668 ^ 1'b0 ;
  assign n38666 = n22951 | n24505 ;
  assign n38667 = n38666 ^ n10393 ^ 1'b0 ;
  assign n38671 = n38670 ^ n38667 ^ n23231 ;
  assign n38672 = n38671 ^ n4443 ^ n2556 ;
  assign n38673 = n25312 ^ n12392 ^ n2491 ;
  assign n38674 = n38673 ^ n532 ^ 1'b0 ;
  assign n38675 = n38672 | n38674 ;
  assign n38676 = n8236 & n27553 ;
  assign n38677 = ~n25730 & n38676 ;
  assign n38679 = n14345 ^ n10761 ^ n2957 ;
  assign n38680 = ( n6426 & n15456 ) | ( n6426 & ~n38679 ) | ( n15456 & ~n38679 ) ;
  assign n38678 = n17359 ^ n14480 ^ n1594 ;
  assign n38681 = n38680 ^ n38678 ^ 1'b0 ;
  assign n38682 = n19760 & n38681 ;
  assign n38683 = ( ~n14739 & n27552 ) | ( ~n14739 & n28670 ) | ( n27552 & n28670 ) ;
  assign n38684 = ( ~n2527 & n24746 ) | ( ~n2527 & n36640 ) | ( n24746 & n36640 ) ;
  assign n38685 = n10431 ^ n5463 ^ n3172 ;
  assign n38686 = n19376 ^ n9316 ^ n1936 ;
  assign n38687 = n38686 ^ n13301 ^ n5026 ;
  assign n38688 = n38687 ^ n7657 ^ 1'b0 ;
  assign n38689 = n36848 ^ n21261 ^ n15826 ;
  assign n38690 = ( n19226 & n23908 ) | ( n19226 & n38689 ) | ( n23908 & n38689 ) ;
  assign n38691 = n11739 & n17660 ;
  assign n38692 = n9091 & n38691 ;
  assign n38693 = n36620 & ~n38692 ;
  assign n38694 = ( n14247 & ~n27397 ) | ( n14247 & n33416 ) | ( ~n27397 & n33416 ) ;
  assign n38695 = n38694 ^ n8232 ^ n8020 ;
  assign n38696 = n7885 & n8051 ;
  assign n38697 = n38696 ^ n27983 ^ n5580 ;
  assign n38698 = n22089 ^ n10186 ^ 1'b0 ;
  assign n38699 = n14088 & ~n17511 ;
  assign n38700 = n38699 ^ n37872 ^ 1'b0 ;
  assign n38701 = n18505 & n30924 ;
  assign n38702 = n38701 ^ n32242 ^ 1'b0 ;
  assign n38703 = n2497 | n33722 ;
  assign n38704 = n38703 ^ n16308 ^ 1'b0 ;
  assign n38705 = n27656 ^ n6553 ^ n4822 ;
  assign n38706 = n1030 ^ n694 ^ 1'b0 ;
  assign n38707 = ~n6602 & n38706 ;
  assign n38708 = ( n21599 & n38705 ) | ( n21599 & n38707 ) | ( n38705 & n38707 ) ;
  assign n38709 = n38708 ^ n22682 ^ n7736 ;
  assign n38710 = n5871 & ~n38709 ;
  assign n38711 = n17948 ^ n910 ^ 1'b0 ;
  assign n38712 = n38711 ^ n24505 ^ n9428 ;
  assign n38713 = n6269 & n20537 ;
  assign n38714 = n38713 ^ n2051 ^ 1'b0 ;
  assign n38715 = ( n1297 & n2455 ) | ( n1297 & n29373 ) | ( n2455 & n29373 ) ;
  assign n38716 = n16263 ^ n11987 ^ n11676 ;
  assign n38717 = n20128 & n38716 ;
  assign n38718 = ( n14567 & n38715 ) | ( n14567 & n38717 ) | ( n38715 & n38717 ) ;
  assign n38719 = ( n6914 & ~n25223 ) | ( n6914 & n38718 ) | ( ~n25223 & n38718 ) ;
  assign n38720 = n14264 | n38719 ;
  assign n38721 = n21990 & ~n38720 ;
  assign n38722 = n2814 ^ n522 ^ 1'b0 ;
  assign n38723 = ~n23447 & n38722 ;
  assign n38724 = n28836 ^ n25960 ^ n17622 ;
  assign n38725 = n38724 ^ n22313 ^ 1'b0 ;
  assign n38726 = n38723 & n38725 ;
  assign n38727 = n30300 ^ n7615 ^ n6344 ;
  assign n38728 = n37876 ^ n7283 ^ n4985 ;
  assign n38732 = n7630 | n21492 ;
  assign n38729 = n28679 & ~n29147 ;
  assign n38730 = n38729 ^ n20240 ^ 1'b0 ;
  assign n38731 = ( n9713 & n14382 ) | ( n9713 & ~n38730 ) | ( n14382 & ~n38730 ) ;
  assign n38733 = n38732 ^ n38731 ^ n22314 ;
  assign n38734 = n3584 ^ n3051 ^ n1074 ;
  assign n38735 = ( n5854 & n16267 ) | ( n5854 & n18325 ) | ( n16267 & n18325 ) ;
  assign n38736 = ( n4015 & n12919 ) | ( n4015 & n23356 ) | ( n12919 & n23356 ) ;
  assign n38737 = ( ~n20675 & n38735 ) | ( ~n20675 & n38736 ) | ( n38735 & n38736 ) ;
  assign n38738 = n38737 ^ n37318 ^ 1'b0 ;
  assign n38739 = ( n14827 & n38734 ) | ( n14827 & n38738 ) | ( n38734 & n38738 ) ;
  assign n38740 = n37882 ^ n12415 ^ n1768 ;
  assign n38741 = n38740 ^ n34910 ^ n15216 ;
  assign n38745 = n9024 ^ n7190 ^ n2090 ;
  assign n38743 = n16958 & n19286 ;
  assign n38744 = n38743 ^ n323 ^ 1'b0 ;
  assign n38742 = n14539 ^ n12881 ^ n12056 ;
  assign n38746 = n38745 ^ n38744 ^ n38742 ;
  assign n38747 = n6213 ^ n2397 ^ 1'b0 ;
  assign n38750 = ( n4328 & n9125 ) | ( n4328 & ~n37050 ) | ( n9125 & ~n37050 ) ;
  assign n38748 = n11365 ^ n4600 ^ 1'b0 ;
  assign n38749 = n38748 ^ n38213 ^ n20583 ;
  assign n38751 = n38750 ^ n38749 ^ n5139 ;
  assign n38752 = n12090 ^ n11598 ^ x135 ;
  assign n38753 = ( n8427 & n23250 ) | ( n8427 & ~n38752 ) | ( n23250 & ~n38752 ) ;
  assign n38754 = n38753 ^ n31583 ^ 1'b0 ;
  assign n38755 = ( n6483 & n8366 ) | ( n6483 & n38754 ) | ( n8366 & n38754 ) ;
  assign n38756 = n25203 ^ n9668 ^ n8230 ;
  assign n38757 = n28284 ^ n15843 ^ n10622 ;
  assign n38758 = ( n27014 & n38756 ) | ( n27014 & n38757 ) | ( n38756 & n38757 ) ;
  assign n38759 = n11156 | n38758 ;
  assign n38760 = n6831 & ~n38759 ;
  assign n38761 = ( n1830 & ~n6162 ) | ( n1830 & n38760 ) | ( ~n6162 & n38760 ) ;
  assign n38763 = ( n3176 & n5317 ) | ( n3176 & n11684 ) | ( n5317 & n11684 ) ;
  assign n38762 = n37411 ^ n4098 ^ 1'b0 ;
  assign n38764 = n38763 ^ n38762 ^ n18785 ;
  assign n38765 = n38764 ^ n31746 ^ n28316 ;
  assign n38766 = n18624 ^ n10865 ^ n8599 ;
  assign n38767 = n38766 ^ n21460 ^ 1'b0 ;
  assign n38768 = n38767 ^ n33436 ^ n18180 ;
  assign n38769 = ( n2471 & n3443 ) | ( n2471 & n18537 ) | ( n3443 & n18537 ) ;
  assign n38770 = n38769 ^ n4113 ^ n2403 ;
  assign n38771 = n38770 ^ n11351 ^ n5546 ;
  assign n38772 = n25630 ^ n15428 ^ n1508 ;
  assign n38773 = ( n19382 & n38771 ) | ( n19382 & n38772 ) | ( n38771 & n38772 ) ;
  assign n38774 = n38773 ^ n20516 ^ 1'b0 ;
  assign n38775 = ( n10722 & ~n23324 ) | ( n10722 & n31500 ) | ( ~n23324 & n31500 ) ;
  assign n38776 = n38775 ^ n24704 ^ 1'b0 ;
  assign n38778 = n36277 ^ n17512 ^ n6537 ;
  assign n38779 = n38778 ^ n12521 ^ n10394 ;
  assign n38777 = ( n10559 & ~n17224 ) | ( n10559 & n21520 ) | ( ~n17224 & n21520 ) ;
  assign n38780 = n38779 ^ n38777 ^ n13796 ;
  assign n38781 = n37793 ^ n37112 ^ 1'b0 ;
  assign n38782 = n14288 & ~n24274 ;
  assign n38783 = n38782 ^ n15011 ^ 1'b0 ;
  assign n38784 = ( ~n12235 & n13295 ) | ( ~n12235 & n27013 ) | ( n13295 & n27013 ) ;
  assign n38785 = ~n3966 & n7323 ;
  assign n38787 = n2612 ^ n1233 ^ 1'b0 ;
  assign n38788 = n38787 ^ n38717 ^ n6718 ;
  assign n38786 = n1941 & n3722 ;
  assign n38789 = n38788 ^ n38786 ^ 1'b0 ;
  assign n38790 = n6610 | n38789 ;
  assign n38791 = n23939 ^ n17655 ^ 1'b0 ;
  assign n38792 = n28739 | n38791 ;
  assign n38793 = n21430 ^ x200 ^ 1'b0 ;
  assign n38794 = n15992 | n38793 ;
  assign n38795 = ( ~n5151 & n24643 ) | ( ~n5151 & n38794 ) | ( n24643 & n38794 ) ;
  assign n38796 = ( ~n3471 & n13813 ) | ( ~n3471 & n17749 ) | ( n13813 & n17749 ) ;
  assign n38797 = n27368 | n38796 ;
  assign n38798 = n38797 ^ n1278 ^ 1'b0 ;
  assign n38799 = ( n11987 & n38795 ) | ( n11987 & n38798 ) | ( n38795 & n38798 ) ;
  assign n38801 = ( ~n2620 & n9633 ) | ( ~n2620 & n11285 ) | ( n9633 & n11285 ) ;
  assign n38802 = n38801 ^ n35635 ^ n3828 ;
  assign n38803 = ( n15257 & n18624 ) | ( n15257 & n38802 ) | ( n18624 & n38802 ) ;
  assign n38800 = n12044 & n17845 ;
  assign n38804 = n38803 ^ n38800 ^ 1'b0 ;
  assign n38805 = n12624 | n37144 ;
  assign n38806 = n15681 ^ n10766 ^ 1'b0 ;
  assign n38807 = n38805 & ~n38806 ;
  assign n38808 = ( n1440 & n8388 ) | ( n1440 & n11403 ) | ( n8388 & n11403 ) ;
  assign n38809 = ( ~n3593 & n15949 ) | ( ~n3593 & n24386 ) | ( n15949 & n24386 ) ;
  assign n38810 = ( ~n11283 & n29949 ) | ( ~n11283 & n38809 ) | ( n29949 & n38809 ) ;
  assign n38811 = n1304 & ~n38810 ;
  assign n38812 = n38808 & n38811 ;
  assign n38813 = n5699 & n28648 ;
  assign n38814 = ( n9296 & ~n22978 ) | ( n9296 & n38813 ) | ( ~n22978 & n38813 ) ;
  assign n38815 = n38814 ^ n22176 ^ n16572 ;
  assign n38816 = ( n8901 & ~n37592 ) | ( n8901 & n38815 ) | ( ~n37592 & n38815 ) ;
  assign n38817 = n30970 ^ n15823 ^ n10467 ;
  assign n38818 = ~n12455 & n14843 ;
  assign n38819 = n34930 ^ n20941 ^ n9653 ;
  assign n38820 = ( n18147 & ~n27913 ) | ( n18147 & n38819 ) | ( ~n27913 & n38819 ) ;
  assign n38821 = ( n282 & ~n31173 ) | ( n282 & n31528 ) | ( ~n31173 & n31528 ) ;
  assign n38822 = n8095 ^ n6185 ^ 1'b0 ;
  assign n38823 = n7796 | n38822 ;
  assign n38824 = n5530 & n38823 ;
  assign n38825 = ( n15144 & n15431 ) | ( n15144 & ~n38824 ) | ( n15431 & ~n38824 ) ;
  assign n38826 = n29158 ^ n20447 ^ n14045 ;
  assign n38827 = n33423 ^ n25892 ^ n17386 ;
  assign n38828 = ~n1274 & n21139 ;
  assign n38829 = ( n8740 & n38242 ) | ( n8740 & n38828 ) | ( n38242 & n38828 ) ;
  assign n38830 = n19360 ^ n7292 ^ n4664 ;
  assign n38832 = n29283 ^ n23088 ^ n16029 ;
  assign n38831 = n8611 | n27548 ;
  assign n38833 = n38832 ^ n38831 ^ 1'b0 ;
  assign n38834 = n14799 & ~n25302 ;
  assign n38835 = ~n9183 & n38834 ;
  assign n38836 = ( ~n25879 & n28212 ) | ( ~n25879 & n32259 ) | ( n28212 & n32259 ) ;
  assign n38837 = n38836 ^ n36717 ^ n2511 ;
  assign n38838 = n22549 ^ n3625 ^ n1091 ;
  assign n38839 = ( n11298 & ~n29398 ) | ( n11298 & n38588 ) | ( ~n29398 & n38588 ) ;
  assign n38840 = ( n1899 & n22174 ) | ( n1899 & ~n30863 ) | ( n22174 & ~n30863 ) ;
  assign n38841 = ( n9530 & ~n38839 ) | ( n9530 & n38840 ) | ( ~n38839 & n38840 ) ;
  assign n38842 = ( n12641 & n21049 ) | ( n12641 & n38841 ) | ( n21049 & n38841 ) ;
  assign n38843 = ~n16099 & n25287 ;
  assign n38844 = n38843 ^ n4008 ^ 1'b0 ;
  assign n38845 = n38844 ^ n24008 ^ n11113 ;
  assign n38846 = ( n2171 & n22903 ) | ( n2171 & n35529 ) | ( n22903 & n35529 ) ;
  assign n38847 = ( n19533 & n28148 ) | ( n19533 & n36256 ) | ( n28148 & n36256 ) ;
  assign n38848 = n630 | n8055 ;
  assign n38849 = n38847 | n38848 ;
  assign n38850 = n22392 & ~n23212 ;
  assign n38851 = n38850 ^ n5490 ^ 1'b0 ;
  assign n38853 = n7906 & ~n26772 ;
  assign n38854 = n5725 & n38853 ;
  assign n38855 = n38854 ^ n7549 ^ n5030 ;
  assign n38852 = n23992 ^ n22564 ^ n11022 ;
  assign n38856 = n38855 ^ n38852 ^ 1'b0 ;
  assign n38857 = n14549 ^ n7080 ^ n6687 ;
  assign n38858 = n38857 ^ n28973 ^ n4072 ;
  assign n38859 = n11969 ^ n5959 ^ 1'b0 ;
  assign n38860 = n19691 ^ n4647 ^ 1'b0 ;
  assign n38861 = n20748 | n38860 ;
  assign n38862 = n26843 ^ n5625 ^ 1'b0 ;
  assign n38863 = ( n29542 & n38861 ) | ( n29542 & n38862 ) | ( n38861 & n38862 ) ;
  assign n38864 = n19465 ^ n16788 ^ n797 ;
  assign n38865 = ( n10111 & n22950 ) | ( n10111 & ~n23390 ) | ( n22950 & ~n23390 ) ;
  assign n38866 = n38865 ^ n30501 ^ 1'b0 ;
  assign n38867 = n7323 & ~n27125 ;
  assign n38868 = n38867 ^ n3267 ^ 1'b0 ;
  assign n38869 = ( n2546 & n8203 ) | ( n2546 & ~n19699 ) | ( n8203 & ~n19699 ) ;
  assign n38870 = n15435 & ~n31529 ;
  assign n38871 = ( n4328 & n5952 ) | ( n4328 & ~n20876 ) | ( n5952 & ~n20876 ) ;
  assign n38872 = n1071 | n3360 ;
  assign n38873 = n38871 & ~n38872 ;
  assign n38874 = n14293 ^ n9968 ^ n4245 ;
  assign n38875 = n11318 ^ n7797 ^ n6100 ;
  assign n38876 = ~n12103 & n28312 ;
  assign n38877 = n38875 & n38876 ;
  assign n38879 = n3617 ^ n1173 ^ 1'b0 ;
  assign n38878 = ( n3096 & n8207 ) | ( n3096 & ~n14290 ) | ( n8207 & ~n14290 ) ;
  assign n38880 = n38879 ^ n38878 ^ n1612 ;
  assign n38881 = n38880 ^ n16363 ^ n16098 ;
  assign n38882 = ( n6525 & n17450 ) | ( n6525 & ~n38881 ) | ( n17450 & ~n38881 ) ;
  assign n38883 = n7351 | n38882 ;
  assign n38884 = n38877 & ~n38883 ;
  assign n38885 = ( n38873 & n38874 ) | ( n38873 & n38884 ) | ( n38874 & n38884 ) ;
  assign n38886 = ( n7061 & n23841 ) | ( n7061 & n38499 ) | ( n23841 & n38499 ) ;
  assign n38887 = ( n7854 & n8845 ) | ( n7854 & n38886 ) | ( n8845 & n38886 ) ;
  assign n38888 = n31297 | n38887 ;
  assign n38889 = n23588 & ~n38888 ;
  assign n38890 = ~n632 & n24069 ;
  assign n38891 = n38890 ^ n33548 ^ 1'b0 ;
  assign n38892 = ( ~n4701 & n9237 ) | ( ~n4701 & n30765 ) | ( n9237 & n30765 ) ;
  assign n38893 = n2407 | n9329 ;
  assign n38894 = n38893 ^ n11487 ^ 1'b0 ;
  assign n38895 = n38894 ^ n12570 ^ n6621 ;
  assign n38896 = ( n981 & n10036 ) | ( n981 & ~n29573 ) | ( n10036 & ~n29573 ) ;
  assign n38899 = ( n4464 & n9326 ) | ( n4464 & ~n11235 ) | ( n9326 & ~n11235 ) ;
  assign n38897 = n18111 | n37555 ;
  assign n38898 = n38897 ^ n7907 ^ 1'b0 ;
  assign n38900 = n38899 ^ n38898 ^ n33458 ;
  assign n38908 = ( x69 & n3350 ) | ( x69 & ~n35118 ) | ( n3350 & ~n35118 ) ;
  assign n38901 = n17109 ^ n15788 ^ n12992 ;
  assign n38902 = n18084 ^ n10961 ^ 1'b0 ;
  assign n38903 = ~n32310 & n38902 ;
  assign n38904 = n38903 ^ n31702 ^ 1'b0 ;
  assign n38905 = n38904 ^ n3306 ^ 1'b0 ;
  assign n38906 = ( ~n35540 & n38901 ) | ( ~n35540 & n38905 ) | ( n38901 & n38905 ) ;
  assign n38907 = ( n8783 & ~n28035 ) | ( n8783 & n38906 ) | ( ~n28035 & n38906 ) ;
  assign n38909 = n38908 ^ n38907 ^ n17309 ;
  assign n38910 = n38909 ^ n17652 ^ n14470 ;
  assign n38911 = n38910 ^ n30109 ^ n12558 ;
  assign n38912 = ( n14255 & n14862 ) | ( n14255 & n25666 ) | ( n14862 & n25666 ) ;
  assign n38913 = ( ~n6726 & n17485 ) | ( ~n6726 & n18417 ) | ( n17485 & n18417 ) ;
  assign n38914 = ( x218 & ~n36286 ) | ( x218 & n38913 ) | ( ~n36286 & n38913 ) ;
  assign n38915 = ( n9981 & n24871 ) | ( n9981 & n38914 ) | ( n24871 & n38914 ) ;
  assign n38918 = ( n1257 & ~n9155 ) | ( n1257 & n14307 ) | ( ~n9155 & n14307 ) ;
  assign n38917 = n15547 ^ n14381 ^ n6328 ;
  assign n38916 = n7450 & ~n11841 ;
  assign n38919 = n38918 ^ n38917 ^ n38916 ;
  assign n38920 = n24327 ^ n10737 ^ 1'b0 ;
  assign n38921 = n3632 & ~n33208 ;
  assign n38922 = n38921 ^ n29405 ^ 1'b0 ;
  assign n38923 = ( n10140 & n21257 ) | ( n10140 & n21602 ) | ( n21257 & n21602 ) ;
  assign n38924 = ( ~n3840 & n25217 ) | ( ~n3840 & n38923 ) | ( n25217 & n38923 ) ;
  assign n38925 = n4642 & ~n7309 ;
  assign n38926 = n38191 ^ n35042 ^ n7837 ;
  assign n38927 = n2363 & n12196 ;
  assign n38932 = n16980 ^ n4564 ^ 1'b0 ;
  assign n38930 = ~n4908 & n25239 ;
  assign n38931 = n17522 & n38930 ;
  assign n38928 = ( ~n3814 & n9551 ) | ( ~n3814 & n32115 ) | ( n9551 & n32115 ) ;
  assign n38929 = ( ~n9818 & n11899 ) | ( ~n9818 & n38928 ) | ( n11899 & n38928 ) ;
  assign n38933 = n38932 ^ n38931 ^ n38929 ;
  assign n38934 = ( n27157 & n30200 ) | ( n27157 & n38933 ) | ( n30200 & n38933 ) ;
  assign n38935 = n28248 ^ n14612 ^ n4078 ;
  assign n38936 = ( n3355 & n24958 ) | ( n3355 & n38935 ) | ( n24958 & n38935 ) ;
  assign n38937 = ( n2528 & n12717 ) | ( n2528 & n24616 ) | ( n12717 & n24616 ) ;
  assign n38938 = n38937 ^ n28772 ^ n7081 ;
  assign n38939 = n38938 ^ n19739 ^ n14543 ;
  assign n38940 = n18193 ^ n15809 ^ n8025 ;
  assign n38941 = n33397 ^ n15265 ^ n11365 ;
  assign n38942 = n8676 | n10359 ;
  assign n38943 = n38942 ^ n10393 ^ 1'b0 ;
  assign n38944 = n13463 ^ n4580 ^ n740 ;
  assign n38945 = n38944 ^ n5590 ^ n416 ;
  assign n38946 = n689 | n3016 ;
  assign n38947 = n38945 & ~n38946 ;
  assign n38948 = ( n35046 & n38943 ) | ( n35046 & ~n38947 ) | ( n38943 & ~n38947 ) ;
  assign n38949 = n38948 ^ n32071 ^ n1557 ;
  assign n38950 = n32973 ^ n21961 ^ 1'b0 ;
  assign n38951 = ( n10484 & n25597 ) | ( n10484 & ~n35939 ) | ( n25597 & ~n35939 ) ;
  assign n38952 = ( n26882 & n29713 ) | ( n26882 & n38951 ) | ( n29713 & n38951 ) ;
  assign n38953 = n38952 ^ n31095 ^ n4423 ;
  assign n38954 = n34367 ^ n13101 ^ n2188 ;
  assign n38955 = n38954 ^ n30623 ^ 1'b0 ;
  assign n38956 = n7065 | n38955 ;
  assign n38957 = ( ~n20640 & n28522 ) | ( ~n20640 & n30107 ) | ( n28522 & n30107 ) ;
  assign n38958 = ( ~n14390 & n17702 ) | ( ~n14390 & n38957 ) | ( n17702 & n38957 ) ;
  assign n38959 = ~n28851 & n38958 ;
  assign n38960 = n5208 | n14485 ;
  assign n38961 = n20419 | n38960 ;
  assign n38962 = n30947 ^ n10430 ^ n6935 ;
  assign n38963 = n38962 ^ n27384 ^ n2698 ;
  assign n38965 = n38769 ^ n6659 ^ 1'b0 ;
  assign n38966 = ~n10289 & n38965 ;
  assign n38967 = ~n3034 & n38966 ;
  assign n38968 = ~n22137 & n38967 ;
  assign n38964 = n21780 ^ n8777 ^ n3848 ;
  assign n38969 = n38968 ^ n38964 ^ n28812 ;
  assign n38975 = ( n581 & n8455 ) | ( n581 & n13222 ) | ( n8455 & n13222 ) ;
  assign n38970 = ( ~n20449 & n32325 ) | ( ~n20449 & n38791 ) | ( n32325 & n38791 ) ;
  assign n38971 = n38707 ^ n9877 ^ n6042 ;
  assign n38972 = ( n4119 & ~n36149 ) | ( n4119 & n38971 ) | ( ~n36149 & n38971 ) ;
  assign n38973 = ( n24741 & ~n30392 ) | ( n24741 & n38972 ) | ( ~n30392 & n38972 ) ;
  assign n38974 = ( n23752 & n38970 ) | ( n23752 & ~n38973 ) | ( n38970 & ~n38973 ) ;
  assign n38976 = n38975 ^ n38974 ^ n2043 ;
  assign n38977 = n37851 ^ n24643 ^ n18797 ;
  assign n38979 = ~n9810 & n15598 ;
  assign n38978 = n30949 ^ n20916 ^ n4520 ;
  assign n38980 = n38979 ^ n38978 ^ n8020 ;
  assign n38981 = n13440 | n20462 ;
  assign n38982 = n10508 ^ n6087 ^ 1'b0 ;
  assign n38983 = ( n8232 & ~n33973 ) | ( n8232 & n38982 ) | ( ~n33973 & n38982 ) ;
  assign n38984 = ( n12944 & ~n38981 ) | ( n12944 & n38983 ) | ( ~n38981 & n38983 ) ;
  assign n38986 = n12042 ^ n7799 ^ n2108 ;
  assign n38985 = n25437 ^ n14070 ^ n2147 ;
  assign n38987 = n38986 ^ n38985 ^ n20936 ;
  assign n38988 = ~n4641 & n38987 ;
  assign n38989 = n35871 ^ n9655 ^ 1'b0 ;
  assign n38990 = ( n11801 & n22016 ) | ( n11801 & n38655 ) | ( n22016 & n38655 ) ;
  assign n38991 = n34693 & n38990 ;
  assign n38992 = ~n38990 & n38991 ;
  assign n38994 = n17345 ^ n12014 ^ 1'b0 ;
  assign n38995 = ( n2241 & n8994 ) | ( n2241 & ~n38994 ) | ( n8994 & ~n38994 ) ;
  assign n38993 = ( n7001 & n23183 ) | ( n7001 & ~n26306 ) | ( n23183 & ~n26306 ) ;
  assign n38996 = n38995 ^ n38993 ^ 1'b0 ;
  assign n38997 = n35811 ^ n27320 ^ n9116 ;
  assign n38998 = ( n9280 & ~n19373 ) | ( n9280 & n23596 ) | ( ~n19373 & n23596 ) ;
  assign n38999 = ( ~n15072 & n17088 ) | ( ~n15072 & n38998 ) | ( n17088 & n38998 ) ;
  assign n39000 = ( n24150 & n34053 ) | ( n24150 & ~n36157 ) | ( n34053 & ~n36157 ) ;
  assign n39001 = n19390 ^ n12817 ^ n12801 ;
  assign n39002 = n27223 ^ n16937 ^ n9086 ;
  assign n39003 = ~n9028 & n39002 ;
  assign n39004 = ~n36058 & n39003 ;
  assign n39005 = ( ~n11801 & n20274 ) | ( ~n11801 & n30594 ) | ( n20274 & n30594 ) ;
  assign n39006 = n13774 & ~n39005 ;
  assign n39007 = n39006 ^ n34684 ^ 1'b0 ;
  assign n39008 = n12970 ^ n9241 ^ n1530 ;
  assign n39009 = n39008 ^ n24933 ^ n15066 ;
  assign n39010 = n17696 ^ n14511 ^ n14123 ;
  assign n39011 = n39010 ^ n27341 ^ n7755 ;
  assign n39012 = n19595 ^ n16180 ^ n5935 ;
  assign n39013 = n39012 ^ n24223 ^ n22959 ;
  assign n39014 = n38270 ^ n14682 ^ 1'b0 ;
  assign n39016 = n20884 ^ n9106 ^ n8213 ;
  assign n39017 = n39016 ^ n14649 ^ n6407 ;
  assign n39015 = n6278 & n19932 ;
  assign n39018 = n39017 ^ n39015 ^ n38463 ;
  assign n39019 = n39018 ^ n5446 ^ 1'b0 ;
  assign n39020 = n36849 ^ n32270 ^ 1'b0 ;
  assign n39021 = n36071 ^ n26500 ^ 1'b0 ;
  assign n39022 = n8720 & ~n39021 ;
  assign n39023 = ( ~n3698 & n6312 ) | ( ~n3698 & n39022 ) | ( n6312 & n39022 ) ;
  assign n39024 = n39023 ^ n20535 ^ 1'b0 ;
  assign n39025 = ~n25803 & n39024 ;
  assign n39026 = n39025 ^ n13771 ^ 1'b0 ;
  assign n39027 = n17703 ^ n9644 ^ n8039 ;
  assign n39028 = n38397 ^ n37778 ^ 1'b0 ;
  assign n39029 = n39027 | n39028 ;
  assign n39030 = n28852 & ~n39029 ;
  assign n39031 = n7066 | n15506 ;
  assign n39032 = n8286 & ~n39031 ;
  assign n39033 = n39032 ^ n4426 ^ 1'b0 ;
  assign n39034 = n39033 ^ n38789 ^ n21628 ;
  assign n39037 = n18481 ^ n16595 ^ 1'b0 ;
  assign n39038 = ~n9713 & n39037 ;
  assign n39035 = ( n19863 & ~n29060 ) | ( n19863 & n37923 ) | ( ~n29060 & n37923 ) ;
  assign n39036 = n3831 & ~n39035 ;
  assign n39039 = n39038 ^ n39036 ^ 1'b0 ;
  assign n39040 = ( ~n12441 & n19719 ) | ( ~n12441 & n39039 ) | ( n19719 & n39039 ) ;
  assign n39041 = n898 & ~n17406 ;
  assign n39042 = ~n13356 & n39041 ;
  assign n39043 = n38390 ^ n7006 ^ 1'b0 ;
  assign n39044 = n39042 & n39043 ;
  assign n39045 = n17446 ^ n10232 ^ n8762 ;
  assign n39046 = n4764 | n6019 ;
  assign n39047 = n1313 & ~n39046 ;
  assign n39048 = ( n2226 & ~n4941 ) | ( n2226 & n5715 ) | ( ~n4941 & n5715 ) ;
  assign n39049 = ( n22525 & n31115 ) | ( n22525 & ~n39048 ) | ( n31115 & ~n39048 ) ;
  assign n39050 = n28318 ^ n5399 ^ n2250 ;
  assign n39054 = n15122 ^ n7132 ^ 1'b0 ;
  assign n39051 = n2838 & n16340 ;
  assign n39052 = n39051 ^ n6243 ^ 1'b0 ;
  assign n39053 = ( n6482 & n27271 ) | ( n6482 & ~n39052 ) | ( n27271 & ~n39052 ) ;
  assign n39055 = n39054 ^ n39053 ^ 1'b0 ;
  assign n39056 = ~n39050 & n39055 ;
  assign n39057 = n14093 ^ n7684 ^ n464 ;
  assign n39058 = ( n9665 & n17821 ) | ( n9665 & n39057 ) | ( n17821 & n39057 ) ;
  assign n39059 = n24108 ^ n15118 ^ n15099 ;
  assign n39060 = ( n16272 & n28344 ) | ( n16272 & n39059 ) | ( n28344 & n39059 ) ;
  assign n39061 = ( n5446 & n21087 ) | ( n5446 & ~n39060 ) | ( n21087 & ~n39060 ) ;
  assign n39062 = n9116 & n32588 ;
  assign n39063 = n39062 ^ n9885 ^ 1'b0 ;
  assign n39064 = n39063 ^ n22166 ^ n20787 ;
  assign n39065 = ( n14448 & n37522 ) | ( n14448 & n39064 ) | ( n37522 & n39064 ) ;
  assign n39067 = ~n20113 & n30643 ;
  assign n39068 = n39067 ^ n19315 ^ 1'b0 ;
  assign n39066 = n31783 & ~n34111 ;
  assign n39069 = n39068 ^ n39066 ^ 1'b0 ;
  assign n39071 = ( n1951 & n14705 ) | ( n1951 & ~n20326 ) | ( n14705 & ~n20326 ) ;
  assign n39072 = n39071 ^ n23580 ^ n4738 ;
  assign n39073 = n31483 ^ n20663 ^ 1'b0 ;
  assign n39074 = n11889 & n39073 ;
  assign n39075 = ( n292 & n14423 ) | ( n292 & ~n39074 ) | ( n14423 & ~n39074 ) ;
  assign n39076 = ( ~n4638 & n39072 ) | ( ~n4638 & n39075 ) | ( n39072 & n39075 ) ;
  assign n39070 = ( n7348 & ~n22344 ) | ( n7348 & n37241 ) | ( ~n22344 & n37241 ) ;
  assign n39077 = n39076 ^ n39070 ^ 1'b0 ;
  assign n39078 = ~n7004 & n39077 ;
  assign n39086 = n27956 ^ n26499 ^ 1'b0 ;
  assign n39084 = ( n16515 & n17681 ) | ( n16515 & ~n38905 ) | ( n17681 & ~n38905 ) ;
  assign n39079 = n4146 & ~n27854 ;
  assign n39080 = ~n26699 & n39079 ;
  assign n39081 = n14185 ^ n6387 ^ n4332 ;
  assign n39082 = n39081 ^ n19737 ^ x50 ;
  assign n39083 = n39080 & ~n39082 ;
  assign n39085 = n39084 ^ n39083 ^ n19895 ;
  assign n39087 = n39086 ^ n39085 ^ n34202 ;
  assign n39088 = ( n5990 & n29260 ) | ( n5990 & ~n38975 ) | ( n29260 & ~n38975 ) ;
  assign n39089 = n25314 ^ n13033 ^ n9476 ;
  assign n39090 = ~n9329 & n39089 ;
  assign n39091 = n20067 ^ n12830 ^ n3315 ;
  assign n39092 = n39091 ^ n26669 ^ n3122 ;
  assign n39093 = n39092 ^ n14785 ^ 1'b0 ;
  assign n39094 = ( n973 & ~n1810 ) | ( n973 & n3528 ) | ( ~n1810 & n3528 ) ;
  assign n39095 = n28802 ^ n6400 ^ 1'b0 ;
  assign n39096 = n39094 | n39095 ;
  assign n39102 = ( ~n12647 & n19310 ) | ( ~n12647 & n20957 ) | ( n19310 & n20957 ) ;
  assign n39103 = ( ~n15019 & n21327 ) | ( ~n15019 & n39102 ) | ( n21327 & n39102 ) ;
  assign n39100 = n27950 ^ n5236 ^ n4151 ;
  assign n39098 = n11287 ^ n8329 ^ 1'b0 ;
  assign n39099 = n13924 & n39098 ;
  assign n39101 = n39100 ^ n39099 ^ n22839 ;
  assign n39104 = n39103 ^ n39101 ^ n38258 ;
  assign n39097 = x231 & ~n22015 ;
  assign n39105 = n39104 ^ n39097 ^ 1'b0 ;
  assign n39106 = n19086 ^ n12809 ^ n10618 ;
  assign n39107 = ~n9796 & n11336 ;
  assign n39108 = n39107 ^ n26186 ^ 1'b0 ;
  assign n39109 = n28871 ^ n4859 ^ n3546 ;
  assign n39110 = n1236 & ~n7540 ;
  assign n39111 = n1147 & n39110 ;
  assign n39112 = n39111 ^ n22825 ^ n1627 ;
  assign n39113 = n39112 ^ n37911 ^ n7385 ;
  assign n39114 = ( n25842 & ~n39109 ) | ( n25842 & n39113 ) | ( ~n39109 & n39113 ) ;
  assign n39116 = ( n518 & n6238 ) | ( n518 & n14545 ) | ( n6238 & n14545 ) ;
  assign n39115 = ~n13282 & n19220 ;
  assign n39117 = n39116 ^ n39115 ^ n15391 ;
  assign n39118 = n39117 ^ n24838 ^ n1424 ;
  assign n39119 = ( n13251 & n18006 ) | ( n13251 & ~n26084 ) | ( n18006 & ~n26084 ) ;
  assign n39120 = n10914 ^ n9364 ^ n5512 ;
  assign n39121 = ~n1211 & n5555 ;
  assign n39122 = ~n39120 & n39121 ;
  assign n39123 = ( x74 & ~n11343 ) | ( x74 & n17627 ) | ( ~n11343 & n17627 ) ;
  assign n39124 = n34476 ^ n16297 ^ 1'b0 ;
  assign n39125 = n39123 & ~n39124 ;
  assign n39126 = ( ~n39119 & n39122 ) | ( ~n39119 & n39125 ) | ( n39122 & n39125 ) ;
  assign n39127 = n11497 ^ n8745 ^ n6769 ;
  assign n39128 = ( n1464 & ~n9129 ) | ( n1464 & n23061 ) | ( ~n9129 & n23061 ) ;
  assign n39129 = n35633 ^ n3631 ^ x19 ;
  assign n39130 = n22324 ^ n4298 ^ n3021 ;
  assign n39131 = ~n39129 & n39130 ;
  assign n39132 = ~n21457 & n39131 ;
  assign n39133 = ~n35588 & n38586 ;
  assign n39134 = ~n29959 & n39133 ;
  assign n39137 = n969 | n2523 ;
  assign n39138 = n13030 | n39137 ;
  assign n39135 = n11820 & ~n20166 ;
  assign n39136 = ~n29057 & n39135 ;
  assign n39139 = n39138 ^ n39136 ^ n815 ;
  assign n39140 = ( n7717 & ~n15628 ) | ( n7717 & n32312 ) | ( ~n15628 & n32312 ) ;
  assign n39141 = n1690 ^ n1686 ^ 1'b0 ;
  assign n39142 = ( ~n9227 & n38263 ) | ( ~n9227 & n39141 ) | ( n38263 & n39141 ) ;
  assign n39143 = n32600 ^ n2983 ^ 1'b0 ;
  assign n39145 = ( n1800 & n8631 ) | ( n1800 & ~n22418 ) | ( n8631 & ~n22418 ) ;
  assign n39144 = n18516 ^ n11349 ^ n7806 ;
  assign n39146 = n39145 ^ n39144 ^ 1'b0 ;
  assign n39147 = n19521 ^ n10010 ^ n9779 ;
  assign n39148 = n30818 ^ n30078 ^ n851 ;
  assign n39149 = n19035 ^ n12611 ^ n4908 ;
  assign n39150 = ( n39147 & n39148 ) | ( n39147 & n39149 ) | ( n39148 & n39149 ) ;
  assign n39151 = n38308 ^ n5744 ^ 1'b0 ;
  assign n39152 = n15298 & ~n39151 ;
  assign n39153 = n26647 ^ n18610 ^ 1'b0 ;
  assign n39154 = n19703 & ~n39153 ;
  assign n39155 = n37469 | n39154 ;
  assign n39156 = n39155 ^ n16764 ^ 1'b0 ;
  assign n39157 = n14712 ^ n5170 ^ n4024 ;
  assign n39158 = n39157 ^ n13073 ^ n2202 ;
  assign n39159 = n38534 ^ n14083 ^ 1'b0 ;
  assign n39167 = ( n916 & n9438 ) | ( n916 & ~n26178 ) | ( n9438 & ~n26178 ) ;
  assign n39168 = n39167 ^ n5799 ^ n2805 ;
  assign n39160 = ( n7056 & ~n26137 ) | ( n7056 & n35746 ) | ( ~n26137 & n35746 ) ;
  assign n39161 = ~n7997 & n9942 ;
  assign n39162 = n12322 ^ n10410 ^ 1'b0 ;
  assign n39163 = n39161 & ~n39162 ;
  assign n39164 = ( n24435 & n39160 ) | ( n24435 & ~n39163 ) | ( n39160 & ~n39163 ) ;
  assign n39165 = n18645 ^ n16027 ^ 1'b0 ;
  assign n39166 = n39164 | n39165 ;
  assign n39169 = n39168 ^ n39166 ^ 1'b0 ;
  assign n39170 = n20040 ^ n12454 ^ n8183 ;
  assign n39171 = ~n24286 & n39170 ;
  assign n39172 = n17383 & n39171 ;
  assign n39173 = ( n7882 & n10606 ) | ( n7882 & n28388 ) | ( n10606 & n28388 ) ;
  assign n39174 = n39173 ^ n5146 ^ 1'b0 ;
  assign n39175 = ( n1958 & n12819 ) | ( n1958 & n26013 ) | ( n12819 & n26013 ) ;
  assign n39177 = n5979 | n6491 ;
  assign n39176 = n35951 ^ n25217 ^ 1'b0 ;
  assign n39178 = n39177 ^ n39176 ^ n38810 ;
  assign n39181 = n3293 | n3493 ;
  assign n39179 = n32660 ^ n25399 ^ n12338 ;
  assign n39180 = n39179 ^ n17059 ^ n5721 ;
  assign n39182 = n39181 ^ n39180 ^ n1505 ;
  assign n39183 = n3756 ^ n1768 ^ 1'b0 ;
  assign n39184 = n39183 ^ n29089 ^ n28597 ;
  assign n39185 = ( n1226 & n23102 ) | ( n1226 & ~n24891 ) | ( n23102 & ~n24891 ) ;
  assign n39186 = n39185 ^ n15055 ^ 1'b0 ;
  assign n39187 = n39186 ^ n32015 ^ n13931 ;
  assign n39188 = ( ~n1263 & n5810 ) | ( ~n1263 & n39187 ) | ( n5810 & n39187 ) ;
  assign n39192 = n20033 ^ n11953 ^ n2658 ;
  assign n39193 = ( n2527 & n4417 ) | ( n2527 & ~n6766 ) | ( n4417 & ~n6766 ) ;
  assign n39194 = n39193 ^ n38279 ^ 1'b0 ;
  assign n39195 = ~n39192 & n39194 ;
  assign n39196 = n39195 ^ n38612 ^ n2244 ;
  assign n39189 = n10271 & ~n26292 ;
  assign n39190 = n39189 ^ n31475 ^ 1'b0 ;
  assign n39191 = ~n4092 & n39190 ;
  assign n39197 = n39196 ^ n39191 ^ 1'b0 ;
  assign n39202 = n19927 ^ n10018 ^ n7050 ;
  assign n39198 = ( x102 & ~n17334 ) | ( x102 & n19405 ) | ( ~n17334 & n19405 ) ;
  assign n39199 = ( n15139 & ~n21341 ) | ( n15139 & n39198 ) | ( ~n21341 & n39198 ) ;
  assign n39200 = ( n19265 & n22593 ) | ( n19265 & ~n24231 ) | ( n22593 & ~n24231 ) ;
  assign n39201 = ( n14510 & n39199 ) | ( n14510 & n39200 ) | ( n39199 & n39200 ) ;
  assign n39203 = n39202 ^ n39201 ^ n17764 ;
  assign n39204 = n19246 ^ n10956 ^ n3616 ;
  assign n39205 = ( n352 & n4597 ) | ( n352 & n26146 ) | ( n4597 & n26146 ) ;
  assign n39206 = ( n2704 & n5766 ) | ( n2704 & ~n35614 ) | ( n5766 & ~n35614 ) ;
  assign n39207 = n20897 & n24356 ;
  assign n39208 = n39207 ^ n13105 ^ 1'b0 ;
  assign n39209 = ( n4834 & n7592 ) | ( n4834 & ~n24620 ) | ( n7592 & ~n24620 ) ;
  assign n39210 = ( ~n6533 & n18435 ) | ( ~n6533 & n39209 ) | ( n18435 & n39209 ) ;
  assign n39211 = n629 & ~n10735 ;
  assign n39212 = n39211 ^ n13105 ^ 1'b0 ;
  assign n39213 = ( n26901 & n31144 ) | ( n26901 & ~n39212 ) | ( n31144 & ~n39212 ) ;
  assign n39214 = n39213 ^ n13442 ^ 1'b0 ;
  assign n39215 = n10768 | n39214 ;
  assign n39216 = ( n21709 & ~n39210 ) | ( n21709 & n39215 ) | ( ~n39210 & n39215 ) ;
  assign n39217 = ( n9803 & ~n17943 ) | ( n9803 & n39216 ) | ( ~n17943 & n39216 ) ;
  assign n39218 = n1408 | n29270 ;
  assign n39219 = n39218 ^ n7080 ^ 1'b0 ;
  assign n39220 = n39219 ^ n20068 ^ n14912 ;
  assign n39221 = n37721 ^ n25117 ^ n9804 ;
  assign n39222 = n1257 | n23210 ;
  assign n39223 = ( n4910 & ~n25486 ) | ( n4910 & n27805 ) | ( ~n25486 & n27805 ) ;
  assign n39224 = ( n4246 & ~n7047 ) | ( n4246 & n24703 ) | ( ~n7047 & n24703 ) ;
  assign n39225 = n7567 & ~n39224 ;
  assign n39226 = n37556 ^ n32280 ^ n4903 ;
  assign n39227 = n28942 | n39226 ;
  assign n39228 = n39227 ^ n18779 ^ 1'b0 ;
  assign n39229 = ( n25512 & n39225 ) | ( n25512 & ~n39228 ) | ( n39225 & ~n39228 ) ;
  assign n39230 = ( n11338 & ~n39223 ) | ( n11338 & n39229 ) | ( ~n39223 & n39229 ) ;
  assign n39231 = n9086 ^ x221 ^ x1 ;
  assign n39232 = n31205 & n39231 ;
  assign n39233 = n39232 ^ n14118 ^ n10835 ;
  assign n39234 = ( n8097 & n8845 ) | ( n8097 & n23555 ) | ( n8845 & n23555 ) ;
  assign n39235 = ( ~n17050 & n21709 ) | ( ~n17050 & n39234 ) | ( n21709 & n39234 ) ;
  assign n39236 = n39235 ^ n28810 ^ n24088 ;
  assign n39237 = n12797 & n33008 ;
  assign n39238 = n39237 ^ n16280 ^ n11684 ;
  assign n39239 = n14787 & ~n24566 ;
  assign n39240 = n39239 ^ n11197 ^ 1'b0 ;
  assign n39241 = ( ~n21399 & n25365 ) | ( ~n21399 & n39240 ) | ( n25365 & n39240 ) ;
  assign n39242 = n39241 ^ n2362 ^ 1'b0 ;
  assign n39243 = ~n39238 & n39242 ;
  assign n39244 = n11301 ^ n9930 ^ n9745 ;
  assign n39245 = n28295 ^ n22736 ^ n18560 ;
  assign n39246 = ( ~n15125 & n31564 ) | ( ~n15125 & n39245 ) | ( n31564 & n39245 ) ;
  assign n39247 = ( n2551 & n14793 ) | ( n2551 & n33014 ) | ( n14793 & n33014 ) ;
  assign n39248 = ( n10453 & n17096 ) | ( n10453 & n39247 ) | ( n17096 & n39247 ) ;
  assign n39249 = n31599 | n35051 ;
  assign n39250 = n39248 | n39249 ;
  assign n39251 = ( n21127 & n39246 ) | ( n21127 & ~n39250 ) | ( n39246 & ~n39250 ) ;
  assign n39252 = ( n10661 & n22834 ) | ( n10661 & ~n31330 ) | ( n22834 & ~n31330 ) ;
  assign n39253 = n20623 ^ n12658 ^ 1'b0 ;
  assign n39254 = n31930 & n39253 ;
  assign n39255 = ( n2799 & n14960 ) | ( n2799 & n39254 ) | ( n14960 & n39254 ) ;
  assign n39256 = n36485 & ~n39255 ;
  assign n39257 = ( n8451 & n17943 ) | ( n8451 & ~n30819 ) | ( n17943 & ~n30819 ) ;
  assign n39258 = ( ~n778 & n1544 ) | ( ~n778 & n28130 ) | ( n1544 & n28130 ) ;
  assign n39261 = n17594 ^ n8534 ^ n7927 ;
  assign n39262 = n39261 ^ n22957 ^ n21870 ;
  assign n39259 = n17651 ^ n8701 ^ n6574 ;
  assign n39260 = n39259 ^ n16774 ^ 1'b0 ;
  assign n39263 = n39262 ^ n39260 ^ n30109 ;
  assign n39264 = n7354 ^ n7227 ^ 1'b0 ;
  assign n39265 = ( n4496 & ~n11204 ) | ( n4496 & n39264 ) | ( ~n11204 & n39264 ) ;
  assign n39266 = n39265 ^ n2587 ^ n1243 ;
  assign n39267 = n2318 & n39266 ;
  assign n39268 = ( ~n2905 & n5030 ) | ( ~n2905 & n39267 ) | ( n5030 & n39267 ) ;
  assign n39269 = n34017 ^ n27297 ^ 1'b0 ;
  assign n39270 = n32975 ^ n2371 ^ 1'b0 ;
  assign n39271 = ~n4408 & n39270 ;
  assign n39272 = n16346 ^ n5200 ^ n585 ;
  assign n39273 = n39272 ^ n25317 ^ n21684 ;
  assign n39274 = ( ~n9352 & n39271 ) | ( ~n9352 & n39273 ) | ( n39271 & n39273 ) ;
  assign n39275 = n30595 ^ n13304 ^ 1'b0 ;
  assign n39276 = n20081 & n39275 ;
  assign n39277 = ( n6617 & n23854 ) | ( n6617 & ~n27142 ) | ( n23854 & ~n27142 ) ;
  assign n39278 = n24266 ^ n13719 ^ n6437 ;
  assign n39279 = n39278 ^ n26612 ^ n15557 ;
  assign n39280 = ( n12871 & n20821 ) | ( n12871 & ~n39279 ) | ( n20821 & ~n39279 ) ;
  assign n39281 = n24983 ^ n5685 ^ 1'b0 ;
  assign n39282 = ~n14185 & n39281 ;
  assign n39283 = n39282 ^ n38431 ^ n9236 ;
  assign n39290 = n16093 & ~n22957 ;
  assign n39291 = n14953 & n39290 ;
  assign n39284 = n7493 ^ n5446 ^ n2655 ;
  assign n39285 = n39284 ^ n38763 ^ n9932 ;
  assign n39286 = n33887 ^ n23518 ^ 1'b0 ;
  assign n39287 = n39285 & ~n39286 ;
  assign n39288 = n39287 ^ n14958 ^ n7211 ;
  assign n39289 = n39288 ^ n28256 ^ n4471 ;
  assign n39292 = n39291 ^ n39289 ^ n38386 ;
  assign n39293 = ( n6535 & n6619 ) | ( n6535 & ~n25253 ) | ( n6619 & ~n25253 ) ;
  assign n39294 = ( n3374 & ~n10661 ) | ( n3374 & n30248 ) | ( ~n10661 & n30248 ) ;
  assign n39295 = n24022 ^ n18658 ^ 1'b0 ;
  assign n39296 = ~n39294 & n39295 ;
  assign n39297 = n21278 & n39296 ;
  assign n39298 = ( n32301 & n39293 ) | ( n32301 & n39297 ) | ( n39293 & n39297 ) ;
  assign n39299 = ~n1457 & n39048 ;
  assign n39300 = ~n28269 & n39299 ;
  assign n39301 = n21990 | n28877 ;
  assign n39302 = n3557 | n39301 ;
  assign n39303 = n33890 ^ n26094 ^ n21353 ;
  assign n39304 = n39303 ^ n26335 ^ n3996 ;
  assign n39305 = n39304 ^ n34382 ^ n26715 ;
  assign n39309 = ( n4427 & ~n6058 ) | ( n4427 & n32449 ) | ( ~n6058 & n32449 ) ;
  assign n39306 = ( n12113 & n12830 ) | ( n12113 & ~n35243 ) | ( n12830 & ~n35243 ) ;
  assign n39307 = ( x209 & n36508 ) | ( x209 & ~n39306 ) | ( n36508 & ~n39306 ) ;
  assign n39308 = ( n2599 & n14984 ) | ( n2599 & ~n39307 ) | ( n14984 & ~n39307 ) ;
  assign n39310 = n39309 ^ n39308 ^ n14257 ;
  assign n39311 = ( n4444 & n29004 ) | ( n4444 & ~n37201 ) | ( n29004 & ~n37201 ) ;
  assign n39312 = n30385 | n39311 ;
  assign n39313 = ( n5901 & n15681 ) | ( n5901 & n25326 ) | ( n15681 & n25326 ) ;
  assign n39314 = n12869 ^ n3695 ^ 1'b0 ;
  assign n39315 = n14420 & ~n39314 ;
  assign n39316 = ~n39313 & n39315 ;
  assign n39317 = n35424 ^ n13996 ^ n7023 ;
  assign n39318 = n39317 ^ n29543 ^ x33 ;
  assign n39319 = n747 & n4066 ;
  assign n39320 = ( n18643 & ~n19079 ) | ( n18643 & n39319 ) | ( ~n19079 & n39319 ) ;
  assign n39321 = n39320 ^ n21632 ^ n8691 ;
  assign n39322 = n3129 | n5615 ;
  assign n39323 = n39322 ^ n9354 ^ 1'b0 ;
  assign n39324 = ( ~n9649 & n24546 ) | ( ~n9649 & n38461 ) | ( n24546 & n38461 ) ;
  assign n39325 = ( n21063 & n39323 ) | ( n21063 & ~n39324 ) | ( n39323 & ~n39324 ) ;
  assign n39326 = n39085 & n39325 ;
  assign n39328 = ( n8786 & ~n24548 ) | ( n8786 & n26250 ) | ( ~n24548 & n26250 ) ;
  assign n39327 = n28794 ^ n19417 ^ 1'b0 ;
  assign n39329 = n39328 ^ n39327 ^ n15176 ;
  assign n39330 = n24117 ^ n22978 ^ n18947 ;
  assign n39331 = n24649 ^ n10141 ^ n5365 ;
  assign n39332 = ( n7262 & ~n8032 ) | ( n7262 & n12815 ) | ( ~n8032 & n12815 ) ;
  assign n39333 = n34482 ^ n25399 ^ n7008 ;
  assign n39336 = n18933 ^ n17751 ^ 1'b0 ;
  assign n39334 = n14533 ^ n9441 ^ 1'b0 ;
  assign n39335 = ~n19120 & n39334 ;
  assign n39337 = n39336 ^ n39335 ^ n29105 ;
  assign n39338 = n39337 ^ n3714 ^ 1'b0 ;
  assign n39339 = n39333 & n39338 ;
  assign n39341 = ( ~n1245 & n21764 ) | ( ~n1245 & n24597 ) | ( n21764 & n24597 ) ;
  assign n39340 = n30011 | n33494 ;
  assign n39342 = n39341 ^ n39340 ^ 1'b0 ;
  assign n39343 = n14989 ^ n12879 ^ n8449 ;
  assign n39344 = n39343 ^ n14790 ^ n11867 ;
  assign n39345 = n39344 ^ n31224 ^ n28178 ;
  assign n39346 = ~n1515 & n2857 ;
  assign n39347 = n39346 ^ n25500 ^ 1'b0 ;
  assign n39348 = n17530 ^ n9415 ^ n4580 ;
  assign n39349 = n26955 & n39348 ;
  assign n39350 = ~x53 & n39349 ;
  assign n39351 = n39350 ^ n39129 ^ n38370 ;
  assign n39352 = n5227 | n14619 ;
  assign n39353 = ( n3104 & ~n11589 ) | ( n3104 & n22727 ) | ( ~n11589 & n22727 ) ;
  assign n39354 = ( n1139 & n21895 ) | ( n1139 & n23112 ) | ( n21895 & n23112 ) ;
  assign n39355 = n16760 & ~n39354 ;
  assign n39356 = n39355 ^ n13202 ^ 1'b0 ;
  assign n39357 = n37912 & ~n39356 ;
  assign n39358 = ~n9691 & n14748 ;
  assign n39359 = ~n39357 & n39358 ;
  assign n39360 = n39359 ^ n10955 ^ n9997 ;
  assign n39361 = ( n418 & n39353 ) | ( n418 & ~n39360 ) | ( n39353 & ~n39360 ) ;
  assign n39362 = n38642 ^ n12893 ^ 1'b0 ;
  assign n39363 = ( n13052 & n28358 ) | ( n13052 & n39362 ) | ( n28358 & n39362 ) ;
  assign n39364 = n36754 ^ n7003 ^ n5998 ;
  assign n39365 = ( ~n11624 & n11781 ) | ( ~n11624 & n39364 ) | ( n11781 & n39364 ) ;
  assign n39366 = ( ~n20251 & n22833 ) | ( ~n20251 & n32573 ) | ( n22833 & n32573 ) ;
  assign n39367 = n39366 ^ n33708 ^ n22772 ;
  assign n39368 = n25464 ^ n13711 ^ 1'b0 ;
  assign n39369 = n39368 ^ n18364 ^ n15526 ;
  assign n39370 = n30345 ^ n22187 ^ n572 ;
  assign n39371 = n22785 ^ n18496 ^ 1'b0 ;
  assign n39372 = n39370 | n39371 ;
  assign n39375 = n29505 ^ n6324 ^ x57 ;
  assign n39376 = n39375 ^ n11274 ^ 1'b0 ;
  assign n39377 = n11742 & ~n39376 ;
  assign n39373 = n9539 & n32457 ;
  assign n39374 = n39373 ^ n21326 ^ 1'b0 ;
  assign n39378 = n39377 ^ n39374 ^ n32926 ;
  assign n39379 = n16222 ^ n15079 ^ n8683 ;
  assign n39380 = ( ~n3347 & n15405 ) | ( ~n3347 & n39379 ) | ( n15405 & n39379 ) ;
  assign n39381 = n6026 ^ n3954 ^ n1595 ;
  assign n39382 = ~n5244 & n19080 ;
  assign n39383 = ~n2550 & n39382 ;
  assign n39384 = ( n17682 & n39381 ) | ( n17682 & n39383 ) | ( n39381 & n39383 ) ;
  assign n39389 = n24613 ^ n12384 ^ n3610 ;
  assign n39385 = ( n4398 & n9517 ) | ( n4398 & n12705 ) | ( n9517 & n12705 ) ;
  assign n39386 = n16459 & ~n22141 ;
  assign n39387 = ~n39385 & n39386 ;
  assign n39388 = n39387 ^ n5699 ^ 1'b0 ;
  assign n39390 = n39389 ^ n39388 ^ n33002 ;
  assign n39393 = x168 & ~n22274 ;
  assign n39394 = n30539 & n39393 ;
  assign n39391 = n8525 | n13677 ;
  assign n39392 = n5673 | n39391 ;
  assign n39395 = n39394 ^ n39392 ^ n10586 ;
  assign n39396 = n18710 | n31445 ;
  assign n39397 = n21016 & n37316 ;
  assign n39398 = n39397 ^ n23613 ^ 1'b0 ;
  assign n39399 = n27157 ^ n13261 ^ n11577 ;
  assign n39400 = n33099 ^ n21471 ^ 1'b0 ;
  assign n39401 = n27024 ^ n11651 ^ 1'b0 ;
  assign n39402 = n10604 ^ n8977 ^ n2686 ;
  assign n39403 = ( n707 & n9642 ) | ( n707 & ~n13905 ) | ( n9642 & ~n13905 ) ;
  assign n39404 = n22358 & n27575 ;
  assign n39405 = ~n7613 & n39404 ;
  assign n39406 = ( n6393 & n10619 ) | ( n6393 & n13345 ) | ( n10619 & n13345 ) ;
  assign n39407 = ( n39403 & n39405 ) | ( n39403 & n39406 ) | ( n39405 & n39406 ) ;
  assign n39408 = n2457 | n18042 ;
  assign n39409 = n23591 | n39408 ;
  assign n39410 = n17059 ^ n6393 ^ n2095 ;
  assign n39411 = n14619 & n39410 ;
  assign n39412 = n39411 ^ n27686 ^ 1'b0 ;
  assign n39413 = n13627 & n14031 ;
  assign n39414 = n39413 ^ n33442 ^ 1'b0 ;
  assign n39415 = n39414 ^ n27826 ^ n8794 ;
  assign n39416 = n6328 | n23875 ;
  assign n39417 = ( ~n4320 & n21635 ) | ( ~n4320 & n30731 ) | ( n21635 & n30731 ) ;
  assign n39418 = ( n17503 & n39416 ) | ( n17503 & ~n39417 ) | ( n39416 & ~n39417 ) ;
  assign n39419 = ( n30667 & ~n32783 ) | ( n30667 & n39418 ) | ( ~n32783 & n39418 ) ;
  assign n39420 = n34148 ^ n13877 ^ n4395 ;
  assign n39423 = ~n20763 & n35909 ;
  assign n39421 = n3142 & ~n19102 ;
  assign n39422 = n39421 ^ n15522 ^ n14315 ;
  assign n39424 = n39423 ^ n39422 ^ n929 ;
  assign n39425 = n18865 | n31048 ;
  assign n39426 = n17496 | n39425 ;
  assign n39427 = n20755 ^ n5328 ^ n4638 ;
  assign n39428 = ( n535 & n9596 ) | ( n535 & ~n39427 ) | ( n9596 & ~n39427 ) ;
  assign n39429 = ( n12701 & ~n14819 ) | ( n12701 & n24791 ) | ( ~n14819 & n24791 ) ;
  assign n39430 = n39429 ^ n5419 ^ n903 ;
  assign n39431 = n39430 ^ n30116 ^ n8845 ;
  assign n39432 = ( n369 & n28006 ) | ( n369 & n39431 ) | ( n28006 & n39431 ) ;
  assign n39433 = ( ~n39426 & n39428 ) | ( ~n39426 & n39432 ) | ( n39428 & n39432 ) ;
  assign n39434 = n39385 ^ n28976 ^ n3983 ;
  assign n39435 = n9645 & ~n25283 ;
  assign n39436 = n15413 | n35036 ;
  assign n39437 = n19910 | n39436 ;
  assign n39438 = n34270 ^ n22033 ^ 1'b0 ;
  assign n39439 = n39438 ^ n30901 ^ n4639 ;
  assign n39440 = ( n26424 & n27778 ) | ( n26424 & n36226 ) | ( n27778 & n36226 ) ;
  assign n39441 = ( n2176 & n8281 ) | ( n2176 & ~n15097 ) | ( n8281 & ~n15097 ) ;
  assign n39442 = n20593 & n39441 ;
  assign n39443 = ( n17329 & ~n21879 ) | ( n17329 & n39442 ) | ( ~n21879 & n39442 ) ;
  assign n39444 = n34254 ^ n18174 ^ n909 ;
  assign n39445 = n26684 ^ n2276 ^ 1'b0 ;
  assign n39446 = n17363 ^ n15086 ^ n9435 ;
  assign n39447 = ( n11064 & n21773 ) | ( n11064 & ~n39446 ) | ( n21773 & ~n39446 ) ;
  assign n39448 = n13050 & n17381 ;
  assign n39449 = ~n19839 & n39448 ;
  assign n39450 = ( n37529 & ~n39447 ) | ( n37529 & n39449 ) | ( ~n39447 & n39449 ) ;
  assign n39451 = n13214 ^ n539 ^ 1'b0 ;
  assign n39452 = n39451 ^ n12704 ^ n864 ;
  assign n39453 = n17813 ^ n14515 ^ 1'b0 ;
  assign n39454 = n32236 ^ n21258 ^ n5693 ;
  assign n39455 = n39454 ^ n22429 ^ n11399 ;
  assign n39456 = n39455 ^ n13339 ^ n11486 ;
  assign n39457 = n23949 ^ n20821 ^ 1'b0 ;
  assign n39458 = n11609 & n39457 ;
  assign n39460 = n9899 ^ n347 ^ 1'b0 ;
  assign n39459 = n14524 | n16829 ;
  assign n39461 = n39460 ^ n39459 ^ n36323 ;
  assign n39462 = n39458 | n39461 ;
  assign n39467 = n33597 ^ n13867 ^ n3509 ;
  assign n39463 = n13983 ^ n10125 ^ n1218 ;
  assign n39464 = ~n12589 & n16952 ;
  assign n39465 = ~n39463 & n39464 ;
  assign n39466 = ( n1007 & ~n1268 ) | ( n1007 & n39465 ) | ( ~n1268 & n39465 ) ;
  assign n39468 = n39467 ^ n39466 ^ 1'b0 ;
  assign n39469 = n39468 ^ n6959 ^ 1'b0 ;
  assign n39470 = n16329 ^ n8127 ^ n1617 ;
  assign n39471 = ( n4002 & n14383 ) | ( n4002 & ~n24048 ) | ( n14383 & ~n24048 ) ;
  assign n39472 = n30849 ^ n10012 ^ x39 ;
  assign n39473 = n39472 ^ n25141 ^ 1'b0 ;
  assign n39474 = ( ~n32098 & n39471 ) | ( ~n32098 & n39473 ) | ( n39471 & n39473 ) ;
  assign n39475 = n21997 ^ n21808 ^ 1'b0 ;
  assign n39476 = n27046 ^ n10900 ^ n10057 ;
  assign n39477 = n22788 ^ n5098 ^ n4934 ;
  assign n39478 = n39477 ^ n20684 ^ n3841 ;
  assign n39479 = ( n20018 & ~n27119 ) | ( n20018 & n39478 ) | ( ~n27119 & n39478 ) ;
  assign n39480 = ( n35597 & ~n39476 ) | ( n35597 & n39479 ) | ( ~n39476 & n39479 ) ;
  assign n39481 = n9401 & ~n33088 ;
  assign n39482 = n4760 | n8990 ;
  assign n39483 = n39482 ^ n16109 ^ 1'b0 ;
  assign n39484 = ( n19412 & n35513 ) | ( n19412 & ~n39483 ) | ( n35513 & ~n39483 ) ;
  assign n39485 = ~n3090 & n36017 ;
  assign n39494 = n12740 ^ n11521 ^ n2114 ;
  assign n39490 = n25442 | n28399 ;
  assign n39491 = n39490 ^ n29400 ^ 1'b0 ;
  assign n39486 = n35831 ^ n13699 ^ n333 ;
  assign n39487 = ( n23258 & ~n31202 ) | ( n23258 & n39486 ) | ( ~n31202 & n39486 ) ;
  assign n39488 = ( x219 & ~n22382 ) | ( x219 & n29639 ) | ( ~n22382 & n29639 ) ;
  assign n39489 = ( ~n8320 & n39487 ) | ( ~n8320 & n39488 ) | ( n39487 & n39488 ) ;
  assign n39492 = n39491 ^ n39489 ^ n23564 ;
  assign n39493 = ~n19912 & n39492 ;
  assign n39495 = n39494 ^ n39493 ^ 1'b0 ;
  assign n39496 = n14278 ^ n14044 ^ n12879 ;
  assign n39497 = n39496 ^ n12551 ^ n9058 ;
  assign n39498 = n27535 ^ n17132 ^ n9352 ;
  assign n39499 = n39498 ^ n9125 ^ n9069 ;
  assign n39500 = n18879 ^ n9805 ^ 1'b0 ;
  assign n39501 = ( n16181 & n17821 ) | ( n16181 & n37455 ) | ( n17821 & n37455 ) ;
  assign n39502 = n16339 ^ n4358 ^ x61 ;
  assign n39503 = ( n16607 & n39501 ) | ( n16607 & n39502 ) | ( n39501 & n39502 ) ;
  assign n39504 = n17898 ^ n13352 ^ 1'b0 ;
  assign n39505 = n17576 & n36848 ;
  assign n39506 = n39505 ^ n7521 ^ 1'b0 ;
  assign n39507 = n39504 & n39506 ;
  assign n39508 = n6172 & n24865 ;
  assign n39509 = n39508 ^ n7692 ^ 1'b0 ;
  assign n39510 = n25401 ^ n8765 ^ 1'b0 ;
  assign n39511 = ~n32533 & n39510 ;
  assign n39512 = ( n4109 & ~n7567 ) | ( n4109 & n39511 ) | ( ~n7567 & n39511 ) ;
  assign n39513 = n28735 ^ n11458 ^ n5787 ;
  assign n39514 = n6572 ^ n5912 ^ n1839 ;
  assign n39515 = n39513 & n39514 ;
  assign n39516 = n36527 & n37595 ;
  assign n39517 = ( n16534 & n27858 ) | ( n16534 & n38058 ) | ( n27858 & n38058 ) ;
  assign n39518 = ( n12491 & n20752 ) | ( n12491 & ~n20812 ) | ( n20752 & ~n20812 ) ;
  assign n39519 = n17873 ^ n2905 ^ 1'b0 ;
  assign n39520 = n25401 ^ n7627 ^ n6454 ;
  assign n39521 = n39519 | n39520 ;
  assign n39522 = ~n11081 & n23292 ;
  assign n39523 = n39522 ^ n21464 ^ 1'b0 ;
  assign n39524 = n3408 ^ n3122 ^ 1'b0 ;
  assign n39525 = n23655 & n39524 ;
  assign n39526 = n15512 | n16148 ;
  assign n39527 = n39526 ^ n2887 ^ 1'b0 ;
  assign n39528 = n8983 | n19252 ;
  assign n39529 = n39527 | n39528 ;
  assign n39530 = ( n6891 & ~n16533 ) | ( n6891 & n23991 ) | ( ~n16533 & n23991 ) ;
  assign n39531 = n22462 ^ n4187 ^ n757 ;
  assign n39532 = n39531 ^ n14649 ^ n9164 ;
  assign n39533 = ( ~n340 & n20052 ) | ( ~n340 & n39532 ) | ( n20052 & n39532 ) ;
  assign n39534 = ( n16170 & n39530 ) | ( n16170 & n39533 ) | ( n39530 & n39533 ) ;
  assign n39535 = n20298 ^ n14677 ^ 1'b0 ;
  assign n39536 = ( x41 & ~n12708 ) | ( x41 & n12830 ) | ( ~n12708 & n12830 ) ;
  assign n39537 = n39536 ^ n28949 ^ 1'b0 ;
  assign n39538 = n1496 & ~n31148 ;
  assign n39539 = ~n14554 & n39538 ;
  assign n39540 = n16616 ^ n11400 ^ n794 ;
  assign n39541 = n8536 & n39540 ;
  assign n39542 = n21967 & n39541 ;
  assign n39544 = n2072 & ~n6740 ;
  assign n39545 = n39544 ^ n8340 ^ 1'b0 ;
  assign n39543 = n13022 ^ n6330 ^ 1'b0 ;
  assign n39546 = n39545 ^ n39543 ^ n7596 ;
  assign n39547 = ( n12683 & n30372 ) | ( n12683 & n34436 ) | ( n30372 & n34436 ) ;
  assign n39548 = n37695 ^ n27432 ^ 1'b0 ;
  assign n39549 = n6570 & n8186 ;
  assign n39550 = n9907 & n39549 ;
  assign n39551 = n39550 ^ n36040 ^ n10831 ;
  assign n39552 = ( n4836 & n6549 ) | ( n4836 & n9040 ) | ( n6549 & n9040 ) ;
  assign n39553 = n39552 ^ n39223 ^ 1'b0 ;
  assign n39554 = ( n23065 & n39551 ) | ( n23065 & n39553 ) | ( n39551 & n39553 ) ;
  assign n39556 = n24172 ^ n12228 ^ n7821 ;
  assign n39555 = n35460 ^ n3112 ^ 1'b0 ;
  assign n39557 = n39556 ^ n39555 ^ n25244 ;
  assign n39558 = n15052 ^ n8953 ^ n1988 ;
  assign n39559 = n21726 | n24723 ;
  assign n39560 = n10666 ^ n7556 ^ n3186 ;
  assign n39561 = ( n7793 & n35599 ) | ( n7793 & ~n39560 ) | ( n35599 & ~n39560 ) ;
  assign n39562 = n39561 ^ n5854 ^ 1'b0 ;
  assign n39563 = n34802 | n39562 ;
  assign n39564 = n39563 ^ n30835 ^ n3242 ;
  assign n39565 = n2003 & ~n3629 ;
  assign n39566 = n39565 ^ n24396 ^ 1'b0 ;
  assign n39567 = n39566 ^ n13473 ^ n2676 ;
  assign n39568 = ( ~n15897 & n16955 ) | ( ~n15897 & n39567 ) | ( n16955 & n39567 ) ;
  assign n39569 = ~n9649 & n32366 ;
  assign n39570 = ~n8034 & n24914 ;
  assign n39571 = ~n39569 & n39570 ;
  assign n39572 = n9523 & n39571 ;
  assign n39573 = n37454 ^ n22137 ^ n10762 ;
  assign n39574 = ( n13796 & ~n16898 ) | ( n13796 & n39573 ) | ( ~n16898 & n39573 ) ;
  assign n39575 = n20615 & n33788 ;
  assign n39576 = n32608 ^ n16309 ^ n4018 ;
  assign n39577 = n19604 ^ n11781 ^ n9283 ;
  assign n39578 = n23469 & ~n39577 ;
  assign n39579 = ~n22608 & n39578 ;
  assign n39580 = n15523 ^ n13902 ^ 1'b0 ;
  assign n39581 = n39580 ^ n12643 ^ n3429 ;
  assign n39582 = n20073 ^ n1986 ^ 1'b0 ;
  assign n39583 = ( n3756 & n12501 ) | ( n3756 & n39582 ) | ( n12501 & n39582 ) ;
  assign n39584 = n39583 ^ n4190 ^ 1'b0 ;
  assign n39585 = ~n39581 & n39584 ;
  assign n39588 = n21464 ^ n11852 ^ n8366 ;
  assign n39589 = ( ~n6665 & n8291 ) | ( ~n6665 & n39588 ) | ( n8291 & n39588 ) ;
  assign n39590 = ( ~n5782 & n10173 ) | ( ~n5782 & n39589 ) | ( n10173 & n39589 ) ;
  assign n39586 = n36206 ^ n3358 ^ 1'b0 ;
  assign n39587 = ( n7395 & n17014 ) | ( n7395 & n39586 ) | ( n17014 & n39586 ) ;
  assign n39591 = n39590 ^ n39587 ^ n25514 ;
  assign n39592 = n20893 & n24689 ;
  assign n39593 = ( ~n1819 & n2420 ) | ( ~n1819 & n35148 ) | ( n2420 & n35148 ) ;
  assign n39594 = ( n9885 & n10011 ) | ( n9885 & n39593 ) | ( n10011 & n39593 ) ;
  assign n39595 = ( n11755 & n39592 ) | ( n11755 & n39594 ) | ( n39592 & n39594 ) ;
  assign n39596 = ( n7667 & n21402 ) | ( n7667 & n32293 ) | ( n21402 & n32293 ) ;
  assign n39597 = ( n7050 & n31438 ) | ( n7050 & n32140 ) | ( n31438 & n32140 ) ;
  assign n39598 = n39597 ^ n28470 ^ n1844 ;
  assign n39599 = n39598 ^ n36545 ^ n23690 ;
  assign n39600 = n19189 ^ n5786 ^ 1'b0 ;
  assign n39601 = ( n3246 & ~n28235 ) | ( n3246 & n39600 ) | ( ~n28235 & n39600 ) ;
  assign n39602 = ( n21759 & ~n24661 ) | ( n21759 & n28625 ) | ( ~n24661 & n28625 ) ;
  assign n39603 = ( n6464 & n33507 ) | ( n6464 & ~n39602 ) | ( n33507 & ~n39602 ) ;
  assign n39604 = n20184 ^ n12022 ^ n8005 ;
  assign n39605 = ~n17520 & n39604 ;
  assign n39606 = ~n38212 & n39605 ;
  assign n39607 = n22010 ^ n8581 ^ n7402 ;
  assign n39610 = ( n9870 & n15482 ) | ( n9870 & n28124 ) | ( n15482 & n28124 ) ;
  assign n39609 = n8333 | n19924 ;
  assign n39608 = n2954 & n9437 ;
  assign n39611 = n39610 ^ n39609 ^ n39608 ;
  assign n39612 = n31455 ^ n25772 ^ 1'b0 ;
  assign n39616 = n5442 | n7728 ;
  assign n39613 = n18390 ^ n18175 ^ n4742 ;
  assign n39614 = ~n14523 & n39613 ;
  assign n39615 = n39614 ^ n17910 ^ 1'b0 ;
  assign n39617 = n39616 ^ n39615 ^ n15401 ;
  assign n39618 = ( n4686 & ~n12353 ) | ( n4686 & n31723 ) | ( ~n12353 & n31723 ) ;
  assign n39619 = n39618 ^ n30020 ^ 1'b0 ;
  assign n39620 = n36765 ^ n23702 ^ n15261 ;
  assign n39621 = n39620 ^ n33394 ^ n14921 ;
  assign n39622 = n19607 ^ n18724 ^ n10440 ;
  assign n39623 = n27638 ^ n4862 ^ n857 ;
  assign n39624 = ( n814 & ~n8785 ) | ( n814 & n39623 ) | ( ~n8785 & n39623 ) ;
  assign n39625 = n25179 ^ n14318 ^ n4020 ;
  assign n39626 = ( n36950 & n39624 ) | ( n36950 & ~n39625 ) | ( n39624 & ~n39625 ) ;
  assign n39627 = n39626 ^ n22821 ^ 1'b0 ;
  assign n39631 = ( n8688 & n8722 ) | ( n8688 & n9164 ) | ( n8722 & n9164 ) ;
  assign n39628 = ~n4070 & n8920 ;
  assign n39629 = n39628 ^ n16600 ^ n5205 ;
  assign n39630 = n39629 ^ n31029 ^ n11383 ;
  assign n39632 = n39631 ^ n39630 ^ n26013 ;
  assign n39633 = n7103 & ~n20540 ;
  assign n39634 = n39633 ^ n36307 ^ 1'b0 ;
  assign n39635 = ~n5624 & n5799 ;
  assign n39636 = n5127 & n39635 ;
  assign n39637 = n21904 & n39636 ;
  assign n39638 = ( n2606 & n9976 ) | ( n2606 & ~n13283 ) | ( n9976 & ~n13283 ) ;
  assign n39639 = n34248 & n39638 ;
  assign n39640 = ( n7542 & n28830 ) | ( n7542 & n34998 ) | ( n28830 & n34998 ) ;
  assign n39642 = ~n1955 & n10224 ;
  assign n39643 = n39642 ^ n31740 ^ 1'b0 ;
  assign n39641 = ~n18503 & n21444 ;
  assign n39644 = n39643 ^ n39641 ^ n17030 ;
  assign n39645 = n39644 ^ n38506 ^ n35708 ;
  assign n39646 = n39645 ^ n28970 ^ n16768 ;
  assign n39647 = ( n7392 & ~n11594 ) | ( n7392 & n37971 ) | ( ~n11594 & n37971 ) ;
  assign n39648 = ( n911 & n7507 ) | ( n911 & n12090 ) | ( n7507 & n12090 ) ;
  assign n39649 = ( n3889 & n4809 ) | ( n3889 & n39648 ) | ( n4809 & n39648 ) ;
  assign n39650 = ( ~n1629 & n11467 ) | ( ~n1629 & n18433 ) | ( n11467 & n18433 ) ;
  assign n39651 = ( n21328 & n39649 ) | ( n21328 & n39650 ) | ( n39649 & n39650 ) ;
  assign n39656 = n2533 & ~n6665 ;
  assign n39654 = ~n3696 & n37201 ;
  assign n39653 = n4321 | n10936 ;
  assign n39652 = n3763 | n25019 ;
  assign n39655 = n39654 ^ n39653 ^ n39652 ;
  assign n39657 = n39656 ^ n39655 ^ 1'b0 ;
  assign n39658 = n31776 ^ n14374 ^ 1'b0 ;
  assign n39659 = n16762 ^ n7618 ^ n7388 ;
  assign n39660 = ~n983 & n39659 ;
  assign n39661 = ( ~n5189 & n10544 ) | ( ~n5189 & n22824 ) | ( n10544 & n22824 ) ;
  assign n39662 = n39661 ^ n14667 ^ 1'b0 ;
  assign n39663 = n12926 ^ n7444 ^ n3399 ;
  assign n39664 = ( ~n3118 & n6942 ) | ( ~n3118 & n30720 ) | ( n6942 & n30720 ) ;
  assign n39665 = ( n4531 & n25844 ) | ( n4531 & n39664 ) | ( n25844 & n39664 ) ;
  assign n39666 = n39665 ^ n29717 ^ n2851 ;
  assign n39667 = n39666 ^ n34587 ^ n24022 ;
  assign n39668 = ( n3064 & ~n4008 ) | ( n3064 & n21341 ) | ( ~n4008 & n21341 ) ;
  assign n39670 = n32649 ^ n24148 ^ n11470 ;
  assign n39669 = ~n14718 & n16667 ;
  assign n39671 = n39670 ^ n39669 ^ 1'b0 ;
  assign n39672 = n10219 ^ n3112 ^ 1'b0 ;
  assign n39673 = n16088 & n39672 ;
  assign n39674 = ( n16780 & n17566 ) | ( n16780 & ~n39673 ) | ( n17566 & ~n39673 ) ;
  assign n39675 = ( ~n1793 & n13558 ) | ( ~n1793 & n31203 ) | ( n13558 & n31203 ) ;
  assign n39676 = n15881 ^ n3777 ^ 1'b0 ;
  assign n39677 = n39676 ^ n22504 ^ 1'b0 ;
  assign n39678 = ( ~n39674 & n39675 ) | ( ~n39674 & n39677 ) | ( n39675 & n39677 ) ;
  assign n39679 = n5461 ^ n4170 ^ n2135 ;
  assign n39680 = ~n2020 & n39679 ;
  assign n39681 = n36692 ^ n8844 ^ 1'b0 ;
  assign n39682 = ( n1642 & ~n18896 ) | ( n1642 & n37603 ) | ( ~n18896 & n37603 ) ;
  assign n39683 = n16270 ^ n12059 ^ n1246 ;
  assign n39684 = ( n749 & n2367 ) | ( n749 & n5694 ) | ( n2367 & n5694 ) ;
  assign n39685 = ( ~n12384 & n39683 ) | ( ~n12384 & n39684 ) | ( n39683 & n39684 ) ;
  assign n39686 = ( ~n29739 & n30380 ) | ( ~n29739 & n39685 ) | ( n30380 & n39685 ) ;
  assign n39687 = ( ~n26222 & n31484 ) | ( ~n26222 & n36890 ) | ( n31484 & n36890 ) ;
  assign n39688 = ( ~n10334 & n16315 ) | ( ~n10334 & n29577 ) | ( n16315 & n29577 ) ;
  assign n39689 = ( n24279 & n39687 ) | ( n24279 & n39688 ) | ( n39687 & n39688 ) ;
  assign n39690 = ~n3165 & n11660 ;
  assign n39691 = n4165 & n39690 ;
  assign n39692 = ( n18896 & n26057 ) | ( n18896 & n39691 ) | ( n26057 & n39691 ) ;
  assign n39693 = ( n12691 & n19426 ) | ( n12691 & n39692 ) | ( n19426 & n39692 ) ;
  assign n39694 = n30186 ^ n18742 ^ n10614 ;
  assign n39695 = ( ~x33 & n17085 ) | ( ~x33 & n32675 ) | ( n17085 & n32675 ) ;
  assign n39696 = ~n7381 & n22907 ;
  assign n39697 = n39696 ^ n5623 ^ 1'b0 ;
  assign n39698 = n7236 & n24660 ;
  assign n39699 = n30727 ^ n13577 ^ 1'b0 ;
  assign n39700 = n30984 & n39699 ;
  assign n39701 = n39700 ^ n33336 ^ n24788 ;
  assign n39702 = ( n4521 & n29496 ) | ( n4521 & n39701 ) | ( n29496 & n39701 ) ;
  assign n39703 = n35066 ^ n9068 ^ x201 ;
  assign n39704 = n11782 & ~n19871 ;
  assign n39705 = n39704 ^ n37705 ^ n16842 ;
  assign n39706 = n39705 ^ n4280 ^ n2161 ;
  assign n39707 = ( n7514 & n20677 ) | ( n7514 & ~n38173 ) | ( n20677 & ~n38173 ) ;
  assign n39708 = n1249 & n6890 ;
  assign n39709 = ~n5168 & n39708 ;
  assign n39710 = ( n8949 & n14914 ) | ( n8949 & n39709 ) | ( n14914 & n39709 ) ;
  assign n39711 = ( n3578 & n6913 ) | ( n3578 & ~n23907 ) | ( n6913 & ~n23907 ) ;
  assign n39712 = ( n39707 & n39710 ) | ( n39707 & n39711 ) | ( n39710 & n39711 ) ;
  assign n39713 = ( x70 & n10031 ) | ( x70 & ~n28087 ) | ( n10031 & ~n28087 ) ;
  assign n39714 = ( n869 & n3207 ) | ( n869 & n10563 ) | ( n3207 & n10563 ) ;
  assign n39715 = n24667 ^ n15526 ^ n2392 ;
  assign n39716 = ( ~n5510 & n33070 ) | ( ~n5510 & n39715 ) | ( n33070 & n39715 ) ;
  assign n39717 = ( ~n39713 & n39714 ) | ( ~n39713 & n39716 ) | ( n39714 & n39716 ) ;
  assign n39718 = n460 | n19207 ;
  assign n39719 = n39718 ^ n17487 ^ 1'b0 ;
  assign n39720 = n4533 | n20138 ;
  assign n39721 = n35386 | n39720 ;
  assign n39722 = n38563 ^ n33272 ^ 1'b0 ;
  assign n39723 = ( n11858 & ~n17351 ) | ( n11858 & n35407 ) | ( ~n17351 & n35407 ) ;
  assign n39724 = n39723 ^ n19043 ^ n441 ;
  assign n39725 = n30027 ^ n27161 ^ n12508 ;
  assign n39726 = n29365 ^ n18672 ^ 1'b0 ;
  assign n39727 = n25128 | n39726 ;
  assign n39728 = n39727 ^ n25989 ^ n25102 ;
  assign n39729 = n39728 ^ n12218 ^ n1195 ;
  assign n39730 = ( n4884 & ~n17295 ) | ( n4884 & n28511 ) | ( ~n17295 & n28511 ) ;
  assign n39731 = ( n3990 & ~n6138 ) | ( n3990 & n11136 ) | ( ~n6138 & n11136 ) ;
  assign n39732 = n39731 ^ n2954 ^ 1'b0 ;
  assign n39737 = n1349 & n8704 ;
  assign n39738 = n17421 & n39737 ;
  assign n39733 = n14895 ^ n10249 ^ n10186 ;
  assign n39734 = ( n18503 & ~n23014 ) | ( n18503 & n39733 ) | ( ~n23014 & n39733 ) ;
  assign n39735 = n39734 ^ n12769 ^ 1'b0 ;
  assign n39736 = n25137 | n39735 ;
  assign n39739 = n39738 ^ n39736 ^ n26328 ;
  assign n39740 = ~n9364 & n11684 ;
  assign n39741 = ( ~n30691 & n30953 ) | ( ~n30691 & n39740 ) | ( n30953 & n39740 ) ;
  assign n39743 = ~n22811 & n39247 ;
  assign n39742 = n5430 & ~n7825 ;
  assign n39744 = n39743 ^ n39742 ^ 1'b0 ;
  assign n39745 = ~n3003 & n7482 ;
  assign n39746 = n39745 ^ n7801 ^ 1'b0 ;
  assign n39747 = n30832 ^ n11053 ^ 1'b0 ;
  assign n39748 = ~n39746 & n39747 ;
  assign n39749 = n11915 & ~n29403 ;
  assign n39750 = n15640 & n18673 ;
  assign n39751 = n39750 ^ n12537 ^ n10643 ;
  assign n39752 = ( ~n8325 & n11353 ) | ( ~n8325 & n24386 ) | ( n11353 & n24386 ) ;
  assign n39753 = ( ~x226 & n13009 ) | ( ~x226 & n25192 ) | ( n13009 & n25192 ) ;
  assign n39754 = ( n4049 & n39752 ) | ( n4049 & ~n39753 ) | ( n39752 & ~n39753 ) ;
  assign n39755 = n22472 & ~n31219 ;
  assign n39756 = n17976 & n39755 ;
  assign n39757 = n9268 & n22165 ;
  assign n39758 = n39757 ^ n26805 ^ 1'b0 ;
  assign n39759 = n11845 & ~n39758 ;
  assign n39760 = ( n14937 & n39756 ) | ( n14937 & ~n39759 ) | ( n39756 & ~n39759 ) ;
  assign n39761 = ~n8581 & n8692 ;
  assign n39762 = n39761 ^ n23311 ^ 1'b0 ;
  assign n39763 = ( n11715 & n28427 ) | ( n11715 & ~n39762 ) | ( n28427 & ~n39762 ) ;
  assign n39764 = ( n1863 & n7636 ) | ( n1863 & ~n21279 ) | ( n7636 & ~n21279 ) ;
  assign n39765 = n39764 ^ n22036 ^ 1'b0 ;
  assign n39766 = n39763 | n39765 ;
  assign n39767 = n8977 & ~n16890 ;
  assign n39768 = n31909 ^ n10254 ^ 1'b0 ;
  assign n39769 = n20909 ^ n12536 ^ n5187 ;
  assign n39770 = n4410 & ~n7708 ;
  assign n39771 = n39770 ^ n27070 ^ 1'b0 ;
  assign n39772 = n11864 & ~n37993 ;
  assign n39773 = n10929 & n39772 ;
  assign n39774 = ( n28410 & n39771 ) | ( n28410 & ~n39773 ) | ( n39771 & ~n39773 ) ;
  assign n39775 = ~n6113 & n12729 ;
  assign n39776 = ~n5824 & n39775 ;
  assign n39777 = ( n26709 & ~n37694 ) | ( n26709 & n39776 ) | ( ~n37694 & n39776 ) ;
  assign n39778 = n39161 ^ n33292 ^ n17466 ;
  assign n39779 = ( n27933 & n32406 ) | ( n27933 & n39778 ) | ( n32406 & n39778 ) ;
  assign n39780 = n13120 | n16040 ;
  assign n39781 = ~n1208 & n10056 ;
  assign n39782 = ~n39780 & n39781 ;
  assign n39783 = ( x54 & ~n32764 ) | ( x54 & n39782 ) | ( ~n32764 & n39782 ) ;
  assign n39784 = n28178 ^ n6673 ^ 1'b0 ;
  assign n39785 = ( ~n35380 & n39248 ) | ( ~n35380 & n39784 ) | ( n39248 & n39784 ) ;
  assign n39786 = n20976 ^ n10425 ^ 1'b0 ;
  assign n39787 = ~n19457 & n39786 ;
  assign n39788 = n807 | n35073 ;
  assign n39789 = n39788 ^ n22201 ^ 1'b0 ;
  assign n39790 = n39787 & ~n39789 ;
  assign n39791 = n39790 ^ n2391 ^ 1'b0 ;
  assign n39792 = n31580 ^ n27692 ^ n8047 ;
  assign n39793 = n24710 ^ n7430 ^ 1'b0 ;
  assign n39794 = n24101 & n39793 ;
  assign n39795 = n39792 & n39794 ;
  assign n39796 = ( n403 & ~n4472 ) | ( n403 & n29558 ) | ( ~n4472 & n29558 ) ;
  assign n39797 = n39796 ^ n30382 ^ n2878 ;
  assign n39798 = ( ~n2647 & n14896 ) | ( ~n2647 & n28498 ) | ( n14896 & n28498 ) ;
  assign n39801 = ( n2676 & ~n4071 ) | ( n2676 & n17549 ) | ( ~n4071 & n17549 ) ;
  assign n39802 = ( ~n18781 & n38905 ) | ( ~n18781 & n39801 ) | ( n38905 & n39801 ) ;
  assign n39799 = ( n1217 & ~n14186 ) | ( n1217 & n38279 ) | ( ~n14186 & n38279 ) ;
  assign n39800 = n39799 ^ n38211 ^ n2005 ;
  assign n39803 = n39802 ^ n39800 ^ n406 ;
  assign n39804 = ( n8117 & ~n22453 ) | ( n8117 & n23859 ) | ( ~n22453 & n23859 ) ;
  assign n39805 = n39804 ^ n11217 ^ n1560 ;
  assign n39806 = n21258 | n26582 ;
  assign n39807 = n39805 | n39806 ;
  assign n39808 = n31081 ^ n13725 ^ n11523 ;
  assign n39810 = ( n3157 & ~n22744 ) | ( n3157 & n22998 ) | ( ~n22744 & n22998 ) ;
  assign n39809 = n38935 ^ n19459 ^ n6955 ;
  assign n39811 = n39810 ^ n39809 ^ n3735 ;
  assign n39812 = n14140 ^ n2705 ^ 1'b0 ;
  assign n39813 = n1935 | n39812 ;
  assign n39814 = ~n7867 & n39813 ;
  assign n39815 = n36031 ^ n21359 ^ 1'b0 ;
  assign n39816 = n13333 ^ n7055 ^ 1'b0 ;
  assign n39817 = n39816 ^ n19256 ^ n13696 ;
  assign n39820 = n7323 ^ n3888 ^ n3058 ;
  assign n39818 = ~n18624 & n30045 ;
  assign n39819 = n39818 ^ n1293 ^ 1'b0 ;
  assign n39821 = n39820 ^ n39819 ^ n8590 ;
  assign n39822 = n39821 ^ n5053 ^ 1'b0 ;
  assign n39823 = n938 | n4463 ;
  assign n39824 = ( n12531 & ~n24179 ) | ( n12531 & n31383 ) | ( ~n24179 & n31383 ) ;
  assign n39825 = ~n11565 & n39527 ;
  assign n39826 = ( n2392 & n13301 ) | ( n2392 & ~n39825 ) | ( n13301 & ~n39825 ) ;
  assign n39827 = ~n39824 & n39826 ;
  assign n39828 = ~n39823 & n39827 ;
  assign n39829 = n16972 ^ n9684 ^ n6232 ;
  assign n39830 = n12050 & n39829 ;
  assign n39831 = ( ~n16375 & n20322 ) | ( ~n16375 & n35648 ) | ( n20322 & n35648 ) ;
  assign n39832 = n39831 ^ n35388 ^ n24177 ;
  assign n39833 = n11683 ^ n3867 ^ 1'b0 ;
  assign n39834 = n37900 & ~n39833 ;
  assign n39835 = n39834 ^ n1114 ^ x196 ;
  assign n39836 = n6621 & ~n28048 ;
  assign n39837 = n12702 | n15270 ;
  assign n39838 = ~n24971 & n39837 ;
  assign n39839 = n39838 ^ n29927 ^ n12868 ;
  assign n39840 = ( n6442 & n13043 ) | ( n6442 & ~n20781 ) | ( n13043 & ~n20781 ) ;
  assign n39841 = ( x161 & n16474 ) | ( x161 & ~n38578 ) | ( n16474 & ~n38578 ) ;
  assign n39842 = n39841 ^ n28478 ^ 1'b0 ;
  assign n39843 = n27945 & n39842 ;
  assign n39844 = n39843 ^ n28363 ^ n17143 ;
  assign n39845 = n2533 & n31526 ;
  assign n39846 = ( n1658 & n5888 ) | ( n1658 & n11740 ) | ( n5888 & n11740 ) ;
  assign n39847 = n39845 & ~n39846 ;
  assign n39848 = n39847 ^ n2680 ^ 1'b0 ;
  assign n39849 = n39848 ^ n31782 ^ n28855 ;
  assign n39850 = n22058 ^ n17685 ^ n2444 ;
  assign n39852 = n23939 ^ n9980 ^ n1296 ;
  assign n39853 = ( x175 & ~n15503 ) | ( x175 & n39852 ) | ( ~n15503 & n39852 ) ;
  assign n39851 = ( n7689 & ~n10904 ) | ( n7689 & n25843 ) | ( ~n10904 & n25843 ) ;
  assign n39854 = n39853 ^ n39851 ^ n12795 ;
  assign n39855 = n34400 & ~n39854 ;
  assign n39856 = n38431 & n39855 ;
  assign n39857 = ( ~n22110 & n39850 ) | ( ~n22110 & n39856 ) | ( n39850 & n39856 ) ;
  assign n39858 = n1496 & n30588 ;
  assign n39859 = n6514 & n39858 ;
  assign n39860 = ~n7406 & n9952 ;
  assign n39861 = ( n20430 & n39859 ) | ( n20430 & ~n39860 ) | ( n39859 & ~n39860 ) ;
  assign n39867 = ( n1099 & ~n3702 ) | ( n1099 & n24350 ) | ( ~n3702 & n24350 ) ;
  assign n39868 = n39867 ^ n23692 ^ n6614 ;
  assign n39862 = n24237 ^ n5007 ^ n4496 ;
  assign n39863 = n39862 ^ n7058 ^ n6934 ;
  assign n39864 = n12062 ^ n11312 ^ n3003 ;
  assign n39865 = n39864 ^ n36304 ^ n24324 ;
  assign n39866 = ( n12494 & ~n39863 ) | ( n12494 & n39865 ) | ( ~n39863 & n39865 ) ;
  assign n39869 = n39868 ^ n39866 ^ n3211 ;
  assign n39870 = n14193 & ~n19057 ;
  assign n39871 = n5451 & n39870 ;
  assign n39872 = ( n1554 & n37911 ) | ( n1554 & ~n39871 ) | ( n37911 & ~n39871 ) ;
  assign n39873 = ( n3871 & ~n6288 ) | ( n3871 & n22430 ) | ( ~n6288 & n22430 ) ;
  assign n39874 = n29389 & n39873 ;
  assign n39875 = ( n9456 & n23187 ) | ( n9456 & n38014 ) | ( n23187 & n38014 ) ;
  assign n39876 = n37122 ^ n6529 ^ n4180 ;
  assign n39877 = n27204 ^ n22995 ^ n797 ;
  assign n39878 = n39877 ^ n6437 ^ 1'b0 ;
  assign n39879 = n39876 & n39878 ;
  assign n39880 = n39879 ^ n32025 ^ n10998 ;
  assign n39881 = n21025 ^ n13066 ^ n10193 ;
  assign n39882 = n39881 ^ n10927 ^ n4919 ;
  assign n39883 = n28737 | n39882 ;
  assign n39884 = ( ~n5591 & n11949 ) | ( ~n5591 & n26280 ) | ( n11949 & n26280 ) ;
  assign n39885 = n34618 ^ n33063 ^ 1'b0 ;
  assign n39886 = ( n1715 & n26647 ) | ( n1715 & n32065 ) | ( n26647 & n32065 ) ;
  assign n39887 = n39886 ^ n25888 ^ n6302 ;
  assign n39888 = ( n19068 & n39885 ) | ( n19068 & n39887 ) | ( n39885 & n39887 ) ;
  assign n39889 = ( n1706 & n4605 ) | ( n1706 & n7595 ) | ( n4605 & n7595 ) ;
  assign n39891 = n28202 ^ n24068 ^ n11155 ;
  assign n39890 = n7101 & n36845 ;
  assign n39892 = n39891 ^ n39890 ^ 1'b0 ;
  assign n39895 = ( n2106 & n6364 ) | ( n2106 & n8618 ) | ( n6364 & n8618 ) ;
  assign n39896 = n5714 ^ n4925 ^ 1'b0 ;
  assign n39897 = n39896 ^ n3392 ^ 1'b0 ;
  assign n39898 = n39895 & n39897 ;
  assign n39893 = n31617 ^ n27613 ^ n19694 ;
  assign n39894 = n24483 | n39893 ;
  assign n39899 = n39898 ^ n39894 ^ 1'b0 ;
  assign n39900 = n31392 ^ n1363 ^ 1'b0 ;
  assign n39902 = n25961 ^ n15301 ^ n15182 ;
  assign n39903 = n39902 ^ n14349 ^ n4624 ;
  assign n39904 = n39903 ^ n25547 ^ n14109 ;
  assign n39901 = n7574 ^ n6452 ^ 1'b0 ;
  assign n39905 = n39904 ^ n39901 ^ n26218 ;
  assign n39906 = n34083 ^ n26004 ^ n21141 ;
  assign n39907 = n16966 ^ n11549 ^ n5199 ;
  assign n39908 = n39907 ^ n25407 ^ n1434 ;
  assign n39909 = n39908 ^ n3478 ^ n2217 ;
  assign n39910 = ~n2608 & n2975 ;
  assign n39911 = n39910 ^ n4583 ^ n1489 ;
  assign n39912 = n36205 ^ n26047 ^ 1'b0 ;
  assign n39913 = ( n12800 & ~n17855 ) | ( n12800 & n22172 ) | ( ~n17855 & n22172 ) ;
  assign n39914 = n19729 ^ n7917 ^ n1627 ;
  assign n39915 = x194 & n39914 ;
  assign n39916 = ~n4896 & n7958 ;
  assign n39917 = n7685 & n39916 ;
  assign n39918 = ( ~n39913 & n39915 ) | ( ~n39913 & n39917 ) | ( n39915 & n39917 ) ;
  assign n39919 = ( n3260 & n19047 ) | ( n3260 & n29392 ) | ( n19047 & n29392 ) ;
  assign n39920 = ( n884 & n13725 ) | ( n884 & n19111 ) | ( n13725 & n19111 ) ;
  assign n39921 = n39920 ^ n25422 ^ n25226 ;
  assign n39922 = ( n2175 & ~n11063 ) | ( n2175 & n39921 ) | ( ~n11063 & n39921 ) ;
  assign n39923 = ( ~n8115 & n39919 ) | ( ~n8115 & n39922 ) | ( n39919 & n39922 ) ;
  assign n39929 = n12725 ^ n10024 ^ n3420 ;
  assign n39930 = n39929 ^ n17756 ^ n14380 ;
  assign n39931 = n31318 & n39930 ;
  assign n39932 = n39931 ^ n23709 ^ 1'b0 ;
  assign n39924 = ~n2850 & n21528 ;
  assign n39925 = n39924 ^ n17022 ^ 1'b0 ;
  assign n39926 = n39925 ^ n34010 ^ n12762 ;
  assign n39927 = n14695 | n39926 ;
  assign n39928 = n25404 | n39927 ;
  assign n39933 = n39932 ^ n39928 ^ 1'b0 ;
  assign n39938 = n27208 ^ n14166 ^ 1'b0 ;
  assign n39939 = ~n788 & n39938 ;
  assign n39934 = ( n2998 & n5215 ) | ( n2998 & n7632 ) | ( n5215 & n7632 ) ;
  assign n39935 = n39934 ^ n28692 ^ 1'b0 ;
  assign n39936 = n39935 ^ n7888 ^ n3929 ;
  assign n39937 = n39936 ^ n8655 ^ x27 ;
  assign n39940 = n39939 ^ n39937 ^ n1873 ;
  assign n39941 = n39940 ^ n37890 ^ n3137 ;
  assign n39942 = n39941 ^ n17500 ^ n9903 ;
  assign n39943 = ( n3957 & n7324 ) | ( n3957 & ~n7337 ) | ( n7324 & ~n7337 ) ;
  assign n39944 = n35310 ^ n33122 ^ n31197 ;
  assign n39945 = ( n18635 & n39943 ) | ( n18635 & n39944 ) | ( n39943 & n39944 ) ;
  assign n39946 = n39945 ^ n24449 ^ n11236 ;
  assign n39947 = n35353 ^ n14782 ^ 1'b0 ;
  assign n39948 = n39947 ^ n37788 ^ n15483 ;
  assign n39949 = n39948 ^ n34240 ^ n31570 ;
  assign n39950 = n28443 | n37433 ;
  assign n39951 = n28938 & ~n39950 ;
  assign n39952 = ( n7352 & ~n31822 ) | ( n7352 & n39951 ) | ( ~n31822 & n39951 ) ;
  assign n39953 = ~n23941 & n23972 ;
  assign n39954 = n39953 ^ n15134 ^ 1'b0 ;
  assign n39955 = n32087 ^ n30505 ^ n7183 ;
  assign n39956 = n38852 ^ n37616 ^ n20390 ;
  assign n39957 = n21801 ^ n18943 ^ n10383 ;
  assign n39958 = n39957 ^ n21857 ^ n11668 ;
  assign n39959 = ( n2976 & n7748 ) | ( n2976 & ~n9432 ) | ( n7748 & ~n9432 ) ;
  assign n39960 = ( n11406 & n39081 ) | ( n11406 & n39959 ) | ( n39081 & n39959 ) ;
  assign n39961 = n39960 ^ n15504 ^ n7997 ;
  assign n39962 = ( n12801 & ~n28339 ) | ( n12801 & n29116 ) | ( ~n28339 & n29116 ) ;
  assign n39963 = ~n26292 & n38568 ;
  assign n39964 = n3584 & n39963 ;
  assign n39965 = ( n5036 & n15506 ) | ( n5036 & ~n39964 ) | ( n15506 & ~n39964 ) ;
  assign n39966 = n27845 ^ n13440 ^ n3701 ;
  assign n39967 = ( n7923 & ~n17119 ) | ( n7923 & n21375 ) | ( ~n17119 & n21375 ) ;
  assign n39968 = n39967 ^ n1865 ^ 1'b0 ;
  assign n39969 = n39519 | n39968 ;
  assign n39970 = n3277 ^ x109 ^ 1'b0 ;
  assign n39975 = n21948 ^ n1374 ^ 1'b0 ;
  assign n39971 = n7522 | n15830 ;
  assign n39972 = n39971 ^ n1448 ^ 1'b0 ;
  assign n39973 = n39972 ^ n26557 ^ 1'b0 ;
  assign n39974 = n8077 & ~n39973 ;
  assign n39976 = n39975 ^ n39974 ^ n1028 ;
  assign n39977 = n39976 ^ n25035 ^ n1968 ;
  assign n39978 = n19085 ^ n18227 ^ n11750 ;
  assign n39979 = ( n17507 & ~n31818 ) | ( n17507 & n38944 ) | ( ~n31818 & n38944 ) ;
  assign n39980 = ( ~n1964 & n16269 ) | ( ~n1964 & n21814 ) | ( n16269 & n21814 ) ;
  assign n39981 = n6202 & n6760 ;
  assign n39982 = n39981 ^ n6484 ^ n4863 ;
  assign n39983 = n9508 & ~n39982 ;
  assign n39984 = n39983 ^ n38087 ^ 1'b0 ;
  assign n39987 = ( n915 & ~n2342 ) | ( n915 & n6245 ) | ( ~n2342 & n6245 ) ;
  assign n39988 = n39987 ^ n20361 ^ n4373 ;
  assign n39985 = n39532 ^ n9682 ^ 1'b0 ;
  assign n39986 = n2477 & ~n39985 ;
  assign n39989 = n39988 ^ n39986 ^ n6649 ;
  assign n39990 = ( n17672 & n27928 ) | ( n17672 & ~n34431 ) | ( n27928 & ~n34431 ) ;
  assign n39991 = ( n4865 & ~n10270 ) | ( n4865 & n35676 ) | ( ~n10270 & n35676 ) ;
  assign n39997 = n504 & ~n16026 ;
  assign n39998 = n11033 & n39997 ;
  assign n39992 = n10585 ^ n6803 ^ n5267 ;
  assign n39993 = n18544 ^ n16383 ^ 1'b0 ;
  assign n39994 = n39992 & ~n39993 ;
  assign n39995 = n39994 ^ n37754 ^ 1'b0 ;
  assign n39996 = ~n13583 & n39995 ;
  assign n39999 = n39998 ^ n39996 ^ n20361 ;
  assign n40000 = ( n12880 & n23004 ) | ( n12880 & ~n26637 ) | ( n23004 & ~n26637 ) ;
  assign n40001 = n40000 ^ n21671 ^ n1497 ;
  assign n40002 = n40001 ^ n39821 ^ n3682 ;
  assign n40003 = n40002 ^ n13874 ^ n5987 ;
  assign n40004 = n1560 & n3802 ;
  assign n40005 = ~n1137 & n40004 ;
  assign n40006 = n9920 & ~n27259 ;
  assign n40007 = n7433 & ~n14534 ;
  assign n40008 = ( n5601 & ~n9855 ) | ( n5601 & n12094 ) | ( ~n9855 & n12094 ) ;
  assign n40009 = n6662 & n28193 ;
  assign n40010 = ( n2294 & n31470 ) | ( n2294 & n40009 ) | ( n31470 & n40009 ) ;
  assign n40011 = n40010 ^ n32668 ^ n7699 ;
  assign n40012 = n31214 ^ n21515 ^ n10177 ;
  assign n40014 = n24675 ^ n17155 ^ n1205 ;
  assign n40015 = ( ~n9529 & n17131 ) | ( ~n9529 & n40014 ) | ( n17131 & n40014 ) ;
  assign n40016 = ( n6155 & n17362 ) | ( n6155 & n40015 ) | ( n17362 & n40015 ) ;
  assign n40013 = n27189 ^ n8549 ^ n531 ;
  assign n40017 = n40016 ^ n40013 ^ n16651 ;
  assign n40018 = ( n3004 & ~n14493 ) | ( n3004 & n40017 ) | ( ~n14493 & n40017 ) ;
  assign n40019 = n40018 ^ n12296 ^ n3123 ;
  assign n40020 = n40019 ^ n20238 ^ 1'b0 ;
  assign n40022 = ( n654 & n7026 ) | ( n654 & n19350 ) | ( n7026 & n19350 ) ;
  assign n40023 = n12877 ^ n12353 ^ n9508 ;
  assign n40024 = ( ~n1168 & n15880 ) | ( ~n1168 & n40023 ) | ( n15880 & n40023 ) ;
  assign n40025 = ( n26142 & n40022 ) | ( n26142 & n40024 ) | ( n40022 & n40024 ) ;
  assign n40021 = ( n1442 & n11227 ) | ( n1442 & ~n22691 ) | ( n11227 & ~n22691 ) ;
  assign n40026 = n40025 ^ n40021 ^ n25273 ;
  assign n40027 = ( ~n19220 & n25737 ) | ( ~n19220 & n30220 ) | ( n25737 & n30220 ) ;
  assign n40028 = ( n15814 & ~n16922 ) | ( n15814 & n26066 ) | ( ~n16922 & n26066 ) ;
  assign n40029 = n40027 & ~n40028 ;
  assign n40031 = n18124 ^ n7764 ^ n4152 ;
  assign n40030 = ~n8881 & n18350 ;
  assign n40032 = n40031 ^ n40030 ^ 1'b0 ;
  assign n40033 = n16471 ^ n12132 ^ 1'b0 ;
  assign n40034 = n35929 ^ n31723 ^ n15852 ;
  assign n40035 = n7474 & ~n18204 ;
  assign n40036 = n40035 ^ n15082 ^ 1'b0 ;
  assign n40037 = ( n1818 & n6917 ) | ( n1818 & ~n40036 ) | ( n6917 & ~n40036 ) ;
  assign n40038 = n34107 ^ n13842 ^ n11852 ;
  assign n40039 = ( n2122 & ~n8924 ) | ( n2122 & n20443 ) | ( ~n8924 & n20443 ) ;
  assign n40040 = n6901 | n9374 ;
  assign n40041 = n33993 ^ n1399 ^ 1'b0 ;
  assign n40042 = n10546 | n40041 ;
  assign n40043 = ( n14200 & ~n33889 ) | ( n14200 & n40042 ) | ( ~n33889 & n40042 ) ;
  assign n40044 = n40043 ^ n8254 ^ 1'b0 ;
  assign n40045 = ( n17256 & n19338 ) | ( n17256 & ~n40044 ) | ( n19338 & ~n40044 ) ;
  assign n40046 = n34766 & n40045 ;
  assign n40047 = ~n25966 & n40046 ;
  assign n40048 = n5552 & n13490 ;
  assign n40049 = ~n31168 & n40048 ;
  assign n40050 = ( n7815 & ~n10282 ) | ( n7815 & n34716 ) | ( ~n10282 & n34716 ) ;
  assign n40053 = n13467 ^ n3552 ^ n2300 ;
  assign n40052 = ~n8627 & n31921 ;
  assign n40054 = n40053 ^ n40052 ^ 1'b0 ;
  assign n40051 = n3216 & ~n9693 ;
  assign n40055 = n40054 ^ n40051 ^ n7143 ;
  assign n40056 = ( n6221 & ~n17463 ) | ( n6221 & n37372 ) | ( ~n17463 & n37372 ) ;
  assign n40057 = n40056 ^ n3678 ^ 1'b0 ;
  assign n40058 = n34725 ^ n30002 ^ n14039 ;
  assign n40059 = n34190 ^ n19344 ^ n2904 ;
  assign n40061 = n11801 ^ n4575 ^ 1'b0 ;
  assign n40060 = ( n11439 & n16627 ) | ( n11439 & n22410 ) | ( n16627 & n22410 ) ;
  assign n40062 = n40061 ^ n40060 ^ n25770 ;
  assign n40063 = ( n29639 & n33303 ) | ( n29639 & ~n40062 ) | ( n33303 & ~n40062 ) ;
  assign n40070 = ( n5987 & n16036 ) | ( n5987 & ~n33765 ) | ( n16036 & ~n33765 ) ;
  assign n40066 = n4961 ^ n4006 ^ 1'b0 ;
  assign n40064 = n7973 | n8086 ;
  assign n40065 = n40064 ^ n17018 ^ 1'b0 ;
  assign n40067 = n40066 ^ n40065 ^ n32307 ;
  assign n40068 = n24214 & n40067 ;
  assign n40069 = ~n21899 & n40068 ;
  assign n40071 = n40070 ^ n40069 ^ 1'b0 ;
  assign n40072 = n35713 ^ n16247 ^ n3375 ;
  assign n40073 = ( ~n10125 & n14426 ) | ( ~n10125 & n28212 ) | ( n14426 & n28212 ) ;
  assign n40074 = n40073 ^ n36362 ^ n18644 ;
  assign n40075 = n18429 & ~n25051 ;
  assign n40076 = n32972 ^ n27817 ^ n19192 ;
  assign n40077 = n40076 ^ n18066 ^ n8708 ;
  assign n40078 = n24110 ^ n5584 ^ n3549 ;
  assign n40079 = n32464 & ~n35229 ;
  assign n40080 = n40078 & n40079 ;
  assign n40081 = n24420 & ~n25122 ;
  assign n40082 = ~n36089 & n40081 ;
  assign n40083 = n13777 ^ n7485 ^ 1'b0 ;
  assign n40084 = ( n17582 & n34048 ) | ( n17582 & n40083 ) | ( n34048 & n40083 ) ;
  assign n40085 = ( n12511 & n18608 ) | ( n12511 & ~n20303 ) | ( n18608 & ~n20303 ) ;
  assign n40086 = n31184 ^ n7175 ^ 1'b0 ;
  assign n40087 = ( ~n24819 & n38943 ) | ( ~n24819 & n40086 ) | ( n38943 & n40086 ) ;
  assign n40088 = n2600 & n22698 ;
  assign n40089 = n40088 ^ n8014 ^ 1'b0 ;
  assign n40090 = n17897 ^ n12382 ^ 1'b0 ;
  assign n40091 = n17809 & n39551 ;
  assign n40092 = n40091 ^ n9612 ^ 1'b0 ;
  assign n40093 = ( n10920 & n40090 ) | ( n10920 & ~n40092 ) | ( n40090 & ~n40092 ) ;
  assign n40094 = ( n11012 & ~n40089 ) | ( n11012 & n40093 ) | ( ~n40089 & n40093 ) ;
  assign n40095 = n33498 ^ n17418 ^ n14094 ;
  assign n40096 = ~n13667 & n23695 ;
  assign n40097 = ~n10515 & n40096 ;
  assign n40098 = ( n4093 & n13845 ) | ( n4093 & n40097 ) | ( n13845 & n40097 ) ;
  assign n40099 = ~n27785 & n40098 ;
  assign n40100 = n6235 ^ n1791 ^ 1'b0 ;
  assign n40101 = n35132 ^ n19207 ^ n1130 ;
  assign n40102 = n40101 ^ n24902 ^ n7481 ;
  assign n40103 = n40102 ^ n2694 ^ 1'b0 ;
  assign n40104 = n40100 & n40103 ;
  assign n40105 = n30535 ^ n7004 ^ 1'b0 ;
  assign n40106 = n20592 | n40105 ;
  assign n40107 = ( n472 & n3087 ) | ( n472 & n4947 ) | ( n3087 & n4947 ) ;
  assign n40108 = n40107 ^ n25937 ^ 1'b0 ;
  assign n40109 = ( n336 & n7157 ) | ( n336 & n10490 ) | ( n7157 & n10490 ) ;
  assign n40110 = ( n16158 & n22986 ) | ( n16158 & n40109 ) | ( n22986 & n40109 ) ;
  assign n40111 = n30792 ^ n13474 ^ n6134 ;
  assign n40112 = n29532 ^ n19633 ^ 1'b0 ;
  assign n40113 = n40112 ^ n27711 ^ n20354 ;
  assign n40114 = n40113 ^ n29706 ^ n18776 ;
  assign n40116 = ( ~n286 & n19484 ) | ( ~n286 & n21607 ) | ( n19484 & n21607 ) ;
  assign n40115 = n34796 ^ n19090 ^ 1'b0 ;
  assign n40117 = n40116 ^ n40115 ^ n19713 ;
  assign n40118 = n14967 & ~n23103 ;
  assign n40119 = n40118 ^ n1038 ^ 1'b0 ;
  assign n40120 = ( n7571 & n23903 ) | ( n7571 & n40119 ) | ( n23903 & n40119 ) ;
  assign n40121 = n40120 ^ n30608 ^ n26891 ;
  assign n40122 = ( n2920 & n30677 ) | ( n2920 & n38342 ) | ( n30677 & n38342 ) ;
  assign n40123 = n21573 ^ n11415 ^ n4437 ;
  assign n40124 = n40123 ^ n18981 ^ 1'b0 ;
  assign n40125 = n30900 & ~n40124 ;
  assign n40126 = n18732 & ~n19511 ;
  assign n40127 = ~n24612 & n40126 ;
  assign n40128 = n13841 | n21081 ;
  assign n40129 = n40128 ^ n35002 ^ 1'b0 ;
  assign n40130 = ~n34503 & n40129 ;
  assign n40131 = ~n30192 & n34216 ;
  assign n40132 = ~n871 & n11770 ;
  assign n40133 = n40132 ^ n17555 ^ 1'b0 ;
  assign n40134 = n5089 & ~n40133 ;
  assign n40135 = n23807 & n40134 ;
  assign n40136 = n9390 | n32702 ;
  assign n40137 = n8320 | n40136 ;
  assign n40138 = n40137 ^ n25879 ^ n23677 ;
  assign n40139 = n19225 ^ n2825 ^ 1'b0 ;
  assign n40140 = n40139 ^ n18723 ^ n8076 ;
  assign n40141 = n2598 | n32331 ;
  assign n40142 = n10234 | n40141 ;
  assign n40143 = n2127 | n19513 ;
  assign n40144 = n40143 ^ n17315 ^ 1'b0 ;
  assign n40145 = n40144 ^ n8070 ^ 1'b0 ;
  assign n40146 = ~n21428 & n40145 ;
  assign n40147 = ~n3420 & n18437 ;
  assign n40148 = n15592 & n35948 ;
  assign n40149 = n40148 ^ n31075 ^ n5458 ;
  assign n40150 = ( n10413 & n12259 ) | ( n10413 & n40149 ) | ( n12259 & n40149 ) ;
  assign n40151 = n18586 ^ n9156 ^ 1'b0 ;
  assign n40152 = n40151 ^ n9465 ^ n7166 ;
  assign n40153 = n37093 ^ n13015 ^ 1'b0 ;
  assign n40154 = n36763 ^ n26140 ^ n1343 ;
  assign n40155 = ( n28059 & ~n40153 ) | ( n28059 & n40154 ) | ( ~n40153 & n40154 ) ;
  assign n40156 = n3200 | n30613 ;
  assign n40157 = n10729 & ~n40156 ;
  assign n40158 = n40157 ^ n311 ^ 1'b0 ;
  assign n40159 = n27679 | n40158 ;
  assign n40160 = x172 & n32736 ;
  assign n40161 = n3120 & n40160 ;
  assign n40162 = ~n388 & n20533 ;
  assign n40163 = n40162 ^ n24735 ^ 1'b0 ;
  assign n40164 = n40163 ^ n10766 ^ 1'b0 ;
  assign n40165 = ( n11182 & n20678 ) | ( n11182 & n23789 ) | ( n20678 & n23789 ) ;
  assign n40167 = n12957 | n26884 ;
  assign n40166 = ( ~n2112 & n10429 ) | ( ~n2112 & n35485 ) | ( n10429 & n35485 ) ;
  assign n40168 = n40167 ^ n40166 ^ 1'b0 ;
  assign n40170 = n32928 ^ n6634 ^ n4088 ;
  assign n40169 = n19605 ^ n16637 ^ n9920 ;
  assign n40171 = n40170 ^ n40169 ^ n1928 ;
  assign n40172 = n13683 ^ n10940 ^ n1911 ;
  assign n40173 = n11589 ^ n7006 ^ n6287 ;
  assign n40174 = ( n11301 & n28183 ) | ( n11301 & n38810 ) | ( n28183 & n38810 ) ;
  assign n40175 = n40174 ^ n15181 ^ 1'b0 ;
  assign n40176 = n11202 ^ n6864 ^ n6487 ;
  assign n40177 = n4864 & n20150 ;
  assign n40178 = n40177 ^ n33911 ^ 1'b0 ;
  assign n40179 = n40178 ^ n34532 ^ n21452 ;
  assign n40180 = n25306 ^ n21656 ^ n9848 ;
  assign n40181 = n24339 & n40180 ;
  assign n40182 = ~n14017 & n40181 ;
  assign n40183 = n34107 ^ n6716 ^ 1'b0 ;
  assign n40184 = n21209 & ~n40183 ;
  assign n40185 = n40184 ^ n6997 ^ n3702 ;
  assign n40186 = n40185 ^ n4166 ^ n1575 ;
  assign n40187 = n888 | n40186 ;
  assign n40188 = n6746 & ~n40187 ;
  assign n40189 = ( n4398 & n20710 ) | ( n4398 & ~n25498 ) | ( n20710 & ~n25498 ) ;
  assign n40190 = n40189 ^ n21776 ^ n7050 ;
  assign n40191 = ( n6933 & n34058 ) | ( n6933 & ~n40190 ) | ( n34058 & ~n40190 ) ;
  assign n40192 = n4423 & ~n18686 ;
  assign n40193 = ( ~n13209 & n16065 ) | ( ~n13209 & n17443 ) | ( n16065 & n17443 ) ;
  assign n40194 = n39070 ^ n6206 ^ 1'b0 ;
  assign n40195 = n8202 & ~n14373 ;
  assign n40196 = ~n4315 & n40195 ;
  assign n40197 = n40196 ^ n28059 ^ n12183 ;
  assign n40198 = n22362 ^ n7547 ^ n867 ;
  assign n40199 = ( ~n5145 & n40197 ) | ( ~n5145 & n40198 ) | ( n40197 & n40198 ) ;
  assign n40200 = n10867 ^ n1954 ^ n824 ;
  assign n40201 = n40200 ^ n22968 ^ n5314 ;
  assign n40202 = n40201 ^ n15933 ^ n7936 ;
  assign n40203 = n17714 ^ n13579 ^ n8867 ;
  assign n40204 = n14196 ^ n10614 ^ 1'b0 ;
  assign n40205 = ( ~n20952 & n40203 ) | ( ~n20952 & n40204 ) | ( n40203 & n40204 ) ;
  assign n40206 = n40205 ^ n13301 ^ n12822 ;
  assign n40207 = ( n11929 & n33324 ) | ( n11929 & n40206 ) | ( n33324 & n40206 ) ;
  assign n40208 = ( ~n2694 & n6381 ) | ( ~n2694 & n9281 ) | ( n6381 & n9281 ) ;
  assign n40209 = n40208 ^ n18153 ^ 1'b0 ;
  assign n40210 = n29878 & n40209 ;
  assign n40211 = n40210 ^ n10357 ^ n7440 ;
  assign n40212 = n33178 ^ n23427 ^ n3394 ;
  assign n40215 = n11881 ^ n1220 ^ 1'b0 ;
  assign n40213 = ( n10266 & n17601 ) | ( n10266 & n31127 ) | ( n17601 & n31127 ) ;
  assign n40214 = n40213 ^ n34192 ^ n8025 ;
  assign n40216 = n40215 ^ n40214 ^ 1'b0 ;
  assign n40217 = n19334 & ~n40216 ;
  assign n40218 = n5173 & ~n34927 ;
  assign n40219 = n31221 ^ n17329 ^ n1857 ;
  assign n40220 = ( ~n1994 & n2714 ) | ( ~n1994 & n4365 ) | ( n2714 & n4365 ) ;
  assign n40221 = ~n33340 & n37225 ;
  assign n40222 = ( n27720 & n40220 ) | ( n27720 & n40221 ) | ( n40220 & n40221 ) ;
  assign n40223 = ( x9 & ~n40219 ) | ( x9 & n40222 ) | ( ~n40219 & n40222 ) ;
  assign n40224 = n19691 ^ n4122 ^ x123 ;
  assign n40228 = n31181 ^ n17117 ^ 1'b0 ;
  assign n40229 = ~n14160 & n40228 ;
  assign n40225 = n20517 & ~n38904 ;
  assign n40226 = n40225 ^ n18243 ^ 1'b0 ;
  assign n40227 = ~n19771 & n40226 ;
  assign n40230 = n40229 ^ n40227 ^ 1'b0 ;
  assign n40231 = n40230 ^ n27591 ^ n18066 ;
  assign n40232 = ( n1987 & ~n8246 ) | ( n1987 & n24755 ) | ( ~n8246 & n24755 ) ;
  assign n40235 = ( n3469 & n14037 ) | ( n3469 & n22530 ) | ( n14037 & n22530 ) ;
  assign n40234 = x0 & ~n14013 ;
  assign n40233 = ( ~n19519 & n25829 ) | ( ~n19519 & n30815 ) | ( n25829 & n30815 ) ;
  assign n40236 = n40235 ^ n40234 ^ n40233 ;
  assign n40237 = n3498 ^ n622 ^ 1'b0 ;
  assign n40238 = ~n16573 & n40237 ;
  assign n40240 = n21187 ^ n6564 ^ n3364 ;
  assign n40239 = ( ~n883 & n13573 ) | ( ~n883 & n17769 ) | ( n13573 & n17769 ) ;
  assign n40241 = n40240 ^ n40239 ^ n25040 ;
  assign n40242 = ( ~n9996 & n10142 ) | ( ~n9996 & n40241 ) | ( n10142 & n40241 ) ;
  assign n40243 = n13653 | n19808 ;
  assign n40244 = n40243 ^ n8756 ^ 1'b0 ;
  assign n40245 = ( n1964 & n27702 ) | ( n1964 & n34031 ) | ( n27702 & n34031 ) ;
  assign n40246 = ( n10854 & n40244 ) | ( n10854 & n40245 ) | ( n40244 & n40245 ) ;
  assign n40247 = n40246 ^ n39498 ^ n37851 ;
  assign n40248 = ~n2592 & n28754 ;
  assign n40249 = ~n5387 & n17740 ;
  assign n40250 = ~n565 & n40249 ;
  assign n40251 = ( ~n5976 & n40248 ) | ( ~n5976 & n40250 ) | ( n40248 & n40250 ) ;
  assign n40252 = n28150 ^ n25565 ^ n11617 ;
  assign n40253 = n40252 ^ n14747 ^ 1'b0 ;
  assign n40254 = n26212 & n34003 ;
  assign n40255 = n10982 & n40254 ;
  assign n40256 = n30818 ^ n28843 ^ n26032 ;
  assign n40257 = n14407 ^ n12030 ^ 1'b0 ;
  assign n40258 = ~n4180 & n40257 ;
  assign n40259 = ( n40255 & ~n40256 ) | ( n40255 & n40258 ) | ( ~n40256 & n40258 ) ;
  assign n40260 = n18499 ^ n4764 ^ 1'b0 ;
  assign n40261 = n33918 & ~n40260 ;
  assign n40262 = n40261 ^ n15122 ^ n14326 ;
  assign n40263 = n2322 & n15535 ;
  assign n40264 = n40263 ^ n25792 ^ 1'b0 ;
  assign n40266 = ( n3118 & n15565 ) | ( n3118 & n26758 ) | ( n15565 & n26758 ) ;
  assign n40265 = ~n1935 & n39999 ;
  assign n40267 = n40266 ^ n40265 ^ 1'b0 ;
  assign n40268 = ( n3690 & n4448 ) | ( n3690 & n7732 ) | ( n4448 & n7732 ) ;
  assign n40269 = n40268 ^ n36872 ^ n16194 ;
  assign n40270 = ( n19006 & n25186 ) | ( n19006 & n38823 ) | ( n25186 & n38823 ) ;
  assign n40272 = ~n22538 & n25001 ;
  assign n40273 = n40272 ^ n3823 ^ 1'b0 ;
  assign n40271 = n18389 ^ n14422 ^ n11732 ;
  assign n40274 = n40273 ^ n40271 ^ n6789 ;
  assign n40275 = ( n22547 & n24465 ) | ( n22547 & ~n40274 ) | ( n24465 & ~n40274 ) ;
  assign n40276 = ( n1781 & n8727 ) | ( n1781 & ~n14307 ) | ( n8727 & ~n14307 ) ;
  assign n40277 = n23293 ^ n8137 ^ n2051 ;
  assign n40278 = n26794 ^ n828 ^ 1'b0 ;
  assign n40279 = n4640 & n17736 ;
  assign n40280 = n40279 ^ n4280 ^ 1'b0 ;
  assign n40281 = n20026 ^ n19240 ^ n4332 ;
  assign n40282 = n40281 ^ n14213 ^ n12871 ;
  assign n40283 = n40282 ^ n23478 ^ n20354 ;
  assign n40284 = n13384 & n18352 ;
  assign n40285 = n32121 & n40284 ;
  assign n40286 = n40285 ^ n5259 ^ n1905 ;
  assign n40287 = ( n2386 & ~n4652 ) | ( n2386 & n11507 ) | ( ~n4652 & n11507 ) ;
  assign n40288 = n16334 ^ n14153 ^ n13638 ;
  assign n40289 = n12385 ^ n6182 ^ n6164 ;
  assign n40290 = n40289 ^ n27733 ^ n16759 ;
  assign n40291 = ( n16756 & ~n18957 ) | ( n16756 & n40290 ) | ( ~n18957 & n40290 ) ;
  assign n40293 = n26421 ^ n24768 ^ 1'b0 ;
  assign n40294 = n40293 ^ n10359 ^ 1'b0 ;
  assign n40292 = ( n258 & n8730 ) | ( n258 & ~n29713 ) | ( n8730 & ~n29713 ) ;
  assign n40295 = n40294 ^ n40292 ^ n1181 ;
  assign n40296 = n11482 & ~n15896 ;
  assign n40297 = n40296 ^ n14409 ^ 1'b0 ;
  assign n40298 = n14535 | n40297 ;
  assign n40299 = n40298 ^ n14977 ^ 1'b0 ;
  assign n40300 = ( ~n2200 & n4549 ) | ( ~n2200 & n23146 ) | ( n4549 & n23146 ) ;
  assign n40305 = n10990 ^ n9769 ^ 1'b0 ;
  assign n40306 = ~n11541 & n40305 ;
  assign n40301 = n30345 ^ n17215 ^ 1'b0 ;
  assign n40302 = n25504 & ~n40301 ;
  assign n40303 = n40302 ^ n10479 ^ n1083 ;
  assign n40304 = ( n25130 & n34047 ) | ( n25130 & n40303 ) | ( n34047 & n40303 ) ;
  assign n40307 = n40306 ^ n40304 ^ 1'b0 ;
  assign n40308 = n40300 | n40307 ;
  assign n40309 = ( n4747 & ~n29603 ) | ( n4747 & n33023 ) | ( ~n29603 & n33023 ) ;
  assign n40310 = ( n10332 & n14909 ) | ( n10332 & ~n19395 ) | ( n14909 & ~n19395 ) ;
  assign n40311 = ( n3221 & n40309 ) | ( n3221 & ~n40310 ) | ( n40309 & ~n40310 ) ;
  assign n40312 = n40311 ^ n5193 ^ 1'b0 ;
  assign n40313 = n3329 & ~n19209 ;
  assign n40314 = n40313 ^ n34515 ^ n31888 ;
  assign n40315 = n40314 ^ n28625 ^ n2607 ;
  assign n40316 = ~n15371 & n16023 ;
  assign n40317 = n14909 & n35764 ;
  assign n40318 = ~n9758 & n40317 ;
  assign n40319 = ( n2963 & n37068 ) | ( n2963 & ~n40318 ) | ( n37068 & ~n40318 ) ;
  assign n40320 = n20254 ^ n16779 ^ 1'b0 ;
  assign n40321 = n21357 & n40320 ;
  assign n40322 = n21608 ^ n19992 ^ 1'b0 ;
  assign n40323 = n34348 | n40322 ;
  assign n40324 = n40323 ^ x187 ^ 1'b0 ;
  assign n40325 = ( n2946 & ~n40321 ) | ( n2946 & n40324 ) | ( ~n40321 & n40324 ) ;
  assign n40326 = n40325 ^ n33592 ^ n5714 ;
  assign n40327 = n18371 ^ n8986 ^ 1'b0 ;
  assign n40328 = n22519 & ~n40327 ;
  assign n40329 = ( ~n37523 & n38067 ) | ( ~n37523 & n40328 ) | ( n38067 & n40328 ) ;
  assign n40330 = n37818 ^ n19258 ^ n2928 ;
  assign n40331 = n3477 & n29454 ;
  assign n40332 = n25700 & n40331 ;
  assign n40334 = ( n8903 & n12664 ) | ( n8903 & ~n34462 ) | ( n12664 & ~n34462 ) ;
  assign n40335 = n40334 ^ n39478 ^ n18575 ;
  assign n40333 = ( n2130 & n13863 ) | ( n2130 & n17635 ) | ( n13863 & n17635 ) ;
  assign n40336 = n40335 ^ n40333 ^ n20940 ;
  assign n40337 = ( ~n2425 & n17173 ) | ( ~n2425 & n28174 ) | ( n17173 & n28174 ) ;
  assign n40338 = n23580 & n40337 ;
  assign n40339 = n22957 | n31547 ;
  assign n40340 = n13417 ^ n9591 ^ 1'b0 ;
  assign n40341 = ( n7511 & n26492 ) | ( n7511 & n34006 ) | ( n26492 & n34006 ) ;
  assign n40342 = ( n26087 & ~n38975 ) | ( n26087 & n40341 ) | ( ~n38975 & n40341 ) ;
  assign n40343 = ~n10776 & n35465 ;
  assign n40344 = ~n23071 & n40343 ;
  assign n40345 = ( n28665 & n34598 ) | ( n28665 & ~n40344 ) | ( n34598 & ~n40344 ) ;
  assign n40346 = n26575 ^ n14649 ^ 1'b0 ;
  assign n40347 = ~n37251 & n40346 ;
  assign n40348 = ( n6435 & n7755 ) | ( n6435 & n32244 ) | ( n7755 & n32244 ) ;
  assign n40349 = n10544 & ~n40348 ;
  assign n40350 = n40349 ^ n35229 ^ 1'b0 ;
  assign n40351 = ( n11301 & n29228 ) | ( n11301 & ~n40350 ) | ( n29228 & ~n40350 ) ;
  assign n40352 = n33673 ^ n19905 ^ n11415 ;
  assign n40354 = n10612 ^ n8020 ^ n3115 ;
  assign n40353 = ~n14003 & n28262 ;
  assign n40355 = n40354 ^ n40353 ^ n23682 ;
  assign n40357 = n623 & n13988 ;
  assign n40358 = ~n7393 & n40357 ;
  assign n40356 = n22960 ^ n10154 ^ n4676 ;
  assign n40359 = n40358 ^ n40356 ^ n19409 ;
  assign n40360 = n37357 ^ n28960 ^ 1'b0 ;
  assign n40361 = n8462 | n40360 ;
  assign n40362 = ( n10521 & n14148 ) | ( n10521 & ~n40361 ) | ( n14148 & ~n40361 ) ;
  assign n40363 = ( n4655 & n38872 ) | ( n4655 & n40362 ) | ( n38872 & n40362 ) ;
  assign n40364 = n17214 ^ n6087 ^ 1'b0 ;
  assign n40365 = n17223 | n40364 ;
  assign n40366 = n40365 ^ n11986 ^ 1'b0 ;
  assign n40367 = n40363 & ~n40366 ;
  assign n40369 = n14391 ^ n9772 ^ 1'b0 ;
  assign n40370 = ~n15376 & n40369 ;
  assign n40368 = n9931 & n24567 ;
  assign n40371 = n40370 ^ n40368 ^ 1'b0 ;
  assign n40372 = n12645 ^ n1690 ^ n474 ;
  assign n40374 = n5541 ^ n3319 ^ n903 ;
  assign n40375 = ( n13290 & n22959 ) | ( n13290 & ~n40374 ) | ( n22959 & ~n40374 ) ;
  assign n40373 = n11236 ^ n6585 ^ 1'b0 ;
  assign n40376 = n40375 ^ n40373 ^ n8801 ;
  assign n40377 = n37942 ^ n19506 ^ n7118 ;
  assign n40378 = n403 & n5890 ;
  assign n40379 = ~n13685 & n40378 ;
  assign n40382 = ( n8234 & ~n17075 ) | ( n8234 & n34443 ) | ( ~n17075 & n34443 ) ;
  assign n40383 = ( ~n4376 & n20931 ) | ( ~n4376 & n40382 ) | ( n20931 & n40382 ) ;
  assign n40380 = n3628 | n7016 ;
  assign n40381 = n40380 ^ n16652 ^ 1'b0 ;
  assign n40384 = n40383 ^ n40381 ^ n9769 ;
  assign n40385 = n22766 ^ n4741 ^ n2704 ;
  assign n40386 = n39925 ^ n7830 ^ 1'b0 ;
  assign n40387 = ( ~n13222 & n28833 ) | ( ~n13222 & n29172 ) | ( n28833 & n29172 ) ;
  assign n40388 = ( n1355 & n7793 ) | ( n1355 & ~n8162 ) | ( n7793 & ~n8162 ) ;
  assign n40389 = ~n14674 & n32464 ;
  assign n40390 = n40389 ^ n22077 ^ n8795 ;
  assign n40391 = n9756 ^ n7178 ^ n3920 ;
  assign n40392 = n28465 & ~n40391 ;
  assign n40393 = ~n40390 & n40392 ;
  assign n40394 = ( n3151 & ~n9504 ) | ( n3151 & n27682 ) | ( ~n9504 & n27682 ) ;
  assign n40395 = n22556 ^ n20009 ^ n10620 ;
  assign n40396 = ( ~n14065 & n34659 ) | ( ~n14065 & n40395 ) | ( n34659 & n40395 ) ;
  assign n40397 = n40396 ^ n31629 ^ 1'b0 ;
  assign n40398 = ~n40394 & n40397 ;
  assign n40399 = n2258 & ~n12617 ;
  assign n40400 = n40399 ^ n4121 ^ 1'b0 ;
  assign n40401 = n40400 ^ n18483 ^ n1677 ;
  assign n40402 = n1487 & ~n6156 ;
  assign n40403 = ~n40401 & n40402 ;
  assign n40404 = n27264 ^ n20115 ^ n4337 ;
  assign n40405 = ( n12800 & n15983 ) | ( n12800 & ~n20741 ) | ( n15983 & ~n20741 ) ;
  assign n40407 = ( n2362 & n10336 ) | ( n2362 & ~n12391 ) | ( n10336 & ~n12391 ) ;
  assign n40406 = ( ~n6305 & n19558 ) | ( ~n6305 & n35493 ) | ( n19558 & n35493 ) ;
  assign n40408 = n40407 ^ n40406 ^ 1'b0 ;
  assign n40409 = n16992 ^ n16206 ^ n6258 ;
  assign n40410 = n40409 ^ n28241 ^ n9250 ;
  assign n40411 = n21257 ^ n9605 ^ n6255 ;
  assign n40412 = n40411 ^ n35256 ^ n26751 ;
  assign n40413 = ( n30955 & ~n36593 ) | ( n30955 & n36616 ) | ( ~n36593 & n36616 ) ;
  assign n40414 = n20363 ^ n12135 ^ 1'b0 ;
  assign n40415 = n23752 & n40414 ;
  assign n40416 = n36275 ^ n36228 ^ n1731 ;
  assign n40417 = n9072 ^ n2358 ^ 1'b0 ;
  assign n40418 = ~n40416 & n40417 ;
  assign n40419 = ( n582 & ~n7649 ) | ( n582 & n15667 ) | ( ~n7649 & n15667 ) ;
  assign n40420 = ( ~n21294 & n30746 ) | ( ~n21294 & n40419 ) | ( n30746 & n40419 ) ;
  assign n40421 = ( n4002 & ~n18180 ) | ( n4002 & n23524 ) | ( ~n18180 & n23524 ) ;
  assign n40422 = ( n4150 & ~n29419 ) | ( n4150 & n40421 ) | ( ~n29419 & n40421 ) ;
  assign n40423 = ( n25850 & ~n30058 ) | ( n25850 & n30801 ) | ( ~n30058 & n30801 ) ;
  assign n40424 = n21477 ^ n19448 ^ 1'b0 ;
  assign n40425 = ( n10233 & ~n37962 ) | ( n10233 & n40424 ) | ( ~n37962 & n40424 ) ;
  assign n40426 = n14185 ^ x234 ^ 1'b0 ;
  assign n40427 = ( ~n26607 & n29285 ) | ( ~n26607 & n40426 ) | ( n29285 & n40426 ) ;
  assign n40430 = ( n7532 & n8340 ) | ( n7532 & ~n11684 ) | ( n8340 & ~n11684 ) ;
  assign n40429 = ( n8909 & n17119 ) | ( n8909 & n32603 ) | ( n17119 & n32603 ) ;
  assign n40428 = n28101 ^ n13564 ^ 1'b0 ;
  assign n40431 = n40430 ^ n40429 ^ n40428 ;
  assign n40432 = n316 | n8776 ;
  assign n40433 = n6989 | n40432 ;
  assign n40434 = n24087 & n40433 ;
  assign n40435 = n3828 | n4894 ;
  assign n40436 = ( n5848 & ~n6113 ) | ( n5848 & n40435 ) | ( ~n6113 & n40435 ) ;
  assign n40437 = n40436 ^ n19193 ^ n17747 ;
  assign n40438 = n28401 ^ n3932 ^ 1'b0 ;
  assign n40439 = n5691 ^ n2590 ^ 1'b0 ;
  assign n40440 = n40439 ^ n8783 ^ n1708 ;
  assign n40441 = n40440 ^ n5178 ^ n3425 ;
  assign n40442 = ( ~n5255 & n7871 ) | ( ~n5255 & n39664 ) | ( n7871 & n39664 ) ;
  assign n40443 = ( n661 & n40441 ) | ( n661 & ~n40442 ) | ( n40441 & ~n40442 ) ;
  assign n40444 = n25448 & n40443 ;
  assign n40445 = ( n6333 & ~n7654 ) | ( n6333 & n36665 ) | ( ~n7654 & n36665 ) ;
  assign n40446 = n40445 ^ n38518 ^ n4663 ;
  assign n40447 = n30862 ^ n4812 ^ n3719 ;
  assign n40448 = ( n13132 & ~n16780 ) | ( n13132 & n40447 ) | ( ~n16780 & n40447 ) ;
  assign n40449 = n18472 ^ n18083 ^ n5510 ;
  assign n40450 = ( n364 & n2043 ) | ( n364 & n12775 ) | ( n2043 & n12775 ) ;
  assign n40451 = n40450 ^ n22191 ^ n6975 ;
  assign n40452 = ( n9425 & n40449 ) | ( n9425 & ~n40451 ) | ( n40449 & ~n40451 ) ;
  assign n40453 = n10245 ^ n6974 ^ 1'b0 ;
  assign n40454 = n1954 & n40453 ;
  assign n40455 = ( n4094 & n10048 ) | ( n4094 & n10560 ) | ( n10048 & n10560 ) ;
  assign n40456 = ( n15923 & n38014 ) | ( n15923 & n40455 ) | ( n38014 & n40455 ) ;
  assign n40457 = ( n4777 & n8130 ) | ( n4777 & n33907 ) | ( n8130 & n33907 ) ;
  assign n40458 = ( n27011 & ~n33357 ) | ( n27011 & n40457 ) | ( ~n33357 & n40457 ) ;
  assign n40459 = n40458 ^ n35217 ^ n32036 ;
  assign n40460 = ( ~n2950 & n6883 ) | ( ~n2950 & n23548 ) | ( n6883 & n23548 ) ;
  assign n40464 = n36077 ^ n25316 ^ n5183 ;
  assign n40461 = n21241 ^ n13062 ^ n7213 ;
  assign n40462 = n40461 ^ n24607 ^ 1'b0 ;
  assign n40463 = n40462 ^ n22540 ^ n12393 ;
  assign n40465 = n40464 ^ n40463 ^ n28597 ;
  assign n40471 = n10690 & ~n34175 ;
  assign n40469 = n34321 ^ n19613 ^ n11720 ;
  assign n40466 = n19205 ^ n13499 ^ n11482 ;
  assign n40467 = n40466 ^ n20277 ^ n13396 ;
  assign n40468 = ( n4543 & ~n21699 ) | ( n4543 & n40467 ) | ( ~n21699 & n40467 ) ;
  assign n40470 = n40469 ^ n40468 ^ n20132 ;
  assign n40472 = n40471 ^ n40470 ^ n23603 ;
  assign n40473 = n23840 | n23964 ;
  assign n40474 = ( n2729 & n21485 ) | ( n2729 & n40473 ) | ( n21485 & n40473 ) ;
  assign n40475 = x132 & n7983 ;
  assign n40476 = n40475 ^ n331 ^ 1'b0 ;
  assign n40477 = ~n14840 & n40476 ;
  assign n40478 = n40477 ^ n19518 ^ n14292 ;
  assign n40481 = ( n13073 & n18453 ) | ( n13073 & ~n19141 ) | ( n18453 & ~n19141 ) ;
  assign n40479 = ~n2333 & n13286 ;
  assign n40480 = n40479 ^ n13100 ^ n4581 ;
  assign n40482 = n40481 ^ n40480 ^ n14862 ;
  assign n40483 = n34398 ^ n10325 ^ 1'b0 ;
  assign n40484 = n4343 & ~n40483 ;
  assign n40485 = ~n21982 & n32371 ;
  assign n40486 = n19715 & n40485 ;
  assign n40487 = ( n14027 & n17182 ) | ( n14027 & n24523 ) | ( n17182 & n24523 ) ;
  assign n40488 = n23941 ^ n954 ^ 1'b0 ;
  assign n40489 = n24377 & n40488 ;
  assign n40490 = n39429 ^ n20595 ^ n1518 ;
  assign n40491 = n40490 ^ n6709 ^ 1'b0 ;
  assign n40492 = ( n18332 & n25836 ) | ( n18332 & ~n39383 ) | ( n25836 & ~n39383 ) ;
  assign n40493 = ( n5878 & n8367 ) | ( n5878 & n10167 ) | ( n8367 & n10167 ) ;
  assign n40494 = n13756 ^ n2004 ^ n1088 ;
  assign n40495 = ( ~n6240 & n8557 ) | ( ~n6240 & n40494 ) | ( n8557 & n40494 ) ;
  assign n40496 = n40495 ^ n27322 ^ 1'b0 ;
  assign n40497 = n9188 & n20761 ;
  assign n40498 = ( ~n13439 & n40496 ) | ( ~n13439 & n40497 ) | ( n40496 & n40497 ) ;
  assign n40499 = n4778 ^ n3353 ^ n690 ;
  assign n40500 = ( n1953 & n14370 ) | ( n1953 & ~n40499 ) | ( n14370 & ~n40499 ) ;
  assign n40501 = n40500 ^ n28976 ^ n14988 ;
  assign n40502 = ( n4772 & n10416 ) | ( n4772 & ~n40501 ) | ( n10416 & ~n40501 ) ;
  assign n40503 = n40502 ^ n27494 ^ n4685 ;
  assign n40504 = n4536 ^ n2682 ^ n2443 ;
  assign n40505 = ( n36416 & n40503 ) | ( n36416 & ~n40504 ) | ( n40503 & ~n40504 ) ;
  assign n40506 = ( n1748 & n8874 ) | ( n1748 & n36380 ) | ( n8874 & n36380 ) ;
  assign n40510 = n1022 & ~n30744 ;
  assign n40511 = n40510 ^ n8006 ^ 1'b0 ;
  assign n40512 = n40511 ^ n33102 ^ n2212 ;
  assign n40507 = n5915 | n8356 ;
  assign n40508 = n40507 ^ n3813 ^ 1'b0 ;
  assign n40509 = n40508 ^ n33662 ^ n4494 ;
  assign n40513 = n40512 ^ n40509 ^ n21679 ;
  assign n40514 = ( n3927 & ~n40506 ) | ( n3927 & n40513 ) | ( ~n40506 & n40513 ) ;
  assign n40515 = n26459 ^ n18298 ^ 1'b0 ;
  assign n40516 = n11179 ^ n7343 ^ 1'b0 ;
  assign n40517 = n29023 | n40516 ;
  assign n40518 = n40517 ^ n6944 ^ 1'b0 ;
  assign n40519 = ( ~n10293 & n15040 ) | ( ~n10293 & n17547 ) | ( n15040 & n17547 ) ;
  assign n40520 = n10635 & ~n14006 ;
  assign n40521 = ~n40519 & n40520 ;
  assign n40522 = n327 & n18353 ;
  assign n40523 = ~x31 & n40522 ;
  assign n40524 = n38947 | n40523 ;
  assign n40525 = n39941 ^ n8837 ^ 1'b0 ;
  assign n40526 = n26270 ^ n8858 ^ n2444 ;
  assign n40527 = ~n1182 & n7408 ;
  assign n40528 = n40527 ^ n21226 ^ 1'b0 ;
  assign n40529 = n13806 ^ n6215 ^ 1'b0 ;
  assign n40530 = n40529 ^ n37562 ^ n9496 ;
  assign n40534 = ( n5340 & n9442 ) | ( n5340 & ~n22660 ) | ( n9442 & ~n22660 ) ;
  assign n40533 = ( n2936 & n5223 ) | ( n2936 & ~n19250 ) | ( n5223 & ~n19250 ) ;
  assign n40531 = n21234 | n32726 ;
  assign n40532 = ( n4256 & n8542 ) | ( n4256 & ~n40531 ) | ( n8542 & ~n40531 ) ;
  assign n40535 = n40534 ^ n40533 ^ n40532 ;
  assign n40536 = ( n9249 & ~n16419 ) | ( n9249 & n22132 ) | ( ~n16419 & n22132 ) ;
  assign n40537 = n40536 ^ n35816 ^ n34495 ;
  assign n40538 = ~n17685 & n40537 ;
  assign n40541 = n24390 | n39982 ;
  assign n40539 = n25122 ^ n9177 ^ 1'b0 ;
  assign n40540 = n40539 ^ n23026 ^ n21381 ;
  assign n40542 = n40541 ^ n40540 ^ n38309 ;
  assign n40543 = n31793 ^ n19035 ^ 1'b0 ;
  assign n40544 = n21168 & ~n22380 ;
  assign n40545 = n40544 ^ n2601 ^ 1'b0 ;
  assign n40546 = x150 & ~n33645 ;
  assign n40547 = x84 | n25766 ;
  assign n40548 = n33379 ^ n19754 ^ n4699 ;
  assign n40550 = n18903 ^ n14443 ^ n8653 ;
  assign n40551 = n40550 ^ n8597 ^ n4664 ;
  assign n40549 = n40044 ^ n27807 ^ n7830 ;
  assign n40552 = n40551 ^ n40549 ^ 1'b0 ;
  assign n40553 = ( n13339 & n13593 ) | ( n13339 & ~n27310 ) | ( n13593 & ~n27310 ) ;
  assign n40554 = n40553 ^ n33173 ^ n7775 ;
  assign n40555 = ~n5707 & n32316 ;
  assign n40556 = ( n8711 & n28577 ) | ( n8711 & ~n37991 ) | ( n28577 & ~n37991 ) ;
  assign n40557 = n21950 & n23122 ;
  assign n40558 = n40557 ^ n8679 ^ 1'b0 ;
  assign n40559 = ( n40555 & n40556 ) | ( n40555 & ~n40558 ) | ( n40556 & ~n40558 ) ;
  assign n40560 = n12792 | n27257 ;
  assign n40561 = n19656 ^ n6197 ^ n4096 ;
  assign n40562 = ( ~n4598 & n40560 ) | ( ~n4598 & n40561 ) | ( n40560 & n40561 ) ;
  assign n40563 = n40562 ^ n16865 ^ n12768 ;
  assign n40564 = n696 & n4581 ;
  assign n40565 = n40564 ^ n30200 ^ 1'b0 ;
  assign n40566 = ~n9801 & n40565 ;
  assign n40567 = n38841 ^ n7059 ^ n4025 ;
  assign n40568 = ( n1352 & ~n28150 ) | ( n1352 & n40567 ) | ( ~n28150 & n40567 ) ;
  assign n40569 = ( n12518 & ~n40566 ) | ( n12518 & n40568 ) | ( ~n40566 & n40568 ) ;
  assign n40570 = n9264 & ~n22080 ;
  assign n40571 = n38416 ^ n9336 ^ 1'b0 ;
  assign n40572 = n40570 | n40571 ;
  assign n40573 = ( n17128 & n29310 ) | ( n17128 & n37589 ) | ( n29310 & n37589 ) ;
  assign n40574 = n38260 ^ n24036 ^ n18480 ;
  assign n40575 = n18236 & ~n40574 ;
  assign n40576 = ( n18041 & n19036 ) | ( n18041 & ~n34084 ) | ( n19036 & ~n34084 ) ;
  assign n40582 = n7392 ^ n5332 ^ 1'b0 ;
  assign n40580 = n22052 | n36704 ;
  assign n40581 = n40580 ^ n21339 ^ 1'b0 ;
  assign n40577 = n25437 ^ n1320 ^ 1'b0 ;
  assign n40578 = n34909 ^ n19692 ^ n17672 ;
  assign n40579 = ( n2046 & n40577 ) | ( n2046 & ~n40578 ) | ( n40577 & ~n40578 ) ;
  assign n40583 = n40582 ^ n40581 ^ n40579 ;
  assign n40584 = n12304 ^ n3579 ^ 1'b0 ;
  assign n40585 = n15092 & ~n40584 ;
  assign n40586 = ( n6959 & n12692 ) | ( n6959 & ~n40585 ) | ( n12692 & ~n40585 ) ;
  assign n40587 = n17798 ^ n12900 ^ x2 ;
  assign n40588 = n40587 ^ n28284 ^ n1107 ;
  assign n40589 = ~n3671 & n30454 ;
  assign n40590 = n40589 ^ n14213 ^ 1'b0 ;
  assign n40591 = ( ~n14576 & n16707 ) | ( ~n14576 & n18498 ) | ( n16707 & n18498 ) ;
  assign n40592 = n40591 ^ n9266 ^ n8176 ;
  assign n40593 = n38879 ^ n20460 ^ n10171 ;
  assign n40594 = ( ~n40590 & n40592 ) | ( ~n40590 & n40593 ) | ( n40592 & n40593 ) ;
  assign n40595 = ( ~x183 & n40534 ) | ( ~x183 & n40594 ) | ( n40534 & n40594 ) ;
  assign n40601 = ( ~n10508 & n14974 ) | ( ~n10508 & n15895 ) | ( n14974 & n15895 ) ;
  assign n40599 = n21080 ^ n12291 ^ 1'b0 ;
  assign n40600 = ~n33697 & n40599 ;
  assign n40596 = n29305 ^ n26374 ^ n16269 ;
  assign n40597 = n40596 ^ n21102 ^ 1'b0 ;
  assign n40598 = n1554 & n40597 ;
  assign n40602 = n40601 ^ n40600 ^ n40598 ;
  assign n40603 = n23935 ^ n19963 ^ 1'b0 ;
  assign n40604 = n40602 & ~n40603 ;
  assign n40605 = n7581 & ~n15036 ;
  assign n40606 = n7136 & n40605 ;
  assign n40607 = n40606 ^ n21548 ^ 1'b0 ;
  assign n40608 = n40607 ^ n25747 ^ n422 ;
  assign n40609 = ( n3057 & ~n23088 ) | ( n3057 & n40608 ) | ( ~n23088 & n40608 ) ;
  assign n40610 = ( n22256 & ~n33346 ) | ( n22256 & n40609 ) | ( ~n33346 & n40609 ) ;
  assign n40611 = ( n23077 & ~n24908 ) | ( n23077 & n30631 ) | ( ~n24908 & n30631 ) ;
  assign n40612 = ( ~n1504 & n16555 ) | ( ~n1504 & n40611 ) | ( n16555 & n40611 ) ;
  assign n40613 = n22873 ^ n10617 ^ n9203 ;
  assign n40614 = n2178 & ~n16790 ;
  assign n40615 = ~n13921 & n40614 ;
  assign n40616 = ( n11417 & ~n12205 ) | ( n11417 & n40615 ) | ( ~n12205 & n40615 ) ;
  assign n40617 = n19640 & ~n29224 ;
  assign n40618 = n37202 | n38099 ;
  assign n40619 = ( n7806 & n35899 ) | ( n7806 & ~n40618 ) | ( n35899 & ~n40618 ) ;
  assign n40622 = n6963 & n33493 ;
  assign n40620 = ( ~n11281 & n17018 ) | ( ~n11281 & n38481 ) | ( n17018 & n38481 ) ;
  assign n40621 = n40620 ^ n13004 ^ 1'b0 ;
  assign n40623 = n40622 ^ n40621 ^ n10669 ;
  assign n40624 = ( ~n8567 & n30059 ) | ( ~n8567 & n40623 ) | ( n30059 & n40623 ) ;
  assign n40626 = ( ~x32 & n4396 ) | ( ~x32 & n13686 ) | ( n4396 & n13686 ) ;
  assign n40625 = n8202 & ~n18804 ;
  assign n40627 = n40626 ^ n40625 ^ 1'b0 ;
  assign n40628 = ( n3637 & n32596 ) | ( n3637 & n40627 ) | ( n32596 & n40627 ) ;
  assign n40629 = n11594 ^ n4716 ^ n2626 ;
  assign n40630 = n40629 ^ n13029 ^ n1770 ;
  assign n40631 = n25561 ^ n9372 ^ n1046 ;
  assign n40632 = n27165 ^ n19301 ^ n13198 ;
  assign n40633 = n9028 ^ n2656 ^ 1'b0 ;
  assign n40634 = n18525 & ~n40633 ;
  assign n40635 = ( n19075 & ~n26718 ) | ( n19075 & n35919 ) | ( ~n26718 & n35919 ) ;
  assign n40636 = ~n36614 & n40635 ;
  assign n40637 = ( ~n40632 & n40634 ) | ( ~n40632 & n40636 ) | ( n40634 & n40636 ) ;
  assign n40638 = n40560 ^ n31143 ^ n3261 ;
  assign n40639 = n40638 ^ n18208 ^ n4913 ;
  assign n40640 = ( n599 & n3652 ) | ( n599 & n16784 ) | ( n3652 & n16784 ) ;
  assign n40641 = ~n21135 & n35843 ;
  assign n40642 = n40640 & n40641 ;
  assign n40643 = n22232 | n35005 ;
  assign n40644 = ~n6766 & n39787 ;
  assign n40645 = n2422 & n15795 ;
  assign n40646 = n40645 ^ n9532 ^ 1'b0 ;
  assign n40647 = n40646 ^ n16725 ^ n1568 ;
  assign n40648 = ( ~n3249 & n10693 ) | ( ~n3249 & n12272 ) | ( n10693 & n12272 ) ;
  assign n40651 = n35543 ^ n5000 ^ n2109 ;
  assign n40649 = n16702 ^ n13169 ^ 1'b0 ;
  assign n40650 = ~n9424 & n40649 ;
  assign n40652 = n40651 ^ n40650 ^ n39947 ;
  assign n40653 = n37704 ^ n20197 ^ n1418 ;
  assign n40654 = n17372 ^ n14151 ^ n10721 ;
  assign n40655 = n40654 ^ n2520 ^ 1'b0 ;
  assign n40656 = ( n31094 & n40653 ) | ( n31094 & n40655 ) | ( n40653 & n40655 ) ;
  assign n40657 = ( x14 & n20818 ) | ( x14 & n40656 ) | ( n20818 & n40656 ) ;
  assign n40662 = n7565 & ~n35300 ;
  assign n40658 = n1889 & ~n8707 ;
  assign n40659 = n40658 ^ n25657 ^ 1'b0 ;
  assign n40660 = n1005 & ~n40659 ;
  assign n40661 = ~n33407 & n40660 ;
  assign n40663 = n40662 ^ n40661 ^ n33989 ;
  assign n40666 = n17992 ^ n3662 ^ n2033 ;
  assign n40667 = n40666 ^ n27251 ^ n6729 ;
  assign n40664 = n15135 ^ n6981 ^ n5184 ;
  assign n40665 = ( n15846 & n33232 ) | ( n15846 & ~n40664 ) | ( n33232 & ~n40664 ) ;
  assign n40668 = n40667 ^ n40665 ^ n38750 ;
  assign n40669 = n29450 ^ n27387 ^ n18160 ;
  assign n40670 = n37048 ^ n30443 ^ n2495 ;
  assign n40671 = n25210 ^ n2460 ^ n1618 ;
  assign n40672 = ( n4043 & ~n4823 ) | ( n4043 & n40671 ) | ( ~n4823 & n40671 ) ;
  assign n40673 = ( ~n3390 & n7668 ) | ( ~n3390 & n28312 ) | ( n7668 & n28312 ) ;
  assign n40674 = n14478 ^ n6851 ^ 1'b0 ;
  assign n40675 = n21191 & ~n40674 ;
  assign n40676 = n19686 ^ n15030 ^ n4674 ;
  assign n40677 = n40676 ^ n3538 ^ 1'b0 ;
  assign n40678 = ~n12403 & n40677 ;
  assign n40679 = n11124 ^ n288 ^ 1'b0 ;
  assign n40680 = n6977 | n40679 ;
  assign n40682 = n30765 ^ n19701 ^ 1'b0 ;
  assign n40683 = n5228 | n40682 ;
  assign n40681 = n5685 ^ n4875 ^ n4762 ;
  assign n40684 = n40683 ^ n40681 ^ n14935 ;
  assign n40685 = n40684 ^ n33476 ^ n6950 ;
  assign n40686 = n40680 | n40685 ;
  assign n40687 = n10607 & n24365 ;
  assign n40688 = n40687 ^ n18412 ^ x150 ;
  assign n40689 = n25609 ^ n11019 ^ n2511 ;
  assign n40690 = ( n2895 & n23956 ) | ( n2895 & ~n40689 ) | ( n23956 & ~n40689 ) ;
  assign n40691 = n26073 ^ n16702 ^ 1'b0 ;
  assign n40692 = n9330 ^ n2593 ^ 1'b0 ;
  assign n40693 = n5330 & n40692 ;
  assign n40694 = ( ~n11212 & n35341 ) | ( ~n11212 & n40693 ) | ( n35341 & n40693 ) ;
  assign n40695 = n40694 ^ n29081 ^ 1'b0 ;
  assign n40696 = n14572 | n40695 ;
  assign n40697 = ( n33010 & n34693 ) | ( n33010 & ~n40696 ) | ( n34693 & ~n40696 ) ;
  assign n40698 = ( n2192 & n6835 ) | ( n2192 & n9735 ) | ( n6835 & n9735 ) ;
  assign n40699 = n40698 ^ n21040 ^ n7006 ;
  assign n40700 = ( x178 & n4512 ) | ( x178 & ~n8949 ) | ( n4512 & ~n8949 ) ;
  assign n40701 = n40700 ^ n13613 ^ n10802 ;
  assign n40702 = ( n20623 & ~n30372 ) | ( n20623 & n40701 ) | ( ~n30372 & n40701 ) ;
  assign n40703 = n40702 ^ n25113 ^ n14344 ;
  assign n40704 = n23222 ^ n15711 ^ 1'b0 ;
  assign n40705 = n40703 & n40704 ;
  assign n40706 = ~n14169 & n40705 ;
  assign n40707 = n40706 ^ n28054 ^ 1'b0 ;
  assign n40708 = n18686 & n21315 ;
  assign n40709 = n40708 ^ n11387 ^ 1'b0 ;
  assign n40713 = n19762 ^ n13828 ^ n12455 ;
  assign n40711 = n3752 | n6660 ;
  assign n40712 = n16914 & ~n40711 ;
  assign n40710 = n915 & ~n27507 ;
  assign n40714 = n40713 ^ n40712 ^ n40710 ;
  assign n40715 = ( n649 & n6049 ) | ( n649 & n22595 ) | ( n6049 & n22595 ) ;
  assign n40716 = ( ~n2453 & n3787 ) | ( ~n2453 & n40715 ) | ( n3787 & n40715 ) ;
  assign n40717 = ( n2302 & n16498 ) | ( n2302 & n25552 ) | ( n16498 & n25552 ) ;
  assign n40718 = ( n6227 & n12774 ) | ( n6227 & n24338 ) | ( n12774 & n24338 ) ;
  assign n40719 = n40718 ^ n27159 ^ n17018 ;
  assign n40720 = n40717 | n40719 ;
  assign n40721 = n3471 | n7852 ;
  assign n40722 = ~n17635 & n39569 ;
  assign n40723 = n40722 ^ n18666 ^ n4311 ;
  assign n40724 = n40204 ^ n28131 ^ n2957 ;
  assign n40725 = n13545 | n20556 ;
  assign n40726 = n36726 ^ n13201 ^ 1'b0 ;
  assign n40727 = n40725 & ~n40726 ;
  assign n40728 = ( n40723 & ~n40724 ) | ( n40723 & n40727 ) | ( ~n40724 & n40727 ) ;
  assign n40729 = n12212 & n29008 ;
  assign n40730 = n40729 ^ n35032 ^ 1'b0 ;
  assign n40731 = n15334 & n40730 ;
  assign n40732 = n32395 ^ n19798 ^ n11019 ;
  assign n40733 = n6255 & n15204 ;
  assign n40734 = n40732 & n40733 ;
  assign n40735 = n28310 ^ n23714 ^ n4778 ;
  assign n40736 = ( n8975 & n34351 ) | ( n8975 & n40735 ) | ( n34351 & n40735 ) ;
  assign n40737 = n8735 & n16141 ;
  assign n40738 = n31872 ^ n9501 ^ n3888 ;
  assign n40739 = ( n19835 & n29353 ) | ( n19835 & n40738 ) | ( n29353 & n40738 ) ;
  assign n40740 = ( ~n11681 & n40725 ) | ( ~n11681 & n40739 ) | ( n40725 & n40739 ) ;
  assign n40741 = n40740 ^ n11355 ^ n4381 ;
  assign n40743 = ~n4795 & n22823 ;
  assign n40744 = n4877 & n40743 ;
  assign n40742 = ( n6537 & ~n15433 ) | ( n6537 & n37018 ) | ( ~n15433 & n37018 ) ;
  assign n40745 = n40744 ^ n40742 ^ n4744 ;
  assign n40746 = ( n2403 & n28694 ) | ( n2403 & n38516 ) | ( n28694 & n38516 ) ;
  assign n40747 = n17362 ^ n471 ^ 1'b0 ;
  assign n40749 = n33723 ^ n16678 ^ n16357 ;
  assign n40750 = ( n11783 & n20961 ) | ( n11783 & ~n40749 ) | ( n20961 & ~n40749 ) ;
  assign n40748 = n16572 & ~n24424 ;
  assign n40751 = n40750 ^ n40748 ^ 1'b0 ;
  assign n40752 = n1169 | n31121 ;
  assign n40753 = n8318 | n40752 ;
  assign n40754 = n31339 ^ n30382 ^ 1'b0 ;
  assign n40755 = ~n40753 & n40754 ;
  assign n40756 = ( n18675 & n26046 ) | ( n18675 & n38497 ) | ( n26046 & n38497 ) ;
  assign n40757 = n22501 ^ n5058 ^ n3885 ;
  assign n40758 = ( n11645 & ~n16171 ) | ( n11645 & n19656 ) | ( ~n16171 & n19656 ) ;
  assign n40759 = ( n7461 & n17424 ) | ( n7461 & n40334 ) | ( n17424 & n40334 ) ;
  assign n40760 = n40759 ^ n18404 ^ 1'b0 ;
  assign n40761 = ( ~n9452 & n20731 ) | ( ~n9452 & n40760 ) | ( n20731 & n40760 ) ;
  assign n40762 = ( ~n8513 & n30056 ) | ( ~n8513 & n40761 ) | ( n30056 & n40761 ) ;
  assign n40763 = n16922 | n38097 ;
  assign n40764 = n12019 ^ n9782 ^ n6750 ;
  assign n40765 = ( n20253 & ~n27127 ) | ( n20253 & n28681 ) | ( ~n27127 & n28681 ) ;
  assign n40766 = ( n1425 & n25889 ) | ( n1425 & ~n31471 ) | ( n25889 & ~n31471 ) ;
  assign n40767 = n1189 & n2020 ;
  assign n40768 = ~n33117 & n40767 ;
  assign n40769 = n40536 ^ n39610 ^ n24374 ;
  assign n40770 = n40768 | n40769 ;
  assign n40771 = n22466 ^ n13019 ^ n11715 ;
  assign n40772 = ( n26613 & ~n29020 ) | ( n26613 & n40771 ) | ( ~n29020 & n40771 ) ;
  assign n40773 = ( n31168 & n36178 ) | ( n31168 & n40772 ) | ( n36178 & n40772 ) ;
  assign n40774 = n29699 ^ n20479 ^ 1'b0 ;
  assign n40775 = ~n5516 & n40774 ;
  assign n40776 = ( ~n4695 & n36500 ) | ( ~n4695 & n40775 ) | ( n36500 & n40775 ) ;
  assign n40777 = ( n21039 & n21193 ) | ( n21039 & n40776 ) | ( n21193 & n40776 ) ;
  assign n40778 = ( ~n592 & n23352 ) | ( ~n592 & n34855 ) | ( n23352 & n34855 ) ;
  assign n40779 = n40778 ^ n28202 ^ n3941 ;
  assign n40780 = n11662 ^ n8730 ^ 1'b0 ;
  assign n40781 = n40780 ^ n24768 ^ 1'b0 ;
  assign n40782 = ( n2920 & n12251 ) | ( n2920 & ~n16681 ) | ( n12251 & ~n16681 ) ;
  assign n40783 = n40782 ^ n20438 ^ n5112 ;
  assign n40784 = n20032 ^ n14227 ^ 1'b0 ;
  assign n40785 = n19264 ^ n14863 ^ 1'b0 ;
  assign n40786 = ~n38917 & n40785 ;
  assign n40795 = n35927 ^ n10881 ^ x19 ;
  assign n40793 = n13427 ^ n1136 ^ n312 ;
  assign n40794 = ( ~n12723 & n17505 ) | ( ~n12723 & n40793 ) | ( n17505 & n40793 ) ;
  assign n40796 = n40795 ^ n40794 ^ n3525 ;
  assign n40797 = ( n20759 & n34863 ) | ( n20759 & n40796 ) | ( n34863 & n40796 ) ;
  assign n40790 = n16496 ^ n3353 ^ 1'b0 ;
  assign n40787 = n16602 ^ n8848 ^ n7820 ;
  assign n40788 = n29573 ^ n11955 ^ 1'b0 ;
  assign n40789 = ~n40787 & n40788 ;
  assign n40791 = n40790 ^ n40789 ^ 1'b0 ;
  assign n40792 = ~n28479 & n40791 ;
  assign n40798 = n40797 ^ n40792 ^ n8829 ;
  assign n40799 = ( n1220 & n9162 ) | ( n1220 & ~n36264 ) | ( n9162 & ~n36264 ) ;
  assign n40800 = n28266 ^ n25725 ^ n23761 ;
  assign n40802 = n9372 ^ n2920 ^ 1'b0 ;
  assign n40801 = n26467 ^ n19880 ^ n9893 ;
  assign n40803 = n40802 ^ n40801 ^ n21420 ;
  assign n40804 = n3367 & ~n25626 ;
  assign n40805 = n40804 ^ n15336 ^ 1'b0 ;
  assign n40806 = ( n10583 & ~n17612 ) | ( n10583 & n29490 ) | ( ~n17612 & n29490 ) ;
  assign n40807 = n40806 ^ n6669 ^ x162 ;
  assign n40808 = n17016 ^ n16062 ^ 1'b0 ;
  assign n40809 = n31542 & n40808 ;
  assign n40810 = n40809 ^ n21027 ^ 1'b0 ;
  assign n40811 = ( n18123 & n40807 ) | ( n18123 & ~n40810 ) | ( n40807 & ~n40810 ) ;
  assign n40812 = ( n4044 & n22145 ) | ( n4044 & n36469 ) | ( n22145 & n36469 ) ;
  assign n40813 = ( ~n2493 & n13469 ) | ( ~n2493 & n19263 ) | ( n13469 & n19263 ) ;
  assign n40814 = n40813 ^ n26065 ^ 1'b0 ;
  assign n40815 = n9833 & ~n12823 ;
  assign n40816 = n40815 ^ n6958 ^ 1'b0 ;
  assign n40817 = ( n1060 & n6337 ) | ( n1060 & n40816 ) | ( n6337 & n40816 ) ;
  assign n40818 = ( n7124 & n12769 ) | ( n7124 & n20050 ) | ( n12769 & n20050 ) ;
  assign n40819 = ~n3482 & n7152 ;
  assign n40820 = n40819 ^ n20526 ^ n9374 ;
  assign n40821 = ( n22609 & n31220 ) | ( n22609 & ~n40820 ) | ( n31220 & ~n40820 ) ;
  assign n40822 = ( n4003 & ~n35810 ) | ( n4003 & n40821 ) | ( ~n35810 & n40821 ) ;
  assign n40823 = ( n13933 & n40818 ) | ( n13933 & n40822 ) | ( n40818 & n40822 ) ;
  assign n40824 = ~n4170 & n20950 ;
  assign n40825 = n40824 ^ n25307 ^ n20805 ;
  assign n40826 = n18582 | n40825 ;
  assign n40827 = ~n11234 & n25856 ;
  assign n40828 = ~n18322 & n40827 ;
  assign n40829 = ( ~n25118 & n28547 ) | ( ~n25118 & n40828 ) | ( n28547 & n40828 ) ;
  assign n40830 = n39192 & n40829 ;
  assign n40831 = ( ~n6968 & n17831 ) | ( ~n6968 & n32864 ) | ( n17831 & n32864 ) ;
  assign n40832 = n40831 ^ n26327 ^ 1'b0 ;
  assign n40833 = n40832 ^ n25463 ^ n11926 ;
  assign n40834 = n40833 ^ n13180 ^ 1'b0 ;
  assign n40835 = n28503 ^ n27089 ^ 1'b0 ;
  assign n40836 = ( n19905 & n27055 ) | ( n19905 & ~n40835 ) | ( n27055 & ~n40835 ) ;
  assign n40837 = ( n8669 & n25314 ) | ( n8669 & n40836 ) | ( n25314 & n40836 ) ;
  assign n40838 = n20723 | n29490 ;
  assign n40839 = n40838 ^ n21300 ^ 1'b0 ;
  assign n40840 = ( n23462 & ~n40038 ) | ( n23462 & n40839 ) | ( ~n40038 & n40839 ) ;
  assign n40841 = ( n1534 & n29803 ) | ( n1534 & n39072 ) | ( n29803 & n39072 ) ;
  assign n40842 = n40841 ^ n40325 ^ n25616 ;
  assign n40843 = ( n34602 & n39501 ) | ( n34602 & n40010 ) | ( n39501 & n40010 ) ;
  assign n40844 = n40457 ^ n14123 ^ n12308 ;
  assign n40845 = n2170 & n21460 ;
  assign n40846 = n16783 | n28588 ;
  assign n40847 = n36884 & ~n40846 ;
  assign n40848 = n1335 | n40847 ;
  assign n40849 = n40845 | n40848 ;
  assign n40850 = ( n8011 & n8714 ) | ( n8011 & n20748 ) | ( n8714 & n20748 ) ;
  assign n40851 = n40850 ^ n11500 ^ 1'b0 ;
  assign n40852 = n4358 & n15951 ;
  assign n40853 = ( n1833 & ~n14569 ) | ( n1833 & n40852 ) | ( ~n14569 & n40852 ) ;
  assign n40854 = n40853 ^ n9935 ^ n2566 ;
  assign n40855 = ( n20779 & n36849 ) | ( n20779 & n40854 ) | ( n36849 & n40854 ) ;
  assign n40856 = n33415 & n37851 ;
  assign n40857 = ( n22984 & ~n32316 ) | ( n22984 & n40856 ) | ( ~n32316 & n40856 ) ;
  assign n40858 = n22468 ^ n21819 ^ n20940 ;
  assign n40859 = ( ~n21585 & n24715 ) | ( ~n21585 & n40858 ) | ( n24715 & n40858 ) ;
  assign n40860 = n37698 ^ n36414 ^ n12196 ;
  assign n40861 = n23400 & ~n40860 ;
  assign n40862 = n40861 ^ n35165 ^ 1'b0 ;
  assign n40863 = ( ~n14238 & n39763 ) | ( ~n14238 & n40862 ) | ( n39763 & n40862 ) ;
  assign n40864 = n10654 & n34302 ;
  assign n40865 = ( n10647 & n19623 ) | ( n10647 & n40864 ) | ( n19623 & n40864 ) ;
  assign n40866 = n28937 | n31297 ;
  assign n40867 = n40865 & ~n40866 ;
  assign n40868 = n21210 ^ n6711 ^ n915 ;
  assign n40869 = ( n11806 & ~n14872 ) | ( n11806 & n40868 ) | ( ~n14872 & n40868 ) ;
  assign n40870 = n23998 ^ n6576 ^ n5055 ;
  assign n40871 = n40870 ^ n29852 ^ n4802 ;
  assign n40879 = ( ~n1779 & n6131 ) | ( ~n1779 & n36461 ) | ( n6131 & n36461 ) ;
  assign n40872 = n2542 | n6443 ;
  assign n40873 = n20897 | n40872 ;
  assign n40874 = ~n10776 & n17306 ;
  assign n40875 = n40874 ^ n34462 ^ 1'b0 ;
  assign n40876 = ( n2225 & n40873 ) | ( n2225 & ~n40875 ) | ( n40873 & ~n40875 ) ;
  assign n40877 = n27504 ^ n22089 ^ 1'b0 ;
  assign n40878 = ( n4131 & n40876 ) | ( n4131 & n40877 ) | ( n40876 & n40877 ) ;
  assign n40880 = n40879 ^ n40878 ^ 1'b0 ;
  assign n40881 = ~n6243 & n10897 ;
  assign n40882 = ( n15336 & n18678 ) | ( n15336 & ~n40881 ) | ( n18678 & ~n40881 ) ;
  assign n40883 = ( n2441 & n7202 ) | ( n2441 & n24770 ) | ( n7202 & n24770 ) ;
  assign n40884 = ( ~n15393 & n34789 ) | ( ~n15393 & n40883 ) | ( n34789 & n40883 ) ;
  assign n40888 = n26693 ^ n12894 ^ n3990 ;
  assign n40889 = ( ~n9523 & n12817 ) | ( ~n9523 & n40888 ) | ( n12817 & n40888 ) ;
  assign n40890 = n40889 ^ n28539 ^ n4559 ;
  assign n40885 = n4670 | n13975 ;
  assign n40886 = ( n5015 & n25197 ) | ( n5015 & ~n40885 ) | ( n25197 & ~n40885 ) ;
  assign n40887 = n40886 ^ n21394 ^ n10241 ;
  assign n40891 = n40890 ^ n40887 ^ n21610 ;
  assign n40892 = n9126 & n10186 ;
  assign n40893 = n23266 ^ n6028 ^ 1'b0 ;
  assign n40894 = n29785 | n40893 ;
  assign n40895 = n8454 & ~n16877 ;
  assign n40896 = ( n17466 & n24669 ) | ( n17466 & ~n32641 ) | ( n24669 & ~n32641 ) ;
  assign n40901 = n9206 & n22158 ;
  assign n40897 = n16228 ^ n7013 ^ 1'b0 ;
  assign n40898 = n7125 & ~n22628 ;
  assign n40899 = n4034 & n40898 ;
  assign n40900 = n40897 | n40899 ;
  assign n40902 = n40901 ^ n40900 ^ n7443 ;
  assign n40903 = n19965 & n40902 ;
  assign n40904 = n40903 ^ n15092 ^ 1'b0 ;
  assign n40905 = n40904 ^ n37553 ^ n22210 ;
  assign n40906 = n36777 ^ n17468 ^ n4840 ;
  assign n40907 = n40906 ^ n32236 ^ n27065 ;
  assign n40908 = n35694 ^ n14323 ^ 1'b0 ;
  assign n40913 = n23633 ^ n3418 ^ 1'b0 ;
  assign n40914 = n5613 | n40913 ;
  assign n40915 = n40914 ^ n29472 ^ 1'b0 ;
  assign n40916 = n40915 ^ n16155 ^ n7079 ;
  assign n40911 = n24668 & n28799 ;
  assign n40909 = ( ~n11937 & n18013 ) | ( ~n11937 & n36567 ) | ( n18013 & n36567 ) ;
  assign n40910 = n40909 ^ n17460 ^ 1'b0 ;
  assign n40912 = n40911 ^ n40910 ^ n14820 ;
  assign n40917 = n40916 ^ n40912 ^ n30801 ;
  assign n40918 = n1872 & n10500 ;
  assign n40919 = ~n21466 & n40918 ;
  assign n40920 = n40919 ^ n36083 ^ n20718 ;
  assign n40921 = n36568 | n38927 ;
  assign n40922 = n18044 & ~n40921 ;
  assign n40924 = n1024 & ~n14595 ;
  assign n40925 = ~n4251 & n40924 ;
  assign n40926 = n40925 ^ n36021 ^ n32180 ;
  assign n40923 = n32543 ^ n14989 ^ n8948 ;
  assign n40927 = n40926 ^ n40923 ^ n36770 ;
  assign n40928 = ~n9653 & n25942 ;
  assign n40929 = n10877 ^ n8210 ^ n6281 ;
  assign n40930 = n27841 ^ n20296 ^ n16786 ;
  assign n40931 = ( n37203 & n40929 ) | ( n37203 & n40930 ) | ( n40929 & n40930 ) ;
  assign n40932 = ( ~n11864 & n40458 ) | ( ~n11864 & n40931 ) | ( n40458 & n40931 ) ;
  assign n40933 = ( ~n31304 & n38380 ) | ( ~n31304 & n40932 ) | ( n38380 & n40932 ) ;
  assign n40934 = ( n687 & n9635 ) | ( n687 & ~n30077 ) | ( n9635 & ~n30077 ) ;
  assign n40935 = n40934 ^ n40651 ^ n26903 ;
  assign n40936 = ( ~n13656 & n16081 ) | ( ~n13656 & n29046 ) | ( n16081 & n29046 ) ;
  assign n40937 = n18732 ^ n2109 ^ 1'b0 ;
  assign n40938 = n18664 & ~n40937 ;
  assign n40939 = ~n35602 & n40938 ;
  assign n40940 = ~n37060 & n40939 ;
  assign n40941 = ~n10882 & n35460 ;
  assign n40942 = n40941 ^ n23290 ^ 1'b0 ;
  assign n40943 = ( n23320 & n26410 ) | ( n23320 & n30198 ) | ( n26410 & n30198 ) ;
  assign n40944 = n25693 ^ n16528 ^ n10844 ;
  assign n40945 = n28743 & ~n38957 ;
  assign n40946 = n9859 ^ n414 ^ 1'b0 ;
  assign n40947 = n22856 ^ n9271 ^ n1398 ;
  assign n40948 = ( n11566 & n17140 ) | ( n11566 & ~n40947 ) | ( n17140 & ~n40947 ) ;
  assign n40949 = ( ~n411 & n10582 ) | ( ~n411 & n22560 ) | ( n10582 & n22560 ) ;
  assign n40950 = n40949 ^ n12259 ^ n1939 ;
  assign n40951 = ~n402 & n40950 ;
  assign n40952 = ~n5182 & n9517 ;
  assign n40953 = n40952 ^ n12641 ^ 1'b0 ;
  assign n40954 = ( n6999 & ~n8270 ) | ( n6999 & n17398 ) | ( ~n8270 & n17398 ) ;
  assign n40955 = n4282 | n32630 ;
  assign n40956 = n40955 ^ n9685 ^ 1'b0 ;
  assign n40957 = n40956 ^ n21676 ^ n11263 ;
  assign n40958 = n23758 ^ n3695 ^ n2467 ;
  assign n40959 = n2840 & ~n6995 ;
  assign n40960 = n36998 & n40959 ;
  assign n40961 = n40960 ^ n34602 ^ n17576 ;
  assign n40962 = ( n9076 & n13319 ) | ( n9076 & n22892 ) | ( n13319 & n22892 ) ;
  assign n40963 = ( n16723 & ~n26745 ) | ( n16723 & n40962 ) | ( ~n26745 & n40962 ) ;
  assign n40964 = ( n12508 & ~n12822 ) | ( n12508 & n37346 ) | ( ~n12822 & n37346 ) ;
  assign n40965 = n32778 ^ n27206 ^ n18376 ;
  assign n40967 = n10462 | n30833 ;
  assign n40966 = n2829 & n8296 ;
  assign n40968 = n40967 ^ n40966 ^ 1'b0 ;
  assign n40969 = n29539 & ~n31779 ;
  assign n40970 = ~n28210 & n40969 ;
  assign n40974 = n29281 ^ n8642 ^ 1'b0 ;
  assign n40975 = n699 & n40974 ;
  assign n40976 = ( n4021 & n28890 ) | ( n4021 & n40975 ) | ( n28890 & n40975 ) ;
  assign n40971 = n9157 ^ n7081 ^ 1'b0 ;
  assign n40972 = n37962 ^ n31252 ^ 1'b0 ;
  assign n40973 = n40971 & n40972 ;
  assign n40977 = n40976 ^ n40973 ^ n13059 ;
  assign n40978 = n17619 ^ n1482 ^ 1'b0 ;
  assign n40979 = n5782 & n9128 ;
  assign n40980 = ( ~n3767 & n40978 ) | ( ~n3767 & n40979 ) | ( n40978 & n40979 ) ;
  assign n40981 = n18021 ^ n12565 ^ 1'b0 ;
  assign n40982 = n9467 & n40981 ;
  assign n40983 = n40982 ^ n24658 ^ n8093 ;
  assign n40984 = ( n7941 & n40980 ) | ( n7941 & ~n40983 ) | ( n40980 & ~n40983 ) ;
  assign n40985 = n40550 ^ n14843 ^ n7648 ;
  assign n40986 = n40985 ^ n19515 ^ n661 ;
  assign n40987 = n36668 ^ n3932 ^ 1'b0 ;
  assign n40988 = ( n353 & ~n6050 ) | ( n353 & n36869 ) | ( ~n6050 & n36869 ) ;
  assign n40989 = ( ~n6733 & n18639 ) | ( ~n6733 & n22158 ) | ( n18639 & n22158 ) ;
  assign n40990 = n32474 | n40989 ;
  assign n40991 = n33494 & ~n40990 ;
  assign n40992 = n40991 ^ n24025 ^ 1'b0 ;
  assign n40994 = ~n9519 & n11946 ;
  assign n40993 = n26956 ^ n23363 ^ n10879 ;
  assign n40995 = n40994 ^ n40993 ^ n17311 ;
  assign n40996 = ( ~n15263 & n40992 ) | ( ~n15263 & n40995 ) | ( n40992 & n40995 ) ;
  assign n40997 = n16456 ^ n2247 ^ 1'b0 ;
  assign n40998 = ~n26853 & n40997 ;
  assign n40999 = n38333 ^ n29690 ^ n14413 ;
  assign n41000 = n40999 ^ n37442 ^ 1'b0 ;
  assign n41001 = n33969 | n41000 ;
  assign n41003 = n30752 ^ n20447 ^ n2392 ;
  assign n41002 = x87 & n35729 ;
  assign n41004 = n41003 ^ n41002 ^ 1'b0 ;
  assign n41005 = n6995 | n8292 ;
  assign n41006 = n8247 | n41005 ;
  assign n41007 = n41006 ^ n35016 ^ 1'b0 ;
  assign n41008 = n15995 | n41007 ;
  assign n41009 = n41008 ^ n23123 ^ n3935 ;
  assign n41010 = ( n11281 & n21799 ) | ( n11281 & ~n40061 ) | ( n21799 & ~n40061 ) ;
  assign n41011 = n28478 & ~n41010 ;
  assign n41012 = n41009 & n41011 ;
  assign n41014 = n16858 ^ n8497 ^ n6282 ;
  assign n41013 = n19327 ^ n9927 ^ 1'b0 ;
  assign n41015 = n41014 ^ n41013 ^ n21632 ;
  assign n41016 = ( n982 & ~n12042 ) | ( n982 & n37808 ) | ( ~n12042 & n37808 ) ;
  assign n41017 = n14359 | n41016 ;
  assign n41018 = ( n11740 & n15061 ) | ( n11740 & ~n30931 ) | ( n15061 & ~n30931 ) ;
  assign n41019 = ( n14945 & n34581 ) | ( n14945 & n41018 ) | ( n34581 & n41018 ) ;
  assign n41020 = ( n26022 & ~n41017 ) | ( n26022 & n41019 ) | ( ~n41017 & n41019 ) ;
  assign n41021 = ( n1370 & n13998 ) | ( n1370 & n25524 ) | ( n13998 & n25524 ) ;
  assign n41022 = n41021 ^ n3224 ^ 1'b0 ;
  assign n41023 = ( n23261 & ~n40220 ) | ( n23261 & n41022 ) | ( ~n40220 & n41022 ) ;
  assign n41024 = ( n6126 & n33738 ) | ( n6126 & ~n41023 ) | ( n33738 & ~n41023 ) ;
  assign n41025 = n41024 ^ n34381 ^ n11164 ;
  assign n41026 = n37014 ^ n22206 ^ n4439 ;
  assign n41027 = ( n3583 & n17237 ) | ( n3583 & ~n17421 ) | ( n17237 & ~n17421 ) ;
  assign n41028 = n41027 ^ n38344 ^ 1'b0 ;
  assign n41029 = ~n41026 & n41028 ;
  assign n41032 = ( n2278 & n7466 ) | ( n2278 & ~n19308 ) | ( n7466 & ~n19308 ) ;
  assign n41030 = ( n2587 & ~n25269 ) | ( n2587 & n25701 ) | ( ~n25269 & n25701 ) ;
  assign n41031 = ( n3573 & ~n24745 ) | ( n3573 & n41030 ) | ( ~n24745 & n41030 ) ;
  assign n41033 = n41032 ^ n41031 ^ n11821 ;
  assign n41034 = n41033 ^ n6712 ^ 1'b0 ;
  assign n41035 = n26452 ^ n5628 ^ n1660 ;
  assign n41036 = ( n968 & ~n23920 ) | ( n968 & n41035 ) | ( ~n23920 & n41035 ) ;
  assign n41037 = n41036 ^ n3004 ^ 1'b0 ;
  assign n41038 = n5460 & n36057 ;
  assign n41039 = ( n4355 & n18162 ) | ( n4355 & n18392 ) | ( n18162 & n18392 ) ;
  assign n41040 = ( n2566 & n22730 ) | ( n2566 & ~n41039 ) | ( n22730 & ~n41039 ) ;
  assign n41041 = ( n7302 & n8686 ) | ( n7302 & ~n15406 ) | ( n8686 & ~n15406 ) ;
  assign n41042 = ( n20019 & n28577 ) | ( n20019 & n41041 ) | ( n28577 & n41041 ) ;
  assign n41043 = ( ~n16958 & n22313 ) | ( ~n16958 & n41042 ) | ( n22313 & n41042 ) ;
  assign n41044 = ( n38514 & n41035 ) | ( n38514 & n41043 ) | ( n41035 & n41043 ) ;
  assign n41045 = n41040 | n41044 ;
  assign n41046 = ( n8711 & n17262 ) | ( n8711 & ~n32398 ) | ( n17262 & ~n32398 ) ;
  assign n41047 = n17809 & n41046 ;
  assign n41048 = n41047 ^ n21006 ^ 1'b0 ;
  assign n41049 = n24061 ^ n14808 ^ n3859 ;
  assign n41050 = n25096 ^ n21680 ^ n13776 ;
  assign n41051 = n34175 ^ n16827 ^ n15860 ;
  assign n41052 = ( n6285 & ~n12068 ) | ( n6285 & n41051 ) | ( ~n12068 & n41051 ) ;
  assign n41053 = ( ~n1279 & n2457 ) | ( ~n1279 & n17619 ) | ( n2457 & n17619 ) ;
  assign n41054 = n41053 ^ n17876 ^ n11269 ;
  assign n41055 = ( ~n16641 & n41052 ) | ( ~n16641 & n41054 ) | ( n41052 & n41054 ) ;
  assign n41056 = ( n6845 & ~n12053 ) | ( n6845 & n33811 ) | ( ~n12053 & n33811 ) ;
  assign n41057 = n41056 ^ n15116 ^ n3490 ;
  assign n41058 = n18857 ^ n4506 ^ n1117 ;
  assign n41059 = n41058 ^ n28617 ^ n8285 ;
  assign n41060 = n6926 ^ n3764 ^ n3146 ;
  assign n41061 = ( n16529 & n23123 ) | ( n16529 & n25903 ) | ( n23123 & n25903 ) ;
  assign n41062 = ( n4465 & ~n41060 ) | ( n4465 & n41061 ) | ( ~n41060 & n41061 ) ;
  assign n41063 = n41062 ^ n37346 ^ 1'b0 ;
  assign n41064 = n25388 ^ n10128 ^ n9953 ;
  assign n41065 = ( ~n33386 & n34959 ) | ( ~n33386 & n41064 ) | ( n34959 & n41064 ) ;
  assign n41066 = n27945 ^ n15167 ^ n1062 ;
  assign n41067 = ( n1242 & n18913 ) | ( n1242 & n41066 ) | ( n18913 & n41066 ) ;
  assign n41068 = n25873 & ~n41067 ;
  assign n41069 = n41068 ^ n36762 ^ 1'b0 ;
  assign n41070 = n41069 ^ n11309 ^ n10500 ;
  assign n41071 = n33589 ^ n4085 ^ 1'b0 ;
  assign n41072 = ( x184 & n5195 ) | ( x184 & n6095 ) | ( n5195 & n6095 ) ;
  assign n41073 = n41072 ^ n20907 ^ n11203 ;
  assign n41074 = ( n5238 & n41071 ) | ( n5238 & ~n41073 ) | ( n41071 & ~n41073 ) ;
  assign n41075 = n19485 ^ n18984 ^ n5941 ;
  assign n41076 = n41075 ^ n11151 ^ n2976 ;
  assign n41077 = ~n35182 & n40219 ;
  assign n41078 = n41076 & n41077 ;
  assign n41079 = n41078 ^ n28101 ^ n17318 ;
  assign n41080 = ( ~n18331 & n21034 ) | ( ~n18331 & n23746 ) | ( n21034 & n23746 ) ;
  assign n41081 = n15060 | n41080 ;
  assign n41085 = ~n8094 & n34073 ;
  assign n41082 = n5413 & ~n17404 ;
  assign n41083 = n41082 ^ n31017 ^ n15181 ;
  assign n41084 = n41083 ^ n19102 ^ n13279 ;
  assign n41086 = n41085 ^ n41084 ^ n1659 ;
  assign n41089 = ( n722 & n6463 ) | ( n722 & n7961 ) | ( n6463 & n7961 ) ;
  assign n41090 = n21188 & ~n41089 ;
  assign n41091 = ~n12797 & n41090 ;
  assign n41092 = n3272 | n41091 ;
  assign n41087 = n24371 & ~n32612 ;
  assign n41088 = n41087 ^ n40787 ^ 1'b0 ;
  assign n41093 = n41092 ^ n41088 ^ 1'b0 ;
  assign n41094 = n8662 ^ n3932 ^ n2973 ;
  assign n41095 = n20509 & n34742 ;
  assign n41096 = ~n41094 & n41095 ;
  assign n41097 = n6884 & n7537 ;
  assign n41098 = n41097 ^ n1889 ^ 1'b0 ;
  assign n41099 = n16951 & ~n41098 ;
  assign n41100 = n41099 ^ n18475 ^ 1'b0 ;
  assign n41101 = ( n3932 & ~n8685 ) | ( n3932 & n18204 ) | ( ~n8685 & n18204 ) ;
  assign n41102 = ( ~n15072 & n34335 ) | ( ~n15072 & n41101 ) | ( n34335 & n41101 ) ;
  assign n41103 = ( n29566 & n41100 ) | ( n29566 & n41102 ) | ( n41100 & n41102 ) ;
  assign n41104 = n41103 ^ n10085 ^ n6876 ;
  assign n41105 = n34944 ^ n13969 ^ n10094 ;
  assign n41106 = n28144 ^ n692 ^ 1'b0 ;
  assign n41107 = n20441 & n41106 ;
  assign n41108 = n41107 ^ n8885 ^ 1'b0 ;
  assign n41109 = ( x143 & n868 ) | ( x143 & n5185 ) | ( n868 & n5185 ) ;
  assign n41110 = ( n7759 & n8151 ) | ( n7759 & ~n41109 ) | ( n8151 & ~n41109 ) ;
  assign n41111 = ( n7023 & ~n16788 ) | ( n7023 & n37931 ) | ( ~n16788 & n37931 ) ;
  assign n41112 = n41111 ^ n37508 ^ n10914 ;
  assign n41113 = n37879 & n41112 ;
  assign n41114 = n35740 ^ n16868 ^ n4676 ;
  assign n41115 = n41114 ^ n29799 ^ n15034 ;
  assign n41116 = ~n19531 & n41115 ;
  assign n41117 = n35834 ^ n35513 ^ n2985 ;
  assign n41118 = ~n16627 & n41006 ;
  assign n41119 = ~n4213 & n41118 ;
  assign n41120 = ( n7245 & ~n17190 ) | ( n7245 & n41119 ) | ( ~n17190 & n41119 ) ;
  assign n41121 = n14364 ^ n12516 ^ 1'b0 ;
  assign n41122 = n41121 ^ n40204 ^ n8082 ;
  assign n41123 = n30226 ^ n16877 ^ n5312 ;
  assign n41127 = n3747 & ~n19849 ;
  assign n41125 = n9189 | n19060 ;
  assign n41126 = n3202 & ~n41125 ;
  assign n41124 = n8836 ^ n7849 ^ n7191 ;
  assign n41128 = n41127 ^ n41126 ^ n41124 ;
  assign n41129 = n7614 | n31554 ;
  assign n41130 = n41129 ^ n11027 ^ 1'b0 ;
  assign n41131 = n41130 ^ n36545 ^ n16435 ;
  assign n41132 = n14315 ^ n323 ^ 1'b0 ;
  assign n41133 = n41132 ^ n31561 ^ n22479 ;
  assign n41134 = n32609 ^ x11 ^ 1'b0 ;
  assign n41135 = ~n22323 & n41134 ;
  assign n41136 = ( n7689 & n12556 ) | ( n7689 & ~n28630 ) | ( n12556 & ~n28630 ) ;
  assign n41137 = ( n6597 & ~n27861 ) | ( n6597 & n41136 ) | ( ~n27861 & n41136 ) ;
  assign n41138 = n9933 & n41137 ;
  assign n41139 = n8545 | n41138 ;
  assign n41140 = n41139 ^ n32150 ^ 1'b0 ;
  assign n41141 = n15592 | n16023 ;
  assign n41142 = ( ~n18394 & n41140 ) | ( ~n18394 & n41141 ) | ( n41140 & n41141 ) ;
  assign n41143 = ( ~n11236 & n27219 ) | ( ~n11236 & n31074 ) | ( n27219 & n31074 ) ;
  assign n41144 = n24316 & ~n32391 ;
  assign n41145 = ( n8577 & n12587 ) | ( n8577 & ~n20366 ) | ( n12587 & ~n20366 ) ;
  assign n41146 = n7292 & n17470 ;
  assign n41147 = n4285 & n41146 ;
  assign n41148 = ( n19117 & n26872 ) | ( n19117 & n41147 ) | ( n26872 & n41147 ) ;
  assign n41149 = ~n17500 & n25401 ;
  assign n41150 = ~n41148 & n41149 ;
  assign n41151 = n30432 ^ n15526 ^ 1'b0 ;
  assign n41152 = n36370 ^ n16323 ^ n15881 ;
  assign n41153 = n30012 ^ n24615 ^ n21831 ;
  assign n41154 = ( n6711 & ~n9343 ) | ( n6711 & n11899 ) | ( ~n9343 & n11899 ) ;
  assign n41155 = ( n365 & ~n20296 ) | ( n365 & n22083 ) | ( ~n20296 & n22083 ) ;
  assign n41156 = n41155 ^ n10550 ^ n2807 ;
  assign n41157 = ( n28188 & ~n41154 ) | ( n28188 & n41156 ) | ( ~n41154 & n41156 ) ;
  assign n41158 = ( n38403 & n41153 ) | ( n38403 & ~n41157 ) | ( n41153 & ~n41157 ) ;
  assign n41159 = ( n19046 & n19883 ) | ( n19046 & ~n21663 ) | ( n19883 & ~n21663 ) ;
  assign n41160 = n26646 | n29260 ;
  assign n41161 = n41160 ^ n28804 ^ 1'b0 ;
  assign n41162 = n41161 ^ n7157 ^ n873 ;
  assign n41163 = ( ~n2676 & n3074 ) | ( ~n2676 & n20416 ) | ( n3074 & n20416 ) ;
  assign n41168 = x31 & n27888 ;
  assign n41169 = n21373 & n41168 ;
  assign n41170 = n41169 ^ n12838 ^ n11447 ;
  assign n41171 = ( n10323 & ~n14862 ) | ( n10323 & n33819 ) | ( ~n14862 & n33819 ) ;
  assign n41172 = n41171 ^ n8007 ^ n3990 ;
  assign n41173 = n41170 & n41172 ;
  assign n41174 = n41173 ^ n23813 ^ n7085 ;
  assign n41164 = n31437 ^ n18524 ^ n4460 ;
  assign n41165 = ( n13690 & n27562 ) | ( n13690 & n41164 ) | ( n27562 & n41164 ) ;
  assign n41166 = n41165 ^ n22083 ^ n12135 ;
  assign n41167 = n8353 & ~n41166 ;
  assign n41175 = n41174 ^ n41167 ^ 1'b0 ;
  assign n41176 = n7944 ^ n4774 ^ 1'b0 ;
  assign n41177 = x102 & ~n41176 ;
  assign n41178 = ~n993 & n13415 ;
  assign n41179 = n17802 & n41178 ;
  assign n41180 = ~n18493 & n18911 ;
  assign n41181 = n41180 ^ n21590 ^ 1'b0 ;
  assign n41182 = n29319 ^ n11261 ^ 1'b0 ;
  assign n41183 = ( n37788 & n41181 ) | ( n37788 & ~n41182 ) | ( n41181 & ~n41182 ) ;
  assign n41186 = ( x127 & ~n3564 ) | ( x127 & n9476 ) | ( ~n3564 & n9476 ) ;
  assign n41184 = n20524 | n24338 ;
  assign n41185 = n13401 & n41184 ;
  assign n41187 = n41186 ^ n41185 ^ 1'b0 ;
  assign n41188 = ( ~n19613 & n41183 ) | ( ~n19613 & n41187 ) | ( n41183 & n41187 ) ;
  assign n41189 = n10893 ^ n4860 ^ n937 ;
  assign n41190 = n18634 & ~n41189 ;
  assign n41191 = ~n873 & n41190 ;
  assign n41192 = n41191 ^ n35970 ^ n13974 ;
  assign n41193 = ( x252 & n33899 ) | ( x252 & n41192 ) | ( n33899 & n41192 ) ;
  assign n41194 = ( n6281 & n13506 ) | ( n6281 & n16128 ) | ( n13506 & n16128 ) ;
  assign n41195 = n6134 & ~n41194 ;
  assign n41196 = ~n7598 & n41195 ;
  assign n41197 = ( n6913 & n19936 ) | ( n6913 & n41196 ) | ( n19936 & n41196 ) ;
  assign n41198 = ( n18721 & n27419 ) | ( n18721 & n41197 ) | ( n27419 & n41197 ) ;
  assign n41208 = n27413 ^ n17985 ^ n9608 ;
  assign n41206 = n8977 | n22468 ;
  assign n41204 = n10369 ^ n4150 ^ n1674 ;
  assign n41199 = n6111 & ~n6368 ;
  assign n41200 = n32015 & n41199 ;
  assign n41201 = n20335 ^ n1188 ^ 1'b0 ;
  assign n41202 = ~n2490 & n41201 ;
  assign n41203 = ( n15488 & n41200 ) | ( n15488 & n41202 ) | ( n41200 & n41202 ) ;
  assign n41205 = n41204 ^ n41203 ^ n40304 ;
  assign n41207 = n41206 ^ n41205 ^ n38737 ;
  assign n41209 = n41208 ^ n41207 ^ n10607 ;
  assign n41210 = n10094 ^ n8497 ^ n2168 ;
  assign n41211 = n41210 ^ n25973 ^ n11612 ;
  assign n41212 = ( n866 & ~n33897 ) | ( n866 & n41211 ) | ( ~n33897 & n41211 ) ;
  assign n41213 = n7431 ^ n4030 ^ n1595 ;
  assign n41214 = n34742 & ~n41213 ;
  assign n41215 = ~x218 & n41214 ;
  assign n41216 = n14156 ^ n8304 ^ 1'b0 ;
  assign n41217 = ~n15101 & n41216 ;
  assign n41219 = ( ~n11804 & n19006 ) | ( ~n11804 & n23393 ) | ( n19006 & n23393 ) ;
  assign n41218 = n10315 | n22227 ;
  assign n41220 = n41219 ^ n41218 ^ 1'b0 ;
  assign n41221 = n41220 ^ n33914 ^ 1'b0 ;
  assign n41222 = n12252 ^ n1128 ^ 1'b0 ;
  assign n41223 = n41222 ^ n25337 ^ n6582 ;
  assign n41224 = n37814 ^ n4834 ^ 1'b0 ;
  assign n41225 = n1304 & ~n41224 ;
  assign n41226 = ( n4035 & n41223 ) | ( n4035 & n41225 ) | ( n41223 & n41225 ) ;
  assign n41227 = ( n11893 & ~n14232 ) | ( n11893 & n41226 ) | ( ~n14232 & n41226 ) ;
  assign n41228 = n35395 ^ n18162 ^ n11304 ;
  assign n41229 = ( n7397 & n18822 ) | ( n7397 & n30588 ) | ( n18822 & n30588 ) ;
  assign n41230 = n9936 & n24904 ;
  assign n41231 = ( n1638 & n4753 ) | ( n1638 & ~n36994 ) | ( n4753 & ~n36994 ) ;
  assign n41232 = n41231 ^ n10207 ^ 1'b0 ;
  assign n41233 = n16659 ^ x69 ^ 1'b0 ;
  assign n41234 = n17857 | n41233 ;
  assign n41235 = ( ~n2323 & n41232 ) | ( ~n2323 & n41234 ) | ( n41232 & n41234 ) ;
  assign n41236 = n34916 ^ n5915 ^ 1'b0 ;
  assign n41237 = n41236 ^ n8203 ^ n7241 ;
  assign n41238 = n32468 ^ n9916 ^ 1'b0 ;
  assign n41239 = ~n41237 & n41238 ;
  assign n41242 = ~n703 & n10492 ;
  assign n41243 = n41242 ^ n33036 ^ 1'b0 ;
  assign n41240 = ( ~n1481 & n26189 ) | ( ~n1481 & n38383 ) | ( n26189 & n38383 ) ;
  assign n41241 = n20895 & ~n41240 ;
  assign n41244 = n41243 ^ n41241 ^ 1'b0 ;
  assign n41245 = n23422 ^ n472 ^ 1'b0 ;
  assign n41246 = ~n15312 & n41245 ;
  assign n41247 = n36425 & n41246 ;
  assign n41248 = n25587 ^ n24634 ^ n11431 ;
  assign n41249 = n41248 ^ n26011 ^ n20902 ;
  assign n41250 = ( ~n21280 & n25472 ) | ( ~n21280 & n41249 ) | ( n25472 & n41249 ) ;
  assign n41251 = ( n33692 & n41247 ) | ( n33692 & n41250 ) | ( n41247 & n41250 ) ;
  assign n41252 = n9686 & n11141 ;
  assign n41253 = ~n36647 & n41252 ;
  assign n41254 = n23839 ^ n12896 ^ n2691 ;
  assign n41255 = n41254 ^ n32501 ^ 1'b0 ;
  assign n41256 = ( n13202 & ~n22023 ) | ( n13202 & n35818 ) | ( ~n22023 & n35818 ) ;
  assign n41257 = ( ~n18932 & n25924 ) | ( ~n18932 & n41256 ) | ( n25924 & n41256 ) ;
  assign n41258 = ( n10982 & n15294 ) | ( n10982 & n37631 ) | ( n15294 & n37631 ) ;
  assign n41259 = n13781 | n41258 ;
  assign n41260 = n13380 ^ n509 ^ x235 ;
  assign n41261 = n3651 & n3882 ;
  assign n41262 = n41260 & n41261 ;
  assign n41263 = ( x234 & n11251 ) | ( x234 & n41262 ) | ( n11251 & n41262 ) ;
  assign n41264 = n41263 ^ n25781 ^ n5924 ;
  assign n41265 = n9382 ^ n7043 ^ n3235 ;
  assign n41266 = n41265 ^ n9289 ^ 1'b0 ;
  assign n41267 = n6421 & n41266 ;
  assign n41268 = ~n39300 & n41267 ;
  assign n41269 = n41268 ^ n20806 ^ 1'b0 ;
  assign n41270 = n7591 ^ n3697 ^ n1733 ;
  assign n41271 = n5774 | n41270 ;
  assign n41272 = n41271 ^ n28655 ^ n26354 ;
  assign n41273 = ( n23355 & n25734 ) | ( n23355 & ~n41272 ) | ( n25734 & ~n41272 ) ;
  assign n41275 = n17081 ^ n15184 ^ n1161 ;
  assign n41276 = ( ~n445 & n9683 ) | ( ~n445 & n41275 ) | ( n9683 & n41275 ) ;
  assign n41274 = n16323 ^ n9385 ^ n8400 ;
  assign n41277 = n41276 ^ n41274 ^ n3447 ;
  assign n41278 = ( n6349 & n6407 ) | ( n6349 & ~n17000 ) | ( n6407 & ~n17000 ) ;
  assign n41279 = n27870 ^ n15536 ^ n926 ;
  assign n41280 = ( ~n6450 & n41278 ) | ( ~n6450 & n41279 ) | ( n41278 & n41279 ) ;
  assign n41281 = n21113 ^ n10819 ^ 1'b0 ;
  assign n41282 = n3883 & ~n41281 ;
  assign n41283 = n18865 ^ n7689 ^ 1'b0 ;
  assign n41284 = ( n5318 & n41282 ) | ( n5318 & n41283 ) | ( n41282 & n41283 ) ;
  assign n41291 = n26913 ^ n11322 ^ 1'b0 ;
  assign n41289 = ( n3767 & n4203 ) | ( n3767 & n24680 ) | ( n4203 & n24680 ) ;
  assign n41287 = n15481 | n30910 ;
  assign n41288 = n41287 ^ n39381 ^ 1'b0 ;
  assign n41285 = n13596 ^ n4573 ^ n2644 ;
  assign n41286 = n41285 ^ n4379 ^ n2088 ;
  assign n41290 = n41289 ^ n41288 ^ n41286 ;
  assign n41292 = n41291 ^ n41290 ^ n12263 ;
  assign n41293 = ( n2688 & n3921 ) | ( n2688 & n5595 ) | ( n3921 & n5595 ) ;
  assign n41294 = n41293 ^ n25286 ^ n11604 ;
  assign n41295 = ( n6535 & ~n32449 ) | ( n6535 & n41294 ) | ( ~n32449 & n41294 ) ;
  assign n41296 = n41295 ^ n23222 ^ 1'b0 ;
  assign n41297 = n29282 | n41296 ;
  assign n41298 = n10006 & n21732 ;
  assign n41299 = n41298 ^ n6323 ^ 1'b0 ;
  assign n41300 = x40 & ~n14612 ;
  assign n41301 = ~n41299 & n41300 ;
  assign n41302 = n41301 ^ n15704 ^ n1559 ;
  assign n41303 = n12746 ^ n7350 ^ n6749 ;
  assign n41304 = ( ~n16408 & n34339 ) | ( ~n16408 & n34890 ) | ( n34339 & n34890 ) ;
  assign n41305 = n4618 | n20611 ;
  assign n41306 = n33073 ^ n9404 ^ n1213 ;
  assign n41307 = n8771 | n31957 ;
  assign n41308 = n13280 | n41307 ;
  assign n41309 = ( n6786 & ~n15191 ) | ( n6786 & n19688 ) | ( ~n15191 & n19688 ) ;
  assign n41310 = ~n3448 & n12894 ;
  assign n41311 = ~n41309 & n41310 ;
  assign n41312 = n29764 ^ n18535 ^ n12313 ;
  assign n41313 = ( ~n34115 & n37558 ) | ( ~n34115 & n41312 ) | ( n37558 & n41312 ) ;
  assign n41314 = ( n4938 & ~n8512 ) | ( n4938 & n24692 ) | ( ~n8512 & n24692 ) ;
  assign n41315 = n41314 ^ n10758 ^ 1'b0 ;
  assign n41316 = ( n3864 & n8806 ) | ( n3864 & n21678 ) | ( n8806 & n21678 ) ;
  assign n41317 = n32856 ^ n26956 ^ n11977 ;
  assign n41318 = n33352 ^ n32073 ^ n29683 ;
  assign n41319 = ( ~n6474 & n12665 ) | ( ~n6474 & n41318 ) | ( n12665 & n41318 ) ;
  assign n41320 = n17329 ^ n9666 ^ n2134 ;
  assign n41321 = ( n25608 & n39455 ) | ( n25608 & n41320 ) | ( n39455 & n41320 ) ;
  assign n41322 = ( n6899 & ~n9561 ) | ( n6899 & n20163 ) | ( ~n9561 & n20163 ) ;
  assign n41323 = n41322 ^ n6011 ^ n5542 ;
  assign n41324 = n33791 ^ n31401 ^ n593 ;
  assign n41325 = ( n4192 & n7250 ) | ( n4192 & ~n14808 ) | ( n7250 & ~n14808 ) ;
  assign n41326 = ( n19316 & ~n41324 ) | ( n19316 & n41325 ) | ( ~n41324 & n41325 ) ;
  assign n41327 = n5340 & n41326 ;
  assign n41328 = ( n10541 & n16142 ) | ( n10541 & ~n20887 ) | ( n16142 & ~n20887 ) ;
  assign n41329 = n41328 ^ n2132 ^ 1'b0 ;
  assign n41330 = n32956 & n41329 ;
  assign n41331 = n27262 ^ n9970 ^ n568 ;
  assign n41332 = n41331 ^ n29357 ^ n24076 ;
  assign n41333 = ( n1907 & n8577 ) | ( n1907 & ~n13574 ) | ( n8577 & ~n13574 ) ;
  assign n41334 = ( ~n4916 & n10010 ) | ( ~n4916 & n41333 ) | ( n10010 & n41333 ) ;
  assign n41335 = ( n20809 & ~n23519 ) | ( n20809 & n25320 ) | ( ~n23519 & n25320 ) ;
  assign n41336 = ( n5448 & n39868 ) | ( n5448 & ~n41335 ) | ( n39868 & ~n41335 ) ;
  assign n41337 = ( n21139 & ~n31777 ) | ( n21139 & n41336 ) | ( ~n31777 & n41336 ) ;
  assign n41338 = ( n36728 & ~n41334 ) | ( n36728 & n41337 ) | ( ~n41334 & n41337 ) ;
  assign n41339 = n11199 | n24505 ;
  assign n41340 = ~n16198 & n23573 ;
  assign n41341 = ( n33062 & n34004 ) | ( n33062 & ~n40442 ) | ( n34004 & ~n40442 ) ;
  assign n41343 = ~n5496 & n15972 ;
  assign n41344 = ~n29188 & n41343 ;
  assign n41342 = n27891 | n30895 ;
  assign n41345 = n41344 ^ n41342 ^ 1'b0 ;
  assign n41346 = n41345 ^ n29893 ^ n29027 ;
  assign n41347 = n5749 & n14864 ;
  assign n41348 = n18359 & n41347 ;
  assign n41349 = ( ~n1891 & n15760 ) | ( ~n1891 & n41348 ) | ( n15760 & n41348 ) ;
  assign n41350 = ( n24108 & ~n29469 ) | ( n24108 & n41349 ) | ( ~n29469 & n41349 ) ;
  assign n41353 = ( n3932 & n5117 ) | ( n3932 & ~n23606 ) | ( n5117 & ~n23606 ) ;
  assign n41351 = n17721 & ~n19675 ;
  assign n41352 = ~n8976 & n41351 ;
  assign n41354 = n41353 ^ n41352 ^ n36413 ;
  assign n41355 = n3938 | n11202 ;
  assign n41356 = n29027 ^ n17501 ^ n1616 ;
  assign n41357 = n41355 & ~n41356 ;
  assign n41358 = ~n30623 & n41357 ;
  assign n41359 = ~n6798 & n41358 ;
  assign n41360 = ( ~x246 & n41354 ) | ( ~x246 & n41359 ) | ( n41354 & n41359 ) ;
  assign n41361 = ( n18665 & n26099 ) | ( n18665 & n29011 ) | ( n26099 & n29011 ) ;
  assign n41362 = ~n11860 & n26394 ;
  assign n41363 = n41362 ^ n17518 ^ n10800 ;
  assign n41364 = ( n669 & n5910 ) | ( n669 & n8065 ) | ( n5910 & n8065 ) ;
  assign n41365 = n41364 ^ n1846 ^ 1'b0 ;
  assign n41366 = n27725 & n41365 ;
  assign n41367 = n41366 ^ n3371 ^ 1'b0 ;
  assign n41368 = ( n1611 & n11237 ) | ( n1611 & ~n12059 ) | ( n11237 & ~n12059 ) ;
  assign n41369 = n41368 ^ n16522 ^ n15904 ;
  assign n41370 = ( n12588 & ~n27433 ) | ( n12588 & n40960 ) | ( ~n27433 & n40960 ) ;
  assign n41371 = ( n4207 & n26641 ) | ( n4207 & ~n41370 ) | ( n26641 & ~n41370 ) ;
  assign n41372 = n11088 ^ n10563 ^ n6594 ;
  assign n41373 = n41372 ^ n23099 ^ n1968 ;
  assign n41374 = n28595 ^ n5897 ^ n3418 ;
  assign n41375 = n3808 & ~n41374 ;
  assign n41376 = n10132 ^ n9887 ^ 1'b0 ;
  assign n41377 = n24077 | n41376 ;
  assign n41378 = ( n2309 & n41375 ) | ( n2309 & n41377 ) | ( n41375 & n41377 ) ;
  assign n41379 = n30746 & ~n36352 ;
  assign n41380 = n41379 ^ n19009 ^ 1'b0 ;
  assign n41381 = n41380 ^ n1803 ^ n1007 ;
  assign n41382 = n7931 & n33913 ;
  assign n41383 = ~n7255 & n41382 ;
  assign n41384 = ( n2850 & n6891 ) | ( n2850 & ~n12884 ) | ( n6891 & ~n12884 ) ;
  assign n41385 = n41384 ^ n13392 ^ n4491 ;
  assign n41386 = n10515 & ~n41385 ;
  assign n41387 = ( n17422 & ~n35618 ) | ( n17422 & n41386 ) | ( ~n35618 & n41386 ) ;
  assign n41388 = n14818 & n30059 ;
  assign n41389 = ( n743 & n17242 ) | ( n743 & n41388 ) | ( n17242 & n41388 ) ;
  assign n41390 = ( ~n3578 & n12953 ) | ( ~n3578 & n15392 ) | ( n12953 & n15392 ) ;
  assign n41391 = n2395 ^ n1579 ^ 1'b0 ;
  assign n41392 = n31493 ^ n10450 ^ n2450 ;
  assign n41393 = n41392 ^ n34307 ^ n2755 ;
  assign n41394 = ( n28591 & n41391 ) | ( n28591 & ~n41393 ) | ( n41391 & ~n41393 ) ;
  assign n41395 = ( n6007 & ~n41390 ) | ( n6007 & n41394 ) | ( ~n41390 & n41394 ) ;
  assign n41396 = n9722 | n13051 ;
  assign n41397 = n7898 | n41396 ;
  assign n41398 = ( n25340 & n25512 ) | ( n25340 & ~n41397 ) | ( n25512 & ~n41397 ) ;
  assign n41399 = ( n11677 & n22576 ) | ( n11677 & n41398 ) | ( n22576 & n41398 ) ;
  assign n41400 = n28181 ^ n861 ^ 1'b0 ;
  assign n41401 = n35654 ^ n33157 ^ 1'b0 ;
  assign n41402 = n41401 ^ n31739 ^ n29064 ;
  assign n41411 = n39868 ^ n11211 ^ n10887 ;
  assign n41405 = n5964 & n38469 ;
  assign n41406 = n568 & n41405 ;
  assign n41407 = n14165 & ~n41406 ;
  assign n41408 = ~n19095 & n41407 ;
  assign n41403 = n37038 ^ n19596 ^ n16351 ;
  assign n41404 = n41403 ^ n17294 ^ n16154 ;
  assign n41409 = n41408 ^ n41404 ^ n2012 ;
  assign n41410 = n41409 ^ n14586 ^ n1967 ;
  assign n41412 = n41411 ^ n41410 ^ n15110 ;
  assign n41413 = ( n8483 & n41402 ) | ( n8483 & ~n41412 ) | ( n41402 & ~n41412 ) ;
  assign n41414 = n8490 ^ n688 ^ 1'b0 ;
  assign n41415 = n7071 & ~n41414 ;
  assign n41416 = n24013 ^ n11392 ^ 1'b0 ;
  assign n41417 = n36294 & ~n41416 ;
  assign n41418 = n18439 ^ n14329 ^ n1190 ;
  assign n41419 = n41418 ^ n29284 ^ n15834 ;
  assign n41420 = n1828 | n12827 ;
  assign n41421 = n14341 | n41420 ;
  assign n41422 = n41421 ^ n39879 ^ n26870 ;
  assign n41423 = n6898 | n14262 ;
  assign n41424 = ( n1562 & n15198 ) | ( n1562 & ~n41423 ) | ( n15198 & ~n41423 ) ;
  assign n41425 = n41424 ^ n32022 ^ n9216 ;
  assign n41426 = ( n4958 & n25211 ) | ( n4958 & ~n41425 ) | ( n25211 & ~n41425 ) ;
  assign n41427 = n1746 & n6581 ;
  assign n41428 = n41427 ^ n3609 ^ 1'b0 ;
  assign n41429 = n23654 ^ n18027 ^ 1'b0 ;
  assign n41430 = ~n19424 & n41429 ;
  assign n41431 = ~n19687 & n23530 ;
  assign n41432 = ( n21927 & n35350 ) | ( n21927 & ~n41431 ) | ( n35350 & ~n41431 ) ;
  assign n41433 = ( n18886 & n25420 ) | ( n18886 & n40381 ) | ( n25420 & n40381 ) ;
  assign n41434 = ( n607 & n12085 ) | ( n607 & n37603 ) | ( n12085 & n37603 ) ;
  assign n41435 = ( n4866 & n6009 ) | ( n4866 & ~n37025 ) | ( n6009 & ~n37025 ) ;
  assign n41436 = n11656 ^ n3354 ^ n1572 ;
  assign n41437 = ( n1431 & n27807 ) | ( n1431 & n41436 ) | ( n27807 & n41436 ) ;
  assign n41438 = ( n13009 & ~n41435 ) | ( n13009 & n41437 ) | ( ~n41435 & n41437 ) ;
  assign n41443 = ( n666 & ~n3067 ) | ( n666 & n8162 ) | ( ~n3067 & n8162 ) ;
  assign n41444 = ( n3735 & n4753 ) | ( n3735 & ~n18281 ) | ( n4753 & ~n18281 ) ;
  assign n41445 = ( n33962 & ~n37930 ) | ( n33962 & n41444 ) | ( ~n37930 & n41444 ) ;
  assign n41446 = ( n10191 & n41443 ) | ( n10191 & n41445 ) | ( n41443 & n41445 ) ;
  assign n41439 = n33528 ^ n17935 ^ n16148 ;
  assign n41440 = n16196 & ~n29717 ;
  assign n41441 = n41439 & n41440 ;
  assign n41442 = n41441 ^ n13929 ^ n267 ;
  assign n41447 = n41446 ^ n41442 ^ n12848 ;
  assign n41448 = ~n11438 & n38314 ;
  assign n41449 = n33760 ^ n23050 ^ 1'b0 ;
  assign n41450 = ~n17691 & n21995 ;
  assign n41451 = n17181 & n41450 ;
  assign n41452 = n19995 ^ n6105 ^ n1953 ;
  assign n41453 = n13414 & ~n41452 ;
  assign n41454 = n41451 & n41453 ;
  assign n41455 = n33647 ^ n32472 ^ n9890 ;
  assign n41456 = n21663 ^ n13037 ^ 1'b0 ;
  assign n41457 = n763 | n20269 ;
  assign n41458 = n41457 ^ n16327 ^ 1'b0 ;
  assign n41459 = ( ~n4315 & n41456 ) | ( ~n4315 & n41458 ) | ( n41456 & n41458 ) ;
  assign n41460 = n41459 ^ n14594 ^ x2 ;
  assign n41466 = ( n4014 & ~n10274 ) | ( n4014 & n15113 ) | ( ~n10274 & n15113 ) ;
  assign n41464 = ( n4744 & ~n8839 ) | ( n4744 & n14371 ) | ( ~n8839 & n14371 ) ;
  assign n41465 = ( n13281 & n28197 ) | ( n13281 & n41464 ) | ( n28197 & n41464 ) ;
  assign n41461 = n24109 ^ n12019 ^ 1'b0 ;
  assign n41462 = ~n14951 & n41461 ;
  assign n41463 = n41462 ^ n27191 ^ n5064 ;
  assign n41467 = n41466 ^ n41465 ^ n41463 ;
  assign n41468 = ( n6542 & ~n12356 ) | ( n6542 & n20316 ) | ( ~n12356 & n20316 ) ;
  assign n41469 = n41468 ^ n5996 ^ 1'b0 ;
  assign n41470 = n16935 & ~n41469 ;
  assign n41471 = n21661 ^ n17957 ^ n14806 ;
  assign n41472 = ( n11532 & ~n41470 ) | ( n11532 & n41471 ) | ( ~n41470 & n41471 ) ;
  assign n41473 = n22087 ^ n19112 ^ 1'b0 ;
  assign n41474 = ( n18911 & n31956 ) | ( n18911 & n37000 ) | ( n31956 & n37000 ) ;
  assign n41475 = n23984 & n33099 ;
  assign n41476 = n18907 & n41475 ;
  assign n41477 = ( ~n4893 & n8448 ) | ( ~n4893 & n12104 ) | ( n8448 & n12104 ) ;
  assign n41478 = n41477 ^ n5526 ^ 1'b0 ;
  assign n41479 = n39229 ^ n38101 ^ n17624 ;
  assign n41480 = ( n5969 & n23936 ) | ( n5969 & ~n32724 ) | ( n23936 & ~n32724 ) ;
  assign n41485 = n2385 & n20097 ;
  assign n41483 = n29105 ^ n7628 ^ n3263 ;
  assign n41481 = n30639 ^ n21161 ^ 1'b0 ;
  assign n41482 = ( n4474 & ~n14886 ) | ( n4474 & n41481 ) | ( ~n14886 & n41481 ) ;
  assign n41484 = n41483 ^ n41482 ^ n512 ;
  assign n41486 = n41485 ^ n41484 ^ n37244 ;
  assign n41487 = n39023 ^ n12071 ^ n10453 ;
  assign n41488 = n41487 ^ n11029 ^ 1'b0 ;
  assign n41489 = ( n5330 & n15861 ) | ( n5330 & n19256 ) | ( n15861 & n19256 ) ;
  assign n41490 = ( ~n788 & n18347 ) | ( ~n788 & n26046 ) | ( n18347 & n26046 ) ;
  assign n41491 = n26963 | n41490 ;
  assign n41492 = ( n22189 & ~n41489 ) | ( n22189 & n41491 ) | ( ~n41489 & n41491 ) ;
  assign n41493 = n5277 & ~n15618 ;
  assign n41494 = n6988 & n41493 ;
  assign n41495 = ~n29126 & n41494 ;
  assign n41496 = n41495 ^ n15336 ^ n4005 ;
  assign n41497 = n30563 ^ n9482 ^ n1225 ;
  assign n41498 = n41497 ^ n10884 ^ n8656 ;
  assign n41499 = ~n17040 & n41498 ;
  assign n41500 = n21894 | n34294 ;
  assign n41501 = ( n4080 & ~n23991 ) | ( n4080 & n30421 ) | ( ~n23991 & n30421 ) ;
  assign n41502 = n41501 ^ n11147 ^ 1'b0 ;
  assign n41503 = n32697 ^ n26526 ^ 1'b0 ;
  assign n41504 = n39102 ^ n25473 ^ n20814 ;
  assign n41505 = ( n6537 & ~n11004 ) | ( n6537 & n41504 ) | ( ~n11004 & n41504 ) ;
  assign n41506 = n41505 ^ n34060 ^ n20173 ;
  assign n41507 = n17824 & ~n41506 ;
  assign n41508 = n41507 ^ n35844 ^ 1'b0 ;
  assign n41509 = ( ~n989 & n13398 ) | ( ~n989 & n14509 ) | ( n13398 & n14509 ) ;
  assign n41510 = n4554 ^ n295 ^ 1'b0 ;
  assign n41511 = n41509 | n41510 ;
  assign n41512 = n31164 ^ n15968 ^ n2018 ;
  assign n41513 = ( n9176 & n19308 ) | ( n9176 & n41512 ) | ( n19308 & n41512 ) ;
  assign n41514 = n26008 ^ n18736 ^ n11266 ;
  assign n41515 = ( n2034 & ~n10339 ) | ( n2034 & n12515 ) | ( ~n10339 & n12515 ) ;
  assign n41516 = n24952 & ~n41515 ;
  assign n41517 = n5429 & n41516 ;
  assign n41518 = n41517 ^ n5962 ^ 1'b0 ;
  assign n41519 = n41518 ^ n29313 ^ n11797 ;
  assign n41520 = n41519 ^ n9147 ^ n6772 ;
  assign n41521 = ( n2176 & ~n4310 ) | ( n2176 & n6207 ) | ( ~n4310 & n6207 ) ;
  assign n41522 = n23474 ^ n10955 ^ n7163 ;
  assign n41523 = ( n33420 & ~n41521 ) | ( n33420 & n41522 ) | ( ~n41521 & n41522 ) ;
  assign n41525 = ( ~n2633 & n3561 ) | ( ~n2633 & n6118 ) | ( n3561 & n6118 ) ;
  assign n41524 = ( n1218 & n9162 ) | ( n1218 & n24877 ) | ( n9162 & n24877 ) ;
  assign n41526 = n41525 ^ n41524 ^ n3153 ;
  assign n41527 = n10596 & ~n28140 ;
  assign n41528 = n41527 ^ n4849 ^ 1'b0 ;
  assign n41529 = n40080 | n41528 ;
  assign n41530 = n5121 & ~n41529 ;
  assign n41531 = n13529 & ~n19800 ;
  assign n41532 = n41531 ^ n32422 ^ 1'b0 ;
  assign n41533 = ( n2430 & ~n31016 ) | ( n2430 & n41532 ) | ( ~n31016 & n41532 ) ;
  assign n41534 = n27909 ^ n19715 ^ 1'b0 ;
  assign n41535 = n41533 & n41534 ;
  assign n41536 = n28203 ^ n17668 ^ n14050 ;
  assign n41537 = ( n6614 & n34883 ) | ( n6614 & n36505 ) | ( n34883 & n36505 ) ;
  assign n41538 = n14026 ^ n10658 ^ n1531 ;
  assign n41539 = n40509 ^ n34492 ^ 1'b0 ;
  assign n41540 = n8594 | n41539 ;
  assign n41541 = n41538 & ~n41540 ;
  assign n41542 = ( n10692 & ~n38349 ) | ( n10692 & n41541 ) | ( ~n38349 & n41541 ) ;
  assign n41543 = n22576 ^ n17348 ^ n15643 ;
  assign n41544 = n41543 ^ n27443 ^ n6426 ;
  assign n41545 = n41544 ^ n34448 ^ n23762 ;
  assign n41546 = n38067 ^ n22898 ^ 1'b0 ;
  assign n41547 = ~n24435 & n37776 ;
  assign n41548 = ~n18537 & n38880 ;
  assign n41549 = n41548 ^ n15592 ^ 1'b0 ;
  assign n41550 = n8284 | n10266 ;
  assign n41551 = ( n41547 & n41549 ) | ( n41547 & ~n41550 ) | ( n41549 & ~n41550 ) ;
  assign n41552 = n20484 ^ n9195 ^ 1'b0 ;
  assign n41553 = n3251 & ~n41552 ;
  assign n41554 = n41553 ^ n39235 ^ n16901 ;
  assign n41557 = ( n2454 & n19050 ) | ( n2454 & n22025 ) | ( n19050 & n22025 ) ;
  assign n41555 = n7135 & ~n24939 ;
  assign n41556 = n41555 ^ n17735 ^ 1'b0 ;
  assign n41558 = n41557 ^ n41556 ^ n12496 ;
  assign n41559 = n39430 ^ n34678 ^ n16955 ;
  assign n41560 = n41559 ^ n26909 ^ n2677 ;
  assign n41561 = n14669 ^ n1031 ^ 1'b0 ;
  assign n41562 = n13308 & n41561 ;
  assign n41563 = n21546 & n33907 ;
  assign n41564 = n7014 & n41563 ;
  assign n41566 = ( n10706 & n23468 ) | ( n10706 & ~n24877 ) | ( n23468 & ~n24877 ) ;
  assign n41565 = n8601 & n32863 ;
  assign n41567 = n41566 ^ n41565 ^ 1'b0 ;
  assign n41568 = n26638 ^ n7547 ^ 1'b0 ;
  assign n41569 = ~n41567 & n41568 ;
  assign n41570 = ( n16820 & n18120 ) | ( n16820 & n24197 ) | ( n18120 & n24197 ) ;
  assign n41571 = n17612 ^ n9881 ^ n4636 ;
  assign n41572 = ( ~n34186 & n35537 ) | ( ~n34186 & n41571 ) | ( n35537 & n41571 ) ;
  assign n41573 = n6732 ^ n4669 ^ n2925 ;
  assign n41574 = ( n7298 & ~n19953 ) | ( n7298 & n41573 ) | ( ~n19953 & n41573 ) ;
  assign n41575 = n24794 ^ n12490 ^ n8401 ;
  assign n41576 = n25711 ^ n19108 ^ n13388 ;
  assign n41577 = n25830 ^ n7763 ^ n5030 ;
  assign n41578 = ~n41576 & n41577 ;
  assign n41579 = ( n41574 & n41575 ) | ( n41574 & n41578 ) | ( n41575 & n41578 ) ;
  assign n41580 = n31965 ^ n4032 ^ n264 ;
  assign n41581 = ( ~n7966 & n21834 ) | ( ~n7966 & n34431 ) | ( n21834 & n34431 ) ;
  assign n41582 = n9360 & ~n41581 ;
  assign n41590 = ~n3927 & n7544 ;
  assign n41591 = n41590 ^ n11706 ^ 1'b0 ;
  assign n41589 = n24819 ^ n16627 ^ n4699 ;
  assign n41583 = n34674 ^ n20158 ^ 1'b0 ;
  assign n41584 = ( n16734 & n25709 ) | ( n16734 & ~n41583 ) | ( n25709 & ~n41583 ) ;
  assign n41585 = n41584 ^ n22623 ^ 1'b0 ;
  assign n41586 = n29946 & ~n41585 ;
  assign n41587 = n18597 | n26167 ;
  assign n41588 = n41586 | n41587 ;
  assign n41592 = n41591 ^ n41589 ^ n41588 ;
  assign n41593 = n38962 ^ n8516 ^ n776 ;
  assign n41594 = ~n13825 & n41593 ;
  assign n41595 = n11114 & n41594 ;
  assign n41596 = n41595 ^ n20239 ^ n9381 ;
  assign n41597 = n5072 & n11197 ;
  assign n41598 = ~n3242 & n41597 ;
  assign n41599 = ( n2946 & n7110 ) | ( n2946 & n15250 ) | ( n7110 & n15250 ) ;
  assign n41600 = n14498 ^ n9195 ^ 1'b0 ;
  assign n41601 = n41600 ^ n38763 ^ n3830 ;
  assign n41602 = n41601 ^ n29535 ^ n20360 ;
  assign n41603 = ( ~n4906 & n7759 ) | ( ~n4906 & n19431 ) | ( n7759 & n19431 ) ;
  assign n41604 = ( n7878 & ~n35684 ) | ( n7878 & n41603 ) | ( ~n35684 & n41603 ) ;
  assign n41605 = n37847 ^ n12582 ^ n6145 ;
  assign n41606 = n41605 ^ n37859 ^ n10262 ;
  assign n41607 = n32525 ^ n31531 ^ n30391 ;
  assign n41608 = n27823 ^ n24200 ^ n22539 ;
  assign n41609 = n41608 ^ n13431 ^ n12090 ;
  assign n41610 = n24419 ^ n13506 ^ 1'b0 ;
  assign n41612 = n12491 | n36990 ;
  assign n41613 = n41612 ^ n11877 ^ 1'b0 ;
  assign n41611 = n30595 ^ n14414 ^ 1'b0 ;
  assign n41614 = n41613 ^ n41611 ^ n38416 ;
  assign n41615 = n19679 ^ n17244 ^ 1'b0 ;
  assign n41616 = n12768 & n33626 ;
  assign n41617 = n41616 ^ n29048 ^ n4677 ;
  assign n41621 = n10074 ^ n8924 ^ 1'b0 ;
  assign n41620 = n13132 & n29293 ;
  assign n41618 = n27441 | n31283 ;
  assign n41619 = n34726 & ~n41618 ;
  assign n41622 = n41621 ^ n41620 ^ n41619 ;
  assign n41623 = n39692 ^ n12671 ^ n10603 ;
  assign n41624 = n41623 ^ n15949 ^ n6759 ;
  assign n41625 = ( n8016 & n22056 ) | ( n8016 & ~n41624 ) | ( n22056 & ~n41624 ) ;
  assign n41626 = n4433 ^ n1654 ^ 1'b0 ;
  assign n41627 = n1114 | n41626 ;
  assign n41628 = n37430 ^ n26909 ^ n12948 ;
  assign n41629 = ~n8453 & n41628 ;
  assign n41630 = n14880 & n41629 ;
  assign n41631 = ( n3019 & n3878 ) | ( n3019 & n7150 ) | ( n3878 & n7150 ) ;
  assign n41632 = n27788 ^ n25864 ^ n3687 ;
  assign n41633 = ( n1569 & n41631 ) | ( n1569 & ~n41632 ) | ( n41631 & ~n41632 ) ;
  assign n41634 = ( n26396 & n41552 ) | ( n26396 & ~n41633 ) | ( n41552 & ~n41633 ) ;
  assign n41635 = n35634 ^ n35065 ^ n4543 ;
  assign n41636 = ( n4130 & n19147 ) | ( n4130 & n22226 ) | ( n19147 & n22226 ) ;
  assign n41637 = n10147 ^ n9914 ^ n3490 ;
  assign n41638 = n36227 ^ n11903 ^ n8925 ;
  assign n41639 = ( n24384 & ~n41637 ) | ( n24384 & n41638 ) | ( ~n41637 & n41638 ) ;
  assign n41640 = ( n24139 & n29742 ) | ( n24139 & ~n41124 ) | ( n29742 & ~n41124 ) ;
  assign n41641 = n25499 ^ n18765 ^ n4541 ;
  assign n41642 = n6010 ^ n5126 ^ 1'b0 ;
  assign n41643 = n41641 | n41642 ;
  assign n41644 = n28026 ^ n17078 ^ n5080 ;
  assign n41645 = ~n41643 & n41644 ;
  assign n41646 = n41645 ^ n7293 ^ 1'b0 ;
  assign n41647 = n4398 & ~n18841 ;
  assign n41648 = ~n17519 & n41647 ;
  assign n41649 = n5211 & ~n23595 ;
  assign n41650 = n41649 ^ n27019 ^ 1'b0 ;
  assign n41651 = ( ~n1889 & n4836 ) | ( ~n1889 & n7764 ) | ( n4836 & n7764 ) ;
  assign n41652 = ( n3994 & n37592 ) | ( n3994 & ~n41651 ) | ( n37592 & ~n41651 ) ;
  assign n41653 = n36731 ^ n33264 ^ n9067 ;
  assign n41654 = ~n41652 & n41653 ;
  assign n41655 = ( n5479 & n23429 ) | ( n5479 & ~n41654 ) | ( n23429 & ~n41654 ) ;
  assign n41656 = ~n14951 & n38390 ;
  assign n41657 = n41656 ^ n8690 ^ 1'b0 ;
  assign n41658 = n41657 ^ n31092 ^ n20507 ;
  assign n41659 = ( ~n23807 & n31686 ) | ( ~n23807 & n41658 ) | ( n31686 & n41658 ) ;
  assign n41660 = n37666 ^ n23919 ^ n5401 ;
  assign n41661 = n18298 ^ n8020 ^ n7627 ;
  assign n41662 = n20426 | n28223 ;
  assign n41663 = n41661 & ~n41662 ;
  assign n41664 = ~n14674 & n22630 ;
  assign n41665 = ~n27513 & n41664 ;
  assign n41666 = n24141 ^ n9996 ^ 1'b0 ;
  assign n41667 = n22823 ^ n21841 ^ n16578 ;
  assign n41668 = n1283 | n35159 ;
  assign n41669 = ( n9735 & ~n14325 ) | ( n9735 & n21580 ) | ( ~n14325 & n21580 ) ;
  assign n41670 = n41669 ^ n15456 ^ n13685 ;
  assign n41671 = ( n3768 & n13778 ) | ( n3768 & ~n14092 ) | ( n13778 & ~n14092 ) ;
  assign n41676 = ( n1282 & n7253 ) | ( n1282 & ~n11521 ) | ( n7253 & ~n11521 ) ;
  assign n41675 = ( n18835 & ~n22685 ) | ( n18835 & n31016 ) | ( ~n22685 & n31016 ) ;
  assign n41677 = n41676 ^ n41675 ^ n28327 ;
  assign n41678 = ( n10824 & n36557 ) | ( n10824 & ~n41677 ) | ( n36557 & ~n41677 ) ;
  assign n41672 = n40407 ^ n23139 ^ 1'b0 ;
  assign n41673 = n18911 & ~n41672 ;
  assign n41674 = n17348 & n41673 ;
  assign n41679 = n41678 ^ n41674 ^ n7136 ;
  assign n41680 = ( n8267 & n31847 ) | ( n8267 & n40258 ) | ( n31847 & n40258 ) ;
  assign n41681 = n39320 ^ n12239 ^ n11560 ;
  assign n41682 = n26198 & ~n26494 ;
  assign n41683 = n16065 ^ n7025 ^ n6173 ;
  assign n41684 = n41683 ^ n17638 ^ x235 ;
  assign n41685 = n41684 ^ n31165 ^ 1'b0 ;
  assign n41686 = n41685 ^ n14935 ^ n2362 ;
  assign n41687 = n27241 ^ n7670 ^ n1366 ;
  assign n41688 = ( n2307 & ~n5041 ) | ( n2307 & n41687 ) | ( ~n5041 & n41687 ) ;
  assign n41689 = n10342 & n12766 ;
  assign n41690 = n6944 & n41689 ;
  assign n41691 = ( n7178 & n11302 ) | ( n7178 & ~n41690 ) | ( n11302 & ~n41690 ) ;
  assign n41692 = ( n15625 & n30113 ) | ( n15625 & ~n41691 ) | ( n30113 & ~n41691 ) ;
  assign n41695 = n31954 ^ n14048 ^ 1'b0 ;
  assign n41693 = n10308 & n30004 ;
  assign n41694 = n41693 ^ n9563 ^ 1'b0 ;
  assign n41696 = n41695 ^ n41694 ^ n5467 ;
  assign n41697 = n41696 ^ n31692 ^ n23226 ;
  assign n41698 = n11497 & n33949 ;
  assign n41699 = n41698 ^ n6676 ^ 1'b0 ;
  assign n41700 = n18012 & n41699 ;
  assign n41701 = ( ~n16036 & n29011 ) | ( ~n16036 & n41700 ) | ( n29011 & n41700 ) ;
  assign n41702 = n20449 ^ n10258 ^ n8102 ;
  assign n41703 = n20273 & ~n41702 ;
  assign n41704 = n41703 ^ n9060 ^ 1'b0 ;
  assign n41705 = n41704 ^ n22983 ^ n633 ;
  assign n41706 = n20743 ^ n6124 ^ n5512 ;
  assign n41707 = n41706 ^ n22813 ^ n1625 ;
  assign n41708 = n24439 ^ n19409 ^ 1'b0 ;
  assign n41709 = n39666 ^ n20170 ^ 1'b0 ;
  assign n41710 = ~n18033 & n41709 ;
  assign n41711 = ( ~n2704 & n6873 ) | ( ~n2704 & n7231 ) | ( n6873 & n7231 ) ;
  assign n41712 = ( ~n8142 & n16233 ) | ( ~n8142 & n41711 ) | ( n16233 & n41711 ) ;
  assign n41713 = ~n6693 & n29460 ;
  assign n41714 = ~n41712 & n41713 ;
  assign n41715 = n41406 ^ n8685 ^ n785 ;
  assign n41716 = n41715 ^ n17970 ^ n4936 ;
  assign n41717 = n6394 | n18446 ;
  assign n41718 = n41717 ^ n5982 ^ 1'b0 ;
  assign n41719 = n41718 ^ n30278 ^ n21495 ;
  assign n41720 = n26178 ^ n658 ^ 1'b0 ;
  assign n41721 = n41720 ^ n22385 ^ 1'b0 ;
  assign n41722 = n38568 ^ n23645 ^ n6931 ;
  assign n41723 = n23910 ^ n15325 ^ 1'b0 ;
  assign n41724 = ~n8909 & n41723 ;
  assign n41725 = ( ~n8879 & n32744 ) | ( ~n8879 & n41724 ) | ( n32744 & n41724 ) ;
  assign n41726 = n41725 ^ n15924 ^ n4159 ;
  assign n41727 = ( n12988 & ~n17157 ) | ( n12988 & n27161 ) | ( ~n17157 & n27161 ) ;
  assign n41730 = n22671 ^ n21856 ^ n19226 ;
  assign n41728 = n9205 ^ n9012 ^ 1'b0 ;
  assign n41729 = n6491 & n41728 ;
  assign n41731 = n41730 ^ n41729 ^ n16033 ;
  assign n41737 = ( ~n11291 & n13514 ) | ( ~n11291 & n29320 ) | ( n13514 & n29320 ) ;
  assign n41735 = n28408 ^ n16445 ^ n15055 ;
  assign n41733 = n6974 & n9750 ;
  assign n41734 = ~n12329 & n41733 ;
  assign n41736 = n41735 ^ n41734 ^ 1'b0 ;
  assign n41732 = ( ~n2141 & n23801 ) | ( ~n2141 & n31219 ) | ( n23801 & n31219 ) ;
  assign n41738 = n41737 ^ n41736 ^ n41732 ;
  assign n41739 = ( n4841 & n31678 ) | ( n4841 & n38600 ) | ( n31678 & n38600 ) ;
  assign n41740 = n36931 ^ n8705 ^ 1'b0 ;
  assign n41741 = n13398 & ~n41740 ;
  assign n41742 = n1588 | n19613 ;
  assign n41743 = n41742 ^ n38880 ^ 1'b0 ;
  assign n41744 = n36134 ^ n10002 ^ n2460 ;
  assign n41750 = ( ~n23205 & n28408 ) | ( ~n23205 & n29700 ) | ( n28408 & n29700 ) ;
  assign n41746 = n17456 ^ n15607 ^ 1'b0 ;
  assign n41747 = n39825 ^ n6650 ^ 1'b0 ;
  assign n41748 = ( n15843 & n41746 ) | ( n15843 & n41747 ) | ( n41746 & n41747 ) ;
  assign n41745 = n34062 ^ n26474 ^ n1946 ;
  assign n41749 = n41748 ^ n41745 ^ n22537 ;
  assign n41751 = n41750 ^ n41749 ^ n16118 ;
  assign n41752 = ( n3464 & n6024 ) | ( n3464 & n14195 ) | ( n6024 & n14195 ) ;
  assign n41753 = ( n9688 & ~n39904 ) | ( n9688 & n41752 ) | ( ~n39904 & n41752 ) ;
  assign n41754 = n24031 ^ n14572 ^ n4042 ;
  assign n41755 = n39895 & n41754 ;
  assign n41756 = n33639 & n41755 ;
  assign n41757 = n5418 & ~n41756 ;
  assign n41758 = n41757 ^ n32106 ^ 1'b0 ;
  assign n41759 = n2593 & n40316 ;
  assign n41760 = ~n10336 & n41759 ;
  assign n41761 = n5175 & n32110 ;
  assign n41762 = n41761 ^ n12226 ^ 1'b0 ;
  assign n41763 = ( n35568 & n39674 ) | ( n35568 & n41762 ) | ( n39674 & n41762 ) ;
  assign n41764 = n2645 & ~n17635 ;
  assign n41765 = n41764 ^ n6981 ^ 1'b0 ;
  assign n41766 = ( ~n1547 & n29563 ) | ( ~n1547 & n41765 ) | ( n29563 & n41765 ) ;
  assign n41767 = n41766 ^ n23489 ^ n21003 ;
  assign n41768 = n32855 ^ n23929 ^ 1'b0 ;
  assign n41769 = n12471 | n41768 ;
  assign n41770 = ( n4767 & ~n5338 ) | ( n4767 & n41769 ) | ( ~n5338 & n41769 ) ;
  assign n41771 = n24442 ^ n3398 ^ 1'b0 ;
  assign n41772 = ( ~n18957 & n41394 ) | ( ~n18957 & n41771 ) | ( n41394 & n41771 ) ;
  assign n41774 = ( n5358 & n20758 ) | ( n5358 & ~n36425 ) | ( n20758 & ~n36425 ) ;
  assign n41775 = ( ~n1541 & n39016 ) | ( ~n1541 & n41774 ) | ( n39016 & n41774 ) ;
  assign n41773 = ( n4869 & n7024 ) | ( n4869 & ~n19102 ) | ( n7024 & ~n19102 ) ;
  assign n41776 = n41775 ^ n41773 ^ 1'b0 ;
  assign n41777 = ( n1060 & n4803 ) | ( n1060 & n9461 ) | ( n4803 & n9461 ) ;
  assign n41778 = n26689 ^ n9074 ^ n1224 ;
  assign n41779 = ( n475 & n41777 ) | ( n475 & ~n41778 ) | ( n41777 & ~n41778 ) ;
  assign n41780 = ( n24751 & n39846 ) | ( n24751 & n41779 ) | ( n39846 & n41779 ) ;
  assign n41784 = n14570 ^ n12030 ^ 1'b0 ;
  assign n41785 = n1363 & n41784 ;
  assign n41782 = ( ~n5237 & n9020 ) | ( ~n5237 & n14116 ) | ( n9020 & n14116 ) ;
  assign n41783 = ( n29663 & ~n34581 ) | ( n29663 & n41782 ) | ( ~n34581 & n41782 ) ;
  assign n41781 = ( n19198 & ~n24905 ) | ( n19198 & n36399 ) | ( ~n24905 & n36399 ) ;
  assign n41786 = n41785 ^ n41783 ^ n41781 ;
  assign n41787 = n41786 ^ n1179 ^ 1'b0 ;
  assign n41788 = n8955 | n41787 ;
  assign n41789 = ( n8145 & n25714 ) | ( n8145 & ~n35394 ) | ( n25714 & ~n35394 ) ;
  assign n41790 = ( ~n5442 & n25729 ) | ( ~n5442 & n35460 ) | ( n25729 & n35460 ) ;
  assign n41791 = n12044 ^ n10871 ^ 1'b0 ;
  assign n41792 = n41791 ^ n29306 ^ n15117 ;
  assign n41793 = ( n18172 & n41790 ) | ( n18172 & n41792 ) | ( n41790 & n41792 ) ;
  assign n41794 = ( ~n20586 & n23026 ) | ( ~n20586 & n37086 ) | ( n23026 & n37086 ) ;
  assign n41795 = n41794 ^ n31495 ^ n12322 ;
  assign n41796 = n12514 & n39935 ;
  assign n41797 = n41796 ^ n20507 ^ 1'b0 ;
  assign n41798 = n41797 ^ n29392 ^ 1'b0 ;
  assign n41799 = ( n6071 & n12622 ) | ( n6071 & ~n26716 ) | ( n12622 & ~n26716 ) ;
  assign n41800 = n41799 ^ n8171 ^ 1'b0 ;
  assign n41801 = n25661 | n41800 ;
  assign n41802 = n25601 | n36453 ;
  assign n41804 = n24771 ^ n9540 ^ n4647 ;
  assign n41803 = n16196 ^ n15318 ^ n3116 ;
  assign n41805 = n41804 ^ n41803 ^ n8901 ;
  assign n41806 = n35844 ^ n22276 ^ n5127 ;
  assign n41807 = ( n938 & n30628 ) | ( n938 & n41806 ) | ( n30628 & n41806 ) ;
  assign n41808 = ( n9029 & ~n37527 ) | ( n9029 & n41807 ) | ( ~n37527 & n41807 ) ;
  assign n41809 = n41808 ^ n33605 ^ n19036 ;
  assign n41810 = n6563 ^ n5045 ^ n2038 ;
  assign n41811 = ( n5909 & n10936 ) | ( n5909 & ~n41810 ) | ( n10936 & ~n41810 ) ;
  assign n41812 = n41811 ^ n36087 ^ n2873 ;
  assign n41813 = n32715 ^ n31783 ^ n29649 ;
  assign n41814 = n41813 ^ n11358 ^ 1'b0 ;
  assign n41815 = n41814 ^ x153 ^ 1'b0 ;
  assign n41816 = n10457 ^ n4894 ^ 1'b0 ;
  assign n41817 = ( n12634 & n17513 ) | ( n12634 & ~n21759 ) | ( n17513 & ~n21759 ) ;
  assign n41818 = ( n4535 & n10948 ) | ( n4535 & ~n41817 ) | ( n10948 & ~n41817 ) ;
  assign n41819 = n41818 ^ n26752 ^ n13479 ;
  assign n41820 = ~n34618 & n34867 ;
  assign n41821 = n41820 ^ n13412 ^ 1'b0 ;
  assign n41822 = n36561 ^ n5700 ^ 1'b0 ;
  assign n41823 = n19795 & n41822 ;
  assign n41824 = ~n899 & n8267 ;
  assign n41825 = n41824 ^ n30607 ^ n7004 ;
  assign n41826 = ( n15316 & n16982 ) | ( n15316 & ~n41825 ) | ( n16982 & ~n41825 ) ;
  assign n41827 = n28861 ^ n24547 ^ n5291 ;
  assign n41828 = ( ~n5233 & n18930 ) | ( ~n5233 & n24207 ) | ( n18930 & n24207 ) ;
  assign n41829 = n12002 ^ n10517 ^ n4698 ;
  assign n41830 = n38624 ^ n27834 ^ n4130 ;
  assign n41831 = n41830 ^ n41278 ^ n24183 ;
  assign n41832 = n10971 | n17075 ;
  assign n41833 = ( n11229 & ~n20884 ) | ( n11229 & n41832 ) | ( ~n20884 & n41832 ) ;
  assign n41834 = n13057 ^ n10326 ^ n2316 ;
  assign n41835 = n41834 ^ n1851 ^ 1'b0 ;
  assign n41836 = ( n12353 & n32004 ) | ( n12353 & ~n41835 ) | ( n32004 & ~n41835 ) ;
  assign n41842 = ( n5689 & n16863 ) | ( n5689 & ~n35831 ) | ( n16863 & ~n35831 ) ;
  assign n41843 = n17478 | n41842 ;
  assign n41837 = n11877 ^ n5834 ^ n362 ;
  assign n41838 = ( n2101 & n5777 ) | ( n2101 & ~n14707 ) | ( n5777 & ~n14707 ) ;
  assign n41839 = n41837 & ~n41838 ;
  assign n41840 = ( ~n13101 & n13496 ) | ( ~n13101 & n41839 ) | ( n13496 & n41839 ) ;
  assign n41841 = n41840 ^ n36557 ^ n8504 ;
  assign n41844 = n41843 ^ n41841 ^ n19043 ;
  assign n41845 = ( ~n2726 & n8910 ) | ( ~n2726 & n31129 ) | ( n8910 & n31129 ) ;
  assign n41846 = n41845 ^ n15940 ^ n2250 ;
  assign n41847 = ( n3359 & n5963 ) | ( n3359 & n15095 ) | ( n5963 & n15095 ) ;
  assign n41848 = n6592 | n24258 ;
  assign n41849 = n41848 ^ n12881 ^ 1'b0 ;
  assign n41850 = ( x8 & n3823 ) | ( x8 & ~n41849 ) | ( n3823 & ~n41849 ) ;
  assign n41851 = ( n1500 & n10023 ) | ( n1500 & ~n12271 ) | ( n10023 & ~n12271 ) ;
  assign n41852 = ( ~n3843 & n31232 ) | ( ~n3843 & n41851 ) | ( n31232 & n41851 ) ;
  assign n41853 = n12810 ^ n1956 ^ 1'b0 ;
  assign n41854 = n41852 & ~n41853 ;
  assign n41855 = n1170 & n32303 ;
  assign n41856 = n12876 & n41855 ;
  assign n41857 = n471 | n41856 ;
  assign n41858 = n7341 & ~n29222 ;
  assign n41859 = n41858 ^ n27343 ^ 1'b0 ;
  assign n41860 = n41859 ^ n38880 ^ 1'b0 ;
  assign n41862 = n1367 | n3503 ;
  assign n41863 = n23430 | n41862 ;
  assign n41861 = ( n17016 & n33887 ) | ( n17016 & n36767 ) | ( n33887 & n36767 ) ;
  assign n41864 = n41863 ^ n41861 ^ n23940 ;
  assign n41865 = ( n14337 & ~n19337 ) | ( n14337 & n41864 ) | ( ~n19337 & n41864 ) ;
  assign n41866 = n30459 ^ n17563 ^ n10226 ;
  assign n41867 = n19652 ^ n7447 ^ n2096 ;
  assign n41868 = ( ~n19857 & n31125 ) | ( ~n19857 & n41867 ) | ( n31125 & n41867 ) ;
  assign n41870 = n4632 & ~n10556 ;
  assign n41871 = ( n14972 & n35810 ) | ( n14972 & n41870 ) | ( n35810 & n41870 ) ;
  assign n41869 = n4012 & n29558 ;
  assign n41872 = n41871 ^ n41869 ^ 1'b0 ;
  assign n41873 = n26070 ^ n24955 ^ 1'b0 ;
  assign n41874 = ~n5536 & n9192 ;
  assign n41875 = ( ~n3383 & n23682 ) | ( ~n3383 & n41874 ) | ( n23682 & n41874 ) ;
  assign n41876 = n41875 ^ n35146 ^ n767 ;
  assign n41882 = ( ~n5584 & n23663 ) | ( ~n5584 & n28920 ) | ( n23663 & n28920 ) ;
  assign n41883 = ( n18423 & n37027 ) | ( n18423 & ~n41882 ) | ( n37027 & ~n41882 ) ;
  assign n41884 = n41883 ^ n25783 ^ n13151 ;
  assign n41877 = n31201 ^ n12269 ^ 1'b0 ;
  assign n41878 = ~n14459 & n41877 ;
  assign n41879 = n12508 | n15232 ;
  assign n41880 = n41879 ^ n8594 ^ 1'b0 ;
  assign n41881 = n41878 & ~n41880 ;
  assign n41885 = n41884 ^ n41881 ^ n4155 ;
  assign n41886 = n19393 ^ n6294 ^ 1'b0 ;
  assign n41887 = n26993 & n41886 ;
  assign n41888 = n41887 ^ n4256 ^ 1'b0 ;
  assign n41889 = ( n11987 & ~n37859 ) | ( n11987 & n41888 ) | ( ~n37859 & n41888 ) ;
  assign n41890 = n22540 ^ n19691 ^ n9352 ;
  assign n41891 = ( n13820 & n38614 ) | ( n13820 & ~n41890 ) | ( n38614 & ~n41890 ) ;
  assign n41892 = n13778 ^ n8091 ^ n1996 ;
  assign n41893 = ( n4806 & n28694 ) | ( n4806 & ~n41892 ) | ( n28694 & ~n41892 ) ;
  assign n41894 = n10965 | n15042 ;
  assign n41895 = n41894 ^ n37225 ^ 1'b0 ;
  assign n41896 = ( ~n5421 & n9000 ) | ( ~n5421 & n39902 ) | ( n9000 & n39902 ) ;
  assign n41897 = n13000 & n28184 ;
  assign n41898 = ~n41896 & n41897 ;
  assign n41899 = n23647 | n41898 ;
  assign n41900 = n41899 ^ n34194 ^ 1'b0 ;
  assign n41901 = n3315 ^ n1564 ^ 1'b0 ;
  assign n41902 = ~n4431 & n41901 ;
  assign n41903 = n19593 & n41902 ;
  assign n41904 = n10073 | n41903 ;
  assign n41908 = ~n18903 & n33662 ;
  assign n41909 = ~n20205 & n41908 ;
  assign n41905 = n18250 ^ n2560 ^ 1'b0 ;
  assign n41906 = n9642 & n41905 ;
  assign n41907 = n41906 ^ n28918 ^ n20865 ;
  assign n41910 = n41909 ^ n41907 ^ n39501 ;
  assign n41911 = ( n11098 & n25745 ) | ( n11098 & ~n29410 ) | ( n25745 & ~n29410 ) ;
  assign n41912 = n11504 & n35592 ;
  assign n41913 = ( n11539 & n37357 ) | ( n11539 & n41912 ) | ( n37357 & n41912 ) ;
  assign n41914 = n41913 ^ n29729 ^ 1'b0 ;
  assign n41915 = ( n10330 & n41911 ) | ( n10330 & ~n41914 ) | ( n41911 & ~n41914 ) ;
  assign n41916 = ( n6847 & n22590 ) | ( n6847 & n36703 ) | ( n22590 & n36703 ) ;
  assign n41917 = ( ~n1782 & n24024 ) | ( ~n1782 & n28341 ) | ( n24024 & n28341 ) ;
  assign n41918 = ( n21373 & n23098 ) | ( n21373 & n41917 ) | ( n23098 & n41917 ) ;
  assign n41919 = ~n10866 & n40314 ;
  assign n41920 = n20833 & n41919 ;
  assign n41921 = n36813 ^ n22253 ^ 1'b0 ;
  assign n41922 = ~n41920 & n41921 ;
  assign n41923 = n29722 ^ n1959 ^ 1'b0 ;
  assign n41924 = ~n3689 & n41923 ;
  assign n41925 = n7125 ^ n4718 ^ 1'b0 ;
  assign n41926 = ~n16905 & n41925 ;
  assign n41927 = ( n5491 & n18720 ) | ( n5491 & ~n22274 ) | ( n18720 & ~n22274 ) ;
  assign n41928 = ( n16488 & ~n41926 ) | ( n16488 & n41927 ) | ( ~n41926 & n41927 ) ;
  assign n41929 = n23544 ^ n16401 ^ 1'b0 ;
  assign n41930 = n10878 | n41929 ;
  assign n41931 = n20940 & ~n41930 ;
  assign n41933 = ( n2797 & n5860 ) | ( n2797 & ~n10485 ) | ( n5860 & ~n10485 ) ;
  assign n41932 = n36557 ^ n30239 ^ n24696 ;
  assign n41934 = n41933 ^ n41932 ^ n2931 ;
  assign n41935 = n19901 ^ n11840 ^ 1'b0 ;
  assign n41936 = n41935 ^ n17182 ^ n4889 ;
  assign n41937 = ( n1695 & n3642 ) | ( n1695 & ~n24739 ) | ( n3642 & ~n24739 ) ;
  assign n41938 = ( n7396 & n33166 ) | ( n7396 & n41937 ) | ( n33166 & n41937 ) ;
  assign n41939 = n41938 ^ n41917 ^ n29234 ;
  assign n41940 = n961 & ~n17233 ;
  assign n41941 = ( n1184 & n16735 ) | ( n1184 & n41940 ) | ( n16735 & n41940 ) ;
  assign n41942 = n32700 ^ n19185 ^ n10999 ;
  assign n41943 = n41942 ^ n9225 ^ 1'b0 ;
  assign n41944 = ~n41941 & n41943 ;
  assign n41945 = n15760 ^ n8453 ^ n2383 ;
  assign n41946 = n11899 ^ n4455 ^ n867 ;
  assign n41947 = n41946 ^ n22328 ^ n16998 ;
  assign n41948 = n41947 ^ n20860 ^ n3608 ;
  assign n41949 = n41948 ^ n3622 ^ 1'b0 ;
  assign n41950 = ~n41945 & n41949 ;
  assign n41951 = n22510 ^ n15631 ^ n13532 ;
  assign n41952 = n7591 & ~n41951 ;
  assign n41953 = n1159 & n20981 ;
  assign n41954 = ~n33198 & n41953 ;
  assign n41955 = n19776 ^ n19148 ^ n2292 ;
  assign n41956 = n7567 | n13737 ;
  assign n41957 = n41955 | n41956 ;
  assign n41958 = ( ~n19843 & n41954 ) | ( ~n19843 & n41957 ) | ( n41954 & n41957 ) ;
  assign n41959 = ( n19327 & n24497 ) | ( n19327 & ~n39665 ) | ( n24497 & ~n39665 ) ;
  assign n41960 = ( n8773 & n32842 ) | ( n8773 & n36041 ) | ( n32842 & n36041 ) ;
  assign n41961 = ( n2782 & ~n11820 ) | ( n2782 & n41960 ) | ( ~n11820 & n41960 ) ;
  assign n41962 = n32195 ^ n28394 ^ n16048 ;
  assign n41963 = n34951 ^ n4675 ^ n1504 ;
  assign n41964 = n9230 ^ n8856 ^ 1'b0 ;
  assign n41965 = n23784 ^ n9583 ^ 1'b0 ;
  assign n41966 = n6018 & ~n35831 ;
  assign n41967 = n4988 | n13658 ;
  assign n41968 = ( x199 & ~n3672 ) | ( x199 & n41967 ) | ( ~n3672 & n41967 ) ;
  assign n41969 = n38036 ^ n1335 ^ 1'b0 ;
  assign n41970 = n2528 & n41969 ;
  assign n41971 = n41970 ^ n28616 ^ n20723 ;
  assign n41972 = ( ~n1866 & n10908 ) | ( ~n1866 & n30169 ) | ( n10908 & n30169 ) ;
  assign n41973 = n1470 & ~n21420 ;
  assign n41974 = n41973 ^ n12847 ^ 1'b0 ;
  assign n41975 = n15749 ^ n13538 ^ n11518 ;
  assign n41976 = n28523 & n41975 ;
  assign n41977 = n39824 & n41976 ;
  assign n41978 = n30521 ^ n16269 ^ n7673 ;
  assign n41979 = n41978 ^ n31575 ^ n1200 ;
  assign n41980 = ( n18646 & n36884 ) | ( n18646 & ~n38636 ) | ( n36884 & ~n38636 ) ;
  assign n41981 = n32206 ^ n16920 ^ n6509 ;
  assign n41982 = n10954 & ~n22466 ;
  assign n41983 = ( n15275 & ~n26901 ) | ( n15275 & n41982 ) | ( ~n26901 & n41982 ) ;
  assign n41984 = n15093 ^ n12741 ^ n8014 ;
  assign n41987 = n9048 ^ n7210 ^ n4640 ;
  assign n41985 = n5247 & n15260 ;
  assign n41986 = ~n6787 & n41985 ;
  assign n41988 = n41987 ^ n41986 ^ 1'b0 ;
  assign n41989 = n1104 & n15666 ;
  assign n41990 = ~n18283 & n41989 ;
  assign n41991 = ( n6593 & ~n11657 ) | ( n6593 & n41990 ) | ( ~n11657 & n41990 ) ;
  assign n41992 = ( n10301 & n23551 ) | ( n10301 & n30890 ) | ( n23551 & n30890 ) ;
  assign n41993 = n41992 ^ n18848 ^ n12141 ;
  assign n41994 = ( ~n14172 & n35460 ) | ( ~n14172 & n41993 ) | ( n35460 & n41993 ) ;
  assign n41995 = ( ~n3054 & n6200 ) | ( ~n3054 & n31313 ) | ( n6200 & n31313 ) ;
  assign n41996 = ( n16599 & ~n29575 ) | ( n16599 & n41995 ) | ( ~n29575 & n41995 ) ;
  assign n41997 = n2319 | n41996 ;
  assign n41998 = n5565 & ~n41997 ;
  assign n41999 = n6598 | n28166 ;
  assign n42000 = ( n22038 & ~n30911 ) | ( n22038 & n32312 ) | ( ~n30911 & n32312 ) ;
  assign n42001 = n42000 ^ n16881 ^ 1'b0 ;
  assign n42002 = ( n1371 & n4825 ) | ( n1371 & ~n25282 ) | ( n4825 & ~n25282 ) ;
  assign n42003 = n17251 ^ n8337 ^ 1'b0 ;
  assign n42004 = ( n29089 & n42002 ) | ( n29089 & n42003 ) | ( n42002 & n42003 ) ;
  assign n42005 = ( n3236 & ~n35672 ) | ( n3236 & n42004 ) | ( ~n35672 & n42004 ) ;
  assign n42006 = n28745 | n31871 ;
  assign n42007 = n455 | n29949 ;
  assign n42008 = n42007 ^ n3612 ^ 1'b0 ;
  assign n42009 = n42008 ^ n33825 ^ n7923 ;
  assign n42010 = n42009 ^ n40464 ^ n30654 ;
  assign n42011 = n22323 ^ n19581 ^ n4057 ;
  assign n42012 = n42011 ^ n18271 ^ n6870 ;
  assign n42013 = n30178 ^ n27939 ^ 1'b0 ;
  assign n42014 = ( n1493 & n23033 ) | ( n1493 & n42013 ) | ( n23033 & n42013 ) ;
  assign n42015 = n31452 ^ n3279 ^ 1'b0 ;
  assign n42016 = n20193 & ~n42015 ;
  assign n42017 = ~n6973 & n31547 ;
  assign n42018 = ~n19110 & n42017 ;
  assign n42019 = n41060 ^ n17802 ^ 1'b0 ;
  assign n42020 = ~n2921 & n42019 ;
  assign n42021 = ( n2897 & ~n16507 ) | ( n2897 & n35795 ) | ( ~n16507 & n35795 ) ;
  assign n42022 = n18071 ^ n13045 ^ n2342 ;
  assign n42023 = n20850 ^ n4529 ^ n1655 ;
  assign n42024 = n42023 ^ n20547 ^ n1425 ;
  assign n42025 = n42024 ^ n13334 ^ n2942 ;
  assign n42029 = n538 & ~n10726 ;
  assign n42026 = ( n9418 & ~n34472 ) | ( n9418 & n36327 ) | ( ~n34472 & n36327 ) ;
  assign n42027 = n42026 ^ n24922 ^ n3453 ;
  assign n42028 = ( n949 & ~n20385 ) | ( n949 & n42027 ) | ( ~n20385 & n42027 ) ;
  assign n42030 = n42029 ^ n42028 ^ 1'b0 ;
  assign n42031 = n31463 ^ n11685 ^ 1'b0 ;
  assign n42032 = ~n30877 & n42031 ;
  assign n42033 = n2343 & n42032 ;
  assign n42034 = n28510 & n42033 ;
  assign n42035 = n11962 ^ n6637 ^ n390 ;
  assign n42036 = n42035 ^ n22166 ^ 1'b0 ;
  assign n42037 = n12787 | n25747 ;
  assign n42038 = ( ~n874 & n6749 ) | ( ~n874 & n17536 ) | ( n6749 & n17536 ) ;
  assign n42041 = ( ~n8865 & n9149 ) | ( ~n8865 & n30877 ) | ( n9149 & n30877 ) ;
  assign n42039 = n22573 & ~n30779 ;
  assign n42040 = ~n4804 & n42039 ;
  assign n42042 = n42041 ^ n42040 ^ x69 ;
  assign n42043 = ( n2585 & n5107 ) | ( n2585 & ~n34923 ) | ( n5107 & ~n34923 ) ;
  assign n42044 = n42043 ^ n38245 ^ n16894 ;
  assign n42045 = ( ~n7176 & n23996 ) | ( ~n7176 & n25161 ) | ( n23996 & n25161 ) ;
  assign n42046 = n17873 | n21636 ;
  assign n42047 = ~n15475 & n39841 ;
  assign n42048 = n42047 ^ n12349 ^ 1'b0 ;
  assign n42049 = n23348 ^ n10005 ^ n9013 ;
  assign n42050 = n18620 & ~n42049 ;
  assign n42051 = n42050 ^ n31291 ^ 1'b0 ;
  assign n42052 = n19188 ^ n11070 ^ 1'b0 ;
  assign n42053 = n15864 & ~n42052 ;
  assign n42054 = ( n2051 & n34294 ) | ( n2051 & n42053 ) | ( n34294 & n42053 ) ;
  assign n42055 = ( n446 & ~n23996 ) | ( n446 & n42054 ) | ( ~n23996 & n42054 ) ;
  assign n42056 = n42055 ^ n40962 ^ 1'b0 ;
  assign n42057 = n42056 ^ n39467 ^ n3738 ;
  assign n42058 = ( n7024 & n7351 ) | ( n7024 & n19114 ) | ( n7351 & n19114 ) ;
  assign n42059 = ( ~n3343 & n26025 ) | ( ~n3343 & n38238 ) | ( n26025 & n38238 ) ;
  assign n42060 = n40862 | n42059 ;
  assign n42061 = n8637 | n42060 ;
  assign n42062 = ( ~n12655 & n42058 ) | ( ~n12655 & n42061 ) | ( n42058 & n42061 ) ;
  assign n42063 = n34505 ^ n6541 ^ 1'b0 ;
  assign n42064 = n22300 & n42063 ;
  assign n42065 = ( n33049 & n33348 ) | ( n33049 & n42064 ) | ( n33348 & n42064 ) ;
  assign n42066 = n16509 ^ n11387 ^ n4404 ;
  assign n42067 = n28712 ^ n20385 ^ n5730 ;
  assign n42068 = n42067 ^ n5531 ^ 1'b0 ;
  assign n42069 = n1959 & n31139 ;
  assign n42070 = n42069 ^ n14730 ^ 1'b0 ;
  assign n42071 = n12658 & n27502 ;
  assign n42072 = n42070 & n42071 ;
  assign n42078 = n34625 ^ n18544 ^ 1'b0 ;
  assign n42075 = n35338 ^ n33338 ^ n6778 ;
  assign n42073 = n6397 & ~n7277 ;
  assign n42074 = n42073 ^ n36970 ^ 1'b0 ;
  assign n42076 = n42075 ^ n42074 ^ 1'b0 ;
  assign n42077 = ~n21234 & n42076 ;
  assign n42079 = n42078 ^ n42077 ^ 1'b0 ;
  assign n42080 = n9569 & n14328 ;
  assign n42081 = ( n14170 & n20493 ) | ( n14170 & ~n42080 ) | ( n20493 & ~n42080 ) ;
  assign n42082 = ( n10973 & n21979 ) | ( n10973 & n42081 ) | ( n21979 & n42081 ) ;
  assign n42083 = n27733 ^ n27267 ^ n20677 ;
  assign n42084 = n42083 ^ n17993 ^ n8010 ;
  assign n42085 = n5978 & n14746 ;
  assign n42086 = n36307 ^ n28694 ^ 1'b0 ;
  assign n42087 = ~n42085 & n42086 ;
  assign n42088 = n42087 ^ n20362 ^ 1'b0 ;
  assign n42089 = ( n31742 & n35066 ) | ( n31742 & n37938 ) | ( n35066 & n37938 ) ;
  assign n42093 = ( n353 & n10451 ) | ( n353 & ~n41810 ) | ( n10451 & ~n41810 ) ;
  assign n42091 = ( n3427 & ~n16757 ) | ( n3427 & n21444 ) | ( ~n16757 & n21444 ) ;
  assign n42092 = n42091 ^ n11881 ^ 1'b0 ;
  assign n42090 = n27573 ^ n21044 ^ n6546 ;
  assign n42094 = n42093 ^ n42092 ^ n42090 ;
  assign n42095 = ( n4803 & ~n15725 ) | ( n4803 & n19832 ) | ( ~n15725 & n19832 ) ;
  assign n42096 = ( n7994 & n13577 ) | ( n7994 & n42095 ) | ( n13577 & n42095 ) ;
  assign n42097 = n41079 & n42096 ;
  assign n42098 = n42097 ^ n24825 ^ 1'b0 ;
  assign n42099 = n2505 ^ n2042 ^ 1'b0 ;
  assign n42100 = ~n36417 & n42099 ;
  assign n42101 = n31170 ^ n30722 ^ n2402 ;
  assign n42102 = n31081 ^ n10760 ^ 1'b0 ;
  assign n42103 = ( n788 & n18084 ) | ( n788 & ~n18730 ) | ( n18084 & ~n18730 ) ;
  assign n42104 = n16828 | n42103 ;
  assign n42105 = ( n12648 & ~n20629 ) | ( n12648 & n31236 ) | ( ~n20629 & n31236 ) ;
  assign n42106 = ( n2535 & ~n2857 ) | ( n2535 & n20086 ) | ( ~n2857 & n20086 ) ;
  assign n42107 = n22616 ^ n3185 ^ n1318 ;
  assign n42108 = ( ~n8858 & n42106 ) | ( ~n8858 & n42107 ) | ( n42106 & n42107 ) ;
  assign n42109 = n4196 & n37592 ;
  assign n42110 = n4873 & n42109 ;
  assign n42111 = n21071 ^ n2654 ^ 1'b0 ;
  assign n42112 = ( ~n13662 & n42110 ) | ( ~n13662 & n42111 ) | ( n42110 & n42111 ) ;
  assign n42115 = ( n5526 & n10515 ) | ( n5526 & n10721 ) | ( n10515 & n10721 ) ;
  assign n42113 = n38527 ^ n35688 ^ n19557 ;
  assign n42114 = n42113 ^ n7044 ^ n3021 ;
  assign n42116 = n42115 ^ n42114 ^ n19000 ;
  assign n42117 = n13436 & ~n36266 ;
  assign n42118 = n42117 ^ n20100 ^ 1'b0 ;
  assign n42119 = n19689 ^ n14798 ^ n11383 ;
  assign n42120 = n42119 ^ x211 ^ 1'b0 ;
  assign n42121 = ~n23481 & n42120 ;
  assign n42122 = n38316 ^ n20491 ^ n4808 ;
  assign n42123 = ( n6065 & n9817 ) | ( n6065 & ~n21252 ) | ( n9817 & ~n21252 ) ;
  assign n42124 = n26121 & ~n42123 ;
  assign n42125 = ~n42122 & n42124 ;
  assign n42126 = n3732 & ~n42125 ;
  assign n42127 = n13498 & n42126 ;
  assign n42128 = n10970 & ~n12333 ;
  assign n42129 = ~n11441 & n42128 ;
  assign n42130 = ( n2331 & n19014 ) | ( n2331 & ~n26942 ) | ( n19014 & ~n26942 ) ;
  assign n42131 = ( n3946 & n42129 ) | ( n3946 & ~n42130 ) | ( n42129 & ~n42130 ) ;
  assign n42132 = n32158 ^ n8922 ^ n7398 ;
  assign n42133 = ( ~x61 & n35603 ) | ( ~x61 & n42132 ) | ( n35603 & n42132 ) ;
  assign n42134 = n33336 ^ n6720 ^ x220 ;
  assign n42135 = n3629 | n42134 ;
  assign n42136 = n42135 ^ n26638 ^ 1'b0 ;
  assign n42137 = n42136 ^ n34566 ^ n3181 ;
  assign n42138 = ( n10424 & n14618 ) | ( n10424 & n35857 ) | ( n14618 & n35857 ) ;
  assign n42139 = ( n2415 & ~n2662 ) | ( n2415 & n18262 ) | ( ~n2662 & n18262 ) ;
  assign n42140 = ( ~n21925 & n28213 ) | ( ~n21925 & n42139 ) | ( n28213 & n42139 ) ;
  assign n42141 = n20583 & ~n42140 ;
  assign n42142 = n42141 ^ n2165 ^ 1'b0 ;
  assign n42143 = n38132 ^ n37803 ^ n22600 ;
  assign n42144 = n37772 ^ n16926 ^ n10743 ;
  assign n42145 = n42144 ^ n40325 ^ n15841 ;
  assign n42146 = n11523 & ~n14770 ;
  assign n42147 = n42146 ^ n4121 ^ 1'b0 ;
  assign n42148 = n40879 ^ n13744 ^ n928 ;
  assign n42149 = ( n2625 & n42147 ) | ( n2625 & ~n42148 ) | ( n42147 & ~n42148 ) ;
  assign n42150 = ( n11597 & n14145 ) | ( n11597 & ~n23498 ) | ( n14145 & ~n23498 ) ;
  assign n42151 = n1120 & n2030 ;
  assign n42152 = ~n42150 & n42151 ;
  assign n42153 = n33858 ^ n13681 ^ n5021 ;
  assign n42154 = n31121 ^ n31054 ^ 1'b0 ;
  assign n42155 = ~n3297 & n42154 ;
  assign n42156 = ~n42153 & n42155 ;
  assign n42159 = ( ~n9346 & n26303 ) | ( ~n9346 & n28236 ) | ( n26303 & n28236 ) ;
  assign n42157 = ( n3357 & n9413 ) | ( n3357 & n35881 ) | ( n9413 & n35881 ) ;
  assign n42158 = n42157 ^ n15755 ^ 1'b0 ;
  assign n42160 = n42159 ^ n42158 ^ n23702 ;
  assign n42161 = n42160 ^ n41803 ^ n13607 ;
  assign n42164 = n25654 ^ n11151 ^ 1'b0 ;
  assign n42162 = ( n6975 & ~n20660 ) | ( n6975 & n41406 ) | ( ~n20660 & n41406 ) ;
  assign n42163 = n42162 ^ n39193 ^ n21552 ;
  assign n42165 = n42164 ^ n42163 ^ n5920 ;
  assign n42166 = ( n10597 & n15642 ) | ( n10597 & n42165 ) | ( n15642 & n42165 ) ;
  assign n42167 = ( n5739 & ~n7485 ) | ( n5739 & n20158 ) | ( ~n7485 & n20158 ) ;
  assign n42168 = n21654 ^ n16862 ^ n6231 ;
  assign n42169 = n42168 ^ n27343 ^ n14588 ;
  assign n42170 = ( n9840 & ~n20013 ) | ( n9840 & n27950 ) | ( ~n20013 & n27950 ) ;
  assign n42171 = n25704 & n27793 ;
  assign n42172 = ( n42169 & n42170 ) | ( n42169 & n42171 ) | ( n42170 & n42171 ) ;
  assign n42173 = ( n953 & n1064 ) | ( n953 & ~n2993 ) | ( n1064 & ~n2993 ) ;
  assign n42174 = ( n25515 & n36611 ) | ( n25515 & ~n42173 ) | ( n36611 & ~n42173 ) ;
  assign n42175 = ( n2491 & n3899 ) | ( n2491 & n34511 ) | ( n3899 & n34511 ) ;
  assign n42176 = ( n8657 & n41204 ) | ( n8657 & ~n42175 ) | ( n41204 & ~n42175 ) ;
  assign n42177 = ( n40824 & n42174 ) | ( n40824 & ~n42176 ) | ( n42174 & ~n42176 ) ;
  assign n42178 = n8765 & ~n10729 ;
  assign n42179 = n42178 ^ n4188 ^ 1'b0 ;
  assign n42180 = n20833 ^ n3536 ^ 1'b0 ;
  assign n42181 = n14231 & ~n42180 ;
  assign n42182 = n4652 & n42181 ;
  assign n42183 = n21765 & n42182 ;
  assign n42184 = n20752 ^ n13969 ^ n13388 ;
  assign n42185 = ( x61 & ~n2876 ) | ( x61 & n22642 ) | ( ~n2876 & n22642 ) ;
  assign n42186 = n19844 & ~n28428 ;
  assign n42187 = n42186 ^ n36900 ^ 1'b0 ;
  assign n42188 = ( ~n25646 & n42185 ) | ( ~n25646 & n42187 ) | ( n42185 & n42187 ) ;
  assign n42189 = ( n14104 & n29136 ) | ( n14104 & ~n42188 ) | ( n29136 & ~n42188 ) ;
  assign n42193 = n15847 ^ n2447 ^ n1651 ;
  assign n42192 = n33775 ^ n8071 ^ 1'b0 ;
  assign n42190 = x159 & ~n7426 ;
  assign n42191 = n42190 ^ n22035 ^ 1'b0 ;
  assign n42194 = n42193 ^ n42192 ^ n42191 ;
  assign n42195 = n31484 ^ n26391 ^ x130 ;
  assign n42196 = n42195 ^ n41811 ^ n29536 ;
  assign n42197 = n5980 ^ n5906 ^ n2402 ;
  assign n42198 = n42197 ^ n25041 ^ 1'b0 ;
  assign n42199 = n42196 | n42198 ;
  assign n42201 = ~n7359 & n28827 ;
  assign n42202 = n42201 ^ n1175 ^ 1'b0 ;
  assign n42200 = ( ~n6935 & n6993 ) | ( ~n6935 & n12386 ) | ( n6993 & n12386 ) ;
  assign n42203 = n42202 ^ n42200 ^ 1'b0 ;
  assign n42204 = n12375 & ~n42203 ;
  assign n42205 = ( n4207 & n6721 ) | ( n4207 & n7746 ) | ( n6721 & n7746 ) ;
  assign n42206 = ( n16194 & n21067 ) | ( n16194 & ~n33460 ) | ( n21067 & ~n33460 ) ;
  assign n42207 = ( ~n12349 & n42205 ) | ( ~n12349 & n42206 ) | ( n42205 & n42206 ) ;
  assign n42208 = ( n22561 & ~n31496 ) | ( n22561 & n42207 ) | ( ~n31496 & n42207 ) ;
  assign n42209 = n19797 ^ n10722 ^ 1'b0 ;
  assign n42210 = n12873 & n21254 ;
  assign n42211 = n42209 & n42210 ;
  assign n42212 = n3060 | n42211 ;
  assign n42213 = ( n2521 & n37628 ) | ( n2521 & n38179 ) | ( n37628 & n38179 ) ;
  assign n42214 = ( n5493 & n9068 ) | ( n5493 & n27925 ) | ( n9068 & n27925 ) ;
  assign n42215 = n27393 ^ n8442 ^ n4746 ;
  assign n42216 = n42215 ^ n10250 ^ 1'b0 ;
  assign n42217 = ( n10803 & n42214 ) | ( n10803 & ~n42216 ) | ( n42214 & ~n42216 ) ;
  assign n42218 = ( ~n7426 & n10270 ) | ( ~n7426 & n27727 ) | ( n10270 & n27727 ) ;
  assign n42219 = ( n1425 & ~n21312 ) | ( n1425 & n42218 ) | ( ~n21312 & n42218 ) ;
  assign n42220 = ~n5950 & n19728 ;
  assign n42221 = n432 & ~n5741 ;
  assign n42222 = ( ~n14269 & n42220 ) | ( ~n14269 & n42221 ) | ( n42220 & n42221 ) ;
  assign n42223 = n42222 ^ n14090 ^ n5998 ;
  assign n42224 = n42223 ^ n1422 ^ n1202 ;
  assign n42225 = ~n2168 & n10293 ;
  assign n42226 = n42225 ^ n29188 ^ 1'b0 ;
  assign n42227 = n2894 & n37870 ;
  assign n42228 = n42227 ^ n18170 ^ 1'b0 ;
  assign n42229 = ~n18714 & n42228 ;
  assign n42230 = n29565 ^ n19491 ^ n16293 ;
  assign n42231 = ( n8412 & n15894 ) | ( n8412 & n17574 ) | ( n15894 & n17574 ) ;
  assign n42232 = ( n15480 & ~n36414 ) | ( n15480 & n42231 ) | ( ~n36414 & n42231 ) ;
  assign n42233 = ( n1329 & ~n6404 ) | ( n1329 & n9307 ) | ( ~n6404 & n9307 ) ;
  assign n42234 = n1981 | n14326 ;
  assign n42235 = n2423 & ~n42234 ;
  assign n42236 = ( n6427 & n12998 ) | ( n6427 & n42235 ) | ( n12998 & n42235 ) ;
  assign n42239 = n4577 & ~n35022 ;
  assign n42237 = ( n9840 & ~n15566 ) | ( n9840 & n27606 ) | ( ~n15566 & n27606 ) ;
  assign n42238 = ~n11612 & n42237 ;
  assign n42240 = n42239 ^ n42238 ^ n37141 ;
  assign n42243 = ( n14534 & n20576 ) | ( n14534 & ~n33843 ) | ( n20576 & ~n33843 ) ;
  assign n42241 = n13776 ^ n8643 ^ 1'b0 ;
  assign n42242 = n22366 | n42241 ;
  assign n42244 = n42243 ^ n42242 ^ 1'b0 ;
  assign n42245 = n42244 ^ n3370 ^ n614 ;
  assign n42247 = n23703 ^ n529 ^ x4 ;
  assign n42246 = n18013 ^ n11193 ^ n3214 ;
  assign n42248 = n42247 ^ n42246 ^ n22341 ;
  assign n42250 = n23066 ^ n2301 ^ n1048 ;
  assign n42252 = ( ~n4678 & n5783 ) | ( ~n4678 & n7114 ) | ( n5783 & n7114 ) ;
  assign n42251 = n17557 ^ n11850 ^ n2240 ;
  assign n42253 = n42252 ^ n42251 ^ 1'b0 ;
  assign n42254 = n42250 & n42253 ;
  assign n42249 = ( ~n11525 & n12702 ) | ( ~n11525 & n36015 ) | ( n12702 & n36015 ) ;
  assign n42255 = n42254 ^ n42249 ^ n39941 ;
  assign n42256 = n8425 ^ n1333 ^ n1146 ;
  assign n42257 = ( n22293 & ~n41173 ) | ( n22293 & n42256 ) | ( ~n41173 & n42256 ) ;
  assign n42258 = n18881 ^ n13190 ^ n5601 ;
  assign n42259 = ( n3697 & n8048 ) | ( n3697 & n22907 ) | ( n8048 & n22907 ) ;
  assign n42260 = ( n17179 & n26411 ) | ( n17179 & n28578 ) | ( n26411 & n28578 ) ;
  assign n42261 = n29045 ^ n19200 ^ 1'b0 ;
  assign n42262 = ( n3739 & ~n7741 ) | ( n3739 & n8274 ) | ( ~n7741 & n8274 ) ;
  assign n42263 = n42262 ^ n37848 ^ n20953 ;
  assign n42264 = n26255 ^ n25931 ^ n1696 ;
  assign n42265 = ~n3011 & n23478 ;
  assign n42266 = ( n28818 & n42264 ) | ( n28818 & n42265 ) | ( n42264 & n42265 ) ;
  assign n42267 = n39620 ^ n37246 ^ n33908 ;
  assign n42272 = ( ~n20517 & n29128 ) | ( ~n20517 & n36169 ) | ( n29128 & n36169 ) ;
  assign n42271 = x192 | n22797 ;
  assign n42269 = n29014 ^ n10785 ^ n10249 ;
  assign n42268 = n9021 ^ x118 ^ x116 ;
  assign n42270 = n42269 ^ n42268 ^ n40353 ;
  assign n42273 = n42272 ^ n42271 ^ n42270 ;
  assign n42274 = n18882 & n31533 ;
  assign n42275 = ( n2009 & ~n6316 ) | ( n2009 & n13630 ) | ( ~n6316 & n13630 ) ;
  assign n42276 = n40014 ^ n26466 ^ n22327 ;
  assign n42277 = n26464 & n29452 ;
  assign n42278 = n29160 & ~n42277 ;
  assign n42279 = n42278 ^ n33324 ^ n30854 ;
  assign n42280 = n335 & n6261 ;
  assign n42281 = n42280 ^ n23444 ^ 1'b0 ;
  assign n42282 = n6130 | n42281 ;
  assign n42283 = ( ~n18532 & n36133 ) | ( ~n18532 & n42282 ) | ( n36133 & n42282 ) ;
  assign n42284 = n36002 ^ n29224 ^ n25126 ;
  assign n42285 = ( n21512 & ~n31881 ) | ( n21512 & n42284 ) | ( ~n31881 & n42284 ) ;
  assign n42286 = n33081 ^ n32338 ^ n8537 ;
  assign n42287 = ( n11408 & n17856 ) | ( n11408 & n42286 ) | ( n17856 & n42286 ) ;
  assign n42288 = n19162 & n25534 ;
  assign n42289 = n42288 ^ n16081 ^ 1'b0 ;
  assign n42290 = ( n2769 & ~n7689 ) | ( n2769 & n42289 ) | ( ~n7689 & n42289 ) ;
  assign n42291 = n21979 ^ n5775 ^ n2535 ;
  assign n42292 = n11260 ^ n9147 ^ n6842 ;
  assign n42293 = n24832 | n42292 ;
  assign n42294 = ( n7575 & ~n42291 ) | ( n7575 & n42293 ) | ( ~n42291 & n42293 ) ;
  assign n42297 = n25313 ^ n10347 ^ n4690 ;
  assign n42296 = ( n14452 & ~n19162 ) | ( n14452 & n36632 ) | ( ~n19162 & n36632 ) ;
  assign n42295 = n35754 ^ n11737 ^ n698 ;
  assign n42298 = n42297 ^ n42296 ^ n42295 ;
  assign n42299 = n20449 ^ n15518 ^ 1'b0 ;
  assign n42300 = n6711 & ~n42299 ;
  assign n42301 = n32960 ^ n25778 ^ 1'b0 ;
  assign n42302 = ~n4598 & n42301 ;
  assign n42303 = n30886 ^ n12767 ^ 1'b0 ;
  assign n42304 = ( n6210 & n14341 ) | ( n6210 & ~n18153 ) | ( n14341 & ~n18153 ) ;
  assign n42305 = ( n34959 & n42303 ) | ( n34959 & n42304 ) | ( n42303 & n42304 ) ;
  assign n42306 = n18384 & ~n42305 ;
  assign n42307 = ~n38753 & n42306 ;
  assign n42308 = n972 | n42307 ;
  assign n42309 = n2834 ^ n1175 ^ n1097 ;
  assign n42310 = n42309 ^ n39359 ^ n1280 ;
  assign n42311 = n37900 ^ n37717 ^ 1'b0 ;
  assign n42312 = n22175 | n42311 ;
  assign n42313 = ( ~n15588 & n37485 ) | ( ~n15588 & n42312 ) | ( n37485 & n42312 ) ;
  assign n42314 = ( ~n619 & n7567 ) | ( ~n619 & n14232 ) | ( n7567 & n14232 ) ;
  assign n42315 = n42314 ^ n36317 ^ n35736 ;
  assign n42316 = n12334 & ~n33590 ;
  assign n42317 = n42316 ^ n35163 ^ 1'b0 ;
  assign n42318 = n3347 | n42317 ;
  assign n42319 = n42318 ^ n16765 ^ 1'b0 ;
  assign n42320 = ( ~n480 & n3996 ) | ( ~n480 & n5008 ) | ( n3996 & n5008 ) ;
  assign n42321 = n42320 ^ n13579 ^ n11541 ;
  assign n42322 = n42321 ^ n36108 ^ 1'b0 ;
  assign n42323 = n42322 ^ n30346 ^ n3873 ;
  assign n42324 = n19897 ^ n1394 ^ 1'b0 ;
  assign n42325 = ~n3799 & n42324 ;
  assign n42326 = ( n8789 & ~n22963 ) | ( n8789 & n42325 ) | ( ~n22963 & n42325 ) ;
  assign n42327 = ( ~n4473 & n13637 ) | ( ~n4473 & n38176 ) | ( n13637 & n38176 ) ;
  assign n42328 = n42327 ^ n8229 ^ n1500 ;
  assign n42329 = n15010 ^ n10174 ^ n6963 ;
  assign n42330 = n31736 | n40101 ;
  assign n42331 = n42330 ^ n33655 ^ n21448 ;
  assign n42332 = n9551 ^ n5984 ^ n4283 ;
  assign n42333 = n42332 ^ n37923 ^ n6145 ;
  assign n42334 = n42333 ^ n34341 ^ n25910 ;
  assign n42335 = n12188 ^ n8116 ^ 1'b0 ;
  assign n42336 = n38871 & ~n42335 ;
  assign n42337 = n11364 ^ n3735 ^ 1'b0 ;
  assign n42338 = n42336 & ~n42337 ;
  assign n42339 = n18195 ^ n11698 ^ n9628 ;
  assign n42340 = ( n3326 & n11260 ) | ( n3326 & ~n13458 ) | ( n11260 & ~n13458 ) ;
  assign n42341 = n42339 | n42340 ;
  assign n42342 = n6741 ^ n4875 ^ n2947 ;
  assign n42343 = ( n20403 & ~n38213 ) | ( n20403 & n42342 ) | ( ~n38213 & n42342 ) ;
  assign n42344 = ( n3900 & ~n28850 ) | ( n3900 & n42343 ) | ( ~n28850 & n42343 ) ;
  assign n42345 = ( n1436 & n2927 ) | ( n1436 & n7951 ) | ( n2927 & n7951 ) ;
  assign n42346 = n42345 ^ n24088 ^ n11903 ;
  assign n42347 = ~n31433 & n42346 ;
  assign n42348 = n42347 ^ n23073 ^ n10514 ;
  assign n42349 = n6128 & n42348 ;
  assign n42350 = n35205 ^ n24925 ^ n24817 ;
  assign n42351 = ( n6048 & ~n6189 ) | ( n6048 & n24778 ) | ( ~n6189 & n24778 ) ;
  assign n42352 = ( ~n12466 & n27389 ) | ( ~n12466 & n42351 ) | ( n27389 & n42351 ) ;
  assign n42353 = n35796 ^ n18192 ^ 1'b0 ;
  assign n42354 = ( n6283 & n42352 ) | ( n6283 & ~n42353 ) | ( n42352 & ~n42353 ) ;
  assign n42355 = ( n3878 & n12600 ) | ( n3878 & ~n17064 ) | ( n12600 & ~n17064 ) ;
  assign n42356 = n8189 & ~n15182 ;
  assign n42357 = n23028 & n42356 ;
  assign n42358 = n38599 ^ n33505 ^ 1'b0 ;
  assign n42359 = n42358 ^ n17548 ^ n15226 ;
  assign n42360 = ( n1188 & n40997 ) | ( n1188 & n42359 ) | ( n40997 & n42359 ) ;
  assign n42361 = ( ~n7977 & n14583 ) | ( ~n7977 & n26437 ) | ( n14583 & n26437 ) ;
  assign n42362 = n1271 | n4581 ;
  assign n42363 = ( n11197 & n11548 ) | ( n11197 & ~n24904 ) | ( n11548 & ~n24904 ) ;
  assign n42364 = n42363 ^ n33703 ^ n26953 ;
  assign n42365 = n40285 ^ n19541 ^ n2595 ;
  assign n42366 = n23329 & ~n42365 ;
  assign n42367 = n42366 ^ n19251 ^ n6064 ;
  assign n42368 = n42367 ^ n9961 ^ n7617 ;
  assign n42369 = n20664 ^ n16209 ^ n3598 ;
  assign n42370 = n42369 ^ n27982 ^ n19306 ;
  assign n42371 = ~n33374 & n37208 ;
  assign n42372 = n24479 ^ n20436 ^ n4921 ;
  assign n42373 = ( ~n14226 & n36852 ) | ( ~n14226 & n42372 ) | ( n36852 & n42372 ) ;
  assign n42374 = n3439 | n38263 ;
  assign n42375 = n8529 | n42374 ;
  assign n42376 = ( n16344 & n21177 ) | ( n16344 & ~n42375 ) | ( n21177 & ~n42375 ) ;
  assign n42377 = ( n15948 & ~n26818 ) | ( n15948 & n42376 ) | ( ~n26818 & n42376 ) ;
  assign n42378 = n42377 ^ n41365 ^ n1749 ;
  assign n42379 = n24343 ^ n4941 ^ n4149 ;
  assign n42380 = ( n13237 & n42332 ) | ( n13237 & n42379 ) | ( n42332 & n42379 ) ;
  assign n42381 = ( ~n2783 & n7546 ) | ( ~n2783 & n7784 ) | ( n7546 & n7784 ) ;
  assign n42382 = n42381 ^ n39083 ^ n15141 ;
  assign n42383 = n6084 & ~n7181 ;
  assign n42384 = n42383 ^ n38642 ^ 1'b0 ;
  assign n42385 = ~n500 & n29784 ;
  assign n42386 = n42385 ^ n20534 ^ 1'b0 ;
  assign n42387 = n7357 & ~n33379 ;
  assign n42388 = n3620 & n42387 ;
  assign n42389 = ( n18791 & n35333 ) | ( n18791 & ~n36512 ) | ( n35333 & ~n36512 ) ;
  assign n42390 = n11680 & n22026 ;
  assign n42391 = n12737 & n42390 ;
  assign n42392 = ( n2544 & n6701 ) | ( n2544 & ~n9850 ) | ( n6701 & ~n9850 ) ;
  assign n42393 = ( ~n1072 & n1528 ) | ( ~n1072 & n42392 ) | ( n1528 & n42392 ) ;
  assign n42394 = ( n31659 & n42391 ) | ( n31659 & ~n42393 ) | ( n42391 & ~n42393 ) ;
  assign n42395 = n38985 ^ n29105 ^ 1'b0 ;
  assign n42396 = ( n2665 & ~n7412 ) | ( n2665 & n15803 ) | ( ~n7412 & n15803 ) ;
  assign n42397 = n42396 ^ n11998 ^ n11648 ;
  assign n42398 = n42397 ^ n34138 ^ n28174 ;
  assign n42399 = n42395 & n42398 ;
  assign n42400 = ( n612 & n28833 ) | ( n612 & ~n30652 ) | ( n28833 & ~n30652 ) ;
  assign n42401 = n3292 | n5839 ;
  assign n42402 = n42401 ^ n37899 ^ n28441 ;
  assign n42403 = n20893 ^ n4642 ^ n2209 ;
  assign n42404 = ( n14532 & n19917 ) | ( n14532 & ~n42403 ) | ( n19917 & ~n42403 ) ;
  assign n42405 = ( n7971 & n36814 ) | ( n7971 & n42404 ) | ( n36814 & n42404 ) ;
  assign n42406 = n42405 ^ n8007 ^ n1487 ;
  assign n42407 = n36869 ^ n33836 ^ n3476 ;
  assign n42408 = n23632 ^ n19340 ^ 1'b0 ;
  assign n42409 = n1463 & n42408 ;
  assign n42410 = ~n31455 & n36710 ;
  assign n42411 = n42410 ^ n36672 ^ 1'b0 ;
  assign n42412 = ( n7344 & n10244 ) | ( n7344 & ~n21130 ) | ( n10244 & ~n21130 ) ;
  assign n42413 = ( ~n5079 & n38258 ) | ( ~n5079 & n42412 ) | ( n38258 & n42412 ) ;
  assign n42414 = ~n8455 & n37667 ;
  assign n42415 = n42414 ^ n10161 ^ 1'b0 ;
  assign n42416 = ( n20631 & ~n38957 ) | ( n20631 & n42415 ) | ( ~n38957 & n42415 ) ;
  assign n42417 = ( n1774 & n25770 ) | ( n1774 & ~n27888 ) | ( n25770 & ~n27888 ) ;
  assign n42418 = ( n8721 & n30178 ) | ( n8721 & n42417 ) | ( n30178 & n42417 ) ;
  assign n42419 = ( ~n14796 & n19369 ) | ( ~n14796 & n42418 ) | ( n19369 & n42418 ) ;
  assign n42420 = ( n3033 & n15593 ) | ( n3033 & n42419 ) | ( n15593 & n42419 ) ;
  assign n42421 = ( n6475 & n13251 ) | ( n6475 & ~n15160 ) | ( n13251 & ~n15160 ) ;
  assign n42422 = n42421 ^ n40203 ^ n23578 ;
  assign n42423 = ~n8234 & n42422 ;
  assign n42425 = n3876 & ~n4755 ;
  assign n42426 = n14845 & n42425 ;
  assign n42427 = n42426 ^ n33002 ^ n8980 ;
  assign n42424 = ( n23466 & n30970 ) | ( n23466 & ~n34012 ) | ( n30970 & ~n34012 ) ;
  assign n42428 = n42427 ^ n42424 ^ n30209 ;
  assign n42429 = n12761 ^ n12039 ^ 1'b0 ;
  assign n42430 = n42429 ^ n35927 ^ n33386 ;
  assign n42431 = n20943 ^ n11280 ^ n8904 ;
  assign n42432 = n42431 ^ n13583 ^ 1'b0 ;
  assign n42433 = n20412 & ~n42432 ;
  assign n42434 = n4343 & ~n36562 ;
  assign n42435 = ~n42433 & n42434 ;
  assign n42436 = ( ~n10620 & n14034 ) | ( ~n10620 & n19485 ) | ( n14034 & n19485 ) ;
  assign n42437 = ( n7630 & ~n31079 ) | ( n7630 & n40989 ) | ( ~n31079 & n40989 ) ;
  assign n42438 = n38518 ^ n15510 ^ n14533 ;
  assign n42440 = n22476 ^ n4064 ^ 1'b0 ;
  assign n42441 = n13673 & ~n42440 ;
  assign n42439 = ( n1956 & n7938 ) | ( n1956 & ~n18182 ) | ( n7938 & ~n18182 ) ;
  assign n42442 = n42441 ^ n42439 ^ n13826 ;
  assign n42444 = n10662 ^ n9753 ^ n6026 ;
  assign n42443 = n30415 ^ n22936 ^ n2601 ;
  assign n42445 = n42444 ^ n42443 ^ n14229 ;
  assign n42446 = n42445 ^ n12872 ^ n7865 ;
  assign n42447 = n5103 | n27908 ;
  assign n42448 = n33595 & ~n42447 ;
  assign n42449 = n36918 ^ n20728 ^ n3625 ;
  assign n42450 = n25197 ^ n22063 ^ n11160 ;
  assign n42451 = n21257 & n37060 ;
  assign n42452 = n6378 & n42451 ;
  assign n42453 = n13782 & n29107 ;
  assign n42454 = n42452 & n42453 ;
  assign n42455 = ( n8945 & n18440 ) | ( n8945 & ~n42454 ) | ( n18440 & ~n42454 ) ;
  assign n42457 = n25314 ^ n11545 ^ 1'b0 ;
  assign n42458 = n16634 | n42457 ;
  assign n42456 = n10514 ^ n3026 ^ 1'b0 ;
  assign n42459 = n42458 ^ n42456 ^ n21448 ;
  assign n42460 = n21419 ^ n7089 ^ 1'b0 ;
  assign n42461 = n32197 ^ n30187 ^ n3917 ;
  assign n42462 = ( n20014 & n42460 ) | ( n20014 & ~n42461 ) | ( n42460 & ~n42461 ) ;
  assign n42463 = n29277 ^ n16145 ^ x251 ;
  assign n42464 = n42463 ^ n19769 ^ 1'b0 ;
  assign n42465 = n7251 | n42464 ;
  assign n42466 = n10611 ^ n8203 ^ 1'b0 ;
  assign n42467 = n21267 & n42466 ;
  assign n42468 = n14008 ^ n7852 ^ 1'b0 ;
  assign n42469 = n30203 | n35036 ;
  assign n42470 = n34945 ^ n28223 ^ 1'b0 ;
  assign n42471 = n26096 ^ n24590 ^ n9510 ;
  assign n42472 = n42471 ^ n15450 ^ n2917 ;
  assign n42473 = n17216 ^ n491 ^ 1'b0 ;
  assign n42474 = ~n32307 & n42473 ;
  assign n42475 = n35262 & n42474 ;
  assign n42476 = n38756 ^ n26062 ^ n9913 ;
  assign n42477 = n25710 | n42476 ;
  assign n42478 = n10853 & ~n42477 ;
  assign n42479 = ( n6779 & n42475 ) | ( n6779 & ~n42478 ) | ( n42475 & ~n42478 ) ;
  assign n42480 = ( n27767 & ~n42472 ) | ( n27767 & n42479 ) | ( ~n42472 & n42479 ) ;
  assign n42481 = n16062 ^ n11691 ^ n994 ;
  assign n42482 = ( ~n406 & n33142 ) | ( ~n406 & n42481 ) | ( n33142 & n42481 ) ;
  assign n42483 = ( n12996 & n17108 ) | ( n12996 & ~n34259 ) | ( n17108 & ~n34259 ) ;
  assign n42484 = n37281 ^ n17691 ^ n5508 ;
  assign n42485 = n42484 ^ n36698 ^ n25516 ;
  assign n42490 = n37693 ^ n30815 ^ n11413 ;
  assign n42486 = n21288 ^ n6674 ^ n1139 ;
  assign n42487 = ( n3334 & ~n11149 ) | ( n3334 & n42486 ) | ( ~n11149 & n42486 ) ;
  assign n42488 = n42487 ^ n38874 ^ 1'b0 ;
  assign n42489 = n30612 & n42488 ;
  assign n42491 = n42490 ^ n42489 ^ n8910 ;
  assign n42492 = ( ~n18523 & n34870 ) | ( ~n18523 & n37493 ) | ( n34870 & n37493 ) ;
  assign n42493 = ( n4319 & n4374 ) | ( n4319 & n5154 ) | ( n4374 & n5154 ) ;
  assign n42494 = n1459 & ~n4520 ;
  assign n42495 = ( n4900 & n42493 ) | ( n4900 & ~n42494 ) | ( n42493 & ~n42494 ) ;
  assign n42496 = ( ~n4799 & n38769 ) | ( ~n4799 & n42495 ) | ( n38769 & n42495 ) ;
  assign n42497 = ( n9317 & n15208 ) | ( n9317 & ~n20296 ) | ( n15208 & ~n20296 ) ;
  assign n42498 = n8337 ^ n7706 ^ n1733 ;
  assign n42499 = n18786 & ~n24670 ;
  assign n42500 = n3189 & n42499 ;
  assign n42501 = ( n42497 & n42498 ) | ( n42497 & n42500 ) | ( n42498 & n42500 ) ;
  assign n42502 = ~n1238 & n7699 ;
  assign n42503 = n42502 ^ n27482 ^ 1'b0 ;
  assign n42504 = ( n8468 & n10428 ) | ( n8468 & n37588 ) | ( n10428 & n37588 ) ;
  assign n42505 = n11847 & n21546 ;
  assign n42506 = n42504 & n42505 ;
  assign n42508 = n18740 ^ n15927 ^ n12448 ;
  assign n42507 = n25461 ^ n21079 ^ n18397 ;
  assign n42509 = n42508 ^ n42507 ^ n2133 ;
  assign n42510 = n42509 ^ n363 ^ 1'b0 ;
  assign n42511 = ~n10357 & n42510 ;
  assign n42512 = ( n27191 & ~n32663 ) | ( n27191 & n37972 ) | ( ~n32663 & n37972 ) ;
  assign n42513 = n22824 ^ n14114 ^ n1436 ;
  assign n42514 = n42513 ^ n40794 ^ 1'b0 ;
  assign n42515 = n31047 ^ n21775 ^ n10828 ;
  assign n42516 = ( n10416 & ~n14307 ) | ( n10416 & n42515 ) | ( ~n14307 & n42515 ) ;
  assign n42517 = ( n2560 & ~n18282 ) | ( n2560 & n22780 ) | ( ~n18282 & n22780 ) ;
  assign n42518 = n9524 & n21421 ;
  assign n42519 = ( n18969 & ~n42517 ) | ( n18969 & n42518 ) | ( ~n42517 & n42518 ) ;
  assign n42520 = n19683 ^ n15760 ^ n6502 ;
  assign n42521 = ( ~n12256 & n22015 ) | ( ~n12256 & n42520 ) | ( n22015 & n42520 ) ;
  assign n42522 = n29168 ^ n23667 ^ 1'b0 ;
  assign n42523 = n40662 ^ n1724 ^ 1'b0 ;
  assign n42524 = n37518 ^ n13918 ^ n9368 ;
  assign n42526 = ( n17299 & n22322 ) | ( n17299 & n24949 ) | ( n22322 & n24949 ) ;
  assign n42525 = n33139 ^ n31000 ^ n12042 ;
  assign n42527 = n42526 ^ n42525 ^ n4099 ;
  assign n42529 = ( n1610 & ~n14184 ) | ( n1610 & n16704 ) | ( ~n14184 & n16704 ) ;
  assign n42528 = n915 & ~n27436 ;
  assign n42530 = n42529 ^ n42528 ^ 1'b0 ;
  assign n42531 = n42530 ^ n38451 ^ n12173 ;
  assign n42532 = n42132 ^ n25358 ^ n6232 ;
  assign n42533 = n42532 ^ n11573 ^ 1'b0 ;
  assign n42534 = n20034 ^ n8784 ^ 1'b0 ;
  assign n42535 = n42534 ^ n36525 ^ n26270 ;
  assign n42536 = n13409 | n18772 ;
  assign n42537 = n40797 ^ n33299 ^ n26719 ;
  assign n42538 = n35180 ^ n28411 ^ n3853 ;
  assign n42539 = n3396 & n16172 ;
  assign n42540 = ~n42538 & n42539 ;
  assign n42541 = n20227 ^ n2223 ^ 1'b0 ;
  assign n42542 = ( n18705 & n36173 ) | ( n18705 & n42541 ) | ( n36173 & n42541 ) ;
  assign n42543 = ~n16315 & n41353 ;
  assign n42544 = ( n21506 & ~n34907 ) | ( n21506 & n42543 ) | ( ~n34907 & n42543 ) ;
  assign n42545 = n32332 ^ n6999 ^ 1'b0 ;
  assign n42546 = ( n21945 & ~n29979 ) | ( n21945 & n42545 ) | ( ~n29979 & n42545 ) ;
  assign n42547 = n20101 ^ n9870 ^ n3495 ;
  assign n42548 = n26662 ^ n11555 ^ 1'b0 ;
  assign n42549 = ( n42546 & n42547 ) | ( n42546 & n42548 ) | ( n42547 & n42548 ) ;
  assign n42556 = n4500 & ~n6083 ;
  assign n42550 = n26811 ^ n15129 ^ 1'b0 ;
  assign n42551 = n10657 | n42550 ;
  assign n42552 = n15115 ^ n4643 ^ n2589 ;
  assign n42553 = ( n29884 & n42551 ) | ( n29884 & ~n42552 ) | ( n42551 & ~n42552 ) ;
  assign n42554 = n42553 ^ n6061 ^ 1'b0 ;
  assign n42555 = n35361 | n42554 ;
  assign n42557 = n42556 ^ n42555 ^ n10505 ;
  assign n42558 = n6886 ^ n1481 ^ 1'b0 ;
  assign n42559 = ( n2363 & n9664 ) | ( n2363 & ~n20892 ) | ( n9664 & ~n20892 ) ;
  assign n42560 = ( n10271 & n42558 ) | ( n10271 & ~n42559 ) | ( n42558 & ~n42559 ) ;
  assign n42561 = n42560 ^ n16244 ^ n3708 ;
  assign n42562 = ( n7884 & ~n15061 ) | ( n7884 & n22704 ) | ( ~n15061 & n22704 ) ;
  assign n42563 = n36357 ^ n28223 ^ n17662 ;
  assign n42564 = n24390 ^ n23439 ^ n8386 ;
  assign n42565 = ( n42562 & n42563 ) | ( n42562 & ~n42564 ) | ( n42563 & ~n42564 ) ;
  assign n42566 = n29014 ^ n15293 ^ n9399 ;
  assign n42567 = n8716 & n36045 ;
  assign n42568 = n42567 ^ n27837 ^ n5761 ;
  assign n42569 = ( n18663 & ~n21733 ) | ( n18663 & n25892 ) | ( ~n21733 & n25892 ) ;
  assign n42570 = n42569 ^ n39588 ^ n7439 ;
  assign n42571 = ( n4637 & ~n13360 ) | ( n4637 & n42570 ) | ( ~n13360 & n42570 ) ;
  assign n42574 = n3941 & n15107 ;
  assign n42575 = n24093 & n42574 ;
  assign n42572 = ( x122 & n14149 ) | ( x122 & n19682 ) | ( n14149 & n19682 ) ;
  assign n42573 = n42572 ^ n13189 ^ 1'b0 ;
  assign n42576 = n42575 ^ n42573 ^ n37111 ;
  assign n42577 = n31971 ^ n6043 ^ n5230 ;
  assign n42578 = n42577 ^ n27916 ^ n23388 ;
  assign n42580 = n15934 | n20517 ;
  assign n42579 = n22755 & ~n37864 ;
  assign n42581 = n42580 ^ n42579 ^ 1'b0 ;
  assign n42582 = ~n19113 & n32129 ;
  assign n42583 = n42582 ^ n30403 ^ 1'b0 ;
  assign n42584 = n36665 ^ n30370 ^ n15346 ;
  assign n42585 = n41643 ^ n3177 ^ 1'b0 ;
  assign n42588 = n18551 ^ n15868 ^ n4448 ;
  assign n42589 = n42588 ^ n26459 ^ n7292 ;
  assign n42586 = ~n3100 & n29738 ;
  assign n42587 = n42586 ^ n29786 ^ 1'b0 ;
  assign n42590 = n42589 ^ n42587 ^ n29282 ;
  assign n42591 = n15112 & ~n26718 ;
  assign n42592 = ( n2938 & ~n23473 ) | ( n2938 & n42591 ) | ( ~n23473 & n42591 ) ;
  assign n42593 = n9624 ^ n3685 ^ 1'b0 ;
  assign n42594 = n12346 ^ n305 ^ 1'b0 ;
  assign n42595 = ( ~n5083 & n31013 ) | ( ~n5083 & n42594 ) | ( n31013 & n42594 ) ;
  assign n42596 = n36226 ^ n22132 ^ 1'b0 ;
  assign n42597 = ~n6809 & n22792 ;
  assign n42598 = ~n9177 & n42597 ;
  assign n42599 = n42598 ^ n14824 ^ 1'b0 ;
  assign n42600 = n42599 ^ n24025 ^ 1'b0 ;
  assign n42601 = n9744 & ~n28347 ;
  assign n42602 = n24827 | n37767 ;
  assign n42603 = ( ~n25935 & n42601 ) | ( ~n25935 & n42602 ) | ( n42601 & n42602 ) ;
  assign n42604 = n42603 ^ n41533 ^ 1'b0 ;
  assign n42605 = n4079 & ~n42604 ;
  assign n42606 = ( n1425 & n7482 ) | ( n1425 & n13393 ) | ( n7482 & n13393 ) ;
  assign n42607 = n42606 ^ n27370 ^ 1'b0 ;
  assign n42608 = n12862 ^ n10400 ^ 1'b0 ;
  assign n42609 = n42607 & n42608 ;
  assign n42610 = n16418 ^ n11750 ^ n4434 ;
  assign n42613 = n18036 ^ n15212 ^ n8463 ;
  assign n42611 = x201 & n4053 ;
  assign n42612 = n3820 & n42611 ;
  assign n42614 = n42613 ^ n42612 ^ n16446 ;
  assign n42615 = ( n28865 & n34307 ) | ( n28865 & ~n42614 ) | ( n34307 & ~n42614 ) ;
  assign n42616 = n42615 ^ n42564 ^ n28291 ;
  assign n42617 = ( n5073 & ~n7615 ) | ( n5073 & n42616 ) | ( ~n7615 & n42616 ) ;
  assign n42618 = n1306 & ~n24443 ;
  assign n42619 = ( n2733 & ~n29079 ) | ( n2733 & n42618 ) | ( ~n29079 & n42618 ) ;
  assign n42620 = n42619 ^ n40790 ^ n2805 ;
  assign n42623 = n39054 ^ n15042 ^ 1'b0 ;
  assign n42621 = n10287 ^ n3204 ^ 1'b0 ;
  assign n42622 = n11739 & ~n42621 ;
  assign n42624 = n42623 ^ n42622 ^ n36057 ;
  assign n42625 = ( n9841 & n20141 ) | ( n9841 & n42624 ) | ( n20141 & n42624 ) ;
  assign n42630 = n23539 ^ n2826 ^ 1'b0 ;
  assign n42631 = n34649 | n42630 ;
  assign n42626 = n8400 ^ n8105 ^ n2523 ;
  assign n42627 = n17124 & ~n19131 ;
  assign n42628 = n42627 ^ n21823 ^ 1'b0 ;
  assign n42629 = ( n2965 & n42626 ) | ( n2965 & ~n42628 ) | ( n42626 & ~n42628 ) ;
  assign n42632 = n42631 ^ n42629 ^ n16511 ;
  assign n42633 = n25437 ^ n6136 ^ 1'b0 ;
  assign n42634 = ~n16579 & n42633 ;
  assign n42635 = n42634 ^ n12320 ^ n4641 ;
  assign n42636 = ( n5921 & n14730 ) | ( n5921 & n29311 ) | ( n14730 & n29311 ) ;
  assign n42637 = ( ~n11809 & n17894 ) | ( ~n11809 & n30142 ) | ( n17894 & n30142 ) ;
  assign n42638 = ( n6981 & n17631 ) | ( n6981 & ~n22583 ) | ( n17631 & ~n22583 ) ;
  assign n42641 = ( n12169 & n13337 ) | ( n12169 & n21525 ) | ( n13337 & n21525 ) ;
  assign n42639 = n14928 & n25089 ;
  assign n42640 = n42639 ^ n28694 ^ n14190 ;
  assign n42642 = n42641 ^ n42640 ^ 1'b0 ;
  assign n42643 = ( n17881 & n32491 ) | ( n17881 & n42642 ) | ( n32491 & n42642 ) ;
  assign n42644 = n21719 ^ n12448 ^ n5797 ;
  assign n42645 = ( ~n6149 & n22761 ) | ( ~n6149 & n42644 ) | ( n22761 & n42644 ) ;
  assign n42646 = ( n8184 & n29817 ) | ( n8184 & ~n42645 ) | ( n29817 & ~n42645 ) ;
  assign n42647 = n37442 ^ n36538 ^ 1'b0 ;
  assign n42648 = ~n29889 & n42647 ;
  assign n42649 = n4044 & n13127 ;
  assign n42650 = ~n2211 & n42649 ;
  assign n42651 = n30203 ^ n12408 ^ 1'b0 ;
  assign n42652 = n1412 & n42651 ;
  assign n42653 = n42652 ^ n35649 ^ n19409 ;
  assign n42654 = n10919 ^ n6327 ^ n747 ;
  assign n42655 = n21694 & ~n42654 ;
  assign n42656 = n42655 ^ n11214 ^ 1'b0 ;
  assign n42657 = ( n4187 & n31127 ) | ( n4187 & n42656 ) | ( n31127 & n42656 ) ;
  assign n42658 = n11252 ^ n9352 ^ n8628 ;
  assign n42659 = n42658 ^ n33505 ^ n32902 ;
  assign n42660 = n3459 & n8040 ;
  assign n42661 = n20863 ^ n10417 ^ 1'b0 ;
  assign n42662 = ~n34877 & n42661 ;
  assign n42663 = n42662 ^ n9524 ^ n5446 ;
  assign n42664 = ( ~n5307 & n8710 ) | ( ~n5307 & n23328 ) | ( n8710 & n23328 ) ;
  assign n42665 = ( n2599 & n9669 ) | ( n2599 & n42664 ) | ( n9669 & n42664 ) ;
  assign n42666 = ( n12882 & ~n35011 ) | ( n12882 & n42665 ) | ( ~n35011 & n42665 ) ;
  assign n42667 = n13938 & n29070 ;
  assign n42668 = n42667 ^ x143 ^ 1'b0 ;
  assign n42669 = n42668 ^ n16248 ^ n6090 ;
  assign n42670 = n7809 & n42669 ;
  assign n42671 = ~n42666 & n42670 ;
  assign n42672 = n26656 ^ n10214 ^ n6824 ;
  assign n42673 = n11190 & ~n27490 ;
  assign n42674 = n42672 & n42673 ;
  assign n42675 = n18195 ^ n7145 ^ n3985 ;
  assign n42676 = ( n796 & ~n1160 ) | ( n796 & n13888 ) | ( ~n1160 & n13888 ) ;
  assign n42677 = ( n19880 & ~n42675 ) | ( n19880 & n42676 ) | ( ~n42675 & n42676 ) ;
  assign n42678 = ( n3701 & n18603 ) | ( n3701 & ~n28241 ) | ( n18603 & ~n28241 ) ;
  assign n42679 = ( n4337 & n4993 ) | ( n4337 & n36307 ) | ( n4993 & n36307 ) ;
  assign n42680 = n42679 ^ n20285 ^ n3259 ;
  assign n42681 = n31530 ^ n11311 ^ 1'b0 ;
  assign n42682 = ( n8279 & n10540 ) | ( n8279 & n12869 ) | ( n10540 & n12869 ) ;
  assign n42683 = ( n11159 & n28333 ) | ( n11159 & ~n42682 ) | ( n28333 & ~n42682 ) ;
  assign n42684 = n42683 ^ n5660 ^ 1'b0 ;
  assign n42685 = n42684 ^ n24834 ^ n18666 ;
  assign n42686 = n11452 | n19235 ;
  assign n42687 = n22060 ^ n10138 ^ n4591 ;
  assign n42688 = ( n1407 & n39241 ) | ( n1407 & ~n42687 ) | ( n39241 & ~n42687 ) ;
  assign n42689 = n33464 | n38886 ;
  assign n42690 = n7140 & ~n42689 ;
  assign n42691 = n42690 ^ n16036 ^ 1'b0 ;
  assign n42692 = n28844 ^ n23728 ^ n7202 ;
  assign n42693 = ( n11270 & n34924 ) | ( n11270 & ~n42692 ) | ( n34924 & ~n42692 ) ;
  assign n42694 = ( n11388 & n28233 ) | ( n11388 & n42693 ) | ( n28233 & n42693 ) ;
  assign n42695 = n18802 & ~n42694 ;
  assign n42696 = ( n7413 & n11270 ) | ( n7413 & ~n18079 ) | ( n11270 & ~n18079 ) ;
  assign n42697 = ( ~n15777 & n36603 ) | ( ~n15777 & n41834 ) | ( n36603 & n41834 ) ;
  assign n42698 = n42697 ^ n25313 ^ 1'b0 ;
  assign n42699 = n20616 ^ n17638 ^ n10658 ;
  assign n42700 = n34812 & n42699 ;
  assign n42701 = ( ~n12624 & n21534 ) | ( ~n12624 & n27347 ) | ( n21534 & n27347 ) ;
  assign n42702 = n38982 ^ n25908 ^ 1'b0 ;
  assign n42703 = n13261 | n42702 ;
  assign n42704 = n42703 ^ n35822 ^ n14055 ;
  assign n42705 = ( n5224 & n5338 ) | ( n5224 & ~n10015 ) | ( n5338 & ~n10015 ) ;
  assign n42706 = n11666 ^ n6677 ^ 1'b0 ;
  assign n42707 = n42705 & ~n42706 ;
  assign n42708 = n12547 ^ x168 ^ 1'b0 ;
  assign n42709 = n40875 ^ n30407 ^ 1'b0 ;
  assign n42710 = n40712 ^ n17629 ^ 1'b0 ;
  assign n42711 = ( ~n24925 & n26702 ) | ( ~n24925 & n30746 ) | ( n26702 & n30746 ) ;
  assign n42712 = n42711 ^ n38233 ^ n10950 ;
  assign n42714 = n14468 ^ n3190 ^ n1769 ;
  assign n42713 = n1483 & ~n29380 ;
  assign n42715 = n42714 ^ n42713 ^ 1'b0 ;
  assign n42717 = ( ~n15266 & n18132 ) | ( ~n15266 & n24702 ) | ( n18132 & n24702 ) ;
  assign n42716 = n27814 ^ n17422 ^ n15139 ;
  assign n42718 = n42717 ^ n42716 ^ n37437 ;
  assign n42719 = ( n13772 & n18532 ) | ( n13772 & n30690 ) | ( n18532 & n30690 ) ;
  assign n42720 = ( n4068 & ~n7440 ) | ( n4068 & n42719 ) | ( ~n7440 & n42719 ) ;
  assign n42721 = n36749 ^ n34828 ^ n30986 ;
  assign n42722 = ~n17854 & n42721 ;
  assign n42723 = n22781 ^ n16096 ^ n9848 ;
  assign n42724 = n42723 ^ n14672 ^ 1'b0 ;
  assign n42725 = n42724 ^ n34306 ^ n9428 ;
  assign n42726 = ( n4699 & n4715 ) | ( n4699 & n13110 ) | ( n4715 & n13110 ) ;
  assign n42727 = n15747 & n34774 ;
  assign n42728 = n42727 ^ n12671 ^ 1'b0 ;
  assign n42729 = ( n1824 & n5857 ) | ( n1824 & n23027 ) | ( n5857 & n23027 ) ;
  assign n42730 = n42729 ^ n29460 ^ n24078 ;
  assign n42731 = n42730 ^ n15169 ^ n7860 ;
  assign n42732 = ( n5016 & ~n11806 ) | ( n5016 & n30936 ) | ( ~n11806 & n30936 ) ;
  assign n42733 = ( n15030 & ~n25343 ) | ( n15030 & n42732 ) | ( ~n25343 & n42732 ) ;
  assign n42734 = ( n1282 & n28300 ) | ( n1282 & ~n37081 ) | ( n28300 & ~n37081 ) ;
  assign n42735 = n25711 | n40761 ;
  assign n42736 = n42735 ^ n4694 ^ 1'b0 ;
  assign n42737 = ( n5721 & n38231 ) | ( n5721 & ~n42736 ) | ( n38231 & ~n42736 ) ;
  assign n42738 = ~n11059 & n42737 ;
  assign n42739 = n33375 ^ n24205 ^ n23776 ;
  assign n42740 = ( ~n1937 & n5590 ) | ( ~n1937 & n10451 ) | ( n5590 & n10451 ) ;
  assign n42741 = n42740 ^ n39764 ^ n11613 ;
  assign n42742 = n10389 & n33117 ;
  assign n42743 = ( n5191 & n10917 ) | ( n5191 & ~n42742 ) | ( n10917 & ~n42742 ) ;
  assign n42744 = ( n958 & n11023 ) | ( n958 & ~n42743 ) | ( n11023 & ~n42743 ) ;
  assign n42745 = n33615 ^ n10039 ^ 1'b0 ;
  assign n42746 = n31699 ^ n17742 ^ 1'b0 ;
  assign n42747 = n13176 & ~n42746 ;
  assign n42748 = ( n477 & n8829 ) | ( n477 & ~n8920 ) | ( n8829 & ~n8920 ) ;
  assign n42749 = n42748 ^ n12733 ^ n11668 ;
  assign n42750 = ~n17252 & n42749 ;
  assign n42751 = ~n18530 & n41863 ;
  assign n42752 = ( n4301 & n42750 ) | ( n4301 & n42751 ) | ( n42750 & n42751 ) ;
  assign n42754 = n41356 ^ n36176 ^ n12980 ;
  assign n42753 = n25844 ^ n11234 ^ n372 ;
  assign n42755 = n42754 ^ n42753 ^ 1'b0 ;
  assign n42756 = n38789 ^ n34389 ^ 1'b0 ;
  assign n42757 = ( n1336 & n22322 ) | ( n1336 & n38947 ) | ( n22322 & n38947 ) ;
  assign n42758 = n12416 & ~n42757 ;
  assign n42759 = n16623 ^ n15703 ^ n6679 ;
  assign n42760 = n42759 ^ n40038 ^ 1'b0 ;
  assign n42761 = n1125 & ~n42760 ;
  assign n42762 = n36291 ^ n12166 ^ 1'b0 ;
  assign n42763 = n42429 ^ n35292 ^ n8826 ;
  assign n42764 = n42763 ^ n5402 ^ 1'b0 ;
  assign n42765 = ~n42762 & n42764 ;
  assign n42766 = n26859 | n37566 ;
  assign n42767 = ( n1707 & n3541 ) | ( n1707 & n11071 ) | ( n3541 & n11071 ) ;
  assign n42768 = n31455 ^ n19232 ^ n2294 ;
  assign n42769 = n31112 ^ n27204 ^ n16582 ;
  assign n42770 = ( n388 & n25745 ) | ( n388 & ~n42769 ) | ( n25745 & ~n42769 ) ;
  assign n42771 = n42770 ^ n40365 ^ n14374 ;
  assign n42772 = n42771 ^ n34254 ^ n11899 ;
  assign n42774 = n27204 ^ n4208 ^ 1'b0 ;
  assign n42773 = n35299 ^ n7174 ^ 1'b0 ;
  assign n42775 = n42774 ^ n42773 ^ n31344 ;
  assign n42776 = ( n20590 & n28871 ) | ( n20590 & n39819 ) | ( n28871 & n39819 ) ;
  assign n42777 = ( n13880 & ~n13942 ) | ( n13880 & n28021 ) | ( ~n13942 & n28021 ) ;
  assign n42778 = n42777 ^ n30393 ^ n25803 ;
  assign n42779 = n42778 ^ n38277 ^ n622 ;
  assign n42780 = n10274 & ~n41890 ;
  assign n42781 = n35852 ^ n12161 ^ 1'b0 ;
  assign n42782 = ~n18262 & n42781 ;
  assign n42783 = n29117 ^ n2311 ^ 1'b0 ;
  assign n42784 = n42783 ^ n11373 ^ n3221 ;
  assign n42785 = n33070 ^ n30403 ^ n9053 ;
  assign n42786 = n5591 ^ n1964 ^ x190 ;
  assign n42787 = ( n12329 & ~n23996 ) | ( n12329 & n42786 ) | ( ~n23996 & n42786 ) ;
  assign n42791 = n5048 & ~n9571 ;
  assign n42792 = n42791 ^ n7977 ^ 1'b0 ;
  assign n42789 = ~n3300 & n17601 ;
  assign n42790 = n6459 & n42789 ;
  assign n42788 = n18854 ^ n10241 ^ n6773 ;
  assign n42793 = n42792 ^ n42790 ^ n42788 ;
  assign n42794 = n41051 ^ n34148 ^ n10002 ;
  assign n42799 = n25428 ^ n14462 ^ n1282 ;
  assign n42800 = ( n20229 & n28382 ) | ( n20229 & ~n33359 ) | ( n28382 & ~n33359 ) ;
  assign n42801 = n42800 ^ n29203 ^ n407 ;
  assign n42802 = ( n12616 & n42799 ) | ( n12616 & ~n42801 ) | ( n42799 & ~n42801 ) ;
  assign n42795 = n4320 ^ n2976 ^ 1'b0 ;
  assign n42796 = n6933 & ~n42795 ;
  assign n42797 = ( ~n5037 & n9609 ) | ( ~n5037 & n19418 ) | ( n9609 & n19418 ) ;
  assign n42798 = ( ~n21003 & n42796 ) | ( ~n21003 & n42797 ) | ( n42796 & n42797 ) ;
  assign n42803 = n42802 ^ n42798 ^ n24316 ;
  assign n42805 = n7614 ^ n4744 ^ n1337 ;
  assign n42804 = ( ~n4025 & n13348 ) | ( ~n4025 & n14944 ) | ( n13348 & n14944 ) ;
  assign n42806 = n42805 ^ n42804 ^ n36751 ;
  assign n42807 = ~n35344 & n42806 ;
  assign n42809 = n24233 ^ n9647 ^ 1'b0 ;
  assign n42808 = n4509 | n30479 ;
  assign n42810 = n42809 ^ n42808 ^ 1'b0 ;
  assign n42811 = ( n7689 & n31333 ) | ( n7689 & n32987 ) | ( n31333 & n32987 ) ;
  assign n42812 = ( n5338 & n15392 ) | ( n5338 & n41463 ) | ( n15392 & n41463 ) ;
  assign n42813 = n29234 ^ n25110 ^ n9608 ;
  assign n42814 = ( n5778 & ~n22663 ) | ( n5778 & n26093 ) | ( ~n22663 & n26093 ) ;
  assign n42815 = ( n8402 & ~n8635 ) | ( n8402 & n40503 ) | ( ~n8635 & n40503 ) ;
  assign n42816 = n11251 ^ n5598 ^ 1'b0 ;
  assign n42817 = n34371 | n42816 ;
  assign n42820 = ( n1463 & n11766 ) | ( n1463 & ~n31092 ) | ( n11766 & ~n31092 ) ;
  assign n42819 = n8017 | n31441 ;
  assign n42821 = n42820 ^ n42819 ^ 1'b0 ;
  assign n42818 = n26130 ^ n24877 ^ n5346 ;
  assign n42822 = n42821 ^ n42818 ^ n13671 ;
  assign n42823 = n32714 | n39471 ;
  assign n42824 = n42822 | n42823 ;
  assign n42825 = n30975 ^ n986 ^ 1'b0 ;
  assign n42826 = n42622 & n42825 ;
  assign n42827 = ( x46 & n3390 ) | ( x46 & ~n27768 ) | ( n3390 & ~n27768 ) ;
  assign n42829 = n13459 ^ n8573 ^ n7454 ;
  assign n42830 = ( n9173 & n24294 ) | ( n9173 & ~n42829 ) | ( n24294 & ~n42829 ) ;
  assign n42828 = n2876 & ~n27955 ;
  assign n42831 = n42830 ^ n42828 ^ n14473 ;
  assign n42832 = n28836 ^ n8968 ^ n2225 ;
  assign n42833 = ( n32252 & ~n41010 ) | ( n32252 & n42832 ) | ( ~n41010 & n42832 ) ;
  assign n42834 = ( n3657 & ~n4544 ) | ( n3657 & n7634 ) | ( ~n4544 & n7634 ) ;
  assign n42835 = n1522 & n8927 ;
  assign n42836 = n16855 ^ n16201 ^ n623 ;
  assign n42837 = n42835 & n42836 ;
  assign n42838 = ( n6788 & n8640 ) | ( n6788 & n42837 ) | ( n8640 & n42837 ) ;
  assign n42839 = x32 & ~n6081 ;
  assign n42840 = n42839 ^ n11782 ^ 1'b0 ;
  assign n42841 = n42840 ^ n20590 ^ n8233 ;
  assign n42847 = ( n7838 & ~n13688 ) | ( n7838 & n30953 ) | ( ~n13688 & n30953 ) ;
  assign n42842 = n30601 ^ n7340 ^ n6958 ;
  assign n42843 = n42842 ^ n28291 ^ n25794 ;
  assign n42844 = ~n1579 & n42843 ;
  assign n42845 = ( n19170 & ~n38500 ) | ( n19170 & n42844 ) | ( ~n38500 & n42844 ) ;
  assign n42846 = n25710 | n42845 ;
  assign n42848 = n42847 ^ n42846 ^ 1'b0 ;
  assign n42849 = x154 & ~n16616 ;
  assign n42850 = n32038 & n42849 ;
  assign n42851 = ( ~n10957 & n11495 ) | ( ~n10957 & n39119 ) | ( n11495 & n39119 ) ;
  assign n42852 = n42851 ^ n31723 ^ 1'b0 ;
  assign n42853 = ~n42850 & n42852 ;
  assign n42854 = n22686 ^ n20431 ^ n16858 ;
  assign n42855 = n13245 & n42854 ;
  assign n42856 = n17989 & n42855 ;
  assign n42857 = ( n6752 & ~n35985 ) | ( n6752 & n42856 ) | ( ~n35985 & n42856 ) ;
  assign n42858 = n14390 ^ n9549 ^ n3414 ;
  assign n42859 = ( n12707 & ~n42857 ) | ( n12707 & n42858 ) | ( ~n42857 & n42858 ) ;
  assign n42860 = n12313 & n26754 ;
  assign n42861 = n32149 ^ n7738 ^ n821 ;
  assign n42862 = n42861 ^ n33926 ^ 1'b0 ;
  assign n42863 = ( n5121 & n6476 ) | ( n5121 & n12520 ) | ( n6476 & n12520 ) ;
  assign n42864 = n42863 ^ n42170 ^ n3976 ;
  assign n42865 = n5803 ^ n805 ^ 1'b0 ;
  assign n42866 = ( n28449 & ~n31226 ) | ( n28449 & n42865 ) | ( ~n31226 & n42865 ) ;
  assign n42867 = ( n2113 & n5658 ) | ( n2113 & ~n22798 ) | ( n5658 & ~n22798 ) ;
  assign n42868 = n38213 ^ n27215 ^ n11591 ;
  assign n42869 = n42867 & n42868 ;
  assign n42870 = n33797 ^ n17471 ^ n11942 ;
  assign n42871 = n42870 ^ n16968 ^ n6312 ;
  assign n42872 = n20843 & n42871 ;
  assign n42873 = n42872 ^ n21774 ^ 1'b0 ;
  assign n42874 = n10928 ^ n8867 ^ 1'b0 ;
  assign n42875 = n35014 ^ n3802 ^ 1'b0 ;
  assign n42876 = n32422 | n42875 ;
  assign n42877 = n25619 ^ n23729 ^ n6592 ;
  assign n42878 = ( n7295 & n10191 ) | ( n7295 & n42877 ) | ( n10191 & n42877 ) ;
  assign n42879 = ( ~n7965 & n41783 ) | ( ~n7965 & n42878 ) | ( n41783 & n42878 ) ;
  assign n42880 = n11319 & ~n27232 ;
  assign n42881 = n648 & n4048 ;
  assign n42882 = n42881 ^ n21321 ^ 1'b0 ;
  assign n42883 = n3908 & ~n13521 ;
  assign n42884 = n35787 & n42883 ;
  assign n42885 = ( n31314 & n42882 ) | ( n31314 & n42884 ) | ( n42882 & n42884 ) ;
  assign n42886 = n31954 ^ n22858 ^ 1'b0 ;
  assign n42887 = ~n7300 & n15356 ;
  assign n42888 = ~n12851 & n42887 ;
  assign n42889 = n42888 ^ n29194 ^ 1'b0 ;
  assign n42890 = n14432 | n28714 ;
  assign n42891 = n3507 & ~n42890 ;
  assign n42892 = ( n16098 & n31637 ) | ( n16098 & n32916 ) | ( n31637 & n32916 ) ;
  assign n42893 = n42891 | n42892 ;
  assign n42894 = n42893 ^ n29578 ^ 1'b0 ;
  assign n42895 = n25775 | n42894 ;
  assign n42896 = n42895 ^ n36316 ^ 1'b0 ;
  assign n42897 = ( n4701 & ~n30021 ) | ( n4701 & n35170 ) | ( ~n30021 & n35170 ) ;
  assign n42898 = n32359 ^ n26265 ^ n9495 ;
  assign n42899 = ( n29150 & n42897 ) | ( n29150 & n42898 ) | ( n42897 & n42898 ) ;
  assign n42902 = ( n21446 & n27690 ) | ( n21446 & ~n36637 ) | ( n27690 & ~n36637 ) ;
  assign n42900 = n6896 & ~n36834 ;
  assign n42901 = ( n653 & n9694 ) | ( n653 & ~n42900 ) | ( n9694 & ~n42900 ) ;
  assign n42903 = n42902 ^ n42901 ^ n39864 ;
  assign n42904 = n20816 ^ n5529 ^ n542 ;
  assign n42905 = n24346 ^ n21799 ^ 1'b0 ;
  assign n42906 = ( n12508 & ~n22441 ) | ( n12508 & n42905 ) | ( ~n22441 & n42905 ) ;
  assign n42907 = n31736 ^ n11383 ^ n2510 ;
  assign n42908 = n42907 ^ n33723 ^ n32035 ;
  assign n42909 = ~n39573 & n42908 ;
  assign n42910 = n36647 ^ n20735 ^ 1'b0 ;
  assign n42911 = n15226 & n42910 ;
  assign n42912 = ( n10109 & n32339 ) | ( n10109 & ~n42911 ) | ( n32339 & ~n42911 ) ;
  assign n42913 = n25130 & ~n30162 ;
  assign n42914 = ( ~n14850 & n38611 ) | ( ~n14850 & n42913 ) | ( n38611 & n42913 ) ;
  assign n42915 = ( n3205 & n42912 ) | ( n3205 & n42914 ) | ( n42912 & n42914 ) ;
  assign n42916 = ( n18924 & n20372 ) | ( n18924 & ~n37262 ) | ( n20372 & ~n37262 ) ;
  assign n42917 = n16616 ^ n15815 ^ n6441 ;
  assign n42918 = n12354 | n21097 ;
  assign n42919 = n42918 ^ n36734 ^ 1'b0 ;
  assign n42920 = n42445 ^ n15755 ^ n5654 ;
  assign n42921 = ( n4883 & n7955 ) | ( n4883 & n17633 ) | ( n7955 & n17633 ) ;
  assign n42923 = n25626 ^ n10999 ^ 1'b0 ;
  assign n42922 = n24421 ^ n18616 ^ n15900 ;
  assign n42924 = n42923 ^ n42922 ^ x202 ;
  assign n42925 = ( n1476 & ~n14915 ) | ( n1476 & n26198 ) | ( ~n14915 & n26198 ) ;
  assign n42926 = n42925 ^ n1184 ^ 1'b0 ;
  assign n42927 = n11565 ^ n1252 ^ 1'b0 ;
  assign n42928 = n2004 | n42927 ;
  assign n42929 = n15058 ^ n5525 ^ 1'b0 ;
  assign n42930 = n42928 | n42929 ;
  assign n42931 = ( n1710 & n20972 ) | ( n1710 & ~n30510 ) | ( n20972 & ~n30510 ) ;
  assign n42932 = ( n31311 & ~n32149 ) | ( n31311 & n42931 ) | ( ~n32149 & n42931 ) ;
  assign n42933 = n42932 ^ n21884 ^ n19380 ;
  assign n42934 = n28299 ^ n6697 ^ 1'b0 ;
  assign n42935 = n24933 & n42934 ;
  assign n42936 = n42935 ^ n17745 ^ 1'b0 ;
  assign n42938 = n22576 ^ n4922 ^ 1'b0 ;
  assign n42939 = n15097 | n42938 ;
  assign n42937 = ( n23378 & n25450 ) | ( n23378 & ~n36957 ) | ( n25450 & ~n36957 ) ;
  assign n42940 = n42939 ^ n42937 ^ n19381 ;
  assign n42941 = ( ~n17127 & n29283 ) | ( ~n17127 & n39483 ) | ( n29283 & n39483 ) ;
  assign n42948 = n16527 ^ n2037 ^ 1'b0 ;
  assign n42944 = n7485 & ~n22977 ;
  assign n42945 = ~n1304 & n42944 ;
  assign n42942 = n8260 & ~n25348 ;
  assign n42943 = n42942 ^ n11972 ^ 1'b0 ;
  assign n42946 = n42945 ^ n42943 ^ n1212 ;
  assign n42947 = ( n916 & n30964 ) | ( n916 & n42946 ) | ( n30964 & n42946 ) ;
  assign n42949 = n42948 ^ n42947 ^ n28238 ;
  assign n42953 = n15944 ^ n5251 ^ x156 ;
  assign n42954 = n42953 ^ n1724 ^ 1'b0 ;
  assign n42952 = n12102 ^ n11114 ^ n7797 ;
  assign n42950 = n14160 ^ n11936 ^ n8881 ;
  assign n42951 = n42950 ^ n18539 ^ n1905 ;
  assign n42955 = n42954 ^ n42952 ^ n42951 ;
  assign n42956 = ( n13887 & n34579 ) | ( n13887 & n34637 ) | ( n34579 & n34637 ) ;
  assign n42957 = n42956 ^ n36096 ^ n10167 ;
  assign n42958 = n21894 & ~n28403 ;
  assign n42959 = n2401 | n42958 ;
  assign n42960 = n10297 ^ n5447 ^ 1'b0 ;
  assign n42961 = n12230 ^ n3794 ^ n3354 ;
  assign n42962 = n20781 & ~n42961 ;
  assign n42963 = n42962 ^ n10959 ^ 1'b0 ;
  assign n42967 = n12273 ^ n5306 ^ n1915 ;
  assign n42968 = n33856 ^ n12482 ^ 1'b0 ;
  assign n42969 = n42967 | n42968 ;
  assign n42964 = n10534 & n19748 ;
  assign n42965 = n12721 & n42964 ;
  assign n42966 = n3335 & ~n42965 ;
  assign n42970 = n42969 ^ n42966 ^ 1'b0 ;
  assign n42971 = ~n42963 & n42970 ;
  assign n42972 = ~n33095 & n42971 ;
  assign n42973 = n42972 ^ n19543 ^ n18752 ;
  assign n42974 = ~n10903 & n31646 ;
  assign n42975 = n3862 & n42974 ;
  assign n42976 = n42975 ^ n13680 ^ n10404 ;
  assign n42977 = n23474 ^ n12221 ^ n6838 ;
  assign n42978 = n14937 & ~n37211 ;
  assign n42979 = n42978 ^ n17623 ^ 1'b0 ;
  assign n42980 = ( n4018 & n14727 ) | ( n4018 & ~n42979 ) | ( n14727 & ~n42979 ) ;
  assign n42981 = n34845 ^ n27989 ^ 1'b0 ;
  assign n42982 = n42981 ^ n26884 ^ n6661 ;
  assign n42992 = n15998 ^ n14910 ^ n1065 ;
  assign n42983 = ( n9472 & n14517 ) | ( n9472 & ~n27250 ) | ( n14517 & ~n27250 ) ;
  assign n42984 = n42983 ^ n27087 ^ n10979 ;
  assign n42985 = n22240 | n42984 ;
  assign n42986 = n2108 & ~n42985 ;
  assign n42987 = n2640 & ~n42986 ;
  assign n42988 = n17944 & n42987 ;
  assign n42989 = n42458 | n42988 ;
  assign n42990 = n2962 | n42989 ;
  assign n42991 = n10959 | n42990 ;
  assign n42993 = n42992 ^ n42991 ^ n17266 ;
  assign n42994 = ( n11968 & ~n12984 ) | ( n11968 & n23602 ) | ( ~n12984 & n23602 ) ;
  assign n42995 = n9659 ^ n6445 ^ 1'b0 ;
  assign n42996 = n42994 | n42995 ;
  assign n42997 = ( n14680 & n36649 ) | ( n14680 & ~n42996 ) | ( n36649 & ~n42996 ) ;
  assign n42998 = n2309 & n3700 ;
  assign n42999 = ~n19528 & n42998 ;
  assign n43000 = n7116 & ~n42999 ;
  assign n43002 = n13568 ^ n6397 ^ x87 ;
  assign n43003 = ( n4426 & n25660 ) | ( n4426 & ~n43002 ) | ( n25660 & ~n43002 ) ;
  assign n43001 = ~n21651 & n30648 ;
  assign n43004 = n43003 ^ n43001 ^ 1'b0 ;
  assign n43005 = ( n30606 & ~n35333 ) | ( n30606 & n42144 ) | ( ~n35333 & n42144 ) ;
  assign n43006 = n20341 ^ n10398 ^ 1'b0 ;
  assign n43007 = n27682 ^ n10977 ^ n7890 ;
  assign n43008 = ( n12620 & n14527 ) | ( n12620 & ~n34306 ) | ( n14527 & ~n34306 ) ;
  assign n43009 = n43008 ^ n12749 ^ n1821 ;
  assign n43010 = n43009 ^ n26919 ^ 1'b0 ;
  assign n43011 = ( ~n6166 & n17551 ) | ( ~n6166 & n27934 ) | ( n17551 & n27934 ) ;
  assign n43012 = ( n7327 & n12693 ) | ( n7327 & ~n41791 ) | ( n12693 & ~n41791 ) ;
  assign n43013 = n26789 & n43012 ;
  assign n43014 = ( n432 & n18283 ) | ( n432 & n28520 ) | ( n18283 & n28520 ) ;
  assign n43015 = n565 & n3167 ;
  assign n43016 = n43014 & n43015 ;
  assign n43017 = n43016 ^ n31790 ^ 1'b0 ;
  assign n43018 = n15865 ^ n2265 ^ 1'b0 ;
  assign n43019 = n43018 ^ n5211 ^ 1'b0 ;
  assign n43020 = n626 & ~n43019 ;
  assign n43021 = ( ~n3825 & n43017 ) | ( ~n3825 & n43020 ) | ( n43017 & n43020 ) ;
  assign n43022 = n14977 ^ n12826 ^ 1'b0 ;
  assign n43023 = n19552 & n43022 ;
  assign n43024 = ~n27386 & n39627 ;
  assign n43025 = ~n43023 & n43024 ;
  assign n43026 = n11370 ^ n7649 ^ 1'b0 ;
  assign n43027 = ( x3 & n19449 ) | ( x3 & ~n34878 ) | ( n19449 & ~n34878 ) ;
  assign n43028 = ( n17862 & ~n43026 ) | ( n17862 & n43027 ) | ( ~n43026 & n43027 ) ;
  assign n43029 = n43028 ^ n23444 ^ n11029 ;
  assign n43030 = n15579 ^ n2286 ^ 1'b0 ;
  assign n43031 = ~n15058 & n43030 ;
  assign n43032 = ( ~n3095 & n23774 ) | ( ~n3095 & n43031 ) | ( n23774 & n43031 ) ;
  assign n43033 = n43029 & n43032 ;
  assign n43034 = n21086 ^ n20437 ^ n16149 ;
  assign n43035 = n43034 ^ n23643 ^ n21829 ;
  assign n43036 = n43035 ^ n24674 ^ n10136 ;
  assign n43037 = n43036 ^ n38164 ^ n30045 ;
  assign n43038 = ~n1560 & n38680 ;
  assign n43039 = n43038 ^ n7510 ^ n5255 ;
  assign n43040 = n4478 ^ n3514 ^ 1'b0 ;
  assign n43041 = ( n23956 & n43039 ) | ( n23956 & ~n43040 ) | ( n43039 & ~n43040 ) ;
  assign n43042 = n4858 & n29573 ;
  assign n43043 = n43042 ^ n26247 ^ 1'b0 ;
  assign n43044 = ( n25429 & n28304 ) | ( n25429 & ~n43043 ) | ( n28304 & ~n43043 ) ;
  assign n43045 = n34625 ^ n3374 ^ 1'b0 ;
  assign n43046 = n3337 | n43045 ;
  assign n43047 = ( n15689 & n42956 ) | ( n15689 & n43046 ) | ( n42956 & n43046 ) ;
  assign n43048 = ~n9875 & n33220 ;
  assign n43049 = n43048 ^ n10562 ^ 1'b0 ;
  assign n43050 = n366 & ~n21582 ;
  assign n43051 = ~n18905 & n43050 ;
  assign n43052 = ( n6999 & ~n15222 ) | ( n6999 & n43051 ) | ( ~n15222 & n43051 ) ;
  assign n43053 = n39952 | n43052 ;
  assign n43054 = n43053 ^ n11324 ^ 1'b0 ;
  assign n43055 = n10328 ^ n5090 ^ n3908 ;
  assign n43056 = n43055 ^ n37627 ^ 1'b0 ;
  assign n43057 = n11114 ^ n1445 ^ 1'b0 ;
  assign n43058 = ( n4009 & n6973 ) | ( n4009 & n36559 ) | ( n6973 & n36559 ) ;
  assign n43059 = ( n1023 & ~n39237 ) | ( n1023 & n43058 ) | ( ~n39237 & n43058 ) ;
  assign n43060 = ( ~n486 & n4196 ) | ( ~n486 & n24947 ) | ( n4196 & n24947 ) ;
  assign n43061 = ( ~n7039 & n7972 ) | ( ~n7039 & n43060 ) | ( n7972 & n43060 ) ;
  assign n43062 = n24847 ^ n12262 ^ n4079 ;
  assign n43063 = ( n1849 & n10310 ) | ( n1849 & ~n43062 ) | ( n10310 & ~n43062 ) ;
  assign n43064 = n42560 ^ n15866 ^ n1857 ;
  assign n43065 = ( n19927 & n20816 ) | ( n19927 & ~n22946 ) | ( n20816 & ~n22946 ) ;
  assign n43066 = n43065 ^ n37803 ^ 1'b0 ;
  assign n43067 = n30957 & ~n43066 ;
  assign n43068 = n41222 ^ n34631 ^ 1'b0 ;
  assign n43069 = n30877 | n43068 ;
  assign n43070 = n43069 ^ n30008 ^ 1'b0 ;
  assign n43077 = n20904 ^ n12480 ^ n3147 ;
  assign n43072 = ( n736 & ~n5601 ) | ( n736 & n12638 ) | ( ~n5601 & n12638 ) ;
  assign n43073 = ( n5077 & ~n26351 ) | ( n5077 & n43072 ) | ( ~n26351 & n43072 ) ;
  assign n43071 = n7064 ^ n4963 ^ 1'b0 ;
  assign n43074 = n43073 ^ n43071 ^ n22724 ;
  assign n43075 = n43074 ^ n10402 ^ 1'b0 ;
  assign n43076 = n26879 & ~n43075 ;
  assign n43078 = n43077 ^ n43076 ^ n26452 ;
  assign n43079 = ( n33593 & n42080 ) | ( n33593 & n43078 ) | ( n42080 & n43078 ) ;
  assign n43080 = n28106 ^ n11455 ^ 1'b0 ;
  assign n43081 = n21916 ^ n18231 ^ n12159 ;
  assign n43082 = n43081 ^ n24377 ^ 1'b0 ;
  assign n43083 = ( ~n43079 & n43080 ) | ( ~n43079 & n43082 ) | ( n43080 & n43082 ) ;
  assign n43084 = ~n14936 & n17431 ;
  assign n43085 = ( n14159 & ~n42024 ) | ( n14159 & n43084 ) | ( ~n42024 & n43084 ) ;
  assign n43086 = ( n5537 & n7849 ) | ( n5537 & ~n31467 ) | ( n7849 & ~n31467 ) ;
  assign n43087 = n43086 ^ n42231 ^ n21768 ;
  assign n43088 = n15834 ^ n15762 ^ n12694 ;
  assign n43089 = n43088 ^ n12853 ^ 1'b0 ;
  assign n43090 = n34004 & n43089 ;
  assign n43091 = ~n4002 & n43090 ;
  assign n43092 = n30250 ^ n10662 ^ 1'b0 ;
  assign n43093 = n25255 | n43092 ;
  assign n43094 = ( n492 & n6345 ) | ( n492 & n22758 ) | ( n6345 & n22758 ) ;
  assign n43095 = ( n14902 & n15592 ) | ( n14902 & ~n30049 ) | ( n15592 & ~n30049 ) ;
  assign n43096 = ( n21448 & ~n30890 ) | ( n21448 & n43095 ) | ( ~n30890 & n43095 ) ;
  assign n43097 = n43096 ^ n5653 ^ 1'b0 ;
  assign n43098 = ( n10274 & n43094 ) | ( n10274 & n43097 ) | ( n43094 & n43097 ) ;
  assign n43099 = n14596 ^ n12066 ^ n5601 ;
  assign n43100 = n43099 ^ n15115 ^ n9966 ;
  assign n43101 = ( n1056 & n4973 ) | ( n1056 & ~n26634 ) | ( n4973 & ~n26634 ) ;
  assign n43102 = n36624 ^ n927 ^ 1'b0 ;
  assign n43107 = n14937 ^ n6252 ^ n348 ;
  assign n43103 = ( ~n970 & n3620 ) | ( ~n970 & n9348 ) | ( n3620 & n9348 ) ;
  assign n43104 = ( n7493 & ~n11865 ) | ( n7493 & n43103 ) | ( ~n11865 & n43103 ) ;
  assign n43105 = n43104 ^ n27345 ^ n26031 ;
  assign n43106 = ~n26749 & n43105 ;
  assign n43108 = n43107 ^ n43106 ^ 1'b0 ;
  assign n43109 = ( n15896 & ~n18438 ) | ( n15896 & n43108 ) | ( ~n18438 & n43108 ) ;
  assign n43110 = ( ~n2239 & n34209 ) | ( ~n2239 & n37616 ) | ( n34209 & n37616 ) ;
  assign n43111 = n29151 ^ n20001 ^ n4117 ;
  assign n43113 = n30033 ^ n9236 ^ n6454 ;
  assign n43112 = ( n7026 & ~n17448 ) | ( n7026 & n18426 ) | ( ~n17448 & n18426 ) ;
  assign n43114 = n43113 ^ n43112 ^ 1'b0 ;
  assign n43115 = ( n36209 & ~n43111 ) | ( n36209 & n43114 ) | ( ~n43111 & n43114 ) ;
  assign n43116 = ( n8020 & n21711 ) | ( n8020 & n41481 ) | ( n21711 & n41481 ) ;
  assign n43117 = n16607 | n43116 ;
  assign n43118 = n43115 | n43117 ;
  assign n43121 = ( n1410 & n2073 ) | ( n1410 & ~n9662 ) | ( n2073 & ~n9662 ) ;
  assign n43119 = n25872 ^ n18361 ^ 1'b0 ;
  assign n43120 = ~n35321 & n43119 ;
  assign n43122 = n43121 ^ n43120 ^ 1'b0 ;
  assign n43123 = n21209 & ~n43122 ;
  assign n43124 = n26322 ^ n18447 ^ n8687 ;
  assign n43125 = ~n6354 & n43124 ;
  assign n43126 = n34014 ^ n1476 ^ 1'b0 ;
  assign n43127 = n20574 & ~n43126 ;
  assign n43128 = n43127 ^ n27890 ^ 1'b0 ;
  assign n43129 = ( ~n26002 & n31912 ) | ( ~n26002 & n43128 ) | ( n31912 & n43128 ) ;
  assign n43130 = n23251 ^ n14791 ^ 1'b0 ;
  assign n43131 = n5496 | n24480 ;
  assign n43132 = n35113 | n43131 ;
  assign n43133 = ( ~n35010 & n43130 ) | ( ~n35010 & n43132 ) | ( n43130 & n43132 ) ;
  assign n43134 = n12694 ^ n8668 ^ n4729 ;
  assign n43135 = n43134 ^ n30869 ^ n22784 ;
  assign n43136 = ( ~n1760 & n4412 ) | ( ~n1760 & n29589 ) | ( n4412 & n29589 ) ;
  assign n43137 = n43136 ^ n40722 ^ n7280 ;
  assign n43138 = n5377 | n6719 ;
  assign n43139 = n43138 ^ n17291 ^ 1'b0 ;
  assign n43140 = n4773 | n19683 ;
  assign n43141 = n10138 | n43140 ;
  assign n43142 = n34256 ^ n14181 ^ n9480 ;
  assign n43143 = n43141 & ~n43142 ;
  assign n43144 = ( ~n3877 & n10378 ) | ( ~n3877 & n12377 ) | ( n10378 & n12377 ) ;
  assign n43145 = n20283 & ~n43144 ;
  assign n43146 = n43145 ^ n12344 ^ 1'b0 ;
  assign n43147 = n11457 ^ n8486 ^ 1'b0 ;
  assign n43148 = n16221 & n43147 ;
  assign n43149 = n43148 ^ n31930 ^ 1'b0 ;
  assign n43150 = n43149 ^ n12376 ^ n4295 ;
  assign n43151 = n43150 ^ n28510 ^ n14133 ;
  assign n43152 = n7398 & n31625 ;
  assign n43153 = n43152 ^ n18055 ^ 1'b0 ;
  assign n43154 = ( n12890 & ~n40620 ) | ( n12890 & n43153 ) | ( ~n40620 & n43153 ) ;
  assign n43155 = n10811 & n11413 ;
  assign n43156 = n43155 ^ n31661 ^ n26891 ;
  assign n43157 = n40374 ^ n36979 ^ 1'b0 ;
  assign n43159 = n17614 ^ n8920 ^ x39 ;
  assign n43158 = ( n4538 & n17553 ) | ( n4538 & n23702 ) | ( n17553 & n23702 ) ;
  assign n43160 = n43159 ^ n43158 ^ n601 ;
  assign n43161 = n43160 ^ n37665 ^ n671 ;
  assign n43162 = n43161 ^ n22987 ^ 1'b0 ;
  assign n43163 = n33748 ^ n4301 ^ n1313 ;
  assign n43164 = n5673 & n42605 ;
  assign n43165 = ~n43163 & n43164 ;
  assign n43166 = n10253 & n34133 ;
  assign n43167 = ( n5482 & n37456 ) | ( n5482 & n43166 ) | ( n37456 & n43166 ) ;
  assign n43168 = ( ~n7089 & n16016 ) | ( ~n7089 & n26880 ) | ( n16016 & n26880 ) ;
  assign n43169 = x22 & n28577 ;
  assign n43170 = ( ~n2711 & n19915 ) | ( ~n2711 & n35793 ) | ( n19915 & n35793 ) ;
  assign n43171 = ( n6824 & ~n17460 ) | ( n6824 & n20317 ) | ( ~n17460 & n20317 ) ;
  assign n43172 = n43171 ^ n20267 ^ n11702 ;
  assign n43177 = n24061 ^ n5660 ^ n2679 ;
  assign n43175 = ( n21065 & n30563 ) | ( n21065 & n35022 ) | ( n30563 & n35022 ) ;
  assign n43176 = n43175 ^ n21158 ^ n10459 ;
  assign n43173 = ( n16493 & n34909 ) | ( n16493 & n36767 ) | ( n34909 & n36767 ) ;
  assign n43174 = n43173 ^ n22436 ^ n19888 ;
  assign n43178 = n43177 ^ n43176 ^ n43174 ;
  assign n43180 = ( ~n2881 & n4599 ) | ( ~n2881 & n21933 ) | ( n4599 & n21933 ) ;
  assign n43181 = ( n4181 & n38590 ) | ( n4181 & n43180 ) | ( n38590 & n43180 ) ;
  assign n43179 = ~n24968 & n36176 ;
  assign n43182 = n43181 ^ n43179 ^ 1'b0 ;
  assign n43183 = n25645 & ~n35009 ;
  assign n43184 = n43183 ^ n22641 ^ 1'b0 ;
  assign n43185 = n28932 ^ n21168 ^ 1'b0 ;
  assign n43186 = n13880 | n43185 ;
  assign n43187 = ( n10785 & ~n21120 ) | ( n10785 & n24523 ) | ( ~n21120 & n24523 ) ;
  assign n43188 = ~n3072 & n30183 ;
  assign n43189 = ( n17604 & ~n28092 ) | ( n17604 & n43188 ) | ( ~n28092 & n43188 ) ;
  assign n43190 = n43189 ^ n25075 ^ n4907 ;
  assign n43191 = n43190 ^ n17611 ^ n12224 ;
  assign n43192 = n22764 ^ n10858 ^ n1796 ;
  assign n43193 = ( n6444 & n21957 ) | ( n6444 & n36559 ) | ( n21957 & n36559 ) ;
  assign n43194 = ( ~n4875 & n43192 ) | ( ~n4875 & n43193 ) | ( n43192 & n43193 ) ;
  assign n43195 = n43194 ^ n18517 ^ n5776 ;
  assign n43196 = n24142 ^ n16149 ^ n9535 ;
  assign n43197 = ( ~n7001 & n14167 ) | ( ~n7001 & n28031 ) | ( n14167 & n28031 ) ;
  assign n43198 = ~n12660 & n19932 ;
  assign n43199 = n43198 ^ n1329 ^ 1'b0 ;
  assign n43200 = ( ~n1483 & n4632 ) | ( ~n1483 & n43199 ) | ( n4632 & n43199 ) ;
  assign n43201 = ( n42509 & n43197 ) | ( n42509 & n43200 ) | ( n43197 & n43200 ) ;
  assign n43202 = ~n2711 & n4167 ;
  assign n43203 = ( ~n4843 & n24259 ) | ( ~n4843 & n43202 ) | ( n24259 & n43202 ) ;
  assign n43205 = n1560 & n42961 ;
  assign n43206 = n17895 & n43205 ;
  assign n43207 = n43206 ^ n28645 ^ n9121 ;
  assign n43204 = ( ~n9944 & n28229 ) | ( ~n9944 & n42935 ) | ( n28229 & n42935 ) ;
  assign n43208 = n43207 ^ n43204 ^ n34903 ;
  assign n43209 = ( n18113 & ~n26176 ) | ( n18113 & n42948 ) | ( ~n26176 & n42948 ) ;
  assign n43210 = n43209 ^ n30400 ^ n30223 ;
  assign n43211 = n41902 ^ n40934 ^ n35481 ;
  assign n43212 = n30093 ^ n15933 ^ 1'b0 ;
  assign n43213 = n11876 | n43212 ;
  assign n43214 = n43213 ^ n4765 ^ 1'b0 ;
  assign n43215 = ( n2538 & n10569 ) | ( n2538 & ~n29918 ) | ( n10569 & ~n29918 ) ;
  assign n43217 = n8743 ^ n7237 ^ n6327 ;
  assign n43218 = ( n13039 & n13908 ) | ( n13039 & n43217 ) | ( n13908 & n43217 ) ;
  assign n43216 = ( n850 & ~n20278 ) | ( n850 & n29501 ) | ( ~n20278 & n29501 ) ;
  assign n43219 = n43218 ^ n43216 ^ n39648 ;
  assign n43220 = ( n5718 & n33978 ) | ( n5718 & n43219 ) | ( n33978 & n43219 ) ;
  assign n43221 = ( n18596 & ~n33324 ) | ( n18596 & n43220 ) | ( ~n33324 & n43220 ) ;
  assign n43222 = n1264 & n40877 ;
  assign n43223 = n19109 & n43222 ;
  assign n43224 = n21315 ^ n13045 ^ 1'b0 ;
  assign n43225 = ( n12538 & ~n26903 ) | ( n12538 & n32443 ) | ( ~n26903 & n32443 ) ;
  assign n43229 = n18784 | n26979 ;
  assign n43230 = n6587 | n25909 ;
  assign n43231 = n18116 | n43230 ;
  assign n43232 = ( n10494 & n19383 ) | ( n10494 & n43231 ) | ( n19383 & n43231 ) ;
  assign n43233 = ( n5098 & n43229 ) | ( n5098 & ~n43232 ) | ( n43229 & ~n43232 ) ;
  assign n43226 = ( n15612 & n18117 ) | ( n15612 & ~n26586 ) | ( n18117 & ~n26586 ) ;
  assign n43227 = n43226 ^ n16847 ^ n7458 ;
  assign n43228 = n36216 & ~n43227 ;
  assign n43234 = n43233 ^ n43228 ^ 1'b0 ;
  assign n43235 = ( n5121 & n16626 ) | ( n5121 & ~n20344 ) | ( n16626 & ~n20344 ) ;
  assign n43236 = ( n13592 & n29234 ) | ( n13592 & ~n43235 ) | ( n29234 & ~n43235 ) ;
  assign n43237 = n10247 & ~n18621 ;
  assign n43238 = n38878 ^ n36738 ^ 1'b0 ;
  assign n43239 = ( ~n9872 & n19000 ) | ( ~n9872 & n43238 ) | ( n19000 & n43238 ) ;
  assign n43240 = ( ~n2176 & n10407 ) | ( ~n2176 & n18260 ) | ( n10407 & n18260 ) ;
  assign n43241 = n43240 ^ n27407 ^ 1'b0 ;
  assign n43242 = n43239 & ~n43241 ;
  assign n43243 = ( n5457 & n12107 ) | ( n5457 & ~n43242 ) | ( n12107 & ~n43242 ) ;
  assign n43244 = ( n6339 & n26877 ) | ( n6339 & ~n31184 ) | ( n26877 & ~n31184 ) ;
  assign n43245 = ~n2260 & n43244 ;
  assign n43246 = ( n3153 & ~n7858 ) | ( n3153 & n14999 ) | ( ~n7858 & n14999 ) ;
  assign n43247 = n12708 ^ n4098 ^ 1'b0 ;
  assign n43248 = ~n1205 & n43247 ;
  assign n43249 = n8378 ^ n6067 ^ 1'b0 ;
  assign n43250 = n27251 | n43249 ;
  assign n43251 = n43250 ^ n13694 ^ n9788 ;
  assign n43252 = n31538 ^ n28891 ^ n9981 ;
  assign n43253 = n11229 & ~n43252 ;
  assign n43254 = n30563 ^ n20398 ^ n19256 ;
  assign n43255 = ( ~n3942 & n13668 ) | ( ~n3942 & n13983 ) | ( n13668 & n13983 ) ;
  assign n43256 = n27611 ^ n8963 ^ n1857 ;
  assign n43257 = ( ~n33775 & n43255 ) | ( ~n33775 & n43256 ) | ( n43255 & n43256 ) ;
  assign n43258 = n43257 ^ n31756 ^ n24945 ;
  assign n43260 = ( n2950 & n12525 ) | ( n2950 & ~n13778 ) | ( n12525 & ~n13778 ) ;
  assign n43259 = n14275 ^ n11634 ^ n7856 ;
  assign n43261 = n43260 ^ n43259 ^ n35438 ;
  assign n43262 = n43261 ^ n7970 ^ n6423 ;
  assign n43263 = n43262 ^ n26424 ^ 1'b0 ;
  assign n43264 = n13909 | n43263 ;
  assign n43265 = ( n7144 & n35957 ) | ( n7144 & ~n43264 ) | ( n35957 & ~n43264 ) ;
  assign n43266 = ( ~n12533 & n17149 ) | ( ~n12533 & n38898 ) | ( n17149 & n38898 ) ;
  assign n43267 = ( ~n3921 & n12532 ) | ( ~n3921 & n43266 ) | ( n12532 & n43266 ) ;
  assign n43268 = ( n3368 & n8919 ) | ( n3368 & n16030 ) | ( n8919 & n16030 ) ;
  assign n43269 = n6489 & ~n24772 ;
  assign n43270 = ~n43268 & n43269 ;
  assign n43271 = ( ~n956 & n21965 ) | ( ~n956 & n43270 ) | ( n21965 & n43270 ) ;
  assign n43272 = n40700 ^ n8925 ^ 1'b0 ;
  assign n43273 = n43271 & ~n43272 ;
  assign n43274 = ( ~n8720 & n41219 ) | ( ~n8720 & n43273 ) | ( n41219 & n43273 ) ;
  assign n43275 = n29000 ^ n1707 ^ 1'b0 ;
  assign n43276 = ~n28318 & n43275 ;
  assign n43277 = n43276 ^ n36779 ^ 1'b0 ;
  assign n43278 = n43274 | n43277 ;
  assign n43279 = ( ~n7141 & n25530 ) | ( ~n7141 & n32209 ) | ( n25530 & n32209 ) ;
  assign n43280 = n10557 & n43279 ;
  assign n43282 = ( n272 & ~n13468 ) | ( n272 & n21049 ) | ( ~n13468 & n21049 ) ;
  assign n43281 = n37721 ^ n31014 ^ n3278 ;
  assign n43283 = n43282 ^ n43281 ^ n17106 ;
  assign n43284 = n5697 ^ n4143 ^ 1'b0 ;
  assign n43285 = n6861 & n43284 ;
  assign n43286 = ( n20811 & n26220 ) | ( n20811 & n43285 ) | ( n26220 & n43285 ) ;
  assign n43287 = ( n2806 & n14449 ) | ( n2806 & ~n22024 ) | ( n14449 & ~n22024 ) ;
  assign n43288 = n1575 & ~n14014 ;
  assign n43289 = n43288 ^ n14253 ^ 1'b0 ;
  assign n43290 = ( n15848 & n43287 ) | ( n15848 & n43289 ) | ( n43287 & n43289 ) ;
  assign n43291 = n43290 ^ n34572 ^ n1216 ;
  assign n43292 = n12899 & ~n29455 ;
  assign n43295 = n17474 ^ n14274 ^ n1871 ;
  assign n43296 = ( n6868 & n17363 ) | ( n6868 & ~n43295 ) | ( n17363 & ~n43295 ) ;
  assign n43293 = n42150 ^ n18490 ^ 1'b0 ;
  assign n43294 = n30519 & ~n43293 ;
  assign n43297 = n43296 ^ n43294 ^ n31226 ;
  assign n43298 = n43297 ^ n8045 ^ 1'b0 ;
  assign n43299 = n16672 & n43298 ;
  assign n43300 = ( ~n5875 & n43292 ) | ( ~n5875 & n43299 ) | ( n43292 & n43299 ) ;
  assign n43301 = n7830 & ~n39103 ;
  assign n43302 = n11548 & n43301 ;
  assign n43303 = ( ~n28766 & n29190 ) | ( ~n28766 & n43302 ) | ( n29190 & n43302 ) ;
  assign n43304 = ( n2721 & ~n9278 ) | ( n2721 & n23635 ) | ( ~n9278 & n23635 ) ;
  assign n43305 = n934 & ~n38139 ;
  assign n43306 = ~n8615 & n43305 ;
  assign n43307 = n29566 ^ n15575 ^ 1'b0 ;
  assign n43308 = ( n17028 & ~n28179 ) | ( n17028 & n32612 ) | ( ~n28179 & n32612 ) ;
  assign n43309 = ~n1663 & n9302 ;
  assign n43310 = ( n11513 & ~n39501 ) | ( n11513 & n43309 ) | ( ~n39501 & n43309 ) ;
  assign n43311 = ( ~n19342 & n35229 ) | ( ~n19342 & n37845 ) | ( n35229 & n37845 ) ;
  assign n43312 = ~n17041 & n43311 ;
  assign n43313 = ( n11624 & n43310 ) | ( n11624 & n43312 ) | ( n43310 & n43312 ) ;
  assign n43314 = n41322 ^ n35386 ^ n16797 ;
  assign n43315 = ( n7204 & n27713 ) | ( n7204 & ~n29619 ) | ( n27713 & ~n29619 ) ;
  assign n43316 = ( n7430 & ~n27777 ) | ( n7430 & n43315 ) | ( ~n27777 & n43315 ) ;
  assign n43317 = n32995 ^ n30391 ^ n27357 ;
  assign n43318 = n22682 ^ n3506 ^ 1'b0 ;
  assign n43319 = n7780 | n43318 ;
  assign n43320 = ( n8858 & ~n10070 ) | ( n8858 & n11251 ) | ( ~n10070 & n11251 ) ;
  assign n43321 = ( n1411 & n13571 ) | ( n1411 & n43320 ) | ( n13571 & n43320 ) ;
  assign n43322 = n43321 ^ n21950 ^ 1'b0 ;
  assign n43323 = ( n8464 & n23017 ) | ( n8464 & ~n43322 ) | ( n23017 & ~n43322 ) ;
  assign n43324 = ( n6482 & n8807 ) | ( n6482 & ~n37976 ) | ( n8807 & ~n37976 ) ;
  assign n43325 = ( x57 & n5660 ) | ( x57 & n13014 ) | ( n5660 & n13014 ) ;
  assign n43326 = ( n7206 & ~n24472 ) | ( n7206 & n43325 ) | ( ~n24472 & n43325 ) ;
  assign n43327 = n12059 ^ n8904 ^ 1'b0 ;
  assign n43328 = ( n335 & n2296 ) | ( n335 & n27221 ) | ( n2296 & n27221 ) ;
  assign n43329 = ( n17025 & n34294 ) | ( n17025 & n43328 ) | ( n34294 & n43328 ) ;
  assign n43330 = ( n38601 & n43327 ) | ( n38601 & n43329 ) | ( n43327 & n43329 ) ;
  assign n43331 = ( ~n1590 & n6013 ) | ( ~n1590 & n7588 ) | ( n6013 & n7588 ) ;
  assign n43332 = ( n7941 & ~n19021 ) | ( n7941 & n43331 ) | ( ~n19021 & n43331 ) ;
  assign n43333 = n32540 & ~n43332 ;
  assign n43335 = ( x190 & n4533 ) | ( x190 & ~n12985 ) | ( n4533 & ~n12985 ) ;
  assign n43334 = n16020 & ~n41294 ;
  assign n43336 = n43335 ^ n43334 ^ n16738 ;
  assign n43337 = n25590 ^ n14133 ^ n11846 ;
  assign n43338 = n3131 & n6106 ;
  assign n43339 = n28393 ^ n21124 ^ 1'b0 ;
  assign n43340 = ~n2000 & n43339 ;
  assign n43341 = n27117 ^ n22854 ^ n14433 ;
  assign n43342 = ( n19451 & n35253 ) | ( n19451 & ~n39467 ) | ( n35253 & ~n39467 ) ;
  assign n43343 = ( n15848 & n19133 ) | ( n15848 & ~n23470 ) | ( n19133 & ~n23470 ) ;
  assign n43344 = n43343 ^ n2912 ^ 1'b0 ;
  assign n43345 = ( n37321 & n39016 ) | ( n37321 & ~n41071 ) | ( n39016 & ~n41071 ) ;
  assign n43346 = ~n13017 & n42244 ;
  assign n43348 = n12883 | n16940 ;
  assign n43349 = n43348 ^ n15708 ^ 1'b0 ;
  assign n43347 = n27355 & ~n27673 ;
  assign n43350 = n43349 ^ n43347 ^ 1'b0 ;
  assign n43351 = n43350 ^ n33055 ^ n15020 ;
  assign n43352 = ( n1471 & ~n3682 ) | ( n1471 & n14048 ) | ( ~n3682 & n14048 ) ;
  assign n43353 = n10307 ^ n9484 ^ n8348 ;
  assign n43354 = n43353 ^ n23808 ^ 1'b0 ;
  assign n43355 = n43352 | n43354 ;
  assign n43356 = ( n869 & n1715 ) | ( n869 & n26362 ) | ( n1715 & n26362 ) ;
  assign n43357 = n19979 | n43356 ;
  assign n43358 = n2517 | n43357 ;
  assign n43360 = n11893 | n12278 ;
  assign n43361 = n43360 ^ n9715 ^ 1'b0 ;
  assign n43359 = n36603 ^ n29264 ^ n2696 ;
  assign n43362 = n43361 ^ n43359 ^ 1'b0 ;
  assign n43363 = n26256 ^ n24795 ^ n828 ;
  assign n43364 = n6502 & n30546 ;
  assign n43365 = n43364 ^ n15010 ^ 1'b0 ;
  assign n43366 = n42954 | n43365 ;
  assign n43367 = n41748 & ~n43366 ;
  assign n43368 = n43367 ^ n27456 ^ n20248 ;
  assign n43369 = ( n10228 & n43363 ) | ( n10228 & ~n43368 ) | ( n43363 & ~n43368 ) ;
  assign n43370 = n27338 ^ n11465 ^ n276 ;
  assign n43371 = ( ~n2474 & n7445 ) | ( ~n2474 & n13938 ) | ( n7445 & n13938 ) ;
  assign n43372 = ( ~n3547 & n12927 ) | ( ~n3547 & n43371 ) | ( n12927 & n43371 ) ;
  assign n43373 = n43372 ^ n30638 ^ 1'b0 ;
  assign n43374 = n36969 ^ n30579 ^ 1'b0 ;
  assign n43376 = n37477 ^ n30462 ^ n9067 ;
  assign n43375 = n23209 & n32377 ;
  assign n43377 = n43376 ^ n43375 ^ 1'b0 ;
  assign n43378 = n2098 & ~n18898 ;
  assign n43379 = n32216 & n43378 ;
  assign n43380 = n41712 & ~n43379 ;
  assign n43381 = ~n33570 & n43380 ;
  assign n43382 = ( ~n19574 & n43377 ) | ( ~n19574 & n43381 ) | ( n43377 & n43381 ) ;
  assign n43383 = n7281 | n26059 ;
  assign n43384 = n43383 ^ n19452 ^ 1'b0 ;
  assign n43385 = n12541 ^ n4784 ^ 1'b0 ;
  assign n43388 = n25283 ^ n17180 ^ n4489 ;
  assign n43386 = n24449 ^ n10476 ^ 1'b0 ;
  assign n43387 = ( ~n850 & n7614 ) | ( ~n850 & n43386 ) | ( n7614 & n43386 ) ;
  assign n43389 = n43388 ^ n43387 ^ n1335 ;
  assign n43390 = ( ~n9942 & n25486 ) | ( ~n9942 & n43389 ) | ( n25486 & n43389 ) ;
  assign n43391 = n43390 ^ n22929 ^ 1'b0 ;
  assign n43392 = ~n43385 & n43391 ;
  assign n43394 = ( n2483 & n7236 ) | ( n2483 & ~n36987 ) | ( n7236 & ~n36987 ) ;
  assign n43395 = n25224 | n43394 ;
  assign n43396 = n43395 ^ n5686 ^ 1'b0 ;
  assign n43393 = n36171 & ~n38292 ;
  assign n43397 = n43396 ^ n43393 ^ 1'b0 ;
  assign n43398 = ~n17631 & n28790 ;
  assign n43399 = ( n5730 & ~n43200 ) | ( n5730 & n43398 ) | ( ~n43200 & n43398 ) ;
  assign n43400 = ( n1405 & ~n26648 ) | ( n1405 & n38054 ) | ( ~n26648 & n38054 ) ;
  assign n43401 = n8338 ^ n7679 ^ n3180 ;
  assign n43402 = n2914 & n43401 ;
  assign n43404 = n26121 ^ n6711 ^ 1'b0 ;
  assign n43405 = ~n7839 & n43404 ;
  assign n43403 = n8880 | n34397 ;
  assign n43406 = n43405 ^ n43403 ^ 1'b0 ;
  assign n43407 = n43406 ^ n14865 ^ 1'b0 ;
  assign n43411 = n12662 ^ n6980 ^ n2956 ;
  assign n43409 = ~n28054 & n33981 ;
  assign n43410 = n43409 ^ n2183 ^ 1'b0 ;
  assign n43408 = n36707 ^ n20800 ^ n15532 ;
  assign n43412 = n43411 ^ n43410 ^ n43408 ;
  assign n43413 = n43412 ^ n3172 ^ 1'b0 ;
  assign n43414 = ( ~n12485 & n15087 ) | ( ~n12485 & n43413 ) | ( n15087 & n43413 ) ;
  assign n43415 = ( n4146 & ~n13175 ) | ( n4146 & n18866 ) | ( ~n13175 & n18866 ) ;
  assign n43416 = n31770 ^ n20873 ^ 1'b0 ;
  assign n43417 = n43415 & n43416 ;
  assign n43418 = n15212 ^ n13364 ^ n3948 ;
  assign n43419 = ( ~n29863 & n43417 ) | ( ~n29863 & n43418 ) | ( n43417 & n43418 ) ;
  assign n43420 = n15510 ^ n4797 ^ 1'b0 ;
  assign n43421 = ~n40430 & n43420 ;
  assign n43422 = ( n21557 & n30838 ) | ( n21557 & n36849 ) | ( n30838 & n36849 ) ;
  assign n43423 = ( ~n18657 & n31334 ) | ( ~n18657 & n34425 ) | ( n31334 & n34425 ) ;
  assign n43424 = n5459 ^ n880 ^ 1'b0 ;
  assign n43425 = n24761 ^ n23142 ^ n3984 ;
  assign n43426 = n7836 & ~n8334 ;
  assign n43427 = n43426 ^ n24268 ^ 1'b0 ;
  assign n43428 = n31785 ^ n30974 ^ 1'b0 ;
  assign n43429 = n43427 & n43428 ;
  assign n43430 = ( n23375 & n43425 ) | ( n23375 & ~n43429 ) | ( n43425 & ~n43429 ) ;
  assign n43431 = ( n5331 & n43424 ) | ( n5331 & ~n43430 ) | ( n43424 & ~n43430 ) ;
  assign n43432 = n267 & ~n11307 ;
  assign n43433 = n43432 ^ n2630 ^ 1'b0 ;
  assign n43434 = n43433 ^ n10386 ^ x214 ;
  assign n43435 = ( n8148 & ~n18867 ) | ( n8148 & n42123 ) | ( ~n18867 & n42123 ) ;
  assign n43436 = n43209 ^ n1868 ^ 1'b0 ;
  assign n43437 = n43436 ^ n37596 ^ n15155 ;
  assign n43438 = n19686 ^ n17794 ^ 1'b0 ;
  assign n43439 = n37329 & ~n43438 ;
  assign n43440 = n43439 ^ n25369 ^ n319 ;
  assign n43444 = ( ~n5008 & n11150 ) | ( ~n5008 & n16758 ) | ( n11150 & n16758 ) ;
  assign n43445 = ( n7143 & ~n28334 ) | ( n7143 & n43444 ) | ( ~n28334 & n43444 ) ;
  assign n43441 = n5201 ^ n1295 ^ 1'b0 ;
  assign n43442 = n43441 ^ n42520 ^ 1'b0 ;
  assign n43443 = n3157 & n43442 ;
  assign n43446 = n43445 ^ n43443 ^ n4841 ;
  assign n43447 = ( n1784 & n9467 ) | ( n1784 & ~n43446 ) | ( n9467 & ~n43446 ) ;
  assign n43448 = ( n2299 & n7159 ) | ( n2299 & ~n9904 ) | ( n7159 & ~n9904 ) ;
  assign n43449 = n4663 & n26687 ;
  assign n43450 = n43448 & n43449 ;
  assign n43451 = n43450 ^ n18013 ^ 1'b0 ;
  assign n43452 = n34389 ^ n20800 ^ n19930 ;
  assign n43453 = n43452 ^ n18579 ^ n5804 ;
  assign n43454 = n40961 & ~n43453 ;
  assign n43455 = n43454 ^ n9478 ^ 1'b0 ;
  assign n43456 = n24316 ^ n17158 ^ 1'b0 ;
  assign n43459 = ( ~n11141 & n20868 ) | ( ~n11141 & n24860 ) | ( n20868 & n24860 ) ;
  assign n43457 = ( n5787 & ~n7224 ) | ( n5787 & n18673 ) | ( ~n7224 & n18673 ) ;
  assign n43458 = n43457 ^ n8506 ^ n2431 ;
  assign n43460 = n43459 ^ n43458 ^ x206 ;
  assign n43461 = ( ~n2472 & n7874 ) | ( ~n2472 & n41243 ) | ( n7874 & n41243 ) ;
  assign n43462 = ( n4657 & n14343 ) | ( n4657 & ~n16071 ) | ( n14343 & ~n16071 ) ;
  assign n43463 = ( n12453 & n16123 ) | ( n12453 & ~n36413 ) | ( n16123 & ~n36413 ) ;
  assign n43464 = n26794 ^ n24350 ^ n567 ;
  assign n43465 = ( n5309 & ~n11838 ) | ( n5309 & n43464 ) | ( ~n11838 & n43464 ) ;
  assign n43466 = ( n12597 & n14840 ) | ( n12597 & n43465 ) | ( n14840 & n43465 ) ;
  assign n43467 = ( ~n42214 & n43463 ) | ( ~n42214 & n43466 ) | ( n43463 & n43466 ) ;
  assign n43468 = n18095 & ~n40361 ;
  assign n43469 = n43468 ^ n8902 ^ 1'b0 ;
  assign n43470 = n40496 ^ n13139 ^ n7468 ;
  assign n43471 = n43470 ^ n10462 ^ 1'b0 ;
  assign n43472 = n11415 & n43471 ;
  assign n43473 = n38067 ^ n18497 ^ 1'b0 ;
  assign n43474 = n22827 & n43473 ;
  assign n43475 = ~n14106 & n43474 ;
  assign n43476 = n43475 ^ n11468 ^ 1'b0 ;
  assign n43477 = n7692 ^ n3495 ^ 1'b0 ;
  assign n43478 = ~n43476 & n43477 ;
  assign n43479 = n43478 ^ n38422 ^ n32777 ;
  assign n43480 = ( n32745 & ~n33319 ) | ( n32745 & n37025 ) | ( ~n33319 & n37025 ) ;
  assign n43481 = n43480 ^ n24171 ^ n22500 ;
  assign n43482 = n6777 & ~n12030 ;
  assign n43485 = n11683 & n13297 ;
  assign n43486 = n43485 ^ n23903 ^ 1'b0 ;
  assign n43483 = n15853 ^ n13865 ^ n13132 ;
  assign n43484 = n43483 ^ n41023 ^ n31811 ;
  assign n43487 = n43486 ^ n43484 ^ n38436 ;
  assign n43488 = n43487 ^ n27785 ^ n5318 ;
  assign n43489 = n718 | n38918 ;
  assign n43490 = n43488 & ~n43489 ;
  assign n43491 = n43490 ^ n18451 ^ 1'b0 ;
  assign n43492 = n21534 & n25544 ;
  assign n43493 = n43492 ^ n39467 ^ 1'b0 ;
  assign n43494 = ( n11924 & n24617 ) | ( n11924 & ~n43493 ) | ( n24617 & ~n43493 ) ;
  assign n43495 = ( x73 & n33917 ) | ( x73 & n42550 ) | ( n33917 & n42550 ) ;
  assign n43496 = ( n8575 & ~n32347 ) | ( n8575 & n38534 ) | ( ~n32347 & n38534 ) ;
  assign n43497 = n43496 ^ n16355 ^ 1'b0 ;
  assign n43498 = ( n18859 & ~n19336 ) | ( n18859 & n26409 ) | ( ~n19336 & n26409 ) ;
  assign n43499 = n43498 ^ n25218 ^ 1'b0 ;
  assign n43500 = ( n3459 & n23145 ) | ( n3459 & ~n43499 ) | ( n23145 & ~n43499 ) ;
  assign n43501 = n43500 ^ n37051 ^ n9451 ;
  assign n43502 = n27511 ^ n23397 ^ 1'b0 ;
  assign n43503 = n35362 & ~n43502 ;
  assign n43504 = n43503 ^ n17059 ^ n4887 ;
  assign n43505 = n31604 ^ n10832 ^ n8938 ;
  assign n43506 = ( ~n5285 & n40638 ) | ( ~n5285 & n43505 ) | ( n40638 & n43505 ) ;
  assign n43507 = n24093 ^ n14155 ^ n10635 ;
  assign n43508 = ( n14279 & n19910 ) | ( n14279 & ~n43507 ) | ( n19910 & ~n43507 ) ;
  assign n43509 = n32073 ^ n23465 ^ n10935 ;
  assign n43510 = n15927 | n23881 ;
  assign n43511 = n8031 & ~n43510 ;
  assign n43512 = ~n7304 & n43511 ;
  assign n43513 = n35310 ^ n962 ^ 1'b0 ;
  assign n43514 = n40310 & ~n43513 ;
  assign n43515 = n10550 & n10658 ;
  assign n43516 = n43515 ^ n22830 ^ n16475 ;
  assign n43517 = n33536 ^ n5135 ^ n1162 ;
  assign n43518 = ( n13787 & n17908 ) | ( n13787 & n43517 ) | ( n17908 & n43517 ) ;
  assign n43519 = n43518 ^ n32438 ^ n6858 ;
  assign n43520 = n27797 ^ n6689 ^ n1614 ;
  assign n43521 = ( n23174 & n38970 ) | ( n23174 & ~n43520 ) | ( n38970 & ~n43520 ) ;
  assign n43522 = n31243 ^ n30195 ^ n23841 ;
  assign n43523 = ~n3436 & n34681 ;
  assign n43524 = n28534 & n43523 ;
  assign n43525 = ( n4995 & n18657 ) | ( n4995 & ~n20978 ) | ( n18657 & ~n20978 ) ;
  assign n43526 = n22602 ^ n21864 ^ x241 ;
  assign n43527 = n43526 ^ n33131 ^ n24338 ;
  assign n43528 = n43527 ^ n39650 ^ n27723 ;
  assign n43533 = ~n994 & n32107 ;
  assign n43534 = n25875 & n43533 ;
  assign n43529 = n37270 ^ n24118 ^ n383 ;
  assign n43530 = ( ~n4765 & n11365 ) | ( ~n4765 & n43529 ) | ( n11365 & n43529 ) ;
  assign n43531 = n43530 ^ n16732 ^ 1'b0 ;
  assign n43532 = ~n18457 & n43531 ;
  assign n43535 = n43534 ^ n43532 ^ n38572 ;
  assign n43536 = n1631 & ~n27560 ;
  assign n43537 = n43536 ^ n30747 ^ n4194 ;
  assign n43538 = n17427 ^ n11048 ^ 1'b0 ;
  assign n43539 = x151 & ~n43538 ;
  assign n43540 = n43539 ^ n20512 ^ n19209 ;
  assign n43541 = n36565 ^ n28705 ^ n3554 ;
  assign n43542 = ( n629 & ~n1023 ) | ( n629 & n26747 ) | ( ~n1023 & n26747 ) ;
  assign n43543 = n16122 | n30195 ;
  assign n43544 = n20689 | n43543 ;
  assign n43545 = ( ~n23821 & n39964 ) | ( ~n23821 & n43544 ) | ( n39964 & n43544 ) ;
  assign n43546 = n43545 ^ n39216 ^ n13884 ;
  assign n43547 = n43546 ^ n2537 ^ 1'b0 ;
  assign n43548 = n28997 | n43547 ;
  assign n43549 = n16185 ^ n14535 ^ n4973 ;
  assign n43550 = ( ~n2042 & n15731 ) | ( ~n2042 & n35705 ) | ( n15731 & n35705 ) ;
  assign n43551 = n32604 & n43550 ;
  assign n43552 = ~n20670 & n43551 ;
  assign n43553 = ( n40062 & n43549 ) | ( n40062 & ~n43552 ) | ( n43549 & ~n43552 ) ;
  assign n43554 = n20577 | n35395 ;
  assign n43555 = n23431 ^ n19718 ^ n827 ;
  assign n43556 = n19974 ^ n16233 ^ 1'b0 ;
  assign n43557 = ~n982 & n23483 ;
  assign n43558 = n9990 ^ n5056 ^ n4588 ;
  assign n43559 = ( n14595 & ~n15615 ) | ( n14595 & n40069 ) | ( ~n15615 & n40069 ) ;
  assign n43560 = n2766 & ~n43559 ;
  assign n43561 = n43560 ^ n6276 ^ 1'b0 ;
  assign n43562 = n43561 ^ n5424 ^ n4354 ;
  assign n43563 = n43562 ^ n30217 ^ n20244 ;
  assign n43564 = n43563 ^ n7332 ^ 1'b0 ;
  assign n43565 = n43558 & ~n43564 ;
  assign n43566 = n35175 ^ x152 ^ 1'b0 ;
  assign n43567 = n14748 & n43566 ;
  assign n43568 = ~n7589 & n8160 ;
  assign n43569 = ~n19737 & n43568 ;
  assign n43570 = ( n31429 & n40326 ) | ( n31429 & n43569 ) | ( n40326 & n43569 ) ;
  assign n43571 = n12616 ^ x237 ^ 1'b0 ;
  assign n43572 = ( ~n2154 & n3183 ) | ( ~n2154 & n43571 ) | ( n3183 & n43571 ) ;
  assign n43573 = ( n1846 & n1925 ) | ( n1846 & n42421 ) | ( n1925 & n42421 ) ;
  assign n43574 = n14164 ^ n7433 ^ n6427 ;
  assign n43575 = n36869 & n43574 ;
  assign n43576 = n43575 ^ n40967 ^ n11409 ;
  assign n43578 = n12366 | n17717 ;
  assign n43577 = n2713 & ~n17807 ;
  assign n43579 = n43578 ^ n43577 ^ 1'b0 ;
  assign n43580 = n6993 ^ n2989 ^ 1'b0 ;
  assign n43581 = n12009 | n43580 ;
  assign n43582 = n11288 & ~n43581 ;
  assign n43583 = ( n6616 & n8140 ) | ( n6616 & ~n8218 ) | ( n8140 & ~n8218 ) ;
  assign n43584 = ( ~n4343 & n16358 ) | ( ~n4343 & n43583 ) | ( n16358 & n43583 ) ;
  assign n43589 = n20206 ^ n1131 ^ 1'b0 ;
  assign n43590 = n5408 & ~n43589 ;
  assign n43591 = ( ~n2636 & n2716 ) | ( ~n2636 & n32701 ) | ( n2716 & n32701 ) ;
  assign n43592 = ( n28438 & n43590 ) | ( n28438 & ~n43591 ) | ( n43590 & ~n43591 ) ;
  assign n43586 = n8239 ^ n3419 ^ 1'b0 ;
  assign n43587 = n12142 & n43586 ;
  assign n43585 = n5242 & ~n41211 ;
  assign n43588 = n43587 ^ n43585 ^ 1'b0 ;
  assign n43593 = n43592 ^ n43588 ^ n13191 ;
  assign n43594 = ( n16607 & ~n43584 ) | ( n16607 & n43593 ) | ( ~n43584 & n43593 ) ;
  assign n43595 = ( n842 & n10703 ) | ( n842 & n13069 ) | ( n10703 & n13069 ) ;
  assign n43596 = n43595 ^ n35359 ^ n31275 ;
  assign n43597 = n21843 ^ n11594 ^ n3855 ;
  assign n43598 = ( ~n10091 & n14133 ) | ( ~n10091 & n25813 ) | ( n14133 & n25813 ) ;
  assign n43599 = n43598 ^ n23945 ^ 1'b0 ;
  assign n43600 = n18435 | n43599 ;
  assign n43601 = n36151 ^ n26318 ^ n9412 ;
  assign n43602 = n19332 ^ n866 ^ 1'b0 ;
  assign n43603 = ( n31577 & n33516 ) | ( n31577 & ~n36352 ) | ( n33516 & ~n36352 ) ;
  assign n43604 = ( n5580 & ~n15955 ) | ( n5580 & n20130 ) | ( ~n15955 & n20130 ) ;
  assign n43605 = n43604 ^ n33554 ^ 1'b0 ;
  assign n43606 = n29446 ^ n18735 ^ 1'b0 ;
  assign n43607 = n6145 | n12731 ;
  assign n43608 = n43607 ^ n11301 ^ 1'b0 ;
  assign n43609 = n43608 ^ n24133 ^ n7688 ;
  assign n43610 = n3798 ^ n1609 ^ n897 ;
  assign n43611 = ~n2832 & n4354 ;
  assign n43612 = n43611 ^ n8310 ^ n1573 ;
  assign n43613 = n43612 ^ n20654 ^ n6353 ;
  assign n43614 = ~n43610 & n43613 ;
  assign n43615 = ( n12147 & n23690 ) | ( n12147 & ~n27583 ) | ( n23690 & ~n27583 ) ;
  assign n43618 = ( n2388 & n4925 ) | ( n2388 & ~n17361 ) | ( n4925 & ~n17361 ) ;
  assign n43616 = n8397 | n34341 ;
  assign n43617 = n5878 | n43616 ;
  assign n43619 = n43618 ^ n43617 ^ 1'b0 ;
  assign n43620 = ( x165 & ~n5215 ) | ( x165 & n32808 ) | ( ~n5215 & n32808 ) ;
  assign n43621 = n43620 ^ n34836 ^ n17454 ;
  assign n43622 = ~n2137 & n43621 ;
  assign n43623 = n13465 & n43622 ;
  assign n43628 = n2517 | n3490 ;
  assign n43624 = ( n519 & n5784 ) | ( n519 & ~n6946 ) | ( n5784 & ~n6946 ) ;
  assign n43625 = n26909 & ~n43624 ;
  assign n43626 = ( n2430 & n13213 ) | ( n2430 & ~n43625 ) | ( n13213 & ~n43625 ) ;
  assign n43627 = n43626 ^ n37707 ^ n26093 ;
  assign n43629 = n43628 ^ n43627 ^ n26420 ;
  assign n43630 = n18527 ^ n11615 ^ 1'b0 ;
  assign n43631 = ~n6357 & n27127 ;
  assign n43632 = ( ~x125 & n4295 ) | ( ~x125 & n43631 ) | ( n4295 & n43631 ) ;
  assign n43633 = n35596 ^ n19035 ^ 1'b0 ;
  assign n43634 = n21433 | n43633 ;
  assign n43635 = n368 | n22930 ;
  assign n43636 = n33587 ^ n8687 ^ n7445 ;
  assign n43639 = ( n13166 & ~n16694 ) | ( n13166 & n21980 ) | ( ~n16694 & n21980 ) ;
  assign n43637 = n12714 & ~n31416 ;
  assign n43638 = ~n14631 & n43637 ;
  assign n43640 = n43639 ^ n43638 ^ n40246 ;
  assign n43642 = ~n5864 & n20201 ;
  assign n43643 = n43642 ^ n23766 ^ 1'b0 ;
  assign n43644 = n43643 ^ n28000 ^ n923 ;
  assign n43641 = ( n4053 & n13548 ) | ( n4053 & n17069 ) | ( n13548 & n17069 ) ;
  assign n43645 = n43644 ^ n43641 ^ n32118 ;
  assign n43646 = n35582 ^ n22251 ^ n1721 ;
  assign n43647 = ( n14076 & n29345 ) | ( n14076 & ~n43646 ) | ( n29345 & ~n43646 ) ;
  assign n43648 = ( ~n24741 & n43645 ) | ( ~n24741 & n43647 ) | ( n43645 & n43647 ) ;
  assign n43649 = ( n2772 & n3865 ) | ( n2772 & ~n6925 ) | ( n3865 & ~n6925 ) ;
  assign n43650 = n5813 | n43649 ;
  assign n43651 = n3651 | n43650 ;
  assign n43652 = ( n11178 & n13146 ) | ( n11178 & ~n35633 ) | ( n13146 & ~n35633 ) ;
  assign n43653 = n31409 & ~n38894 ;
  assign n43654 = ~n24795 & n43653 ;
  assign n43655 = ( n31293 & n43652 ) | ( n31293 & n43654 ) | ( n43652 & n43654 ) ;
  assign n43656 = n25693 ^ n1301 ^ 1'b0 ;
  assign n43657 = ( n4324 & n11833 ) | ( n4324 & ~n37017 ) | ( n11833 & ~n37017 ) ;
  assign n43658 = ( n34639 & n43656 ) | ( n34639 & ~n43657 ) | ( n43656 & ~n43657 ) ;
  assign n43659 = ( n7075 & ~n7969 ) | ( n7075 & n31667 ) | ( ~n7969 & n31667 ) ;
  assign n43660 = n10155 & n43659 ;
  assign n43661 = n26400 ^ n12682 ^ n6516 ;
  assign n43662 = ~n4605 & n43661 ;
  assign n43663 = n43662 ^ n23998 ^ n4252 ;
  assign n43664 = n30049 ^ n13776 ^ 1'b0 ;
  assign n43665 = n43664 ^ n31833 ^ 1'b0 ;
  assign n43666 = n43665 ^ n32246 ^ n11012 ;
  assign n43667 = n31234 ^ n25666 ^ n14821 ;
  assign n43668 = ( n23655 & n43588 ) | ( n23655 & n43667 ) | ( n43588 & n43667 ) ;
  assign n43669 = ( n5852 & n19241 ) | ( n5852 & n43668 ) | ( n19241 & n43668 ) ;
  assign n43674 = ( ~n4655 & n9688 ) | ( ~n4655 & n12986 ) | ( n9688 & n12986 ) ;
  assign n43675 = ( n4322 & n4754 ) | ( n4322 & ~n43674 ) | ( n4754 & ~n43674 ) ;
  assign n43676 = ( n5829 & n8472 ) | ( n5829 & ~n43675 ) | ( n8472 & ~n43675 ) ;
  assign n43677 = ( n9419 & n27858 ) | ( n9419 & n43676 ) | ( n27858 & n43676 ) ;
  assign n43670 = ( ~n3383 & n17007 ) | ( ~n3383 & n24733 ) | ( n17007 & n24733 ) ;
  assign n43671 = ~n7242 & n43670 ;
  assign n43672 = ~n11364 & n43671 ;
  assign n43673 = ( n1335 & n18180 ) | ( n1335 & ~n43672 ) | ( n18180 & ~n43672 ) ;
  assign n43678 = n43677 ^ n43673 ^ 1'b0 ;
  assign n43679 = n10712 & n31873 ;
  assign n43680 = n43679 ^ n23717 ^ 1'b0 ;
  assign n43681 = ( n3102 & n3257 ) | ( n3102 & n8882 ) | ( n3257 & n8882 ) ;
  assign n43682 = n16805 | n43681 ;
  assign n43683 = n21394 | n43682 ;
  assign n43684 = n12628 ^ n4737 ^ n1456 ;
  assign n43685 = ( ~n22749 & n25788 ) | ( ~n22749 & n39337 ) | ( n25788 & n39337 ) ;
  assign n43686 = ~n15843 & n18710 ;
  assign n43687 = n43686 ^ n18088 ^ 1'b0 ;
  assign n43688 = n34608 ^ n17851 ^ n8434 ;
  assign n43689 = ( n43685 & ~n43687 ) | ( n43685 & n43688 ) | ( ~n43687 & n43688 ) ;
  assign n43690 = ( ~n4347 & n7386 ) | ( ~n4347 & n8491 ) | ( n7386 & n8491 ) ;
  assign n43694 = n34337 ^ n20067 ^ n2394 ;
  assign n43692 = n25611 ^ n15905 ^ n1807 ;
  assign n43693 = n43692 ^ n24029 ^ n8852 ;
  assign n43691 = n23001 ^ n18281 ^ n5661 ;
  assign n43695 = n43694 ^ n43693 ^ n43691 ;
  assign n43696 = n21935 ^ n21233 ^ 1'b0 ;
  assign n43697 = n25801 & n43696 ;
  assign n43698 = n30625 ^ n19399 ^ n5591 ;
  assign n43700 = n15170 ^ n13470 ^ n11900 ;
  assign n43699 = n7580 & ~n26296 ;
  assign n43701 = n43700 ^ n43699 ^ 1'b0 ;
  assign n43702 = n35110 ^ n17555 ^ n6316 ;
  assign n43703 = ( n10952 & n11278 ) | ( n10952 & n43077 ) | ( n11278 & n43077 ) ;
  assign n43704 = n14921 ^ n13394 ^ n12532 ;
  assign n43705 = n24552 ^ n13161 ^ 1'b0 ;
  assign n43706 = n43704 & n43705 ;
  assign n43707 = ~n16706 & n43706 ;
  assign n43708 = n43707 ^ n38861 ^ n26554 ;
  assign n43709 = n43708 ^ n38226 ^ 1'b0 ;
  assign n43710 = n43709 ^ n40852 ^ 1'b0 ;
  assign n43711 = ( n2699 & ~n3726 ) | ( n2699 & n26749 ) | ( ~n3726 & n26749 ) ;
  assign n43712 = n41253 ^ n8881 ^ 1'b0 ;
  assign n43713 = n43711 & n43712 ;
  assign n43714 = n3216 & ~n10796 ;
  assign n43715 = n41386 ^ n41115 ^ n20826 ;
  assign n43716 = n17727 ^ n9184 ^ 1'b0 ;
  assign n43717 = ~n43715 & n43716 ;
  assign n43718 = n16098 ^ n8808 ^ n1371 ;
  assign n43719 = ( n6495 & n27343 ) | ( n6495 & n33436 ) | ( n27343 & n33436 ) ;
  assign n43720 = ( n7618 & ~n43718 ) | ( n7618 & n43719 ) | ( ~n43718 & n43719 ) ;
  assign n43721 = n18912 & n24723 ;
  assign n43722 = ~n18441 & n43721 ;
  assign n43723 = ( n2818 & ~n21310 ) | ( n2818 & n43722 ) | ( ~n21310 & n43722 ) ;
  assign n43724 = ( n37264 & n43720 ) | ( n37264 & n43723 ) | ( n43720 & n43723 ) ;
  assign n43725 = ( n26779 & n42619 ) | ( n26779 & n43724 ) | ( n42619 & n43724 ) ;
  assign n43726 = n3333 | n21171 ;
  assign n43727 = n8214 | n43726 ;
  assign n43728 = ( n14473 & n26339 ) | ( n14473 & ~n35658 ) | ( n26339 & ~n35658 ) ;
  assign n43729 = ( n12908 & n43727 ) | ( n12908 & n43728 ) | ( n43727 & n43728 ) ;
  assign n43730 = n43729 ^ n26156 ^ n6858 ;
  assign n43731 = n24944 ^ n5574 ^ 1'b0 ;
  assign n43732 = n7284 & ~n43731 ;
  assign n43733 = n43732 ^ n13400 ^ n8932 ;
  assign n43734 = ( ~n1641 & n5698 ) | ( ~n1641 & n32827 ) | ( n5698 & n32827 ) ;
  assign n43735 = n40186 ^ n30205 ^ n12393 ;
  assign n43738 = n24619 ^ n5269 ^ 1'b0 ;
  assign n43736 = n19491 ^ n11173 ^ n561 ;
  assign n43737 = ( n9064 & n22285 ) | ( n9064 & n43736 ) | ( n22285 & n43736 ) ;
  assign n43739 = n43738 ^ n43737 ^ n33193 ;
  assign n43740 = ( n13639 & n37938 ) | ( n13639 & ~n43739 ) | ( n37938 & ~n43739 ) ;
  assign n43741 = n28882 ^ n24974 ^ n2925 ;
  assign n43742 = n4580 & ~n6655 ;
  assign n43743 = ( n2374 & n19348 ) | ( n2374 & n43742 ) | ( n19348 & n43742 ) ;
  assign n43744 = ~n282 & n43743 ;
  assign n43745 = ~n5422 & n43744 ;
  assign n43746 = n16069 ^ n15949 ^ n15797 ;
  assign n43747 = n3872 | n43746 ;
  assign n43748 = n43747 ^ n28997 ^ 1'b0 ;
  assign n43750 = ( ~n11123 & n22287 ) | ( ~n11123 & n23870 ) | ( n22287 & n23870 ) ;
  assign n43749 = ( n311 & n21219 ) | ( n311 & n27280 ) | ( n21219 & n27280 ) ;
  assign n43751 = n43750 ^ n43749 ^ 1'b0 ;
  assign n43752 = n18665 ^ n10957 ^ 1'b0 ;
  assign n43753 = n15097 & ~n43752 ;
  assign n43754 = ( n22583 & n27420 ) | ( n22583 & n40439 ) | ( n27420 & n40439 ) ;
  assign n43755 = ~n36689 & n39935 ;
  assign n43756 = n43755 ^ n31460 ^ n22219 ;
  assign n43757 = ( n8840 & ~n10119 ) | ( n8840 & n22220 ) | ( ~n10119 & n22220 ) ;
  assign n43758 = ( ~n9776 & n17285 ) | ( ~n9776 & n34307 ) | ( n17285 & n34307 ) ;
  assign n43759 = ( n30978 & n43757 ) | ( n30978 & ~n43758 ) | ( n43757 & ~n43758 ) ;
  assign n43760 = ( n43754 & ~n43756 ) | ( n43754 & n43759 ) | ( ~n43756 & n43759 ) ;
  assign n43761 = n8251 | n24581 ;
  assign n43762 = n43761 ^ n41384 ^ n18110 ;
  assign n43763 = ( n769 & ~n2744 ) | ( n769 & n16295 ) | ( ~n2744 & n16295 ) ;
  assign n43764 = n43763 ^ n24895 ^ n19673 ;
  assign n43765 = n43764 ^ n11557 ^ 1'b0 ;
  assign n43766 = n43765 ^ n28807 ^ n26282 ;
  assign n43767 = ( n26884 & n32716 ) | ( n26884 & ~n40925 ) | ( n32716 & ~n40925 ) ;
  assign n43768 = ~n23842 & n43767 ;
  assign n43769 = ( n5281 & n21002 ) | ( n5281 & n25954 ) | ( n21002 & n25954 ) ;
  assign n43770 = n41586 & n43769 ;
  assign n43771 = ~n30820 & n43770 ;
  assign n43772 = n21860 ^ n4626 ^ n2167 ;
  assign n43773 = n43772 ^ n26160 ^ n7227 ;
  assign n43775 = ( n9479 & ~n16031 ) | ( n9479 & n16242 ) | ( ~n16031 & n16242 ) ;
  assign n43774 = ~n11204 & n21617 ;
  assign n43776 = n43775 ^ n43774 ^ 1'b0 ;
  assign n43777 = ( n5311 & n11824 ) | ( n5311 & n14785 ) | ( n11824 & n14785 ) ;
  assign n43778 = ( n10855 & ~n43776 ) | ( n10855 & n43777 ) | ( ~n43776 & n43777 ) ;
  assign n43779 = n16725 | n31236 ;
  assign n43780 = n43779 ^ n2197 ^ 1'b0 ;
  assign n43781 = n43780 ^ n10498 ^ n8376 ;
  assign n43782 = ( ~n28693 & n43778 ) | ( ~n28693 & n43781 ) | ( n43778 & n43781 ) ;
  assign n43783 = n15151 ^ n13753 ^ n11677 ;
  assign n43784 = n43783 ^ n17583 ^ n7567 ;
  assign n43785 = ( ~n665 & n10509 ) | ( ~n665 & n36723 ) | ( n10509 & n36723 ) ;
  assign n43786 = n43785 ^ n33391 ^ n13340 ;
  assign n43787 = n28452 ^ n7020 ^ n2322 ;
  assign n43788 = n43787 ^ n38777 ^ n2295 ;
  assign n43789 = ( n1442 & ~n33780 ) | ( n1442 & n39479 ) | ( ~n33780 & n39479 ) ;
  assign n43790 = n22515 & ~n28131 ;
  assign n43791 = ( n3349 & n14281 ) | ( n3349 & ~n15841 ) | ( n14281 & ~n15841 ) ;
  assign n43792 = ( ~n8786 & n10106 ) | ( ~n8786 & n43791 ) | ( n10106 & n43791 ) ;
  assign n43793 = n34069 ^ n17366 ^ 1'b0 ;
  assign n43794 = n40991 | n43793 ;
  assign n43795 = ( n4215 & n5228 ) | ( n4215 & ~n5779 ) | ( n5228 & ~n5779 ) ;
  assign n43796 = ( n11322 & n15038 ) | ( n11322 & n43795 ) | ( n15038 & n43795 ) ;
  assign n43797 = n43796 ^ n37381 ^ n635 ;
  assign n43798 = ( n931 & ~n1692 ) | ( n931 & n10301 ) | ( ~n1692 & n10301 ) ;
  assign n43799 = n43798 ^ n29031 ^ n16224 ;
  assign n43800 = ( n8210 & n18311 ) | ( n8210 & n18828 ) | ( n18311 & n18828 ) ;
  assign n43801 = ( n19267 & ~n28721 ) | ( n19267 & n43800 ) | ( ~n28721 & n43800 ) ;
  assign n43802 = n37647 ^ n35654 ^ n2819 ;
  assign n43803 = ( n14770 & ~n18842 ) | ( n14770 & n27292 ) | ( ~n18842 & n27292 ) ;
  assign n43804 = n29198 & n43803 ;
  assign n43805 = ( n23921 & ~n43802 ) | ( n23921 & n43804 ) | ( ~n43802 & n43804 ) ;
  assign n43806 = ( ~n2801 & n11521 ) | ( ~n2801 & n11812 ) | ( n11521 & n11812 ) ;
  assign n43807 = ( n11281 & n21470 ) | ( n11281 & n33035 ) | ( n21470 & n33035 ) ;
  assign n43808 = ( n15943 & n26575 ) | ( n15943 & n39826 ) | ( n26575 & n39826 ) ;
  assign n43809 = n43808 ^ n38044 ^ n25066 ;
  assign n43810 = ( n43806 & ~n43807 ) | ( n43806 & n43809 ) | ( ~n43807 & n43809 ) ;
  assign n43811 = n42572 ^ n13136 ^ 1'b0 ;
  assign n43812 = ( n27410 & n27458 ) | ( n27410 & ~n29312 ) | ( n27458 & ~n29312 ) ;
  assign n43813 = n1577 | n43812 ;
  assign n43814 = n29651 ^ n464 ^ x61 ;
  assign n43815 = ( n24949 & n43813 ) | ( n24949 & ~n43814 ) | ( n43813 & ~n43814 ) ;
  assign n43816 = n39675 ^ n32868 ^ 1'b0 ;
  assign n43817 = n43266 | n43816 ;
  assign n43818 = n287 & ~n38122 ;
  assign n43819 = n43818 ^ n21375 ^ 1'b0 ;
  assign n43820 = n17035 & ~n43819 ;
  assign n43821 = n8980 | n36723 ;
  assign n43822 = n43820 & n43821 ;
  assign n43823 = n13403 & ~n29004 ;
  assign n43824 = n43823 ^ n17820 ^ 1'b0 ;
  assign n43825 = ( n4020 & ~n29785 ) | ( n4020 & n43824 ) | ( ~n29785 & n43824 ) ;
  assign n43826 = n34681 ^ n22339 ^ x37 ;
  assign n43827 = ( n5007 & n23397 ) | ( n5007 & ~n43826 ) | ( n23397 & ~n43826 ) ;
  assign n43829 = ( n2641 & n5233 ) | ( n2641 & ~n23896 ) | ( n5233 & ~n23896 ) ;
  assign n43828 = ( n576 & n14319 ) | ( n576 & ~n37401 ) | ( n14319 & ~n37401 ) ;
  assign n43830 = n43829 ^ n43828 ^ n14936 ;
  assign n43833 = ( n1363 & n1586 ) | ( n1363 & n32933 ) | ( n1586 & n32933 ) ;
  assign n43834 = n43833 ^ n16270 ^ n10661 ;
  assign n43831 = ( ~n2462 & n33697 ) | ( ~n2462 & n34627 ) | ( n33697 & n34627 ) ;
  assign n43832 = ( ~n8497 & n22394 ) | ( ~n8497 & n43831 ) | ( n22394 & n43831 ) ;
  assign n43835 = n43834 ^ n43832 ^ n16184 ;
  assign n43836 = n43835 ^ n1988 ^ 1'b0 ;
  assign n43837 = ~n43498 & n43836 ;
  assign n43840 = n8483 | n27695 ;
  assign n43841 = n43840 ^ n29049 ^ 1'b0 ;
  assign n43838 = n7496 & ~n29580 ;
  assign n43839 = n35583 & n43838 ;
  assign n43842 = n43841 ^ n43839 ^ n9612 ;
  assign n43843 = n635 | n43842 ;
  assign n43845 = ( n5543 & ~n10480 ) | ( n5543 & n25608 ) | ( ~n10480 & n25608 ) ;
  assign n43844 = n17951 ^ n7216 ^ n7169 ;
  assign n43846 = n43845 ^ n43844 ^ n2505 ;
  assign n43847 = ( n17609 & n18703 ) | ( n17609 & n24152 ) | ( n18703 & n24152 ) ;
  assign n43848 = n43847 ^ n15562 ^ n3027 ;
  assign n43849 = n19397 ^ n15867 ^ n4739 ;
  assign n43850 = n35014 ^ n34830 ^ n19852 ;
  assign n43851 = n27105 & ~n42928 ;
  assign n43852 = n20420 & n43851 ;
  assign n43853 = n11963 & n22012 ;
  assign n43854 = n24850 & n43853 ;
  assign n43855 = n43854 ^ n7165 ^ 1'b0 ;
  assign n43856 = n12344 & ~n43855 ;
  assign n43857 = n22339 & n31243 ;
  assign n43858 = n43857 ^ n10996 ^ 1'b0 ;
  assign n43859 = n43856 | n43858 ;
  assign n43860 = ~n9666 & n25013 ;
  assign n43861 = n38588 ^ n23459 ^ 1'b0 ;
  assign n43862 = ~n43860 & n43861 ;
  assign n43863 = ( ~n25784 & n42304 ) | ( ~n25784 & n43862 ) | ( n42304 & n43862 ) ;
  assign n43864 = n19608 ^ n14452 ^ n553 ;
  assign n43865 = ( n16477 & n25272 ) | ( n16477 & n27748 ) | ( n25272 & n27748 ) ;
  assign n43866 = n31855 ^ n29072 ^ n13317 ;
  assign n43867 = n29548 ^ n20140 ^ n13237 ;
  assign n43868 = ( ~n34382 & n43401 ) | ( ~n34382 & n43867 ) | ( n43401 & n43867 ) ;
  assign n43869 = ( n6074 & ~n24648 ) | ( n6074 & n43868 ) | ( ~n24648 & n43868 ) ;
  assign n43870 = n43869 ^ n10728 ^ n6566 ;
  assign n43871 = n42460 ^ n32720 ^ n16220 ;
  assign n43872 = n43871 ^ n7051 ^ 1'b0 ;
  assign n43873 = n10735 ^ n4932 ^ 1'b0 ;
  assign n43874 = n7756 & n43873 ;
  assign n43875 = ~n6779 & n40256 ;
  assign n43876 = n43875 ^ n34800 ^ 1'b0 ;
  assign n43877 = n43876 ^ n13189 ^ 1'b0 ;
  assign n43880 = n38169 ^ n38028 ^ 1'b0 ;
  assign n43881 = n11172 & ~n43880 ;
  assign n43878 = ( n5669 & ~n11648 ) | ( n5669 & n14305 ) | ( ~n11648 & n14305 ) ;
  assign n43879 = n33948 & n43878 ;
  assign n43882 = n43881 ^ n43879 ^ 1'b0 ;
  assign n43883 = ( ~n4869 & n38431 ) | ( ~n4869 & n43882 ) | ( n38431 & n43882 ) ;
  assign n43884 = ( ~n4460 & n17676 ) | ( ~n4460 & n34469 ) | ( n17676 & n34469 ) ;
  assign n43885 = ( ~n8075 & n31362 ) | ( ~n8075 & n33604 ) | ( n31362 & n33604 ) ;
  assign n43886 = n43885 ^ n19806 ^ n11108 ;
  assign n43887 = n15765 | n36596 ;
  assign n43888 = n18396 ^ n7492 ^ 1'b0 ;
  assign n43889 = n43888 ^ n35902 ^ n4910 ;
  assign n43890 = n19519 ^ n16833 ^ 1'b0 ;
  assign n43891 = n23034 ^ n15567 ^ 1'b0 ;
  assign n43892 = n8324 & n43891 ;
  assign n43893 = x235 & ~n7249 ;
  assign n43894 = ~n31854 & n43893 ;
  assign n43895 = n17491 ^ n8412 ^ n4536 ;
  assign n43896 = n14272 & n42096 ;
  assign n43897 = ( n1520 & n28365 ) | ( n1520 & ~n30238 ) | ( n28365 & ~n30238 ) ;
  assign n43898 = ( n7431 & ~n13777 ) | ( n7431 & n30720 ) | ( ~n13777 & n30720 ) ;
  assign n43904 = n39213 ^ n24786 ^ n11099 ;
  assign n43905 = n43904 ^ n27858 ^ n11567 ;
  assign n43899 = n19466 ^ n5628 ^ 1'b0 ;
  assign n43900 = n25727 ^ n4603 ^ 1'b0 ;
  assign n43901 = n23705 & n43900 ;
  assign n43902 = ( n4068 & n39479 ) | ( n4068 & ~n43901 ) | ( n39479 & ~n43901 ) ;
  assign n43903 = ( n23199 & n43899 ) | ( n23199 & ~n43902 ) | ( n43899 & ~n43902 ) ;
  assign n43906 = n43905 ^ n43903 ^ n9787 ;
  assign n43907 = ( n12274 & n15163 ) | ( n12274 & ~n31264 ) | ( n15163 & ~n31264 ) ;
  assign n43908 = n39303 ^ n11056 ^ 1'b0 ;
  assign n43909 = ~n43907 & n43908 ;
  assign n43910 = ( ~x200 & n19275 ) | ( ~x200 & n21109 ) | ( n19275 & n21109 ) ;
  assign n43911 = n31696 | n38035 ;
  assign n43912 = n43910 & ~n43911 ;
  assign n43913 = n22941 ^ n5415 ^ 1'b0 ;
  assign n43914 = n8778 ^ n7774 ^ 1'b0 ;
  assign n43915 = n2687 & ~n43914 ;
  assign n43916 = n43915 ^ n37143 ^ n11236 ;
  assign n43917 = n43916 ^ n43327 ^ n1866 ;
  assign n43918 = ( n10736 & n27151 ) | ( n10736 & n30451 ) | ( n27151 & n30451 ) ;
  assign n43919 = n43918 ^ n18560 ^ n12102 ;
  assign n43920 = n43919 ^ n7230 ^ n1301 ;
  assign n43924 = n4034 & ~n18223 ;
  assign n43925 = n43924 ^ n1038 ^ 1'b0 ;
  assign n43921 = ( n11545 & ~n17943 ) | ( n11545 & n21246 ) | ( ~n17943 & n21246 ) ;
  assign n43922 = n43921 ^ n32275 ^ n19233 ;
  assign n43923 = ( ~n7863 & n25316 ) | ( ~n7863 & n43922 ) | ( n25316 & n43922 ) ;
  assign n43926 = n43925 ^ n43923 ^ n34347 ;
  assign n43927 = ( n10752 & n22813 ) | ( n10752 & ~n27267 ) | ( n22813 & ~n27267 ) ;
  assign n43928 = n43927 ^ n39145 ^ n16324 ;
  assign n43929 = n14307 ^ n5890 ^ 1'b0 ;
  assign n43930 = ( n31866 & n36595 ) | ( n31866 & n43929 ) | ( n36595 & n43929 ) ;
  assign n43931 = n36247 ^ n395 ^ 1'b0 ;
  assign n43932 = n39761 ^ n37011 ^ n9012 ;
  assign n43933 = n14068 ^ n3416 ^ 1'b0 ;
  assign n43934 = n17175 & ~n43933 ;
  assign n43935 = n6116 & n18097 ;
  assign n43936 = n43935 ^ n7808 ^ 1'b0 ;
  assign n43937 = ( n1973 & n5498 ) | ( n1973 & ~n31179 ) | ( n5498 & ~n31179 ) ;
  assign n43938 = n10359 | n20265 ;
  assign n43939 = n43937 & ~n43938 ;
  assign n43940 = n43939 ^ n34176 ^ 1'b0 ;
  assign n43941 = n17271 ^ n11681 ^ n8336 ;
  assign n43942 = ( n9518 & ~n23083 ) | ( n9518 & n31762 ) | ( ~n23083 & n31762 ) ;
  assign n43943 = ( n23143 & n29454 ) | ( n23143 & ~n43942 ) | ( n29454 & ~n43942 ) ;
  assign n43944 = ( n16815 & ~n38438 ) | ( n16815 & n43943 ) | ( ~n38438 & n43943 ) ;
  assign n43945 = n43944 ^ n34737 ^ n3501 ;
  assign n43947 = ( n549 & n2680 ) | ( n549 & n35736 ) | ( n2680 & n35736 ) ;
  assign n43946 = ( n18076 & n32573 ) | ( n18076 & n42697 ) | ( n32573 & n42697 ) ;
  assign n43948 = n43947 ^ n43946 ^ n14261 ;
  assign n43949 = ( n4712 & n36046 ) | ( n4712 & n43948 ) | ( n36046 & n43948 ) ;
  assign n43950 = ( n1471 & n3486 ) | ( n1471 & n41947 ) | ( n3486 & n41947 ) ;
  assign n43951 = n37455 ^ n31570 ^ n15430 ;
  assign n43952 = n14830 ^ n10744 ^ x61 ;
  assign n43953 = n43952 ^ n35170 ^ n11907 ;
  assign n43954 = n14660 & ~n32058 ;
  assign n43955 = n20710 & n43954 ;
  assign n43956 = n31833 ^ n3741 ^ 1'b0 ;
  assign n43957 = n19139 & ~n19939 ;
  assign n43958 = ( n31137 & n34426 ) | ( n31137 & ~n39071 ) | ( n34426 & ~n39071 ) ;
  assign n43959 = ~n16730 & n29743 ;
  assign n43960 = n17549 & n43959 ;
  assign n43961 = n43960 ^ x13 ^ 1'b0 ;
  assign n43962 = n20401 ^ n18442 ^ n11041 ;
  assign n43963 = n43635 ^ n12226 ^ n2403 ;
  assign n43964 = n34841 ^ n16976 ^ n12341 ;
  assign n43965 = ( n1411 & ~n4437 ) | ( n1411 & n37353 ) | ( ~n4437 & n37353 ) ;
  assign n43966 = n43965 ^ n37486 ^ 1'b0 ;
  assign n43967 = n6038 & ~n43966 ;
  assign n43968 = n20621 | n35089 ;
  assign n43969 = n38311 ^ n21567 ^ n13482 ;
  assign n43973 = ( n5359 & n6285 ) | ( n5359 & n30410 ) | ( n6285 & n30410 ) ;
  assign n43974 = n23324 ^ n19599 ^ 1'b0 ;
  assign n43975 = ~n43973 & n43974 ;
  assign n43976 = n43975 ^ n17913 ^ n12737 ;
  assign n43977 = n43976 ^ n21567 ^ n3246 ;
  assign n43970 = n38195 ^ n24723 ^ n3495 ;
  assign n43971 = ( ~n8899 & n24865 ) | ( ~n8899 & n43970 ) | ( n24865 & n43970 ) ;
  assign n43972 = n43971 ^ n33979 ^ n11466 ;
  assign n43978 = n43977 ^ n43972 ^ n16013 ;
  assign n43979 = n42152 ^ n37990 ^ n25041 ;
  assign n43980 = n33972 ^ n26265 ^ n14496 ;
  assign n43981 = n43980 ^ n33353 ^ 1'b0 ;
  assign n43982 = ( ~n12027 & n41794 ) | ( ~n12027 & n43981 ) | ( n41794 & n43981 ) ;
  assign n43983 = n41182 ^ n26824 ^ n10819 ;
  assign n43984 = n43983 ^ n39426 ^ 1'b0 ;
  assign n43985 = n7632 ^ n4701 ^ n272 ;
  assign n43986 = n43985 ^ n22950 ^ n12452 ;
  assign n43987 = ( n4035 & ~n4538 ) | ( n4035 & n41711 ) | ( ~n4538 & n41711 ) ;
  assign n43988 = n41806 ^ n30990 ^ n5664 ;
  assign n43989 = ( n3911 & ~n43987 ) | ( n3911 & n43988 ) | ( ~n43987 & n43988 ) ;
  assign n43990 = ( n807 & ~n9278 ) | ( n807 & n34046 ) | ( ~n9278 & n34046 ) ;
  assign n43991 = ( n799 & n9209 ) | ( n799 & n43990 ) | ( n9209 & n43990 ) ;
  assign n43992 = n17194 & ~n42426 ;
  assign n43993 = n43991 & n43992 ;
  assign n43994 = n19929 ^ n7409 ^ 1'b0 ;
  assign n43995 = n9938 | n43994 ;
  assign n43996 = n27650 ^ n15331 ^ 1'b0 ;
  assign n43997 = ~n13558 & n43996 ;
  assign n43998 = ( ~n1072 & n1363 ) | ( ~n1072 & n16607 ) | ( n1363 & n16607 ) ;
  assign n43999 = ( n9319 & ~n33589 ) | ( n9319 & n43998 ) | ( ~n33589 & n43998 ) ;
  assign n44000 = n23920 ^ n23638 ^ 1'b0 ;
  assign n44001 = n42059 ^ n6890 ^ n6131 ;
  assign n44002 = n44001 ^ n16023 ^ 1'b0 ;
  assign n44003 = n44002 ^ n23758 ^ n4657 ;
  assign n44004 = n30606 ^ n20619 ^ n12105 ;
  assign n44006 = ( n8379 & ~n11698 ) | ( n8379 & n13994 ) | ( ~n11698 & n13994 ) ;
  assign n44005 = ( ~n5276 & n6294 ) | ( ~n5276 & n11021 ) | ( n6294 & n11021 ) ;
  assign n44007 = n44006 ^ n44005 ^ n2982 ;
  assign n44008 = ( n20911 & n22208 ) | ( n20911 & n26055 ) | ( n22208 & n26055 ) ;
  assign n44009 = ( ~n8751 & n9230 ) | ( ~n8751 & n18930 ) | ( n9230 & n18930 ) ;
  assign n44010 = ( ~n958 & n27989 ) | ( ~n958 & n44009 ) | ( n27989 & n44009 ) ;
  assign n44011 = ( n3364 & n5385 ) | ( n3364 & n44010 ) | ( n5385 & n44010 ) ;
  assign n44016 = n24181 ^ n15674 ^ n5059 ;
  assign n44012 = ~n2212 & n9566 ;
  assign n44013 = n44012 ^ n1071 ^ 1'b0 ;
  assign n44014 = ( n3921 & ~n34409 ) | ( n3921 & n44013 ) | ( ~n34409 & n44013 ) ;
  assign n44015 = n44014 ^ n41440 ^ n4403 ;
  assign n44017 = n44016 ^ n44015 ^ n31282 ;
  assign n44018 = ( n10875 & n18773 ) | ( n10875 & ~n27750 ) | ( n18773 & ~n27750 ) ;
  assign n44019 = ( n33988 & n43486 ) | ( n33988 & ~n44018 ) | ( n43486 & ~n44018 ) ;
  assign n44020 = n44019 ^ n4032 ^ 1'b0 ;
  assign n44023 = n4008 | n30559 ;
  assign n44024 = n44023 ^ n42309 ^ 1'b0 ;
  assign n44021 = ( n1784 & n7386 ) | ( n1784 & ~n37608 ) | ( n7386 & ~n37608 ) ;
  assign n44022 = ( n4252 & n36683 ) | ( n4252 & ~n44021 ) | ( n36683 & ~n44021 ) ;
  assign n44025 = n44024 ^ n44022 ^ 1'b0 ;
  assign n44026 = n44020 & ~n44025 ;
  assign n44027 = n4245 ^ n3732 ^ n3608 ;
  assign n44028 = ( n29818 & ~n39636 ) | ( n29818 & n44027 ) | ( ~n39636 & n44027 ) ;
  assign n44029 = n31402 ^ n12055 ^ n1808 ;
  assign n44030 = ~n42937 & n44029 ;
  assign n44031 = ( n14697 & ~n15244 ) | ( n14697 & n26795 ) | ( ~n15244 & n26795 ) ;
  assign n44032 = n44031 ^ n1021 ^ 1'b0 ;
  assign n44033 = ( n1621 & ~n5401 ) | ( n1621 & n29488 ) | ( ~n5401 & n29488 ) ;
  assign n44034 = n44033 ^ n39454 ^ 1'b0 ;
  assign n44035 = n14588 & n25702 ;
  assign n44036 = ( n24127 & ~n35450 ) | ( n24127 & n44035 ) | ( ~n35450 & n44035 ) ;
  assign n44037 = n41272 ^ n34004 ^ n27988 ;
  assign n44038 = n9755 & n44037 ;
  assign n44039 = n44038 ^ n29745 ^ 1'b0 ;
  assign n44040 = ( n8769 & n9668 ) | ( n8769 & n42935 ) | ( n9668 & n42935 ) ;
  assign n44041 = ~n22889 & n43309 ;
  assign n44042 = n15874 ^ n4130 ^ n1910 ;
  assign n44043 = n44042 ^ n24728 ^ n4354 ;
  assign n44044 = ( n1294 & ~n35118 ) | ( n1294 & n35450 ) | ( ~n35118 & n35450 ) ;
  assign n44045 = n44044 ^ n20437 ^ 1'b0 ;
  assign n44046 = n18920 & ~n44045 ;
  assign n44047 = n40128 ^ n39219 ^ n24499 ;
  assign n44048 = n23313 ^ n14796 ^ n10600 ;
  assign n44049 = n3947 ^ n853 ^ n760 ;
  assign n44050 = n44049 ^ n4853 ^ n1684 ;
  assign n44051 = n44050 ^ n35252 ^ n33065 ;
  assign n44052 = ( n17443 & ~n44048 ) | ( n17443 & n44051 ) | ( ~n44048 & n44051 ) ;
  assign n44053 = ( ~x204 & n6767 ) | ( ~x204 & n7542 ) | ( n6767 & n7542 ) ;
  assign n44054 = n26250 & n44053 ;
  assign n44055 = ( n11131 & ~n19346 ) | ( n11131 & n24266 ) | ( ~n19346 & n24266 ) ;
  assign n44056 = n44055 ^ n6143 ^ n5981 ;
  assign n44057 = n24420 ^ n5117 ^ n2039 ;
  assign n44058 = ( n23026 & n44056 ) | ( n23026 & n44057 ) | ( n44056 & n44057 ) ;
  assign n44059 = n647 & ~n33403 ;
  assign n44060 = n44059 ^ n16297 ^ 1'b0 ;
  assign n44061 = n44060 ^ n885 ^ 1'b0 ;
  assign n44062 = n44061 ^ n29821 ^ n26619 ;
  assign n44063 = n12897 ^ n5724 ^ n3826 ;
  assign n44064 = n28333 ^ n17235 ^ 1'b0 ;
  assign n44065 = ( n32578 & n44063 ) | ( n32578 & ~n44064 ) | ( n44063 & ~n44064 ) ;
  assign n44066 = n23708 ^ n23017 ^ 1'b0 ;
  assign n44067 = ~n2592 & n44066 ;
  assign n44068 = n28449 & n44060 ;
  assign n44069 = n44068 ^ n23908 ^ 1'b0 ;
  assign n44070 = n32770 ^ n6057 ^ n1485 ;
  assign n44071 = ( n6500 & n20186 ) | ( n6500 & ~n28655 ) | ( n20186 & ~n28655 ) ;
  assign n44072 = n44070 & ~n44071 ;
  assign n44079 = n26204 ^ n16027 ^ n2440 ;
  assign n44076 = ( n7499 & n11602 ) | ( n7499 & n29396 ) | ( n11602 & n29396 ) ;
  assign n44077 = n1378 & n11009 ;
  assign n44078 = ~n44076 & n44077 ;
  assign n44080 = n44079 ^ n44078 ^ n7748 ;
  assign n44073 = n1899 | n6051 ;
  assign n44074 = n44073 ^ n37721 ^ n25061 ;
  assign n44075 = n33957 & ~n44074 ;
  assign n44081 = n44080 ^ n44075 ^ n11281 ;
  assign n44082 = n14220 ^ n11203 ^ n5517 ;
  assign n44083 = n44082 ^ n14153 ^ n12974 ;
  assign n44084 = n2066 & ~n7098 ;
  assign n44085 = n44084 ^ n28178 ^ 1'b0 ;
  assign n44090 = ( ~n13025 & n19999 ) | ( ~n13025 & n21060 ) | ( n19999 & n21060 ) ;
  assign n44086 = n17477 ^ n15833 ^ n4143 ;
  assign n44087 = n7406 & n33426 ;
  assign n44088 = n44087 ^ n22939 ^ n15309 ;
  assign n44089 = ( ~n43458 & n44086 ) | ( ~n43458 & n44088 ) | ( n44086 & n44088 ) ;
  assign n44091 = n44090 ^ n44089 ^ n14770 ;
  assign n44092 = ( n32828 & n39998 ) | ( n32828 & n40889 ) | ( n39998 & n40889 ) ;
  assign n44093 = ( n11424 & n12868 ) | ( n11424 & n33244 ) | ( n12868 & n33244 ) ;
  assign n44094 = n24899 | n30818 ;
  assign n44095 = n29078 & ~n44094 ;
  assign n44096 = ( n33582 & n43985 ) | ( n33582 & ~n44095 ) | ( n43985 & ~n44095 ) ;
  assign n44097 = ( ~n44092 & n44093 ) | ( ~n44092 & n44096 ) | ( n44093 & n44096 ) ;
  assign n44098 = n9450 ^ x217 ^ 1'b0 ;
  assign n44099 = n13251 & ~n37111 ;
  assign n44100 = n3874 & n44099 ;
  assign n44101 = ~n33800 & n37069 ;
  assign n44102 = n31063 & n44101 ;
  assign n44103 = n36809 ^ n5555 ^ 1'b0 ;
  assign n44104 = ( n27713 & n31816 ) | ( n27713 & ~n41766 ) | ( n31816 & ~n41766 ) ;
  assign n44105 = ( ~n6681 & n10927 ) | ( ~n6681 & n38579 ) | ( n10927 & n38579 ) ;
  assign n44106 = ( ~n5700 & n16517 ) | ( ~n5700 & n38212 ) | ( n16517 & n38212 ) ;
  assign n44107 = n44106 ^ n17215 ^ n6874 ;
  assign n44109 = n5192 ^ n2206 ^ 1'b0 ;
  assign n44108 = n29142 ^ n9998 ^ n6632 ;
  assign n44110 = n44109 ^ n44108 ^ n21578 ;
  assign n44111 = ~n7008 & n30114 ;
  assign n44112 = n44111 ^ n39677 ^ n11261 ;
  assign n44113 = n27070 ^ n10091 ^ n4415 ;
  assign n44114 = ( n7468 & n26715 ) | ( n7468 & n44113 ) | ( n26715 & n44113 ) ;
  assign n44115 = ( n13292 & n21595 ) | ( n13292 & ~n39854 ) | ( n21595 & ~n39854 ) ;
  assign n44116 = n35621 | n35697 ;
  assign n44117 = n44116 ^ n27432 ^ 1'b0 ;
  assign n44118 = ( ~n19251 & n27586 ) | ( ~n19251 & n37566 ) | ( n27586 & n37566 ) ;
  assign n44119 = ( n3892 & n4684 ) | ( n3892 & n14275 ) | ( n4684 & n14275 ) ;
  assign n44120 = n40470 & ~n44119 ;
  assign n44121 = n13374 ^ n6570 ^ 1'b0 ;
  assign n44122 = ~n28706 & n44121 ;
  assign n44123 = ( n6990 & ~n24685 ) | ( n6990 & n44122 ) | ( ~n24685 & n44122 ) ;
  assign n44124 = n33270 ^ n27262 ^ n11288 ;
  assign n44125 = ( n21049 & n32302 ) | ( n21049 & ~n44124 ) | ( n32302 & ~n44124 ) ;
  assign n44126 = n29934 ^ n13291 ^ 1'b0 ;
  assign n44127 = ~n1385 & n44126 ;
  assign n44128 = n44127 ^ n21458 ^ 1'b0 ;
  assign n44129 = n19278 ^ n11361 ^ 1'b0 ;
  assign n44130 = n4560 & n44129 ;
  assign n44131 = n8112 ^ n2931 ^ n1879 ;
  assign n44132 = ( ~n14322 & n25995 ) | ( ~n14322 & n44131 ) | ( n25995 & n44131 ) ;
  assign n44133 = n44132 ^ n11841 ^ n11051 ;
  assign n44134 = ( n12273 & n34736 ) | ( n12273 & ~n44133 ) | ( n34736 & ~n44133 ) ;
  assign n44135 = n28792 ^ n13079 ^ n3834 ;
  assign n44136 = n44135 ^ n10253 ^ n1141 ;
  assign n44137 = n40556 ^ n9220 ^ 1'b0 ;
  assign n44138 = n39789 | n44137 ;
  assign n44139 = n25255 ^ n3915 ^ n3645 ;
  assign n44140 = ( n29400 & n38707 ) | ( n29400 & ~n44139 ) | ( n38707 & ~n44139 ) ;
  assign n44141 = n8123 & ~n9829 ;
  assign n44142 = n44141 ^ n6948 ^ n2780 ;
  assign n44143 = n36247 ^ n31955 ^ n12676 ;
  assign n44144 = ( n14070 & ~n44142 ) | ( n14070 & n44143 ) | ( ~n44142 & n44143 ) ;
  assign n44145 = n17496 ^ n3915 ^ n2815 ;
  assign n44146 = n27407 ^ n16717 ^ n12979 ;
  assign n44147 = n44146 ^ n23924 ^ n5035 ;
  assign n44148 = n5867 | n17226 ;
  assign n44149 = n10350 | n44148 ;
  assign n44150 = n24270 ^ n13460 ^ 1'b0 ;
  assign n44151 = n10557 & ~n44150 ;
  assign n44152 = ( n28260 & n44149 ) | ( n28260 & ~n44151 ) | ( n44149 & ~n44151 ) ;
  assign n44153 = n21993 ^ n15426 ^ 1'b0 ;
  assign n44154 = n37908 & n44153 ;
  assign n44155 = n31260 ^ n17609 ^ n14490 ;
  assign n44156 = ~n9598 & n44155 ;
  assign n44157 = ( n28448 & n29183 ) | ( n28448 & n43918 ) | ( n29183 & n43918 ) ;
  assign n44158 = n44157 ^ n36536 ^ n7412 ;
  assign n44159 = n21542 ^ n5840 ^ 1'b0 ;
  assign n44160 = n25848 ^ n24087 ^ n7394 ;
  assign n44161 = n32651 ^ n18073 ^ n13781 ;
  assign n44162 = n15324 | n15401 ;
  assign n44163 = n964 & ~n44162 ;
  assign n44164 = n1384 | n18042 ;
  assign n44165 = n44164 ^ n15642 ^ 1'b0 ;
  assign n44166 = n9841 ^ n3649 ^ n3004 ;
  assign n44167 = n44166 ^ n13778 ^ n8051 ;
  assign n44168 = ( ~n4245 & n42195 ) | ( ~n4245 & n44167 ) | ( n42195 & n44167 ) ;
  assign n44170 = n13513 ^ n5591 ^ n4197 ;
  assign n44169 = n41652 ^ n20258 ^ n7639 ;
  assign n44171 = n44170 ^ n44169 ^ n6995 ;
  assign n44172 = ( n32304 & n43009 ) | ( n32304 & n44171 ) | ( n43009 & n44171 ) ;
  assign n44173 = ( n31613 & ~n31762 ) | ( n31613 & n42905 ) | ( ~n31762 & n42905 ) ;
  assign n44174 = ( ~n3894 & n31455 ) | ( ~n3894 & n44173 ) | ( n31455 & n44173 ) ;
  assign n44175 = n25935 ^ n15481 ^ n3568 ;
  assign n44176 = n19193 ^ n18429 ^ n2303 ;
  assign n44177 = ( n39381 & n44175 ) | ( n39381 & n44176 ) | ( n44175 & n44176 ) ;
  assign n44178 = n44177 ^ n24164 ^ n14057 ;
  assign n44180 = n11699 ^ n4286 ^ 1'b0 ;
  assign n44179 = ( ~n3165 & n6113 ) | ( ~n3165 & n13274 ) | ( n6113 & n13274 ) ;
  assign n44181 = n44180 ^ n44179 ^ n6414 ;
  assign n44182 = ( ~n20087 & n23843 ) | ( ~n20087 & n44181 ) | ( n23843 & n44181 ) ;
  assign n44183 = n38782 | n40561 ;
  assign n44184 = n42049 ^ n10544 ^ 1'b0 ;
  assign n44185 = n3937 | n44184 ;
  assign n44186 = n3105 & n44185 ;
  assign n44187 = ( n11299 & n30953 ) | ( n11299 & n32242 ) | ( n30953 & n32242 ) ;
  assign n44189 = n19818 ^ n5446 ^ 1'b0 ;
  assign n44190 = ~n9057 & n44189 ;
  assign n44188 = n19360 ^ n12419 ^ n7658 ;
  assign n44191 = n44190 ^ n44188 ^ n6213 ;
  assign n44192 = ( n22628 & ~n34418 ) | ( n22628 & n39216 ) | ( ~n34418 & n39216 ) ;
  assign n44193 = n36513 ^ n22727 ^ 1'b0 ;
  assign n44194 = ( n23705 & n39477 ) | ( n23705 & ~n44193 ) | ( n39477 & ~n44193 ) ;
  assign n44195 = n13844 ^ n11056 ^ 1'b0 ;
  assign n44196 = ( ~n6297 & n9253 ) | ( ~n6297 & n27932 ) | ( n9253 & n27932 ) ;
  assign n44197 = n44196 ^ n32185 ^ n26468 ;
  assign n44198 = n44197 ^ n21193 ^ n2137 ;
  assign n44199 = n44198 ^ n42119 ^ 1'b0 ;
  assign n44200 = n26925 | n44199 ;
  assign n44201 = n44200 ^ n24004 ^ n19494 ;
  assign n44202 = ( n1907 & n11915 ) | ( n1907 & ~n16859 ) | ( n11915 & ~n16859 ) ;
  assign n44203 = n44202 ^ n16990 ^ 1'b0 ;
  assign n44204 = ( ~n44195 & n44201 ) | ( ~n44195 & n44203 ) | ( n44201 & n44203 ) ;
  assign n44205 = n16671 ^ n8298 ^ x16 ;
  assign n44206 = n5357 & ~n8359 ;
  assign n44207 = n44206 ^ n11468 ^ 1'b0 ;
  assign n44208 = ( n16811 & n44205 ) | ( n16811 & n44207 ) | ( n44205 & n44207 ) ;
  assign n44209 = ( ~n11307 & n16101 ) | ( ~n11307 & n44208 ) | ( n16101 & n44208 ) ;
  assign n44210 = n17743 ^ n17179 ^ n13136 ;
  assign n44211 = ( n569 & n12405 ) | ( n569 & ~n21337 ) | ( n12405 & ~n21337 ) ;
  assign n44212 = ( n12836 & n42074 ) | ( n12836 & ~n44211 ) | ( n42074 & ~n44211 ) ;
  assign n44213 = n19502 ^ n3565 ^ 1'b0 ;
  assign n44214 = ( n9954 & n17360 ) | ( n9954 & n44213 ) | ( n17360 & n44213 ) ;
  assign n44215 = ( n1704 & n9975 ) | ( n1704 & ~n44214 ) | ( n9975 & ~n44214 ) ;
  assign n44216 = n25676 ^ n4206 ^ 1'b0 ;
  assign n44217 = n30797 ^ n12871 ^ n2809 ;
  assign n44218 = ( n26438 & n43804 ) | ( n26438 & ~n44217 ) | ( n43804 & ~n44217 ) ;
  assign n44219 = n4824 ^ n4440 ^ 1'b0 ;
  assign n44222 = n23819 ^ n17689 ^ n3366 ;
  assign n44220 = x81 & n11565 ;
  assign n44221 = n11040 & n44220 ;
  assign n44223 = n44222 ^ n44221 ^ 1'b0 ;
  assign n44224 = n42961 & n44223 ;
  assign n44225 = ~n2162 & n14406 ;
  assign n44226 = n44225 ^ n19201 ^ 1'b0 ;
  assign n44234 = ( n4612 & n14669 ) | ( n4612 & n19953 ) | ( n14669 & n19953 ) ;
  assign n44229 = n39654 ^ n11443 ^ n9913 ;
  assign n44230 = n36284 & ~n44229 ;
  assign n44227 = n15163 ^ n5869 ^ n5296 ;
  assign n44228 = n3631 & ~n44227 ;
  assign n44231 = n44230 ^ n44228 ^ 1'b0 ;
  assign n44232 = n44231 ^ n34157 ^ n28365 ;
  assign n44233 = ( n3687 & n24367 ) | ( n3687 & ~n44232 ) | ( n24367 & ~n44232 ) ;
  assign n44235 = n44234 ^ n44233 ^ n13829 ;
  assign n44236 = n36979 ^ n11105 ^ n4599 ;
  assign n44237 = ( n11370 & ~n30609 ) | ( n11370 & n44236 ) | ( ~n30609 & n44236 ) ;
  assign n44238 = n25069 ^ n10243 ^ 1'b0 ;
  assign n44239 = n6945 & n44238 ;
  assign n44240 = ( ~n10961 & n43991 ) | ( ~n10961 & n44239 ) | ( n43991 & n44239 ) ;
  assign n44241 = n33993 | n44240 ;
  assign n44242 = n44241 ^ n35549 ^ n12471 ;
  assign n44243 = n19816 ^ n14787 ^ 1'b0 ;
  assign n44244 = ~n31222 & n44243 ;
  assign n44245 = n44244 ^ n33064 ^ 1'b0 ;
  assign n44246 = ( n3130 & ~n29357 ) | ( n3130 & n37274 ) | ( ~n29357 & n37274 ) ;
  assign n44247 = n25368 ^ n6905 ^ 1'b0 ;
  assign n44248 = n12147 | n41509 ;
  assign n44249 = n44248 ^ n17149 ^ 1'b0 ;
  assign n44250 = ( n17022 & n23734 ) | ( n17022 & n26001 ) | ( n23734 & n26001 ) ;
  assign n44251 = n44250 ^ n43294 ^ n36298 ;
  assign n44252 = n28721 ^ n25208 ^ n24753 ;
  assign n44253 = ( n3248 & n11922 ) | ( n3248 & n44252 ) | ( n11922 & n44252 ) ;
  assign n44254 = n44253 ^ n22849 ^ n9328 ;
  assign n44255 = n18648 & ~n25771 ;
  assign n44256 = ( n10672 & n30141 ) | ( n10672 & ~n41355 ) | ( n30141 & ~n41355 ) ;
  assign n44257 = n27740 ^ n16406 ^ n6247 ;
  assign n44258 = n44257 ^ n694 ^ 1'b0 ;
  assign n44259 = n20077 & ~n44258 ;
  assign n44260 = n5792 & n14275 ;
  assign n44261 = n44260 ^ n12809 ^ 1'b0 ;
  assign n44262 = n8869 ^ n688 ^ 1'b0 ;
  assign n44263 = ~n40042 & n44262 ;
  assign n44264 = n44263 ^ n9922 ^ 1'b0 ;
  assign n44265 = n16376 ^ n4280 ^ 1'b0 ;
  assign n44266 = ( n3672 & n19971 ) | ( n3672 & ~n35014 ) | ( n19971 & ~n35014 ) ;
  assign n44267 = n14534 ^ n10607 ^ n4392 ;
  assign n44268 = ( ~n1831 & n4007 ) | ( ~n1831 & n30437 ) | ( n4007 & n30437 ) ;
  assign n44269 = n44267 | n44268 ;
  assign n44270 = ( n14674 & ~n20078 ) | ( n14674 & n36415 ) | ( ~n20078 & n36415 ) ;
  assign n44271 = n2056 ^ n405 ^ 1'b0 ;
  assign n44272 = ( ~n9309 & n44270 ) | ( ~n9309 & n44271 ) | ( n44270 & n44271 ) ;
  assign n44273 = n33992 ^ n10230 ^ n7593 ;
  assign n44274 = n44273 ^ n23451 ^ 1'b0 ;
  assign n44275 = n27492 ^ n17825 ^ n10656 ;
  assign n44276 = n20130 | n33481 ;
  assign n44277 = n44276 ^ n41370 ^ 1'b0 ;
  assign n44278 = x118 & ~n34401 ;
  assign n44279 = ~n20448 & n44278 ;
  assign n44280 = n21960 ^ n1169 ^ 1'b0 ;
  assign n44281 = n8980 | n33282 ;
  assign n44282 = n34769 & ~n44281 ;
  assign n44283 = ( n21210 & n44280 ) | ( n21210 & n44282 ) | ( n44280 & n44282 ) ;
  assign n44284 = ( n1553 & ~n5502 ) | ( n1553 & n7496 ) | ( ~n5502 & n7496 ) ;
  assign n44285 = n466 & ~n12477 ;
  assign n44286 = ~n10166 & n44285 ;
  assign n44287 = n44286 ^ n4687 ^ 1'b0 ;
  assign n44288 = n9905 & n44287 ;
  assign n44289 = ( n778 & ~n35969 ) | ( n778 & n44288 ) | ( ~n35969 & n44288 ) ;
  assign n44290 = n44289 ^ n7119 ^ n3034 ;
  assign n44291 = ( n7546 & n44284 ) | ( n7546 & n44290 ) | ( n44284 & n44290 ) ;
  assign n44292 = n8095 & ~n35315 ;
  assign n44293 = n9246 ^ n8748 ^ 1'b0 ;
  assign n44294 = n3482 & n44293 ;
  assign n44295 = n44294 ^ n27696 ^ n4006 ;
  assign n44296 = n17812 | n27730 ;
  assign n44297 = n44295 & ~n44296 ;
  assign n44298 = n22121 ^ n12396 ^ 1'b0 ;
  assign n44299 = n44298 ^ n41286 ^ n4405 ;
  assign n44300 = ( n43532 & n44297 ) | ( n43532 & ~n44299 ) | ( n44297 & ~n44299 ) ;
  assign n44301 = n22650 ^ n577 ^ 1'b0 ;
  assign n44302 = ( n1693 & n21816 ) | ( n1693 & n44301 ) | ( n21816 & n44301 ) ;
  assign n44303 = n9481 ^ n9286 ^ n8502 ;
  assign n44304 = n13884 | n16676 ;
  assign n44305 = ~n778 & n16598 ;
  assign n44306 = ( n13100 & n15232 ) | ( n13100 & ~n18738 ) | ( n15232 & ~n18738 ) ;
  assign n44307 = n31397 ^ n22438 ^ n19997 ;
  assign n44308 = ( n28703 & n44306 ) | ( n28703 & n44307 ) | ( n44306 & n44307 ) ;
  assign n44309 = n29209 & n29829 ;
  assign n44310 = n9557 & n44309 ;
  assign n44311 = ( n37473 & ~n40093 ) | ( n37473 & n44310 ) | ( ~n40093 & n44310 ) ;
  assign n44312 = n14238 ^ n6603 ^ n1422 ;
  assign n44313 = n39511 & ~n44312 ;
  assign n44314 = ( n970 & n30660 ) | ( n970 & ~n34112 ) | ( n30660 & ~n34112 ) ;
  assign n44315 = n44314 ^ n40738 ^ n38832 ;
  assign n44316 = ( n21457 & n26298 ) | ( n21457 & n35859 ) | ( n26298 & n35859 ) ;
  assign n44317 = n6378 ^ n4341 ^ n2156 ;
  assign n44318 = n5354 ^ n4641 ^ n4126 ;
  assign n44319 = n44318 ^ n21757 ^ n16955 ;
  assign n44320 = ( n23477 & n44317 ) | ( n23477 & n44319 ) | ( n44317 & n44319 ) ;
  assign n44321 = n44320 ^ n12034 ^ 1'b0 ;
  assign n44322 = ( n26539 & ~n28040 ) | ( n26539 & n44321 ) | ( ~n28040 & n44321 ) ;
  assign n44323 = ~n18278 & n42925 ;
  assign n44324 = n44323 ^ n41482 ^ 1'b0 ;
  assign n44325 = ( n7364 & ~n10857 ) | ( n7364 & n17787 ) | ( ~n10857 & n17787 ) ;
  assign n44326 = n44325 ^ n19260 ^ 1'b0 ;
  assign n44327 = n29891 & n44326 ;
  assign n44328 = ( n418 & ~n1749 ) | ( n418 & n5616 ) | ( ~n1749 & n5616 ) ;
  assign n44329 = n32275 ^ n14033 ^ n8246 ;
  assign n44330 = ( n4496 & n13867 ) | ( n4496 & ~n44329 ) | ( n13867 & ~n44329 ) ;
  assign n44331 = n5335 & n44330 ;
  assign n44332 = n44331 ^ n37112 ^ n25655 ;
  assign n44333 = ( n17356 & ~n29661 ) | ( n17356 & n30854 ) | ( ~n29661 & n30854 ) ;
  assign n44334 = ( n13209 & n24420 ) | ( n13209 & n44333 ) | ( n24420 & n44333 ) ;
  assign n44337 = n37970 ^ n32195 ^ n20270 ;
  assign n44335 = n461 & n20460 ;
  assign n44336 = ( ~n7662 & n14564 ) | ( ~n7662 & n44335 ) | ( n14564 & n44335 ) ;
  assign n44338 = n44337 ^ n44336 ^ n922 ;
  assign n44339 = ( ~n6337 & n12581 ) | ( ~n6337 & n29583 ) | ( n12581 & n29583 ) ;
  assign n44340 = n44339 ^ n36343 ^ n28675 ;
  assign n44341 = ~x87 & n37695 ;
  assign n44342 = n2140 | n28285 ;
  assign n44343 = n14755 | n44342 ;
  assign n44344 = ( n2937 & n17449 ) | ( n2937 & n44343 ) | ( n17449 & n44343 ) ;
  assign n44345 = n29531 ^ n16806 ^ n1659 ;
  assign n44346 = n7890 & n40620 ;
  assign n44347 = ~n44345 & n44346 ;
  assign n44348 = n44347 ^ n32096 ^ n25013 ;
  assign n44349 = n37189 ^ n10690 ^ n6308 ;
  assign n44351 = n25814 ^ n11528 ^ 1'b0 ;
  assign n44352 = ~n32471 & n44351 ;
  assign n44350 = n30974 ^ n30619 ^ n29355 ;
  assign n44353 = n44352 ^ n44350 ^ 1'b0 ;
  assign n44354 = n42078 ^ n8946 ^ n8233 ;
  assign n44355 = n26998 ^ n11234 ^ 1'b0 ;
  assign n44356 = ~n44354 & n44355 ;
  assign n44357 = ( n7088 & ~n19826 ) | ( n7088 & n39074 ) | ( ~n19826 & n39074 ) ;
  assign n44358 = n22171 | n44357 ;
  assign n44359 = n17103 & ~n44358 ;
  assign n44360 = ( ~n15334 & n22665 ) | ( ~n15334 & n44359 ) | ( n22665 & n44359 ) ;
  assign n44361 = n33573 ^ n31045 ^ n6650 ;
  assign n44362 = n44361 ^ n13750 ^ n7726 ;
  assign n44363 = ( n987 & ~n1363 ) | ( n987 & n24511 ) | ( ~n1363 & n24511 ) ;
  assign n44364 = ( ~n561 & n28354 ) | ( ~n561 & n38162 ) | ( n28354 & n38162 ) ;
  assign n44365 = ( ~n25863 & n30350 ) | ( ~n25863 & n44364 ) | ( n30350 & n44364 ) ;
  assign n44371 = n13160 | n44166 ;
  assign n44372 = n44371 ^ n23227 ^ 1'b0 ;
  assign n44366 = n39284 ^ n23808 ^ n21091 ;
  assign n44367 = n44366 ^ n16209 ^ n7801 ;
  assign n44368 = n44367 ^ n16488 ^ 1'b0 ;
  assign n44369 = n11050 & n44368 ;
  assign n44370 = n44369 ^ n40531 ^ 1'b0 ;
  assign n44373 = n44372 ^ n44370 ^ n19896 ;
  assign n44374 = ( n14287 & ~n26146 ) | ( n14287 & n42202 ) | ( ~n26146 & n42202 ) ;
  assign n44375 = n15336 & ~n23668 ;
  assign n44376 = ~n16154 & n44375 ;
  assign n44377 = n9484 & n44376 ;
  assign n44378 = n37755 ^ n19509 ^ 1'b0 ;
  assign n44379 = n9106 ^ n5052 ^ n2816 ;
  assign n44380 = n18376 ^ n11951 ^ 1'b0 ;
  assign n44381 = x103 & n44380 ;
  assign n44382 = ( n2154 & n34947 ) | ( n2154 & ~n44381 ) | ( n34947 & ~n44381 ) ;
  assign n44383 = n38928 ^ n28062 ^ n26567 ;
  assign n44384 = n44383 ^ n43071 ^ n34389 ;
  assign n44385 = ( n44379 & n44382 ) | ( n44379 & ~n44384 ) | ( n44382 & ~n44384 ) ;
  assign n44386 = n5310 & ~n22764 ;
  assign n44387 = n44386 ^ n24981 ^ 1'b0 ;
  assign n44388 = n7797 | n12617 ;
  assign n44389 = n17184 ^ n2815 ^ 1'b0 ;
  assign n44390 = n44389 ^ n26475 ^ n7231 ;
  assign n44391 = n44388 & ~n44390 ;
  assign n44392 = ~n6766 & n44391 ;
  assign n44393 = n44392 ^ n5917 ^ 1'b0 ;
  assign n44394 = ( n16629 & n44387 ) | ( n16629 & n44393 ) | ( n44387 & n44393 ) ;
  assign n44395 = n38998 ^ n21700 ^ 1'b0 ;
  assign n44396 = ( n8640 & n35026 ) | ( n8640 & n35144 ) | ( n35026 & n35144 ) ;
  assign n44398 = ( n874 & n4141 ) | ( n874 & n16542 ) | ( n4141 & n16542 ) ;
  assign n44397 = n862 & n1128 ;
  assign n44399 = n44398 ^ n44397 ^ 1'b0 ;
  assign n44400 = n44399 ^ n27719 ^ 1'b0 ;
  assign n44402 = n22191 ^ n21976 ^ n1006 ;
  assign n44401 = n33913 ^ n14520 ^ n10429 ;
  assign n44403 = n44402 ^ n44401 ^ n6983 ;
  assign n44404 = n42317 ^ n25559 ^ 1'b0 ;
  assign n44405 = ( n1631 & n5322 ) | ( n1631 & n7157 ) | ( n5322 & n7157 ) ;
  assign n44406 = ~n23820 & n44405 ;
  assign n44407 = n44406 ^ n27582 ^ 1'b0 ;
  assign n44408 = n24716 ^ n2580 ^ 1'b0 ;
  assign n44409 = n19477 & n44408 ;
  assign n44410 = ( n6811 & n14800 ) | ( n6811 & n23348 ) | ( n14800 & n23348 ) ;
  assign n44411 = n44410 ^ n30616 ^ 1'b0 ;
  assign n44412 = ( n6529 & n27910 ) | ( n6529 & n36755 ) | ( n27910 & n36755 ) ;
  assign n44415 = n11706 ^ x147 ^ 1'b0 ;
  assign n44416 = n26732 | n44415 ;
  assign n44413 = n18648 ^ n1915 ^ 1'b0 ;
  assign n44414 = n44413 ^ n33436 ^ n2996 ;
  assign n44417 = n44416 ^ n44414 ^ n22741 ;
  assign n44418 = n41490 ^ n30820 ^ n30308 ;
  assign n44419 = ( ~n830 & n39756 ) | ( ~n830 & n39877 ) | ( n39756 & n39877 ) ;
  assign n44420 = ( n33360 & ~n37329 ) | ( n33360 & n44419 ) | ( ~n37329 & n44419 ) ;
  assign n44421 = n39149 ^ n14348 ^ n5156 ;
  assign n44424 = ( n15977 & ~n22911 ) | ( n15977 & n42369 ) | ( ~n22911 & n42369 ) ;
  assign n44422 = n6338 | n40555 ;
  assign n44423 = ~n11923 & n44422 ;
  assign n44425 = n44424 ^ n44423 ^ n10292 ;
  assign n44426 = n44425 ^ n30808 ^ 1'b0 ;
  assign n44427 = n24811 & ~n44426 ;
  assign n44428 = n36809 ^ n34063 ^ n21172 ;
  assign n44429 = n27201 ^ n23143 ^ n4059 ;
  assign n44430 = ~x172 & n44429 ;
  assign n44431 = n5385 | n44430 ;
  assign n44432 = n44428 & ~n44431 ;
  assign n44433 = n37923 ^ n11957 ^ n4922 ;
  assign n44434 = n21282 | n44433 ;
  assign n44435 = n42556 ^ n40858 ^ n16646 ;
  assign n44436 = n6404 | n44435 ;
  assign n44437 = n44436 ^ n40527 ^ n24011 ;
  assign n44438 = n22692 & ~n32608 ;
  assign n44439 = n44438 ^ n14301 ^ n6805 ;
  assign n44440 = ( n9853 & n17648 ) | ( n9853 & ~n35991 ) | ( n17648 & ~n35991 ) ;
  assign n44441 = ( n5978 & n21960 ) | ( n5978 & n33766 ) | ( n21960 & n33766 ) ;
  assign n44442 = ( n23403 & ~n26160 ) | ( n23403 & n44441 ) | ( ~n26160 & n44441 ) ;
  assign n44443 = n31446 ^ n14881 ^ n7842 ;
  assign n44444 = n1435 & ~n8945 ;
  assign n44445 = n44444 ^ n9517 ^ 1'b0 ;
  assign n44446 = ( ~n937 & n3190 ) | ( ~n937 & n30696 ) | ( n3190 & n30696 ) ;
  assign n44447 = ( ~x185 & n1138 ) | ( ~x185 & n8431 ) | ( n1138 & n8431 ) ;
  assign n44448 = n44447 ^ n43282 ^ n7100 ;
  assign n44449 = ( n2322 & n10328 ) | ( n2322 & n44448 ) | ( n10328 & n44448 ) ;
  assign n44450 = ( n44445 & n44446 ) | ( n44445 & n44449 ) | ( n44446 & n44449 ) ;
  assign n44451 = ( n5246 & ~n22604 ) | ( n5246 & n35107 ) | ( ~n22604 & n35107 ) ;
  assign n44452 = n44451 ^ n30845 ^ 1'b0 ;
  assign n44453 = n31865 ^ n14286 ^ 1'b0 ;
  assign n44454 = ( x223 & n20026 ) | ( x223 & ~n44453 ) | ( n20026 & ~n44453 ) ;
  assign n44455 = ( ~n13059 & n16336 ) | ( ~n13059 & n16968 ) | ( n16336 & n16968 ) ;
  assign n44456 = n44455 ^ n9795 ^ 1'b0 ;
  assign n44457 = n44454 & n44456 ;
  assign n44458 = n41211 ^ n17537 ^ n536 ;
  assign n44459 = ( n25730 & ~n26281 ) | ( n25730 & n41191 ) | ( ~n26281 & n41191 ) ;
  assign n44460 = n44459 ^ n28833 ^ 1'b0 ;
  assign n44461 = n14684 & ~n26655 ;
  assign n44462 = n44461 ^ n43250 ^ n40875 ;
  assign n44463 = ( n11203 & n15230 ) | ( n11203 & ~n40015 ) | ( n15230 & ~n40015 ) ;
  assign n44464 = n44463 ^ n2668 ^ 1'b0 ;
  assign n44465 = ( n2344 & ~n10768 ) | ( n2344 & n39819 ) | ( ~n10768 & n39819 ) ;
  assign n44466 = ~n5595 & n16974 ;
  assign n44467 = n44466 ^ n13462 ^ 1'b0 ;
  assign n44471 = ( x31 & n8221 ) | ( x31 & ~n10860 ) | ( n8221 & ~n10860 ) ;
  assign n44470 = n32926 ^ n18437 ^ n14130 ;
  assign n44468 = ( n10787 & n10809 ) | ( n10787 & n28429 ) | ( n10809 & n28429 ) ;
  assign n44469 = n44468 ^ n28577 ^ n25915 ;
  assign n44472 = n44471 ^ n44470 ^ n44469 ;
  assign n44473 = n36209 ^ n19871 ^ 1'b0 ;
  assign n44474 = n44472 & n44473 ;
  assign n44476 = ( n6452 & n19776 ) | ( n6452 & n25650 ) | ( n19776 & n25650 ) ;
  assign n44475 = ~n29612 & n41849 ;
  assign n44477 = n44476 ^ n44475 ^ 1'b0 ;
  assign n44478 = ( n7023 & ~n17965 ) | ( n7023 & n33507 ) | ( ~n17965 & n33507 ) ;
  assign n44479 = n35129 ^ n29439 ^ n9683 ;
  assign n44480 = n18023 ^ n4841 ^ 1'b0 ;
  assign n44481 = n17191 ^ n3146 ^ 1'b0 ;
  assign n44484 = ( n1340 & n5214 ) | ( n1340 & ~n13249 ) | ( n5214 & ~n13249 ) ;
  assign n44485 = n44484 ^ n32809 ^ n28054 ;
  assign n44482 = n13677 ^ n6983 ^ 1'b0 ;
  assign n44483 = n41745 | n44482 ;
  assign n44486 = n44485 ^ n44483 ^ n31553 ;
  assign n44487 = n9123 ^ n5615 ^ n835 ;
  assign n44488 = ( n36816 & n41874 ) | ( n36816 & ~n44487 ) | ( n41874 & ~n44487 ) ;
  assign n44489 = n20386 ^ n16954 ^ n12397 ;
  assign n44490 = ( n2492 & n4271 ) | ( n2492 & ~n11890 ) | ( n4271 & ~n11890 ) ;
  assign n44491 = ( n17379 & n20318 ) | ( n17379 & n44490 ) | ( n20318 & n44490 ) ;
  assign n44492 = n17127 | n44491 ;
  assign n44493 = n44492 ^ n3348 ^ 1'b0 ;
  assign n44494 = n14359 ^ n4162 ^ 1'b0 ;
  assign n44495 = n44494 ^ n23026 ^ n12556 ;
  assign n44496 = ( n2217 & ~n3556 ) | ( n2217 & n44495 ) | ( ~n3556 & n44495 ) ;
  assign n44497 = ~n10853 & n44496 ;
  assign n44498 = n44497 ^ x16 ^ 1'b0 ;
  assign n44499 = n25668 & n28935 ;
  assign n44500 = n44499 ^ n33927 ^ 1'b0 ;
  assign n44501 = n44483 ^ n39838 ^ n19297 ;
  assign n44502 = ( n11348 & ~n26146 ) | ( n11348 & n43919 ) | ( ~n26146 & n43919 ) ;
  assign n44503 = ( n7341 & n7851 ) | ( n7341 & ~n44502 ) | ( n7851 & ~n44502 ) ;
  assign n44504 = n34409 ^ n33949 ^ n5046 ;
  assign n44505 = ( n18791 & n20609 ) | ( n18791 & n37535 ) | ( n20609 & n37535 ) ;
  assign n44506 = n29922 ^ n26273 ^ n5084 ;
  assign n44507 = n12803 & n39502 ;
  assign n44508 = ~n44506 & n44507 ;
  assign n44509 = n40326 ^ n39700 ^ 1'b0 ;
  assign n44510 = n32464 & n44509 ;
  assign n44511 = n29319 ^ n11564 ^ n706 ;
  assign n44512 = ( n547 & n8436 ) | ( n547 & ~n44511 ) | ( n8436 & ~n44511 ) ;
  assign n44513 = ( n3131 & n17171 ) | ( n3131 & ~n37567 ) | ( n17171 & ~n37567 ) ;
  assign n44514 = ( ~n44074 & n44512 ) | ( ~n44074 & n44513 ) | ( n44512 & n44513 ) ;
  assign n44520 = n2105 ^ n1020 ^ 1'b0 ;
  assign n44521 = n44520 ^ n35978 ^ n20898 ;
  assign n44517 = ( x154 & n2967 ) | ( x154 & ~n3917 ) | ( n2967 & ~n3917 ) ;
  assign n44518 = ( n14924 & ~n28663 ) | ( n14924 & n44517 ) | ( ~n28663 & n44517 ) ;
  assign n44515 = n11581 ^ n10992 ^ n8255 ;
  assign n44516 = n44515 ^ n41832 ^ 1'b0 ;
  assign n44519 = n44518 ^ n44516 ^ n24887 ;
  assign n44522 = n44521 ^ n44519 ^ n20013 ;
  assign n44531 = ( n1180 & ~n2271 ) | ( n1180 & n16245 ) | ( ~n2271 & n16245 ) ;
  assign n44523 = n2304 | n5414 ;
  assign n44524 = n44523 ^ n25917 ^ 1'b0 ;
  assign n44526 = n20019 ^ n3927 ^ x43 ;
  assign n44525 = n26112 ^ n25498 ^ n22126 ;
  assign n44527 = n44526 ^ n44525 ^ 1'b0 ;
  assign n44528 = n21070 & n44527 ;
  assign n44529 = n44528 ^ n17625 ^ 1'b0 ;
  assign n44530 = ( ~n11746 & n44524 ) | ( ~n11746 & n44529 ) | ( n44524 & n44529 ) ;
  assign n44532 = n44531 ^ n44530 ^ n4701 ;
  assign n44533 = n9714 ^ n3670 ^ n2653 ;
  assign n44534 = n19429 & ~n44533 ;
  assign n44535 = n44534 ^ n13285 ^ 1'b0 ;
  assign n44536 = ( n10043 & n18212 ) | ( n10043 & ~n44535 ) | ( n18212 & ~n44535 ) ;
  assign n44537 = n44536 ^ n22415 ^ n16910 ;
  assign n44538 = ( n13940 & ~n43474 ) | ( n13940 & n44537 ) | ( ~n43474 & n44537 ) ;
  assign n44541 = ( n2255 & n8006 ) | ( n2255 & n10214 ) | ( n8006 & n10214 ) ;
  assign n44539 = n41091 ^ n40634 ^ n16567 ;
  assign n44540 = n20525 & n44539 ;
  assign n44542 = n44541 ^ n44540 ^ 1'b0 ;
  assign n44553 = n35139 & n39654 ;
  assign n44554 = n44553 ^ n8553 ^ 1'b0 ;
  assign n44549 = ( n5875 & ~n12769 ) | ( n5875 & n42452 ) | ( ~n12769 & n42452 ) ;
  assign n44550 = ( ~n3185 & n36094 ) | ( ~n3185 & n40070 ) | ( n36094 & n40070 ) ;
  assign n44551 = n44550 ^ n41031 ^ n13613 ;
  assign n44552 = ( n14773 & n44549 ) | ( n14773 & ~n44551 ) | ( n44549 & ~n44551 ) ;
  assign n44543 = n11609 ^ n6575 ^ n6482 ;
  assign n44544 = n44543 ^ n32872 ^ n4757 ;
  assign n44545 = n9810 | n36142 ;
  assign n44546 = n44544 & ~n44545 ;
  assign n44547 = n44546 ^ n4341 ^ 1'b0 ;
  assign n44548 = n44547 ^ n21279 ^ n4460 ;
  assign n44555 = n44554 ^ n44552 ^ n44548 ;
  assign n44556 = n36987 ^ n20432 ^ n9116 ;
  assign n44557 = n28363 ^ n11874 ^ 1'b0 ;
  assign n44558 = n19511 | n44557 ;
  assign n44559 = ( n10136 & n41439 ) | ( n10136 & n44558 ) | ( n41439 & n44558 ) ;
  assign n44560 = n21256 & n25297 ;
  assign n44561 = n37615 ^ n10390 ^ 1'b0 ;
  assign n44562 = ~n16776 & n44561 ;
  assign n44563 = n44562 ^ n3887 ^ n468 ;
  assign n44564 = ( ~n40461 & n44560 ) | ( ~n40461 & n44563 ) | ( n44560 & n44563 ) ;
  assign n44565 = ( ~n5222 & n40374 ) | ( ~n5222 & n41549 ) | ( n40374 & n41549 ) ;
  assign n44566 = ( ~n7464 & n40365 ) | ( ~n7464 & n44565 ) | ( n40365 & n44565 ) ;
  assign n44567 = n14434 & n44566 ;
  assign n44568 = n44567 ^ n33356 ^ 1'b0 ;
  assign n44569 = n23677 ^ n14702 ^ n4311 ;
  assign n44570 = ( x211 & ~n4012 ) | ( x211 & n36198 ) | ( ~n4012 & n36198 ) ;
  assign n44575 = n14965 ^ n13508 ^ 1'b0 ;
  assign n44576 = n6166 & n44575 ;
  assign n44577 = n44576 ^ n28597 ^ n27710 ;
  assign n44574 = ~n13813 & n14366 ;
  assign n44578 = n44577 ^ n44574 ^ n17541 ;
  assign n44579 = n44578 ^ n41695 ^ n25176 ;
  assign n44571 = n16342 ^ n9496 ^ n7973 ;
  assign n44572 = n44571 ^ n39816 ^ 1'b0 ;
  assign n44573 = n2632 & n44572 ;
  assign n44580 = n44579 ^ n44573 ^ n28954 ;
  assign n44581 = n44447 ^ n37615 ^ n1876 ;
  assign n44582 = n22862 ^ n3866 ^ 1'b0 ;
  assign n44583 = ~n11418 & n44582 ;
  assign n44584 = n44583 ^ n18376 ^ 1'b0 ;
  assign n44585 = n44584 ^ n12470 ^ n7467 ;
  assign n44588 = n40916 ^ n28650 ^ n23655 ;
  assign n44586 = n23959 ^ n2947 ^ 1'b0 ;
  assign n44587 = n8856 & n44586 ;
  assign n44589 = n44588 ^ n44587 ^ n8147 ;
  assign n44590 = n24653 ^ n10835 ^ 1'b0 ;
  assign n44591 = n22359 & n44590 ;
  assign n44592 = n33555 & n44591 ;
  assign n44593 = n37918 | n39998 ;
  assign n44594 = n44593 ^ n16785 ^ 1'b0 ;
  assign n44595 = ( n6446 & ~n16889 ) | ( n6446 & n18228 ) | ( ~n16889 & n18228 ) ;
  assign n44596 = ( n2498 & ~n26747 ) | ( n2498 & n44595 ) | ( ~n26747 & n44595 ) ;
  assign n44597 = n12256 ^ n11847 ^ n4832 ;
  assign n44598 = ( n5653 & n9270 ) | ( n5653 & ~n44597 ) | ( n9270 & ~n44597 ) ;
  assign n44599 = n44598 ^ n14847 ^ n10688 ;
  assign n44600 = n44599 ^ n14409 ^ 1'b0 ;
  assign n44601 = ~n44596 & n44600 ;
  assign n44602 = ( n11814 & n12868 ) | ( n11814 & ~n33082 ) | ( n12868 & ~n33082 ) ;
  assign n44603 = ( n1072 & n2509 ) | ( n1072 & n24969 ) | ( n2509 & n24969 ) ;
  assign n44604 = ( x188 & n21606 ) | ( x188 & ~n44603 ) | ( n21606 & ~n44603 ) ;
  assign n44605 = n41574 ^ n30351 ^ n20139 ;
  assign n44606 = n29643 ^ n13128 ^ n2541 ;
  assign n44607 = ( n21382 & n44605 ) | ( n21382 & n44606 ) | ( n44605 & n44606 ) ;
  assign n44608 = n13269 ^ n12253 ^ n1545 ;
  assign n44609 = n44608 ^ n10663 ^ n4287 ;
  assign n44610 = ( n1262 & ~n8736 ) | ( n1262 & n44609 ) | ( ~n8736 & n44609 ) ;
  assign n44611 = n13345 & ~n44610 ;
  assign n44612 = n36702 & n44611 ;
  assign n44613 = ( n8325 & n42419 ) | ( n8325 & n44612 ) | ( n42419 & n44612 ) ;
  assign n44615 = n17287 ^ n6364 ^ n2691 ;
  assign n44614 = n6720 & n24029 ;
  assign n44616 = n44615 ^ n44614 ^ n15750 ;
  assign n44617 = ( n28931 & n34615 ) | ( n28931 & n42391 ) | ( n34615 & n42391 ) ;
  assign n44618 = n44617 ^ n16256 ^ n10467 ;
  assign n44619 = n13011 & ~n31277 ;
  assign n44620 = n44619 ^ n8808 ^ 1'b0 ;
  assign n44621 = n43051 ^ n1953 ^ 1'b0 ;
  assign n44622 = n36707 & n44621 ;
  assign n44623 = ( n2311 & n24826 ) | ( n2311 & n27970 ) | ( n24826 & n27970 ) ;
  assign n44625 = ( n9009 & ~n9680 ) | ( n9009 & n27711 ) | ( ~n9680 & n27711 ) ;
  assign n44624 = n8856 & n37341 ;
  assign n44626 = n44625 ^ n44624 ^ n42658 ;
  assign n44627 = ( n5528 & n5602 ) | ( n5528 & ~n18735 ) | ( n5602 & ~n18735 ) ;
  assign n44628 = n44627 ^ n14206 ^ n3037 ;
  assign n44629 = n7953 & ~n26681 ;
  assign n44630 = n44629 ^ n36107 ^ n17757 ;
  assign n44632 = n22488 ^ n10429 ^ n5797 ;
  assign n44631 = n29128 ^ n5123 ^ n2620 ;
  assign n44633 = n44632 ^ n44631 ^ n3739 ;
  assign n44634 = n40822 ^ n26083 ^ n1527 ;
  assign n44635 = n1067 | n17278 ;
  assign n44636 = ( ~x6 & n31712 ) | ( ~x6 & n44635 ) | ( n31712 & n44635 ) ;
  assign n44637 = n44636 ^ n19153 ^ n8732 ;
  assign n44638 = n44637 ^ n40426 ^ n27130 ;
  assign n44639 = n13489 & ~n44638 ;
  assign n44640 = n44639 ^ n27888 ^ 1'b0 ;
  assign n44644 = n11965 ^ n7572 ^ n3483 ;
  assign n44645 = n17595 ^ n16122 ^ 1'b0 ;
  assign n44646 = ~n44644 & n44645 ;
  assign n44641 = n15557 ^ n8020 ^ 1'b0 ;
  assign n44642 = ~n17641 & n44641 ;
  assign n44643 = ~n17108 & n44642 ;
  assign n44647 = n44646 ^ n44643 ^ 1'b0 ;
  assign n44652 = ~n10728 & n12818 ;
  assign n44653 = n44652 ^ n41240 ^ 1'b0 ;
  assign n44648 = n432 & n4322 ;
  assign n44649 = n44648 ^ n5780 ^ 1'b0 ;
  assign n44650 = ( ~n6964 & n25510 ) | ( ~n6964 & n44649 ) | ( n25510 & n44649 ) ;
  assign n44651 = n44650 ^ n17591 ^ n15588 ;
  assign n44654 = n44653 ^ n44651 ^ n20892 ;
  assign n44655 = n40778 ^ n21884 ^ n19396 ;
  assign n44656 = ( n15484 & ~n36328 ) | ( n15484 & n44655 ) | ( ~n36328 & n44655 ) ;
  assign n44657 = n27040 ^ n20077 ^ 1'b0 ;
  assign n44658 = ~n2871 & n44657 ;
  assign n44659 = ( ~n2228 & n20990 ) | ( ~n2228 & n44658 ) | ( n20990 & n44658 ) ;
  assign n44660 = n26473 ^ n8609 ^ n1428 ;
  assign n44661 = ( n3965 & ~n4303 ) | ( n3965 & n5983 ) | ( ~n4303 & n5983 ) ;
  assign n44662 = n19541 ^ n9123 ^ 1'b0 ;
  assign n44663 = ( n5458 & ~n44661 ) | ( n5458 & n44662 ) | ( ~n44661 & n44662 ) ;
  assign n44665 = ( n15200 & n17555 ) | ( n15200 & ~n33872 ) | ( n17555 & ~n33872 ) ;
  assign n44666 = ( n23786 & n30943 ) | ( n23786 & ~n44665 ) | ( n30943 & ~n44665 ) ;
  assign n44667 = n44666 ^ n23367 ^ n2662 ;
  assign n44664 = ( n2686 & n22291 ) | ( n2686 & n37300 ) | ( n22291 & n37300 ) ;
  assign n44668 = n44667 ^ n44664 ^ n26887 ;
  assign n44669 = n44668 ^ n16058 ^ 1'b0 ;
  assign n44670 = ( n6762 & ~n31187 ) | ( n6762 & n31939 ) | ( ~n31187 & n31939 ) ;
  assign n44671 = ( n23494 & ~n26885 ) | ( n23494 & n44670 ) | ( ~n26885 & n44670 ) ;
  assign n44672 = n32845 ^ n11632 ^ n7999 ;
  assign n44673 = n1238 | n44672 ;
  assign n44674 = n44671 | n44673 ;
  assign n44675 = n36892 ^ n11405 ^ n7742 ;
  assign n44676 = n18665 & ~n44675 ;
  assign n44677 = n7668 & n44676 ;
  assign n44678 = n15272 ^ n3488 ^ n452 ;
  assign n44679 = n33899 & n44678 ;
  assign n44680 = ( n10443 & n23424 ) | ( n10443 & ~n42641 ) | ( n23424 & ~n42641 ) ;
  assign n44681 = n37477 ^ n17513 ^ n4883 ;
  assign n44682 = n4184 & n18699 ;
  assign n44683 = n25073 ^ n20731 ^ n8546 ;
  assign n44684 = n9318 & ~n44683 ;
  assign n44685 = n28917 ^ n6861 ^ 1'b0 ;
  assign n44686 = n17142 ^ n12213 ^ n6888 ;
  assign n44687 = n44686 ^ n6775 ^ 1'b0 ;
  assign n44688 = ~n19173 & n44687 ;
  assign n44689 = ~n5205 & n44688 ;
  assign n44690 = n17268 ^ n13997 ^ n6995 ;
  assign n44691 = n43942 ^ n23593 ^ n10215 ;
  assign n44692 = n44691 ^ n42439 ^ n28808 ;
  assign n44693 = n33620 ^ n20797 ^ n7514 ;
  assign n44694 = n44693 ^ n11779 ^ n9108 ;
  assign n44695 = ( n5511 & ~n16373 ) | ( n5511 & n44694 ) | ( ~n16373 & n44694 ) ;
  assign n44696 = ( n16513 & n31399 ) | ( n16513 & n43064 ) | ( n31399 & n43064 ) ;
  assign n44697 = n11796 & ~n31705 ;
  assign n44698 = ( n16184 & n22771 ) | ( n16184 & ~n27443 ) | ( n22771 & ~n27443 ) ;
  assign n44699 = ( n4134 & n7521 ) | ( n4134 & ~n16858 ) | ( n7521 & ~n16858 ) ;
  assign n44700 = ( n18392 & n21204 ) | ( n18392 & ~n28706 ) | ( n21204 & ~n28706 ) ;
  assign n44701 = n37130 | n44700 ;
  assign n44702 = n44701 ^ n7816 ^ 1'b0 ;
  assign n44707 = ( n2842 & n8501 ) | ( n2842 & n17922 ) | ( n8501 & n17922 ) ;
  assign n44708 = ( n12723 & n21225 ) | ( n12723 & ~n44707 ) | ( n21225 & ~n44707 ) ;
  assign n44705 = n623 & ~n12115 ;
  assign n44706 = ( n40778 & n41591 ) | ( n40778 & ~n44705 ) | ( n41591 & ~n44705 ) ;
  assign n44709 = n44708 ^ n44706 ^ n21951 ;
  assign n44703 = ~n19885 & n34449 ;
  assign n44704 = ~n28959 & n44703 ;
  assign n44710 = n44709 ^ n44704 ^ n10254 ;
  assign n44711 = n4407 & ~n44710 ;
  assign n44712 = n44711 ^ n27423 ^ 1'b0 ;
  assign n44713 = n37833 ^ n14240 ^ n8728 ;
  assign n44714 = ( n4890 & n9874 ) | ( n4890 & ~n44713 ) | ( n9874 & ~n44713 ) ;
  assign n44715 = n8199 ^ n1306 ^ 1'b0 ;
  assign n44716 = n18312 ^ n4934 ^ n2585 ;
  assign n44717 = ( n35751 & ~n44715 ) | ( n35751 & n44716 ) | ( ~n44715 & n44716 ) ;
  assign n44718 = ( n18290 & n27286 ) | ( n18290 & ~n33612 ) | ( n27286 & ~n33612 ) ;
  assign n44719 = n44718 ^ n26183 ^ n16578 ;
  assign n44720 = ( n11876 & ~n13732 ) | ( n11876 & n28804 ) | ( ~n13732 & n28804 ) ;
  assign n44721 = n16126 & ~n27417 ;
  assign n44722 = ( n9203 & n44720 ) | ( n9203 & n44721 ) | ( n44720 & n44721 ) ;
  assign n44723 = n2803 ^ n1912 ^ 1'b0 ;
  assign n44724 = n27218 ^ n3074 ^ 1'b0 ;
  assign n44725 = n44724 ^ n14430 ^ n8368 ;
  assign n44726 = n44723 & n44725 ;
  assign n44727 = n9466 & ~n33536 ;
  assign n44728 = ( n4853 & ~n6587 ) | ( n4853 & n14947 ) | ( ~n6587 & n14947 ) ;
  assign n44729 = n13091 | n44728 ;
  assign n44730 = n17276 ^ n9581 ^ n2036 ;
  assign n44731 = n2213 & n5461 ;
  assign n44732 = n44731 ^ n26586 ^ 1'b0 ;
  assign n44733 = n22537 & ~n44732 ;
  assign n44734 = n26469 ^ n7090 ^ 1'b0 ;
  assign n44735 = n40481 ^ n27298 ^ n1069 ;
  assign n44736 = ( n26806 & n44031 ) | ( n26806 & ~n44735 ) | ( n44031 & ~n44735 ) ;
  assign n44737 = ( n7484 & n15708 ) | ( n7484 & ~n17344 ) | ( n15708 & ~n17344 ) ;
  assign n44738 = n27116 ^ n18660 ^ n2599 ;
  assign n44739 = n11619 & ~n27878 ;
  assign n44740 = n44739 ^ n44595 ^ 1'b0 ;
  assign n44741 = ( n25232 & n31963 ) | ( n25232 & n44740 ) | ( n31963 & n44740 ) ;
  assign n44742 = n12929 ^ n10359 ^ x7 ;
  assign n44743 = ~n13865 & n16055 ;
  assign n44744 = n44743 ^ n8686 ^ 1'b0 ;
  assign n44745 = ( ~n17814 & n17987 ) | ( ~n17814 & n27010 ) | ( n17987 & n27010 ) ;
  assign n44746 = n31141 ^ n2372 ^ n1405 ;
  assign n44747 = ( ~n410 & n4768 ) | ( ~n410 & n37920 ) | ( n4768 & n37920 ) ;
  assign n44748 = ( ~x236 & n6546 ) | ( ~x236 & n44747 ) | ( n6546 & n44747 ) ;
  assign n44751 = n10272 | n37496 ;
  assign n44752 = n44751 ^ n19302 ^ n14630 ;
  assign n44749 = ( n10435 & ~n19815 ) | ( n10435 & n28286 ) | ( ~n19815 & n28286 ) ;
  assign n44750 = ( n5670 & n39375 ) | ( n5670 & n44749 ) | ( n39375 & n44749 ) ;
  assign n44753 = n44752 ^ n44750 ^ n10344 ;
  assign n44754 = ( n17877 & n29354 ) | ( n17877 & ~n44753 ) | ( n29354 & ~n44753 ) ;
  assign n44755 = n25940 ^ n7902 ^ x152 ;
  assign n44756 = n44755 ^ n35352 ^ n31315 ;
  assign n44757 = n44756 ^ n19305 ^ n12296 ;
  assign n44758 = n44757 ^ n40440 ^ n29958 ;
  assign n44759 = n3337 | n4914 ;
  assign n44760 = n11079 | n44759 ;
  assign n44761 = n5427 & ~n23998 ;
  assign n44762 = n3300 & n44761 ;
  assign n44763 = n44762 ^ n28216 ^ n23136 ;
  assign n44764 = n28442 ^ n21858 ^ n16858 ;
  assign n44765 = n11067 | n44764 ;
  assign n44770 = ( n2507 & ~n4683 ) | ( n2507 & n6619 ) | ( ~n4683 & n6619 ) ;
  assign n44771 = ( ~n5195 & n38215 ) | ( ~n5195 & n44770 ) | ( n38215 & n44770 ) ;
  assign n44768 = n26012 ^ n17203 ^ n12560 ;
  assign n44766 = ( n6931 & ~n8142 ) | ( n6931 & n18695 ) | ( ~n8142 & n18695 ) ;
  assign n44767 = ( n1606 & n32226 ) | ( n1606 & n44766 ) | ( n32226 & n44766 ) ;
  assign n44769 = n44768 ^ n44767 ^ n30285 ;
  assign n44772 = n44771 ^ n44769 ^ n34498 ;
  assign n44773 = ( n29175 & ~n34018 ) | ( n29175 & n36734 ) | ( ~n34018 & n36734 ) ;
  assign n44774 = n29108 ^ n13387 ^ n12926 ;
  assign n44775 = n44774 ^ n33203 ^ n14981 ;
  assign n44776 = ( ~n13524 & n34774 ) | ( ~n13524 & n40664 ) | ( n34774 & n40664 ) ;
  assign n44777 = ( n17372 & n20744 ) | ( n17372 & ~n32702 ) | ( n20744 & ~n32702 ) ;
  assign n44778 = ( ~n1470 & n14849 ) | ( ~n1470 & n33226 ) | ( n14849 & n33226 ) ;
  assign n44779 = ( n13176 & n35375 ) | ( n13176 & n44778 ) | ( n35375 & n44778 ) ;
  assign n44780 = n44779 ^ n799 ^ 1'b0 ;
  assign n44781 = n7306 & ~n44780 ;
  assign n44782 = n44777 & n44781 ;
  assign n44783 = n32476 ^ n19962 ^ n15277 ;
  assign n44784 = n9060 | n22432 ;
  assign n44785 = n44784 ^ n41835 ^ 1'b0 ;
  assign n44786 = n30366 ^ n11980 ^ n5029 ;
  assign n44787 = ( n5716 & ~n8593 ) | ( n5716 & n40281 ) | ( ~n8593 & n40281 ) ;
  assign n44788 = n10110 & n44787 ;
  assign n44789 = ~n44786 & n44788 ;
  assign n44790 = ( n2469 & n2582 ) | ( n2469 & ~n8635 ) | ( n2582 & ~n8635 ) ;
  assign n44791 = ( n13994 & n14317 ) | ( n13994 & n14406 ) | ( n14317 & n14406 ) ;
  assign n44792 = ( n29935 & n44790 ) | ( n29935 & n44791 ) | ( n44790 & n44791 ) ;
  assign n44793 = ~n1958 & n23189 ;
  assign n44794 = ~n44792 & n44793 ;
  assign n44795 = ( x197 & ~n1092 ) | ( x197 & n4513 ) | ( ~n1092 & n4513 ) ;
  assign n44796 = n44795 ^ n26533 ^ n18325 ;
  assign n44797 = n44796 ^ n10465 ^ 1'b0 ;
  assign n44798 = ( n15500 & ~n25684 ) | ( n15500 & n37325 ) | ( ~n25684 & n37325 ) ;
  assign n44799 = n38236 ^ n10580 ^ 1'b0 ;
  assign n44800 = n5554 | n7037 ;
  assign n44801 = ( n8523 & n15876 ) | ( n8523 & ~n44800 ) | ( n15876 & ~n44800 ) ;
  assign n44802 = ( ~n2447 & n5860 ) | ( ~n2447 & n10900 ) | ( n5860 & n10900 ) ;
  assign n44803 = n16003 & n44802 ;
  assign n44804 = n44803 ^ n33119 ^ 1'b0 ;
  assign n44805 = n18424 & n19894 ;
  assign n44806 = n44805 ^ n35643 ^ n16966 ;
  assign n44807 = n5922 & ~n19765 ;
  assign n44808 = n44807 ^ n28872 ^ 1'b0 ;
  assign n44809 = n9519 ^ n4520 ^ 1'b0 ;
  assign n44810 = ( ~n5491 & n24858 ) | ( ~n5491 & n34596 ) | ( n24858 & n34596 ) ;
  assign n44811 = n2391 | n5522 ;
  assign n44812 = ( n7513 & n34899 ) | ( n7513 & n36239 ) | ( n34899 & n36239 ) ;
  assign n44813 = n40266 ^ n28359 ^ n16471 ;
  assign n44814 = ( n6383 & ~n10467 ) | ( n6383 & n11360 ) | ( ~n10467 & n11360 ) ;
  assign n44815 = n44814 ^ n38023 ^ n14468 ;
  assign n44816 = ( n6330 & n44813 ) | ( n6330 & n44815 ) | ( n44813 & n44815 ) ;
  assign n44817 = n23538 ^ n17768 ^ n12897 ;
  assign n44818 = n25023 ^ n20762 ^ 1'b0 ;
  assign n44819 = n21850 & ~n44818 ;
  assign n44820 = n36046 ^ n32849 ^ n18952 ;
  assign n44821 = ( n5733 & ~n44819 ) | ( n5733 & n44820 ) | ( ~n44819 & n44820 ) ;
  assign n44822 = ( ~n2135 & n4694 ) | ( ~n2135 & n37556 ) | ( n4694 & n37556 ) ;
  assign n44823 = ( n2877 & n12103 ) | ( n2877 & n24846 ) | ( n12103 & n24846 ) ;
  assign n44824 = n10915 & ~n44823 ;
  assign n44825 = n44824 ^ n37095 ^ 1'b0 ;
  assign n44826 = n33807 ^ n20132 ^ 1'b0 ;
  assign n44827 = n44825 & n44826 ;
  assign n44828 = n4218 & n9474 ;
  assign n44829 = ~n44079 & n44828 ;
  assign n44830 = ( n10558 & n17306 ) | ( n10558 & n17621 ) | ( n17306 & n17621 ) ;
  assign n44831 = ( n5303 & n13385 ) | ( n5303 & ~n44830 ) | ( n13385 & ~n44830 ) ;
  assign n44832 = n22645 & n28751 ;
  assign n44833 = ~n44831 & n44832 ;
  assign n44834 = ( n26164 & ~n26748 ) | ( n26164 & n37925 ) | ( ~n26748 & n37925 ) ;
  assign n44835 = n44834 ^ n34431 ^ n1294 ;
  assign n44836 = n44835 ^ n37670 ^ n2825 ;
  assign n44837 = n41431 ^ n38594 ^ n2830 ;
  assign n44838 = ( n11269 & n11654 ) | ( n11269 & n18537 ) | ( n11654 & n18537 ) ;
  assign n44839 = n41285 ^ n4385 ^ 1'b0 ;
  assign n44840 = n18699 & ~n30204 ;
  assign n44841 = n44840 ^ n43983 ^ 1'b0 ;
  assign n44842 = n2504 & ~n4689 ;
  assign n44843 = n44842 ^ n15180 ^ 1'b0 ;
  assign n44844 = ( n10308 & n28270 ) | ( n10308 & ~n42122 ) | ( n28270 & ~n42122 ) ;
  assign n44845 = n44844 ^ n41621 ^ n7169 ;
  assign n44846 = n26000 ^ n12193 ^ 1'b0 ;
  assign n44847 = ( ~n12101 & n16152 ) | ( ~n12101 & n34913 ) | ( n16152 & n34913 ) ;
  assign n44848 = ( n25326 & ~n30731 ) | ( n25326 & n37550 ) | ( ~n30731 & n37550 ) ;
  assign n44849 = n23254 ^ n704 ^ 1'b0 ;
  assign n44850 = n12113 | n16556 ;
  assign n44851 = n41157 & ~n44850 ;
  assign n44852 = n27343 ^ n17406 ^ n10439 ;
  assign n44853 = n15804 ^ n14274 ^ 1'b0 ;
  assign n44854 = ( n22697 & n29700 ) | ( n22697 & ~n39428 ) | ( n29700 & ~n39428 ) ;
  assign n44855 = ( ~n8432 & n8688 ) | ( ~n8432 & n26682 ) | ( n8688 & n26682 ) ;
  assign n44856 = ( ~n21515 & n32621 ) | ( ~n21515 & n44855 ) | ( n32621 & n44855 ) ;
  assign n44857 = ( ~n402 & n4420 ) | ( ~n402 & n6001 ) | ( n4420 & n6001 ) ;
  assign n44858 = ~n5199 & n24634 ;
  assign n44859 = ~n44857 & n44858 ;
  assign n44860 = n29350 & n42714 ;
  assign n44861 = n44860 ^ n4628 ^ 1'b0 ;
  assign n44862 = ( n27246 & n30412 ) | ( n27246 & n44366 ) | ( n30412 & n44366 ) ;
  assign n44863 = n44862 ^ n20232 ^ n8538 ;
  assign n44864 = ( n9270 & n21346 ) | ( n9270 & n24243 ) | ( n21346 & n24243 ) ;
  assign n44865 = ( n4117 & n39459 ) | ( n4117 & n44864 ) | ( n39459 & n44864 ) ;
  assign n44867 = n36486 ^ n25907 ^ n4229 ;
  assign n44868 = ( ~n3509 & n3980 ) | ( ~n3509 & n44867 ) | ( n3980 & n44867 ) ;
  assign n44866 = n42393 ^ n26235 ^ n19357 ;
  assign n44869 = n44868 ^ n44866 ^ n16838 ;
  assign n44870 = ( n1534 & ~n17208 ) | ( n1534 & n34928 ) | ( ~n17208 & n34928 ) ;
  assign n44871 = ( n1501 & n10919 ) | ( n1501 & ~n11400 ) | ( n10919 & ~n11400 ) ;
  assign n44872 = n41691 ^ n13881 ^ n932 ;
  assign n44873 = n44872 ^ n20092 ^ n15426 ;
  assign n44874 = n39273 ^ n24391 ^ n23041 ;
  assign n44875 = n44874 ^ n25711 ^ n9944 ;
  assign n44876 = n23149 ^ n3206 ^ n977 ;
  assign n44877 = n44876 ^ n44709 ^ n27265 ;
  assign n44878 = n17244 & n37687 ;
  assign n44879 = ~n22656 & n44878 ;
  assign n44880 = ( n258 & n30035 ) | ( n258 & ~n39267 ) | ( n30035 & ~n39267 ) ;
  assign n44881 = ~n16494 & n26747 ;
  assign n44882 = n44880 & n44881 ;
  assign n44883 = n522 & ~n10706 ;
  assign n44884 = n41421 & ~n44883 ;
  assign n44885 = n38020 & n44884 ;
  assign n44886 = n44885 ^ n4079 ^ 1'b0 ;
  assign n44889 = n16374 ^ n15399 ^ n294 ;
  assign n44887 = n23102 & n24881 ;
  assign n44888 = n44887 ^ n20747 ^ 1'b0 ;
  assign n44890 = n44889 ^ n44888 ^ n32729 ;
  assign n44891 = ~n8390 & n20780 ;
  assign n44892 = n15977 & n44891 ;
  assign n44893 = n14922 & n44892 ;
  assign n44894 = n38243 ^ n28536 ^ n6454 ;
  assign n44895 = n44894 ^ n19222 ^ n9036 ;
  assign n44897 = ( n16725 & n31385 ) | ( n16725 & n32556 ) | ( n31385 & n32556 ) ;
  assign n44896 = n32259 ^ n12987 ^ n3384 ;
  assign n44898 = n44897 ^ n44896 ^ n34948 ;
  assign n44899 = ( n4585 & n29561 ) | ( n4585 & n44898 ) | ( n29561 & n44898 ) ;
  assign n44900 = ( ~n10833 & n11145 ) | ( ~n10833 & n17831 ) | ( n11145 & n17831 ) ;
  assign n44901 = n21892 ^ n2946 ^ 1'b0 ;
  assign n44902 = n44901 ^ n32524 ^ n12419 ;
  assign n44903 = n977 & n44902 ;
  assign n44904 = n44903 ^ n38840 ^ 1'b0 ;
  assign n44905 = ( n6026 & ~n16161 ) | ( n6026 & n44904 ) | ( ~n16161 & n44904 ) ;
  assign n44906 = n26051 & ~n44905 ;
  assign n44907 = ( n10830 & ~n11942 ) | ( n10830 & n24125 ) | ( ~n11942 & n24125 ) ;
  assign n44908 = ~n34253 & n44907 ;
  assign n44909 = n44908 ^ n25796 ^ 1'b0 ;
  assign n44910 = n29803 ^ n18129 ^ 1'b0 ;
  assign n44911 = ( n9022 & n10225 ) | ( n9022 & n19927 ) | ( n10225 & n19927 ) ;
  assign n44912 = ( ~x170 & n361 ) | ( ~x170 & n21702 ) | ( n361 & n21702 ) ;
  assign n44913 = n44912 ^ n14584 ^ n475 ;
  assign n44914 = ( n4775 & ~n23348 ) | ( n4775 & n23891 ) | ( ~n23348 & n23891 ) ;
  assign n44915 = n6169 ^ n2871 ^ n1104 ;
  assign n44916 = ( ~n3157 & n23375 ) | ( ~n3157 & n44915 ) | ( n23375 & n44915 ) ;
  assign n44917 = n18091 | n39896 ;
  assign n44918 = n44917 ^ n4628 ^ n4034 ;
  assign n44919 = n588 | n28311 ;
  assign n44920 = n22709 | n44919 ;
  assign n44922 = ( n1726 & n4301 ) | ( n1726 & n6857 ) | ( n4301 & n6857 ) ;
  assign n44923 = n5371 & n44922 ;
  assign n44921 = n2428 & ~n25087 ;
  assign n44924 = n44923 ^ n44921 ^ 1'b0 ;
  assign n44925 = ~n28868 & n31763 ;
  assign n44926 = n44925 ^ n34949 ^ n27782 ;
  assign n44927 = ( n18065 & n25338 ) | ( n18065 & ~n44022 ) | ( n25338 & ~n44022 ) ;
  assign n44928 = n31380 ^ n13013 ^ n11301 ;
  assign n44929 = n11525 ^ n11309 ^ n7656 ;
  assign n44930 = n44929 ^ n26652 ^ 1'b0 ;
  assign n44931 = ~n26994 & n44930 ;
  assign n44932 = ( ~n4830 & n36022 ) | ( ~n4830 & n38211 ) | ( n36022 & n38211 ) ;
  assign n44933 = n19408 ^ n3254 ^ 1'b0 ;
  assign n44934 = n18840 ^ n18403 ^ 1'b0 ;
  assign n44935 = ( n10728 & n44933 ) | ( n10728 & n44934 ) | ( n44933 & n44934 ) ;
  assign n44936 = ( n1501 & n1547 ) | ( n1501 & n24356 ) | ( n1547 & n24356 ) ;
  assign n44937 = n44936 ^ n21663 ^ n3678 ;
  assign n44938 = ( n7836 & n8481 ) | ( n7836 & ~n39659 ) | ( n8481 & ~n39659 ) ;
  assign n44939 = n23808 ^ n14695 ^ n2171 ;
  assign n44940 = n39060 ^ n17541 ^ 1'b0 ;
  assign n44943 = ( n1175 & n3835 ) | ( n1175 & n8797 ) | ( n3835 & n8797 ) ;
  assign n44941 = n7755 & n11684 ;
  assign n44942 = n44941 ^ n3049 ^ 1'b0 ;
  assign n44944 = n44943 ^ n44942 ^ n24351 ;
  assign n44945 = n44944 ^ n24033 ^ 1'b0 ;
  assign n44946 = n24910 | n37101 ;
  assign n44947 = n44946 ^ n33093 ^ n32091 ;
  assign n44948 = n44310 ^ n26903 ^ n9749 ;
  assign n44949 = n5041 & ~n17470 ;
  assign n44950 = x175 & n22056 ;
  assign n44951 = ~n43834 & n44950 ;
  assign n44952 = ( n6965 & ~n17454 ) | ( n6965 & n44951 ) | ( ~n17454 & n44951 ) ;
  assign n44953 = ( n2150 & n36902 ) | ( n2150 & ~n44952 ) | ( n36902 & ~n44952 ) ;
  assign n44954 = n24087 ^ n17721 ^ n10901 ;
  assign n44955 = n14511 & ~n44954 ;
  assign n44956 = ( n8025 & n8638 ) | ( n8025 & n44955 ) | ( n8638 & n44955 ) ;
  assign n44957 = ( n14239 & ~n14956 ) | ( n14239 & n23513 ) | ( ~n14956 & n23513 ) ;
  assign n44958 = ( n794 & ~n5310 ) | ( n794 & n41616 ) | ( ~n5310 & n41616 ) ;
  assign n44959 = ( n16202 & n23398 ) | ( n16202 & n44958 ) | ( n23398 & n44958 ) ;
  assign n44960 = n27506 ^ n4607 ^ 1'b0 ;
  assign n44961 = n18104 & ~n44960 ;
  assign n44962 = x59 & n1623 ;
  assign n44963 = ( n32169 & n39688 ) | ( n32169 & n44962 ) | ( n39688 & n44962 ) ;
  assign n44970 = ( n6645 & n8390 ) | ( n6645 & n23036 ) | ( n8390 & n23036 ) ;
  assign n44969 = ( n2565 & n5754 ) | ( n2565 & ~n9945 ) | ( n5754 & ~n9945 ) ;
  assign n44964 = n19564 ^ n16750 ^ n12985 ;
  assign n44965 = n10216 | n13161 ;
  assign n44966 = n2586 & ~n44965 ;
  assign n44967 = n6434 & ~n44966 ;
  assign n44968 = n44964 & n44967 ;
  assign n44971 = n44970 ^ n44969 ^ n44968 ;
  assign n44972 = n44971 ^ n12801 ^ 1'b0 ;
  assign n44973 = n44972 ^ n33361 ^ n13474 ;
  assign n44974 = n2906 & ~n43539 ;
  assign n44975 = n2830 & n44974 ;
  assign n44976 = ( n1879 & ~n6746 ) | ( n1879 & n28997 ) | ( ~n6746 & n28997 ) ;
  assign n44977 = n44976 ^ n18492 ^ 1'b0 ;
  assign n44978 = ~n44975 & n44977 ;
  assign n44979 = n44978 ^ n44605 ^ n810 ;
  assign n44980 = n34550 ^ n23637 ^ n2589 ;
  assign n44981 = n44980 ^ n34612 ^ n11292 ;
  assign n44982 = ( n18585 & n35677 ) | ( n18585 & ~n44981 ) | ( n35677 & ~n44981 ) ;
  assign n44983 = n19633 ^ n10642 ^ n5814 ;
  assign n44987 = n10541 & ~n14832 ;
  assign n44988 = n44987 ^ n33748 ^ 1'b0 ;
  assign n44984 = ( n5430 & ~n24539 ) | ( n5430 & n39845 ) | ( ~n24539 & n39845 ) ;
  assign n44985 = n44984 ^ n20944 ^ 1'b0 ;
  assign n44986 = ( ~n26187 & n39496 ) | ( ~n26187 & n44985 ) | ( n39496 & n44985 ) ;
  assign n44989 = n44988 ^ n44986 ^ n25851 ;
  assign n44990 = n37677 | n43889 ;
  assign n44991 = n44990 ^ n25644 ^ 1'b0 ;
  assign n44992 = n7139 & n12199 ;
  assign n44993 = n5542 & ~n44992 ;
  assign n44994 = n18802 ^ n2688 ^ 1'b0 ;
  assign n44995 = n10952 & ~n44994 ;
  assign n44996 = n44995 ^ n19795 ^ n15391 ;
  assign n44997 = ( ~n11458 & n44993 ) | ( ~n11458 & n44996 ) | ( n44993 & n44996 ) ;
  assign n44998 = ( ~n15419 & n22870 ) | ( ~n15419 & n42115 ) | ( n22870 & n42115 ) ;
  assign n44999 = ( n556 & n39910 ) | ( n556 & n44998 ) | ( n39910 & n44998 ) ;
  assign n45000 = n32678 ^ n11754 ^ 1'b0 ;
  assign n45002 = n36576 ^ n24269 ^ n5010 ;
  assign n45001 = n37767 ^ n18223 ^ n5522 ;
  assign n45003 = n45002 ^ n45001 ^ n29618 ;
  assign n45004 = n42445 ^ n41746 ^ n16380 ;
  assign n45005 = n12064 ^ n11660 ^ n1106 ;
  assign n45006 = n45005 ^ n43470 ^ n4692 ;
  assign n45007 = n38584 ^ n2481 ^ 1'b0 ;
  assign n45008 = n1446 & n45007 ;
  assign n45009 = ( n22428 & n23191 ) | ( n22428 & n37824 ) | ( n23191 & n37824 ) ;
  assign n45010 = n45009 ^ n24917 ^ 1'b0 ;
  assign n45011 = n354 & ~n45010 ;
  assign n45012 = ( n7054 & ~n10882 ) | ( n7054 & n16466 ) | ( ~n10882 & n16466 ) ;
  assign n45013 = n45012 ^ n12412 ^ 1'b0 ;
  assign n45014 = n45013 ^ n37736 ^ n34948 ;
  assign n45015 = ~n5178 & n41468 ;
  assign n45016 = n15179 ^ n4708 ^ n2258 ;
  assign n45017 = n39762 ^ n36937 ^ 1'b0 ;
  assign n45018 = n7877 | n45017 ;
  assign n45019 = ( n19823 & n25714 ) | ( n19823 & ~n45018 ) | ( n25714 & ~n45018 ) ;
  assign n45020 = n45019 ^ n18780 ^ n711 ;
  assign n45023 = n29962 ^ n20123 ^ n5993 ;
  assign n45024 = ( n14667 & n15677 ) | ( n14667 & ~n45023 ) | ( n15677 & ~n45023 ) ;
  assign n45021 = n4904 & ~n29643 ;
  assign n45022 = n10877 & ~n45021 ;
  assign n45025 = n45024 ^ n45022 ^ n10326 ;
  assign n45026 = ~n20797 & n31072 ;
  assign n45027 = ( n19507 & ~n41285 ) | ( n19507 & n45026 ) | ( ~n41285 & n45026 ) ;
  assign n45028 = n45027 ^ n25595 ^ n16379 ;
  assign n45029 = n39235 ^ n29596 ^ n970 ;
  assign n45031 = n14795 ^ n7292 ^ n3480 ;
  assign n45030 = n18024 ^ n6541 ^ 1'b0 ;
  assign n45032 = n45031 ^ n45030 ^ n1870 ;
  assign n45035 = n11345 ^ n597 ^ x247 ;
  assign n45036 = n45035 ^ n32363 ^ n23495 ;
  assign n45033 = n38198 ^ n6744 ^ 1'b0 ;
  assign n45034 = n26539 | n45033 ;
  assign n45037 = n45036 ^ n45034 ^ 1'b0 ;
  assign n45038 = n33219 ^ n8808 ^ 1'b0 ;
  assign n45039 = n15917 & ~n45038 ;
  assign n45040 = ( n1182 & n26777 ) | ( n1182 & n44830 ) | ( n26777 & n44830 ) ;
  assign n45041 = n45040 ^ n9176 ^ n2511 ;
  assign n45042 = n20244 & n37500 ;
  assign n45043 = n45041 & n45042 ;
  assign n45044 = ( ~x26 & n19953 ) | ( ~x26 & n30043 ) | ( n19953 & n30043 ) ;
  assign n45045 = ( n17899 & ~n45043 ) | ( n17899 & n45044 ) | ( ~n45043 & n45044 ) ;
  assign n45046 = ( ~n11061 & n17492 ) | ( ~n11061 & n45045 ) | ( n17492 & n45045 ) ;
  assign n45047 = ( n12463 & n30565 ) | ( n12463 & ~n44290 ) | ( n30565 & ~n44290 ) ;
  assign n45048 = n7959 | n10067 ;
  assign n45049 = n25576 & ~n45048 ;
  assign n45050 = ( ~n31402 & n42095 ) | ( ~n31402 & n45049 ) | ( n42095 & n45049 ) ;
  assign n45051 = ( n587 & n22561 ) | ( n587 & n32267 ) | ( n22561 & n32267 ) ;
  assign n45052 = n45051 ^ n39267 ^ n3713 ;
  assign n45053 = ( n7384 & n12474 ) | ( n7384 & ~n29769 ) | ( n12474 & ~n29769 ) ;
  assign n45054 = ( n1195 & ~n4873 ) | ( n1195 & n7544 ) | ( ~n4873 & n7544 ) ;
  assign n45055 = n44610 ^ n35540 ^ n2476 ;
  assign n45056 = ( n4441 & n4837 ) | ( n4441 & ~n27757 ) | ( n4837 & ~n27757 ) ;
  assign n45057 = n45056 ^ n43088 ^ n33814 ;
  assign n45058 = n10882 ^ n1496 ^ x70 ;
  assign n45059 = ( n2388 & n13394 ) | ( n2388 & n25813 ) | ( n13394 & n25813 ) ;
  assign n45060 = n45059 ^ n28054 ^ 1'b0 ;
  assign n45061 = n18477 & n45060 ;
  assign n45062 = n31236 ^ n17117 ^ 1'b0 ;
  assign n45063 = n45061 & ~n45062 ;
  assign n45064 = n1246 & n7860 ;
  assign n45065 = n32564 & n45064 ;
  assign n45066 = n7750 & n13503 ;
  assign n45067 = n45066 ^ n29372 ^ 1'b0 ;
  assign n45068 = n33372 | n42433 ;
  assign n45069 = n14893 ^ n6579 ^ 1'b0 ;
  assign n45070 = n45069 ^ n41538 ^ n19359 ;
  assign n45071 = n45070 ^ n18917 ^ n3910 ;
  assign n45072 = n19552 ^ n12897 ^ n10688 ;
  assign n45073 = n45072 ^ n22597 ^ n18811 ;
  assign n45074 = n35292 ^ n2110 ^ 1'b0 ;
  assign n45075 = n31634 | n45074 ;
  assign n45076 = ( ~n1435 & n5739 ) | ( ~n1435 & n45075 ) | ( n5739 & n45075 ) ;
  assign n45077 = ( ~n1144 & n44713 ) | ( ~n1144 & n45076 ) | ( n44713 & n45076 ) ;
  assign n45078 = n28552 ^ n6125 ^ n6027 ;
  assign n45079 = n39063 ^ n11038 ^ n6951 ;
  assign n45080 = n16182 ^ n5523 ^ 1'b0 ;
  assign n45081 = n45079 | n45080 ;
  assign n45082 = n44024 ^ n32778 ^ n7689 ;
  assign n45083 = ( n7232 & n7419 ) | ( n7232 & n13671 ) | ( n7419 & n13671 ) ;
  assign n45084 = ( n15742 & n38036 ) | ( n15742 & n45083 ) | ( n38036 & n45083 ) ;
  assign n45085 = n45084 ^ n11508 ^ n5036 ;
  assign n45086 = ( n32987 & ~n45082 ) | ( n32987 & n45085 ) | ( ~n45082 & n45085 ) ;
  assign n45087 = ( n3642 & n9816 ) | ( n3642 & n18236 ) | ( n9816 & n18236 ) ;
  assign n45088 = ( ~n19355 & n35822 ) | ( ~n19355 & n39465 ) | ( n35822 & n39465 ) ;
  assign n45089 = ( ~n8296 & n28128 ) | ( ~n8296 & n41824 ) | ( n28128 & n41824 ) ;
  assign n45091 = n3370 & n4130 ;
  assign n45090 = ( n13481 & n21245 ) | ( n13481 & n27016 ) | ( n21245 & n27016 ) ;
  assign n45092 = n45091 ^ n45090 ^ n9479 ;
  assign n45093 = n38150 ^ n7980 ^ 1'b0 ;
  assign n45094 = ( n761 & n5634 ) | ( n761 & ~n30984 ) | ( n5634 & ~n30984 ) ;
  assign n45095 = ( n8368 & n14716 ) | ( n8368 & ~n45094 ) | ( n14716 & ~n45094 ) ;
  assign n45096 = n45095 ^ n26083 ^ 1'b0 ;
  assign n45097 = n29829 ^ n18280 ^ n14282 ;
  assign n45098 = n34899 ^ n9951 ^ n861 ;
  assign n45099 = n45098 ^ n26925 ^ n12746 ;
  assign n45100 = n45097 & n45099 ;
  assign n45101 = n42788 ^ n32474 ^ n26200 ;
  assign n45102 = ~n3018 & n12838 ;
  assign n45103 = ~n45101 & n45102 ;
  assign n45104 = ~n2688 & n31547 ;
  assign n45105 = n45104 ^ n3786 ^ 1'b0 ;
  assign n45106 = n12314 ^ n2036 ^ n1511 ;
  assign n45107 = n45106 ^ n3402 ^ n3384 ;
  assign n45108 = ( n4859 & n11249 ) | ( n4859 & ~n45107 ) | ( n11249 & ~n45107 ) ;
  assign n45109 = n45105 & n45108 ;
  assign n45110 = n45109 ^ n23259 ^ n20580 ;
  assign n45111 = n13380 & ~n24029 ;
  assign n45112 = n7489 & n23049 ;
  assign n45113 = n45112 ^ n5346 ^ 1'b0 ;
  assign n45114 = n33904 ^ n16995 ^ 1'b0 ;
  assign n45115 = ( n10726 & n45113 ) | ( n10726 & n45114 ) | ( n45113 & n45114 ) ;
  assign n45116 = n31320 ^ n29603 ^ n7075 ;
  assign n45117 = ( ~n24014 & n29445 ) | ( ~n24014 & n45116 ) | ( n29445 & n45116 ) ;
  assign n45118 = ( n6358 & ~n45115 ) | ( n6358 & n45117 ) | ( ~n45115 & n45117 ) ;
  assign n45119 = n270 & ~n16712 ;
  assign n45120 = n45119 ^ n15574 ^ 1'b0 ;
  assign n45121 = n8241 & ~n45120 ;
  assign n45122 = n32608 ^ n30204 ^ n743 ;
  assign n45123 = n45122 ^ n27603 ^ n22199 ;
  assign n45124 = n45123 ^ n25013 ^ n17792 ;
  assign n45125 = n39685 ^ n10590 ^ n10457 ;
  assign n45126 = n33166 | n45125 ;
  assign n45127 = ( ~n8097 & n43220 ) | ( ~n8097 & n45126 ) | ( n43220 & n45126 ) ;
  assign n45128 = ( n6140 & n24180 ) | ( n6140 & n39901 ) | ( n24180 & n39901 ) ;
  assign n45129 = n21840 ^ n19833 ^ n14481 ;
  assign n45130 = n9056 & ~n45129 ;
  assign n45131 = ~n941 & n45130 ;
  assign n45132 = n21357 & ~n43088 ;
  assign n45133 = ( n3451 & n8353 ) | ( n3451 & n29613 ) | ( n8353 & n29613 ) ;
  assign n45134 = n45133 ^ n38206 ^ 1'b0 ;
  assign n45135 = n25772 & n45134 ;
  assign n45136 = n7722 ^ n3277 ^ 1'b0 ;
  assign n45137 = n20322 & n45136 ;
  assign n45138 = n45137 ^ n29616 ^ n3797 ;
  assign n45144 = n32521 ^ n29796 ^ 1'b0 ;
  assign n45145 = ( ~n4478 & n24669 ) | ( ~n4478 & n45144 ) | ( n24669 & n45144 ) ;
  assign n45139 = n40664 ^ n16889 ^ n16833 ;
  assign n45140 = ( ~n20176 & n25684 ) | ( ~n20176 & n40148 ) | ( n25684 & n40148 ) ;
  assign n45141 = n29971 ^ n4231 ^ 1'b0 ;
  assign n45142 = ( n13593 & ~n35751 ) | ( n13593 & n45141 ) | ( ~n35751 & n45141 ) ;
  assign n45143 = ( ~n45139 & n45140 ) | ( ~n45139 & n45142 ) | ( n45140 & n45142 ) ;
  assign n45146 = n45145 ^ n45143 ^ n41425 ;
  assign n45147 = n9153 ^ n593 ^ 1'b0 ;
  assign n45148 = ( ~n8247 & n31914 ) | ( ~n8247 & n45147 ) | ( n31914 & n45147 ) ;
  assign n45149 = ( n4673 & ~n11274 ) | ( n4673 & n26911 ) | ( ~n11274 & n26911 ) ;
  assign n45150 = ( n15727 & n45148 ) | ( n15727 & n45149 ) | ( n45148 & n45149 ) ;
  assign n45151 = n5971 | n19717 ;
  assign n45152 = n9535 & ~n45151 ;
  assign n45153 = n45152 ^ n11118 ^ 1'b0 ;
  assign n45154 = n15435 | n45153 ;
  assign n45155 = n9875 ^ n6594 ^ n5008 ;
  assign n45156 = n12106 & n45155 ;
  assign n45157 = n45156 ^ n13133 ^ 1'b0 ;
  assign n45158 = ( n12885 & ~n45154 ) | ( n12885 & n45157 ) | ( ~n45154 & n45157 ) ;
  assign n45159 = ( n10154 & ~n20144 ) | ( n10154 & n29713 ) | ( ~n20144 & n29713 ) ;
  assign n45160 = n18100 ^ n15906 ^ n10864 ;
  assign n45161 = n2862 & ~n45160 ;
  assign n45162 = ( ~n2583 & n32300 ) | ( ~n2583 & n45161 ) | ( n32300 & n45161 ) ;
  assign n45163 = n28744 ^ n5745 ^ n3537 ;
  assign n45164 = n27470 & ~n45163 ;
  assign n45165 = n1081 | n32589 ;
  assign n45166 = n3115 & ~n45165 ;
  assign n45167 = n22393 ^ n21440 ^ 1'b0 ;
  assign n45168 = n29668 ^ n7081 ^ 1'b0 ;
  assign n45169 = n45167 | n45168 ;
  assign n45170 = n30433 ^ n1751 ^ 1'b0 ;
  assign n45171 = n29732 & n45170 ;
  assign n45172 = n43575 ^ n2374 ^ 1'b0 ;
  assign n45173 = n45026 ^ n40978 ^ n19776 ;
  assign n45174 = n19438 & ~n23563 ;
  assign n45175 = n38754 ^ n17774 ^ n2821 ;
  assign n45179 = n20991 ^ n7458 ^ 1'b0 ;
  assign n45180 = ~n7630 & n45179 ;
  assign n45178 = ( ~n18328 & n26702 ) | ( ~n18328 & n34677 ) | ( n26702 & n34677 ) ;
  assign n45176 = ( ~n2309 & n10044 ) | ( ~n2309 & n12213 ) | ( n10044 & n12213 ) ;
  assign n45177 = n45176 ^ n29692 ^ n2671 ;
  assign n45181 = n45180 ^ n45178 ^ n45177 ;
  assign n45182 = n45181 ^ n36559 ^ n20002 ;
  assign n45183 = n10324 ^ n7781 ^ n596 ;
  assign n45184 = n45183 ^ n41147 ^ n14566 ;
  assign n45185 = ( ~n7281 & n20505 ) | ( ~n7281 & n26664 ) | ( n20505 & n26664 ) ;
  assign n45186 = n20987 ^ n6604 ^ n2829 ;
  assign n45187 = n45186 ^ n32713 ^ n4318 ;
  assign n45188 = ( n5010 & n45185 ) | ( n5010 & n45187 ) | ( n45185 & n45187 ) ;
  assign n45189 = ~n43504 & n45188 ;
  assign n45190 = n24329 & n45189 ;
  assign n45191 = ( n5265 & n36364 ) | ( n5265 & ~n43353 ) | ( n36364 & ~n43353 ) ;
  assign n45192 = n29005 ^ n15336 ^ n14581 ;
  assign n45193 = n34798 ^ n27582 ^ n2493 ;
  assign n45194 = n32254 ^ n6624 ^ 1'b0 ;
  assign n45195 = n13842 | n27141 ;
  assign n45196 = n11646 ^ n6404 ^ n6154 ;
  assign n45197 = ~n1492 & n5578 ;
  assign n45198 = n45197 ^ n18776 ^ 1'b0 ;
  assign n45199 = ( x127 & ~n22436 ) | ( x127 & n45198 ) | ( ~n22436 & n45198 ) ;
  assign n45200 = ( ~n7071 & n45196 ) | ( ~n7071 & n45199 ) | ( n45196 & n45199 ) ;
  assign n45201 = n45200 ^ n19037 ^ 1'b0 ;
  assign n45202 = n9734 | n45201 ;
  assign n45203 = ( n38422 & n44922 ) | ( n38422 & n45202 ) | ( n44922 & n45202 ) ;
  assign n45204 = n31593 ^ n19062 ^ n14531 ;
  assign n45205 = n8130 ^ n4987 ^ n341 ;
  assign n45206 = n45205 ^ n26255 ^ n5214 ;
  assign n45207 = n5648 & ~n20585 ;
  assign n45208 = ~n16732 & n45207 ;
  assign n45209 = n41470 ^ n25349 ^ 1'b0 ;
  assign n45210 = ~n23408 & n45209 ;
  assign n45211 = ( n42024 & ~n45208 ) | ( n42024 & n45210 ) | ( ~n45208 & n45210 ) ;
  assign n45212 = ( n4403 & n37455 ) | ( n4403 & n45211 ) | ( n37455 & n45211 ) ;
  assign n45213 = n9053 | n21461 ;
  assign n45214 = n12507 ^ n2604 ^ x28 ;
  assign n45215 = n45214 ^ n39343 ^ 1'b0 ;
  assign n45216 = n12669 ^ n8161 ^ n3548 ;
  assign n45217 = n23934 & ~n45216 ;
  assign n45218 = n45215 & n45217 ;
  assign n45219 = n45218 ^ n20427 ^ n17096 ;
  assign n45220 = ( ~n1727 & n21044 ) | ( ~n1727 & n21205 ) | ( n21044 & n21205 ) ;
  assign n45221 = n45220 ^ n23059 ^ n413 ;
  assign n45222 = n34999 ^ n14853 ^ n9735 ;
  assign n45223 = n17431 & ~n23637 ;
  assign n45224 = n45223 ^ n40213 ^ n25925 ;
  assign n45226 = ( n13173 & ~n17423 ) | ( n13173 & n17551 ) | ( ~n17423 & n17551 ) ;
  assign n45227 = ~n2202 & n25253 ;
  assign n45228 = n45227 ^ n18460 ^ 1'b0 ;
  assign n45229 = ( n44027 & n45226 ) | ( n44027 & n45228 ) | ( n45226 & n45228 ) ;
  assign n45225 = ( n6262 & n12757 ) | ( n6262 & n27024 ) | ( n12757 & n27024 ) ;
  assign n45230 = n45229 ^ n45225 ^ n23019 ;
  assign n45231 = x226 & ~n13005 ;
  assign n45232 = n16728 | n28022 ;
  assign n45233 = n35789 | n45232 ;
  assign n45234 = n37022 | n44476 ;
  assign n45235 = ( x224 & n6218 ) | ( x224 & n37658 ) | ( n6218 & n37658 ) ;
  assign n45236 = ~n35257 & n45235 ;
  assign n45237 = n45234 & n45236 ;
  assign n45238 = ( n1125 & n6094 ) | ( n1125 & n15460 ) | ( n6094 & n15460 ) ;
  assign n45239 = ( x105 & n15318 ) | ( x105 & n33682 ) | ( n15318 & n33682 ) ;
  assign n45240 = n24612 ^ n19353 ^ 1'b0 ;
  assign n45241 = n3292 | n45240 ;
  assign n45242 = n45241 ^ n20144 ^ 1'b0 ;
  assign n45243 = n40226 & n45242 ;
  assign n45244 = ( n964 & ~n45239 ) | ( n964 & n45243 ) | ( ~n45239 & n45243 ) ;
  assign n45245 = n45244 ^ n10208 ^ 1'b0 ;
  assign n45246 = n20327 & n45245 ;
  assign n45247 = ( n6584 & n45238 ) | ( n6584 & ~n45246 ) | ( n45238 & ~n45246 ) ;
  assign n45248 = n29142 & ~n41528 ;
  assign n45249 = n18226 & n45248 ;
  assign n45250 = ( n27084 & ~n41903 ) | ( n27084 & n45249 ) | ( ~n41903 & n45249 ) ;
  assign n45252 = n9807 ^ n2581 ^ x84 ;
  assign n45251 = n27549 ^ n15918 ^ n2819 ;
  assign n45253 = n45252 ^ n45251 ^ n20514 ;
  assign n45254 = ( n31293 & n32438 ) | ( n31293 & n42754 ) | ( n32438 & n42754 ) ;
  assign n45255 = n13099 | n15014 ;
  assign n45256 = ( n31045 & n33172 ) | ( n31045 & n45255 ) | ( n33172 & n45255 ) ;
  assign n45257 = n15736 | n17237 ;
  assign n45258 = n45257 ^ n44728 ^ 1'b0 ;
  assign n45259 = n13916 & n33288 ;
  assign n45260 = n45259 ^ n29351 ^ 1'b0 ;
  assign n45261 = ( n15282 & ~n22815 ) | ( n15282 & n38247 ) | ( ~n22815 & n38247 ) ;
  assign n45262 = ( n17157 & ~n28782 ) | ( n17157 & n45261 ) | ( ~n28782 & n45261 ) ;
  assign n45263 = n45262 ^ n13335 ^ n10327 ;
  assign n45264 = ( n3097 & ~n10882 ) | ( n3097 & n45263 ) | ( ~n10882 & n45263 ) ;
  assign n45265 = n6797 ^ n5337 ^ 1'b0 ;
  assign n45266 = n45265 ^ n39685 ^ n11911 ;
  assign n45267 = n45264 | n45266 ;
  assign n45268 = n45267 ^ n42525 ^ 1'b0 ;
  assign n45269 = n3888 & n18237 ;
  assign n45270 = ~n31370 & n45269 ;
  assign n45271 = n45270 ^ n19188 ^ n7464 ;
  assign n45272 = n45271 ^ n21150 ^ n20816 ;
  assign n45273 = n42699 ^ n26930 ^ n26365 ;
  assign n45274 = n33636 ^ n18439 ^ n15425 ;
  assign n45275 = ( ~n9044 & n9634 ) | ( ~n9044 & n15402 ) | ( n9634 & n15402 ) ;
  assign n45276 = n45275 ^ n4105 ^ 1'b0 ;
  assign n45277 = n45274 & n45276 ;
  assign n45278 = n45277 ^ n39057 ^ n15803 ;
  assign n45279 = n910 & n24904 ;
  assign n45280 = n45279 ^ n43769 ^ n31314 ;
  assign n45281 = n30217 ^ n2898 ^ 1'b0 ;
  assign n45282 = ~n25584 & n45281 ;
  assign n45283 = n39306 ^ n38238 ^ x31 ;
  assign n45284 = ( ~n4793 & n19560 ) | ( ~n4793 & n24079 ) | ( n19560 & n24079 ) ;
  assign n45285 = n33356 ^ n7913 ^ n4007 ;
  assign n45286 = n27796 ^ n23106 ^ x97 ;
  assign n45287 = n45286 ^ n14172 ^ n13884 ;
  assign n45288 = n39181 ^ n6202 ^ 1'b0 ;
  assign n45289 = n45288 ^ n44082 ^ 1'b0 ;
  assign n45290 = ( n30418 & n32653 ) | ( n30418 & n45289 ) | ( n32653 & n45289 ) ;
  assign n45291 = n11042 ^ n4189 ^ 1'b0 ;
  assign n45292 = n40354 | n45291 ;
  assign n45293 = ( n11888 & ~n20380 ) | ( n11888 & n45292 ) | ( ~n20380 & n45292 ) ;
  assign n45294 = n13731 & n44913 ;
  assign n45295 = n45293 & ~n45294 ;
  assign n45296 = ( n13316 & n26106 ) | ( n13316 & n34319 ) | ( n26106 & n34319 ) ;
  assign n45297 = n2765 ^ n2077 ^ 1'b0 ;
  assign n45298 = n8773 & n45297 ;
  assign n45299 = ~n12879 & n45298 ;
  assign n45300 = n14808 & n45299 ;
  assign n45307 = x89 & n8825 ;
  assign n45308 = n45307 ^ n29349 ^ 1'b0 ;
  assign n45309 = ~n30603 & n45308 ;
  assign n45310 = n45309 ^ n39816 ^ 1'b0 ;
  assign n45301 = n655 & n25837 ;
  assign n45302 = ( n1459 & n8049 ) | ( n1459 & ~n45301 ) | ( n8049 & ~n45301 ) ;
  assign n45304 = ( n929 & ~n3394 ) | ( n929 & n3646 ) | ( ~n3394 & n3646 ) ;
  assign n45303 = ( ~n14240 & n19395 ) | ( ~n14240 & n41170 ) | ( n19395 & n41170 ) ;
  assign n45305 = n45304 ^ n45303 ^ 1'b0 ;
  assign n45306 = n45302 & ~n45305 ;
  assign n45311 = n45310 ^ n45306 ^ n28847 ;
  assign n45312 = ~n10963 & n38791 ;
  assign n45313 = n45312 ^ n23275 ^ 1'b0 ;
  assign n45314 = n35109 ^ n13806 ^ n1082 ;
  assign n45315 = n21259 ^ n20624 ^ n13493 ;
  assign n45316 = ( ~n39845 & n45314 ) | ( ~n39845 & n45315 ) | ( n45314 & n45315 ) ;
  assign n45317 = n33491 ^ n31553 ^ n4994 ;
  assign n45318 = ( ~n4577 & n35110 ) | ( ~n4577 & n45317 ) | ( n35110 & n45317 ) ;
  assign n45319 = ( ~n12800 & n27510 ) | ( ~n12800 & n45069 ) | ( n27510 & n45069 ) ;
  assign n45320 = n34101 ^ n21026 ^ 1'b0 ;
  assign n45321 = ~n45319 & n45320 ;
  assign n45322 = ( ~n4717 & n17747 ) | ( ~n4717 & n31745 ) | ( n17747 & n31745 ) ;
  assign n45323 = ( n10224 & ~n45321 ) | ( n10224 & n45322 ) | ( ~n45321 & n45322 ) ;
  assign n45324 = n6723 & ~n11924 ;
  assign n45325 = n31695 & n45324 ;
  assign n45326 = n37851 ^ n27845 ^ n10463 ;
  assign n45327 = ( n29692 & n40226 ) | ( n29692 & ~n45326 ) | ( n40226 & ~n45326 ) ;
  assign n45328 = ( n20726 & ~n44331 ) | ( n20726 & n45327 ) | ( ~n44331 & n45327 ) ;
  assign n45329 = ( n4325 & n11224 ) | ( n4325 & n13334 ) | ( n11224 & n13334 ) ;
  assign n45330 = ( ~n11983 & n19544 ) | ( ~n11983 & n45329 ) | ( n19544 & n45329 ) ;
  assign n45331 = ( n6649 & ~n11325 ) | ( n6649 & n12656 ) | ( ~n11325 & n12656 ) ;
  assign n45332 = ( n4211 & ~n10545 ) | ( n4211 & n45331 ) | ( ~n10545 & n45331 ) ;
  assign n45333 = ( n2215 & n26223 ) | ( n2215 & n32417 ) | ( n26223 & n32417 ) ;
  assign n45334 = n409 | n7734 ;
  assign n45335 = n45334 ^ n15992 ^ 1'b0 ;
  assign n45336 = n22589 ^ n2462 ^ 1'b0 ;
  assign n45337 = ~n45335 & n45336 ;
  assign n45338 = ( ~n353 & n15849 ) | ( ~n353 & n45337 ) | ( n15849 & n45337 ) ;
  assign n45339 = n3597 & n29079 ;
  assign n45340 = ~n29477 & n45339 ;
  assign n45341 = n19369 & n45340 ;
  assign n45342 = x193 & ~n17182 ;
  assign n45343 = n45342 ^ n972 ^ 1'b0 ;
  assign n45344 = n27595 ^ n15919 ^ n8744 ;
  assign n45345 = n45344 ^ n33955 ^ n19063 ;
  assign n45346 = ( ~n1624 & n14610 ) | ( ~n1624 & n45345 ) | ( n14610 & n45345 ) ;
  assign n45347 = n24940 ^ n1357 ^ 1'b0 ;
  assign n45348 = n45347 ^ n38789 ^ n31196 ;
  assign n45353 = ( ~n20936 & n27231 ) | ( ~n20936 & n32140 ) | ( n27231 & n32140 ) ;
  assign n45350 = n3660 ^ n2704 ^ 1'b0 ;
  assign n45351 = n3340 & n45350 ;
  assign n45352 = n45351 ^ n18507 ^ n13703 ;
  assign n45354 = n45353 ^ n45352 ^ n23318 ;
  assign n45349 = ( n8842 & ~n9583 ) | ( n8842 & n28915 ) | ( ~n9583 & n28915 ) ;
  assign n45355 = n45354 ^ n45349 ^ n20344 ;
  assign n45356 = ~n3808 & n29444 ;
  assign n45357 = ~n27834 & n45356 ;
  assign n45358 = ( n11291 & ~n33773 ) | ( n11291 & n45357 ) | ( ~n33773 & n45357 ) ;
  assign n45359 = ( x118 & n2337 ) | ( x118 & ~n33683 ) | ( n2337 & ~n33683 ) ;
  assign n45360 = ~n9359 & n22355 ;
  assign n45361 = n45360 ^ n16030 ^ 1'b0 ;
  assign n45362 = n23106 ^ n16281 ^ 1'b0 ;
  assign n45363 = n45361 & n45362 ;
  assign n45364 = ~n9708 & n45363 ;
  assign n45365 = ~n20972 & n45364 ;
  assign n45366 = ( ~n20073 & n28048 ) | ( ~n20073 & n35070 ) | ( n28048 & n35070 ) ;
  assign n45367 = n45366 ^ n15043 ^ n8207 ;
  assign n45368 = n45367 ^ n28810 ^ n9575 ;
  assign n45369 = n13369 | n45368 ;
  assign n45370 = n33393 | n45369 ;
  assign n45371 = n12881 & n15281 ;
  assign n45372 = ( n1798 & n24452 ) | ( n1798 & n45371 ) | ( n24452 & n45371 ) ;
  assign n45373 = ( n2443 & n39410 ) | ( n2443 & ~n45372 ) | ( n39410 & ~n45372 ) ;
  assign n45378 = n9235 ^ n5931 ^ n4406 ;
  assign n45374 = n37333 ^ n30006 ^ 1'b0 ;
  assign n45375 = n20042 ^ n13755 ^ n3258 ;
  assign n45376 = n45375 ^ n13159 ^ 1'b0 ;
  assign n45377 = ~n45374 & n45376 ;
  assign n45379 = n45378 ^ n45377 ^ n35638 ;
  assign n45380 = n40590 ^ n20180 ^ n549 ;
  assign n45381 = ( n45373 & n45379 ) | ( n45373 & ~n45380 ) | ( n45379 & ~n45380 ) ;
  assign n45382 = n13629 ^ n12624 ^ n4674 ;
  assign n45384 = ( ~n1080 & n21846 ) | ( ~n1080 & n28345 ) | ( n21846 & n28345 ) ;
  assign n45383 = ( n8333 & n8914 ) | ( n8333 & ~n9852 ) | ( n8914 & ~n9852 ) ;
  assign n45385 = n45384 ^ n45383 ^ n8895 ;
  assign n45386 = ( ~n14273 & n18588 ) | ( ~n14273 & n39540 ) | ( n18588 & n39540 ) ;
  assign n45387 = n4993 & ~n39198 ;
  assign n45388 = n45387 ^ n25304 ^ 1'b0 ;
  assign n45389 = n45388 ^ n11099 ^ n6793 ;
  assign n45390 = n7368 ^ n5684 ^ 1'b0 ;
  assign n45391 = n27652 | n41861 ;
  assign n45392 = n45390 | n45391 ;
  assign n45393 = ( n5556 & ~n8886 ) | ( n5556 & n14253 ) | ( ~n8886 & n14253 ) ;
  assign n45394 = ~n1716 & n17734 ;
  assign n45395 = n45393 & n45394 ;
  assign n45396 = n32897 & n34152 ;
  assign n45397 = n45396 ^ n20742 ^ 1'b0 ;
  assign n45398 = ( n11539 & n16676 ) | ( n11539 & n16734 ) | ( n16676 & n16734 ) ;
  assign n45399 = n13405 ^ n8103 ^ n6649 ;
  assign n45400 = n21455 ^ n18237 ^ n12964 ;
  assign n45401 = ( n1212 & n45399 ) | ( n1212 & ~n45400 ) | ( n45399 & ~n45400 ) ;
  assign n45402 = n18580 ^ n17574 ^ n12388 ;
  assign n45404 = ( n18262 & n21586 ) | ( n18262 & n25684 ) | ( n21586 & n25684 ) ;
  assign n45403 = n33219 ^ n18854 ^ n10361 ;
  assign n45405 = n45404 ^ n45403 ^ n29491 ;
  assign n45406 = n9160 ^ n2708 ^ n2241 ;
  assign n45407 = ( ~n1470 & n21357 ) | ( ~n1470 & n45406 ) | ( n21357 & n45406 ) ;
  assign n45408 = ( n637 & n12879 ) | ( n637 & n45407 ) | ( n12879 & n45407 ) ;
  assign n45409 = ( x162 & ~n7767 ) | ( x162 & n9452 ) | ( ~n7767 & n9452 ) ;
  assign n45410 = n45409 ^ n9789 ^ n7042 ;
  assign n45411 = ( n10015 & ~n21016 ) | ( n10015 & n45410 ) | ( ~n21016 & n45410 ) ;
  assign n45412 = n45411 ^ n41211 ^ n39600 ;
  assign n45413 = ( ~n16676 & n21963 ) | ( ~n16676 & n38882 ) | ( n21963 & n38882 ) ;
  assign n45414 = n11230 & ~n30116 ;
  assign n45415 = n45414 ^ n24037 ^ 1'b0 ;
  assign n45416 = ~n9555 & n35217 ;
  assign n45417 = n45416 ^ n11449 ^ 1'b0 ;
  assign n45418 = n31283 ^ n13721 ^ 1'b0 ;
  assign n45419 = n17734 & n45418 ;
  assign n45420 = n45419 ^ n23301 ^ 1'b0 ;
  assign n45421 = n43171 ^ n31207 ^ n2707 ;
  assign n45422 = n24189 ^ n3604 ^ n690 ;
  assign n45423 = n2572 & ~n24195 ;
  assign n45424 = n45423 ^ n42282 ^ 1'b0 ;
  assign n45425 = ~n11193 & n45424 ;
  assign n45426 = n45425 ^ n43413 ^ n1959 ;
  assign n45427 = n28326 ^ n13500 ^ n12073 ;
  assign n45428 = ( n9378 & ~n17957 ) | ( n9378 & n22455 ) | ( ~n17957 & n22455 ) ;
  assign n45429 = n6029 | n45428 ;
  assign n45430 = ( n11784 & n11830 ) | ( n11784 & ~n45429 ) | ( n11830 & ~n45429 ) ;
  assign n45431 = ( n4278 & ~n6686 ) | ( n4278 & n19089 ) | ( ~n6686 & n19089 ) ;
  assign n45432 = ( ~n1585 & n14631 ) | ( ~n1585 & n20074 ) | ( n14631 & n20074 ) ;
  assign n45433 = n14090 & n31528 ;
  assign n45434 = n45433 ^ n39972 ^ 1'b0 ;
  assign n45435 = n45434 ^ n15000 ^ n7713 ;
  assign n45436 = n45432 & ~n45435 ;
  assign n45437 = n45436 ^ n14379 ^ 1'b0 ;
  assign n45438 = n3720 & ~n45437 ;
  assign n45439 = n24046 ^ n19516 ^ n1376 ;
  assign n45440 = n17249 ^ n15829 ^ 1'b0 ;
  assign n45441 = n45439 & ~n45440 ;
  assign n45442 = ~n1157 & n20919 ;
  assign n45443 = n1262 & ~n45442 ;
  assign n45444 = n45443 ^ n29328 ^ 1'b0 ;
  assign n45445 = ( n7436 & n11820 ) | ( n7436 & n13087 ) | ( n11820 & n13087 ) ;
  assign n45446 = n44383 ^ n30612 ^ n14629 ;
  assign n45447 = ( ~n4227 & n8721 ) | ( ~n4227 & n20448 ) | ( n8721 & n20448 ) ;
  assign n45448 = n13891 & n31547 ;
  assign n45449 = n45448 ^ n9160 ^ n6284 ;
  assign n45450 = n7596 & n42937 ;
  assign n45451 = n35420 ^ n21161 ^ n8720 ;
  assign n45452 = ( ~n45449 & n45450 ) | ( ~n45449 & n45451 ) | ( n45450 & n45451 ) ;
  assign n45453 = ( ~n34671 & n45447 ) | ( ~n34671 & n45452 ) | ( n45447 & n45452 ) ;
  assign n45454 = ( ~n10717 & n31234 ) | ( ~n10717 & n39496 ) | ( n31234 & n39496 ) ;
  assign n45455 = n18548 | n27127 ;
  assign n45456 = n22438 ^ n19359 ^ n8167 ;
  assign n45457 = n5167 & n45456 ;
  assign n45458 = ~n1204 & n45457 ;
  assign n45459 = n43878 ^ n23384 ^ n18784 ;
  assign n45460 = n45459 ^ n45436 ^ n5241 ;
  assign n45462 = n32763 ^ n19697 ^ x78 ;
  assign n45461 = n15217 | n33827 ;
  assign n45463 = n45462 ^ n45461 ^ n14200 ;
  assign n45464 = n18853 ^ n1059 ^ 1'b0 ;
  assign n45465 = n13138 ^ n8201 ^ 1'b0 ;
  assign n45466 = n45465 ^ n7202 ^ n3882 ;
  assign n45467 = n26458 ^ n16951 ^ 1'b0 ;
  assign n45468 = ~n33299 & n45467 ;
  assign n45469 = n38857 & n45468 ;
  assign n45470 = n29588 ^ n18342 ^ 1'b0 ;
  assign n45471 = n18609 ^ n9496 ^ 1'b0 ;
  assign n45472 = n45470 & ~n45471 ;
  assign n45473 = n45472 ^ n13631 ^ 1'b0 ;
  assign n45474 = ~n32313 & n45473 ;
  assign n45475 = n45474 ^ n33237 ^ 1'b0 ;
  assign n45476 = n28764 & n45475 ;
  assign n45477 = ( n9179 & ~n13579 ) | ( n9179 & n24033 ) | ( ~n13579 & n24033 ) ;
  assign n45478 = n45477 ^ n12229 ^ 1'b0 ;
  assign n45479 = n6351 ^ n2797 ^ n1760 ;
  assign n45480 = ~n4203 & n45479 ;
  assign n45481 = n14258 & n45480 ;
  assign n45482 = n29811 ^ n23402 ^ n13138 ;
  assign n45483 = n25837 ^ n1875 ^ 1'b0 ;
  assign n45484 = ( n8882 & n45482 ) | ( n8882 & ~n45483 ) | ( n45482 & ~n45483 ) ;
  assign n45485 = n5193 | n12738 ;
  assign n45486 = n45485 ^ n39655 ^ n30179 ;
  assign n45487 = ~n21109 & n31004 ;
  assign n45488 = n45487 ^ n22102 ^ n5638 ;
  assign n45489 = n2290 & ~n25627 ;
  assign n45490 = n45489 ^ n5588 ^ 1'b0 ;
  assign n45491 = n4304 & ~n16134 ;
  assign n45492 = n45491 ^ n8271 ^ 1'b0 ;
  assign n45493 = n1064 ^ n928 ^ 1'b0 ;
  assign n45494 = ~n16923 & n38494 ;
  assign n45495 = n25618 ^ n13673 ^ n8980 ;
  assign n45496 = n45495 ^ n8243 ^ n5373 ;
  assign n45497 = n17802 & n40795 ;
  assign n45498 = n25600 ^ n5790 ^ 1'b0 ;
  assign n45499 = ( n12919 & n32471 ) | ( n12919 & ~n45498 ) | ( n32471 & ~n45498 ) ;
  assign n45500 = n45499 ^ n23156 ^ 1'b0 ;
  assign n45501 = n33973 & n45500 ;
  assign n45502 = n45497 | n45501 ;
  assign n45504 = ~n25765 & n29890 ;
  assign n45503 = ~n7109 & n23414 ;
  assign n45505 = n45504 ^ n45503 ^ n8220 ;
  assign n45506 = n16351 & ~n20834 ;
  assign n45507 = n17110 ^ n1814 ^ 1'b0 ;
  assign n45508 = n20258 & ~n45507 ;
  assign n45509 = n1329 & n45508 ;
  assign n45510 = ~n16329 & n45509 ;
  assign n45511 = n45510 ^ n31406 ^ n24634 ;
  assign n45512 = n3331 & ~n37683 ;
  assign n45513 = ( n24339 & n43975 ) | ( n24339 & ~n45512 ) | ( n43975 & ~n45512 ) ;
  assign n45514 = n45513 ^ n6269 ^ n6184 ;
  assign n45515 = n18107 ^ n3839 ^ n3116 ;
  assign n45516 = ( n11242 & n30881 ) | ( n11242 & ~n32388 ) | ( n30881 & ~n32388 ) ;
  assign n45517 = ( n829 & n883 ) | ( n829 & ~n11836 ) | ( n883 & ~n11836 ) ;
  assign n45518 = n37855 ^ n37619 ^ n3008 ;
  assign n45519 = n45518 ^ n362 ^ x97 ;
  assign n45520 = ( n7763 & n45517 ) | ( n7763 & ~n45519 ) | ( n45517 & ~n45519 ) ;
  assign n45521 = n36144 ^ n28146 ^ n23703 ;
  assign n45522 = n18569 & n18582 ;
  assign n45523 = n45522 ^ n6179 ^ 1'b0 ;
  assign n45524 = n45523 ^ n27827 ^ 1'b0 ;
  assign n45525 = n18442 & n45524 ;
  assign n45526 = n12767 ^ n3552 ^ 1'b0 ;
  assign n45527 = ( ~n19679 & n45525 ) | ( ~n19679 & n45526 ) | ( n45525 & n45526 ) ;
  assign n45528 = n24252 & n25015 ;
  assign n45529 = ~n45527 & n45528 ;
  assign n45530 = n10136 & n39446 ;
  assign n45531 = n3501 | n19182 ;
  assign n45532 = ( n14595 & ~n31239 ) | ( n14595 & n45531 ) | ( ~n31239 & n45531 ) ;
  assign n45533 = n12443 ^ n5357 ^ n1258 ;
  assign n45534 = n20142 & n45533 ;
  assign n45535 = n6297 & ~n45534 ;
  assign n45536 = ( n15390 & n18921 ) | ( n15390 & n35088 ) | ( n18921 & n35088 ) ;
  assign n45537 = n35356 ^ n28130 ^ n2254 ;
  assign n45538 = ( ~n6656 & n33804 ) | ( ~n6656 & n34190 ) | ( n33804 & n34190 ) ;
  assign n45539 = n45538 ^ n38401 ^ n6108 ;
  assign n45540 = ( n2518 & n11493 ) | ( n2518 & ~n45539 ) | ( n11493 & ~n45539 ) ;
  assign n45544 = n31634 ^ n18903 ^ n4079 ;
  assign n45541 = ( n4813 & n9029 ) | ( n4813 & n17474 ) | ( n9029 & n17474 ) ;
  assign n45542 = n37225 ^ n8606 ^ 1'b0 ;
  assign n45543 = n45541 & ~n45542 ;
  assign n45545 = n45544 ^ n45543 ^ n16062 ;
  assign n45546 = n37493 ^ n15164 ^ n5711 ;
  assign n45547 = n19290 ^ n13205 ^ n7067 ;
  assign n45548 = ( n17531 & ~n45546 ) | ( n17531 & n45547 ) | ( ~n45546 & n45547 ) ;
  assign n45549 = n14540 | n21648 ;
  assign n45550 = n13946 & ~n45549 ;
  assign n45551 = ( n1424 & n13151 ) | ( n1424 & ~n41466 ) | ( n13151 & ~n41466 ) ;
  assign n45553 = n15704 ^ n7122 ^ n6666 ;
  assign n45554 = n45553 ^ n31182 ^ n26863 ;
  assign n45552 = n9060 | n14727 ;
  assign n45555 = n45554 ^ n45552 ^ 1'b0 ;
  assign n45556 = n38724 & n45555 ;
  assign n45557 = ~n45551 & n45556 ;
  assign n45558 = n38591 ^ n6401 ^ 1'b0 ;
  assign n45559 = n34594 & ~n45558 ;
  assign n45560 = n45559 ^ n23655 ^ n9970 ;
  assign n45561 = n31767 | n45560 ;
  assign n45563 = n14057 ^ n10990 ^ n9824 ;
  assign n45564 = n45563 ^ n18302 ^ n6856 ;
  assign n45562 = n27177 ^ n21100 ^ n8057 ;
  assign n45565 = n45564 ^ n45562 ^ n2366 ;
  assign n45566 = n15777 ^ n14572 ^ n784 ;
  assign n45568 = n42346 ^ n29506 ^ n22501 ;
  assign n45567 = ~n24839 & n43574 ;
  assign n45569 = n45568 ^ n45567 ^ n28154 ;
  assign n45570 = n4332 & ~n22189 ;
  assign n45571 = n45570 ^ n24355 ^ n8869 ;
  assign n45572 = n45571 ^ n3265 ^ n352 ;
  assign n45573 = n45572 ^ n36150 ^ 1'b0 ;
  assign n45574 = ~n13635 & n26719 ;
  assign n45575 = n31822 & n45574 ;
  assign n45576 = n12008 & ~n27827 ;
  assign n45577 = ( n5491 & n20800 ) | ( n5491 & ~n45576 ) | ( n20800 & ~n45576 ) ;
  assign n45578 = ( n604 & n42658 ) | ( n604 & ~n45577 ) | ( n42658 & ~n45577 ) ;
  assign n45579 = ( n2587 & n2700 ) | ( n2587 & ~n15516 ) | ( n2700 & ~n15516 ) ;
  assign n45580 = n27276 & n45579 ;
  assign n45581 = n26745 & n45580 ;
  assign n45582 = n45581 ^ n44390 ^ n4104 ;
  assign n45584 = n38527 ^ n15871 ^ 1'b0 ;
  assign n45583 = n1938 & ~n4823 ;
  assign n45585 = n45584 ^ n45583 ^ n32586 ;
  assign n45586 = n41254 ^ n33445 ^ n30963 ;
  assign n45587 = n8878 ^ n6086 ^ x142 ;
  assign n45588 = n1083 & n35286 ;
  assign n45589 = n45588 ^ n42830 ^ n21648 ;
  assign n45590 = ~n19580 & n35545 ;
  assign n45591 = n45590 ^ n6001 ^ 1'b0 ;
  assign n45592 = n25017 ^ n15848 ^ 1'b0 ;
  assign n45593 = n39876 & n45592 ;
  assign n45594 = n34247 & ~n45533 ;
  assign n45596 = n27121 ^ n22734 ^ 1'b0 ;
  assign n45597 = n39649 | n45596 ;
  assign n45595 = ~n1263 & n23205 ;
  assign n45598 = n45597 ^ n45595 ^ n28480 ;
  assign n45599 = n13529 ^ n11873 ^ 1'b0 ;
  assign n45600 = n1475 | n45599 ;
  assign n45601 = n45600 ^ n25069 ^ n21090 ;
  assign n45602 = ( n12750 & n18897 ) | ( n12750 & ~n44214 ) | ( n18897 & ~n44214 ) ;
  assign n45603 = n5890 | n16141 ;
  assign n45604 = ( n14942 & n30014 ) | ( n14942 & n45603 ) | ( n30014 & n45603 ) ;
  assign n45605 = n20870 & ~n39771 ;
  assign n45606 = n3995 & n45605 ;
  assign n45607 = ~n36990 & n45606 ;
  assign n45608 = n17903 ^ n5857 ^ 1'b0 ;
  assign n45609 = n10131 & ~n45608 ;
  assign n45610 = ( n3443 & n3820 ) | ( n3443 & n14039 ) | ( n3820 & n14039 ) ;
  assign n45611 = ( n27837 & n33239 ) | ( n27837 & ~n45610 ) | ( n33239 & ~n45610 ) ;
  assign n45612 = n45611 ^ n8093 ^ 1'b0 ;
  assign n45613 = ~n29949 & n45612 ;
  assign n45614 = ( n12020 & n18172 ) | ( n12020 & n18250 ) | ( n18172 & n18250 ) ;
  assign n45615 = n16677 ^ x100 ^ 1'b0 ;
  assign n45616 = n45615 ^ n27910 ^ n15133 ;
  assign n45617 = n45616 ^ n8953 ^ n4636 ;
  assign n45618 = ( n15288 & n15512 ) | ( n15288 & ~n28333 ) | ( n15512 & ~n28333 ) ;
  assign n45619 = ( n12185 & n13975 ) | ( n12185 & ~n21368 ) | ( n13975 & ~n21368 ) ;
  assign n45620 = ( n33689 & n45618 ) | ( n33689 & n45619 ) | ( n45618 & n45619 ) ;
  assign n45621 = ( ~n2643 & n17918 ) | ( ~n2643 & n34738 ) | ( n17918 & n34738 ) ;
  assign n45622 = n45621 ^ n14959 ^ 1'b0 ;
  assign n45623 = n33419 ^ n6879 ^ n5785 ;
  assign n45624 = n30732 ^ n22280 ^ n6195 ;
  assign n45625 = n4335 & ~n34993 ;
  assign n45626 = ( n932 & n18136 ) | ( n932 & n23647 ) | ( n18136 & n23647 ) ;
  assign n45627 = ( ~n6965 & n8486 ) | ( ~n6965 & n12651 ) | ( n8486 & n12651 ) ;
  assign n45630 = n13812 ^ x58 ^ 1'b0 ;
  assign n45628 = n1161 | n19205 ;
  assign n45629 = n9217 | n45628 ;
  assign n45631 = n45630 ^ n45629 ^ n4430 ;
  assign n45632 = n17155 ^ n7869 ^ n1979 ;
  assign n45633 = n45632 ^ n36635 ^ n22237 ;
  assign n45634 = ~n3320 & n27549 ;
  assign n45635 = n45634 ^ n11528 ^ 1'b0 ;
  assign n45636 = n45635 ^ n21278 ^ n7080 ;
  assign n45637 = n30201 ^ n24682 ^ n17120 ;
  assign n45638 = n13170 & n31854 ;
  assign n45639 = ~n45637 & n45638 ;
  assign n45640 = n17382 ^ n8888 ^ n687 ;
  assign n45641 = n11711 & n45640 ;
  assign n45642 = n17211 ^ n2815 ^ n2491 ;
  assign n45643 = n1030 | n45642 ;
  assign n45644 = n45643 ^ n40759 ^ 1'b0 ;
  assign n45645 = n14747 & n44713 ;
  assign n45646 = ~n45644 & n45645 ;
  assign n45647 = ( n25465 & n36160 ) | ( n25465 & n41191 ) | ( n36160 & n41191 ) ;
  assign n45648 = n28382 ^ n19118 ^ 1'b0 ;
  assign n45649 = n29444 ^ n18867 ^ n16093 ;
  assign n45650 = ( ~n37737 & n45648 ) | ( ~n37737 & n45649 ) | ( n45648 & n45649 ) ;
  assign n45651 = n19377 ^ n19267 ^ n4038 ;
  assign n45652 = n33473 & ~n45651 ;
  assign n45653 = n45652 ^ n37862 ^ 1'b0 ;
  assign n45654 = n45653 ^ n4217 ^ n2691 ;
  assign n45655 = ~n1822 & n17492 ;
  assign n45656 = n6881 ^ n6278 ^ n3892 ;
  assign n45657 = ( n4045 & n14381 ) | ( n4045 & n45656 ) | ( n14381 & n45656 ) ;
  assign n45658 = ( n1286 & n36203 ) | ( n1286 & n45657 ) | ( n36203 & n45657 ) ;
  assign n45660 = n44074 ^ n42891 ^ n25461 ;
  assign n45659 = n10770 & n40015 ;
  assign n45661 = n45660 ^ n45659 ^ 1'b0 ;
  assign n45663 = n35657 ^ n21430 ^ n10410 ;
  assign n45662 = ( n3935 & n20840 ) | ( n3935 & n31982 ) | ( n20840 & n31982 ) ;
  assign n45664 = n45663 ^ n45662 ^ n21241 ;
  assign n45665 = n30929 & n45664 ;
  assign n45667 = ( n4746 & n17412 ) | ( n4746 & n33435 ) | ( n17412 & n33435 ) ;
  assign n45668 = n22515 & ~n45667 ;
  assign n45666 = n21730 ^ n13415 ^ n3332 ;
  assign n45669 = n45668 ^ n45666 ^ n13025 ;
  assign n45670 = n29618 ^ n11341 ^ n10516 ;
  assign n45671 = n17309 | n34636 ;
  assign n45677 = n33825 ^ n7292 ^ n5117 ;
  assign n45678 = n24932 ^ n16743 ^ 1'b0 ;
  assign n45679 = ~n45677 & n45678 ;
  assign n45672 = n21937 ^ n19699 ^ x27 ;
  assign n45673 = n11732 ^ n4446 ^ n2362 ;
  assign n45674 = ( n2505 & ~n28277 ) | ( n2505 & n45673 ) | ( ~n28277 & n45673 ) ;
  assign n45675 = n45674 ^ n23126 ^ n2953 ;
  assign n45676 = ( ~n7635 & n45672 ) | ( ~n7635 & n45675 ) | ( n45672 & n45675 ) ;
  assign n45680 = n45679 ^ n45676 ^ 1'b0 ;
  assign n45681 = n12143 ^ n10537 ^ n10367 ;
  assign n45682 = ( n25627 & n30486 ) | ( n25627 & n35990 ) | ( n30486 & n35990 ) ;
  assign n45683 = n37216 ^ n29089 ^ 1'b0 ;
  assign n45684 = n45683 ^ n41072 ^ n12047 ;
  assign n45686 = n32568 ^ n15013 ^ n3110 ;
  assign n45687 = n45686 ^ n31981 ^ x179 ;
  assign n45685 = ~n2300 & n33462 ;
  assign n45688 = n45687 ^ n45685 ^ 1'b0 ;
  assign n45689 = n35252 & n35334 ;
  assign n45690 = n44286 & n45689 ;
  assign n45691 = ~n19131 & n27938 ;
  assign n45692 = ~n35866 & n45691 ;
  assign n45693 = ~n12409 & n28041 ;
  assign n45694 = n45693 ^ n21529 ^ 1'b0 ;
  assign n45695 = ( ~n4378 & n28026 ) | ( ~n4378 & n45694 ) | ( n28026 & n45694 ) ;
  assign n45696 = n3536 & ~n41006 ;
  assign n45697 = n30221 ^ n15244 ^ 1'b0 ;
  assign n45698 = n25714 ^ n23066 ^ n16696 ;
  assign n45699 = ( n13727 & n25004 ) | ( n13727 & ~n45698 ) | ( n25004 & ~n45698 ) ;
  assign n45700 = ( ~n7334 & n28099 ) | ( ~n7334 & n43213 ) | ( n28099 & n43213 ) ;
  assign n45701 = n25113 & n45700 ;
  assign n45702 = ( n25073 & n36765 ) | ( n25073 & n45701 ) | ( n36765 & n45701 ) ;
  assign n45703 = n36390 ^ n8806 ^ n5771 ;
  assign n45704 = ( n9696 & n45163 ) | ( n9696 & n45703 ) | ( n45163 & n45703 ) ;
  assign n45705 = n30412 & ~n37742 ;
  assign n45706 = ~n6958 & n43515 ;
  assign n45707 = n45706 ^ n15609 ^ 1'b0 ;
  assign n45708 = ~n4468 & n45707 ;
  assign n45709 = n45708 ^ n19525 ^ 1'b0 ;
  assign n45710 = n11829 | n37162 ;
  assign n45711 = ( n27519 & ~n31437 ) | ( n27519 & n45710 ) | ( ~n31437 & n45710 ) ;
  assign n45712 = n45711 ^ n7703 ^ 1'b0 ;
  assign n45713 = n20811 | n45712 ;
  assign n45714 = n1802 & n16273 ;
  assign n45715 = ( n8905 & ~n13160 ) | ( n8905 & n45714 ) | ( ~n13160 & n45714 ) ;
  assign n45716 = n28043 ^ n10318 ^ 1'b0 ;
  assign n45717 = n14683 | n45716 ;
  assign n45718 = n37301 ^ n28567 ^ n10229 ;
  assign n45719 = ( n28836 & ~n42907 ) | ( n28836 & n45718 ) | ( ~n42907 & n45718 ) ;
  assign n45720 = n45719 ^ n39085 ^ 1'b0 ;
  assign n45721 = ( n26632 & n45717 ) | ( n26632 & ~n45720 ) | ( n45717 & ~n45720 ) ;
  assign n45722 = n8150 & ~n20450 ;
  assign n45723 = n45722 ^ n14563 ^ n8667 ;
  assign n45724 = n45723 ^ n43071 ^ n26121 ;
  assign n45725 = ( n3852 & n5929 ) | ( n3852 & n13724 ) | ( n5929 & n13724 ) ;
  assign n45726 = ( n9026 & n29094 ) | ( n9026 & n45725 ) | ( n29094 & n45725 ) ;
  assign n45727 = n7535 & ~n21642 ;
  assign n45728 = ( n2980 & n4295 ) | ( n2980 & ~n26724 ) | ( n4295 & ~n26724 ) ;
  assign n45729 = ~n13346 & n45728 ;
  assign n45730 = n45729 ^ n4861 ^ 1'b0 ;
  assign n45731 = n20070 ^ n16843 ^ n2338 ;
  assign n45732 = n45731 ^ n31770 ^ n3541 ;
  assign n45733 = n6284 & n41355 ;
  assign n45734 = n45733 ^ n14290 ^ 1'b0 ;
  assign n45735 = n45734 ^ n43181 ^ n36171 ;
  assign n45736 = n5930 & ~n44750 ;
  assign n45737 = ( n293 & n1883 ) | ( n293 & n4465 ) | ( n1883 & n4465 ) ;
  assign n45738 = ( n13783 & n14571 ) | ( n13783 & ~n45737 ) | ( n14571 & ~n45737 ) ;
  assign n45739 = n25755 ^ n24884 ^ 1'b0 ;
  assign n45740 = ( x114 & n17336 ) | ( x114 & n45739 ) | ( n17336 & n45739 ) ;
  assign n45741 = ( n511 & n13970 ) | ( n511 & ~n24183 ) | ( n13970 & ~n24183 ) ;
  assign n45742 = ~n21452 & n45741 ;
  assign n45743 = n12697 ^ n3940 ^ 1'b0 ;
  assign n45744 = ~n19905 & n45743 ;
  assign n45745 = ( n14172 & n15008 ) | ( n14172 & n17218 ) | ( n15008 & n17218 ) ;
  assign n45746 = ( ~n15830 & n17568 ) | ( ~n15830 & n19832 ) | ( n17568 & n19832 ) ;
  assign n45748 = ( n884 & n20133 ) | ( n884 & ~n45728 ) | ( n20133 & ~n45728 ) ;
  assign n45749 = n881 & ~n10948 ;
  assign n45750 = n45748 & ~n45749 ;
  assign n45751 = n45750 ^ n27112 ^ 1'b0 ;
  assign n45747 = ~n14896 & n22581 ;
  assign n45752 = n45751 ^ n45747 ^ 1'b0 ;
  assign n45753 = n31634 ^ n8909 ^ n3063 ;
  assign n45754 = n37721 ^ n23741 ^ 1'b0 ;
  assign n45755 = n45753 | n45754 ;
  assign n45756 = ( n43584 & n45752 ) | ( n43584 & ~n45755 ) | ( n45752 & ~n45755 ) ;
  assign n45757 = ( n5278 & n24102 ) | ( n5278 & ~n38649 ) | ( n24102 & ~n38649 ) ;
  assign n45758 = n20710 ^ n5681 ^ n719 ;
  assign n45759 = n45758 ^ n19169 ^ n788 ;
  assign n45760 = n36439 ^ n18180 ^ n2408 ;
  assign n45761 = ( ~n5772 & n10733 ) | ( ~n5772 & n11232 ) | ( n10733 & n11232 ) ;
  assign n45762 = ( ~n31011 & n40590 ) | ( ~n31011 & n45761 ) | ( n40590 & n45761 ) ;
  assign n45763 = n2626 | n3188 ;
  assign n45764 = ( n14172 & ~n27953 ) | ( n14172 & n45763 ) | ( ~n27953 & n45763 ) ;
  assign n45765 = n5060 ^ n4646 ^ n1399 ;
  assign n45766 = n9000 ^ n8485 ^ 1'b0 ;
  assign n45767 = n4352 & ~n45766 ;
  assign n45768 = ( ~n22356 & n22595 ) | ( ~n22356 & n35233 ) | ( n22595 & n35233 ) ;
  assign n45769 = ( n25346 & n28299 ) | ( n25346 & n35051 ) | ( n28299 & n35051 ) ;
  assign n45770 = ( n45767 & n45768 ) | ( n45767 & n45769 ) | ( n45768 & n45769 ) ;
  assign n45776 = ( n5724 & n6296 ) | ( n5724 & ~n9980 ) | ( n6296 & ~n9980 ) ;
  assign n45775 = n40458 ^ n29314 ^ n4781 ;
  assign n45771 = n12533 ^ n10822 ^ n7580 ;
  assign n45772 = ( ~n21451 & n29435 ) | ( ~n21451 & n45771 ) | ( n29435 & n45771 ) ;
  assign n45773 = n45772 ^ n29683 ^ 1'b0 ;
  assign n45774 = ( n25761 & n40725 ) | ( n25761 & ~n45773 ) | ( n40725 & ~n45773 ) ;
  assign n45777 = n45776 ^ n45775 ^ n45774 ;
  assign n45778 = n28300 ^ n8434 ^ 1'b0 ;
  assign n45779 = ( n3695 & ~n25078 ) | ( n3695 & n28651 ) | ( ~n25078 & n28651 ) ;
  assign n45780 = ( n13112 & ~n21120 ) | ( n13112 & n45779 ) | ( ~n21120 & n45779 ) ;
  assign n45781 = n37788 ^ n12030 ^ n4473 ;
  assign n45782 = n45781 ^ n16649 ^ 1'b0 ;
  assign n45783 = n16346 | n37991 ;
  assign n45784 = n15383 ^ n2397 ^ 1'b0 ;
  assign n45785 = n13138 | n45784 ;
  assign n45786 = n45785 ^ n22126 ^ n14083 ;
  assign n45787 = n18180 | n45786 ;
  assign n45788 = n15270 | n33041 ;
  assign n45789 = ~n2891 & n45788 ;
  assign n45790 = n45789 ^ n3997 ^ 1'b0 ;
  assign n45791 = ( ~n8984 & n32643 ) | ( ~n8984 & n45790 ) | ( n32643 & n45790 ) ;
  assign n45792 = n37459 ^ n7598 ^ 1'b0 ;
  assign n45793 = n16671 & ~n43882 ;
  assign n45794 = n26009 ^ n16868 ^ n16036 ;
  assign n45795 = n36800 ^ n16828 ^ n10759 ;
  assign n45796 = ( n3651 & ~n24685 ) | ( n3651 & n35852 ) | ( ~n24685 & n35852 ) ;
  assign n45797 = n45796 ^ n44933 ^ 1'b0 ;
  assign n45798 = ( n7820 & n31948 ) | ( n7820 & n35195 ) | ( n31948 & n35195 ) ;
  assign n45799 = n45798 ^ n42888 ^ n399 ;
  assign n45800 = n2637 & ~n33516 ;
  assign n45801 = ~n44233 & n45800 ;
  assign n45802 = n30297 ^ n9677 ^ 1'b0 ;
  assign n45803 = ~n10731 & n45802 ;
  assign n45804 = ( n22229 & ~n26086 ) | ( n22229 & n34242 ) | ( ~n26086 & n34242 ) ;
  assign n45806 = n26535 ^ n24621 ^ n4375 ;
  assign n45807 = n45806 ^ n40025 ^ n16783 ;
  assign n45805 = ( ~n15608 & n23250 ) | ( ~n15608 & n41153 ) | ( n23250 & n41153 ) ;
  assign n45808 = n45807 ^ n45805 ^ n10636 ;
  assign n45809 = n45808 ^ n10326 ^ 1'b0 ;
  assign n45810 = n23080 ^ n20176 ^ n2248 ;
  assign n45811 = n45810 ^ n23575 ^ 1'b0 ;
  assign n45812 = n5400 & n6475 ;
  assign n45813 = n5138 & n45812 ;
  assign n45814 = ( n31936 & n32280 ) | ( n31936 & ~n45813 ) | ( n32280 & ~n45813 ) ;
  assign n45815 = ( n1893 & n12116 ) | ( n1893 & ~n40382 ) | ( n12116 & ~n40382 ) ;
  assign n45816 = n19746 & ~n45815 ;
  assign n45817 = ( n22038 & n45814 ) | ( n22038 & ~n45816 ) | ( n45814 & ~n45816 ) ;
  assign n45818 = ( n14782 & n27252 ) | ( n14782 & n45817 ) | ( n27252 & n45817 ) ;
  assign n45819 = ( n2059 & n3417 ) | ( n2059 & ~n15864 ) | ( n3417 & ~n15864 ) ;
  assign n45820 = n45819 ^ n14029 ^ n6407 ;
  assign n45821 = n45820 ^ n34258 ^ n3427 ;
  assign n45822 = n42963 ^ n18854 ^ 1'b0 ;
  assign n45823 = n43617 & ~n45822 ;
  assign n45824 = n28604 ^ n22646 ^ 1'b0 ;
  assign n45826 = ( ~n3102 & n5872 ) | ( ~n3102 & n16205 ) | ( n5872 & n16205 ) ;
  assign n45825 = n10740 ^ n7548 ^ 1'b0 ;
  assign n45827 = n45826 ^ n45825 ^ n19506 ;
  assign n45828 = n43260 ^ n37323 ^ n31742 ;
  assign n45829 = n45828 ^ n13607 ^ n4590 ;
  assign n45830 = n38559 & ~n45829 ;
  assign n45831 = ( n8634 & ~n11474 ) | ( n8634 & n15198 ) | ( ~n11474 & n15198 ) ;
  assign n45832 = n45831 ^ n20841 ^ n12343 ;
  assign n45833 = n19350 ^ n11411 ^ n6785 ;
  assign n45834 = ( n15008 & n15528 ) | ( n15008 & n45833 ) | ( n15528 & n45833 ) ;
  assign n45835 = n277 & ~n16161 ;
  assign n45836 = n45835 ^ n24454 ^ 1'b0 ;
  assign n45837 = ~n11960 & n27456 ;
  assign n45838 = n45837 ^ n38709 ^ 1'b0 ;
  assign n45839 = n1554 & n2436 ;
  assign n45840 = n3326 & ~n45839 ;
  assign n45841 = n10849 ^ n9235 ^ n9223 ;
  assign n45842 = ( ~n18435 & n19193 ) | ( ~n18435 & n45841 ) | ( n19193 & n45841 ) ;
  assign n45843 = x125 | n45842 ;
  assign n45844 = ~n33836 & n45843 ;
  assign n45845 = ( n7973 & n25831 ) | ( n7973 & ~n36177 ) | ( n25831 & ~n36177 ) ;
  assign n45846 = n21575 ^ n6258 ^ n5132 ;
  assign n45847 = n45846 ^ n9537 ^ n1528 ;
  assign n45848 = n45847 ^ n18523 ^ 1'b0 ;
  assign n45849 = n45200 ^ n20434 ^ n16667 ;
  assign n45850 = ( n2658 & n7115 ) | ( n2658 & ~n27918 ) | ( n7115 & ~n27918 ) ;
  assign n45851 = n31907 ^ n19488 ^ n2018 ;
  assign n45852 = n45851 ^ n22180 ^ n9711 ;
  assign n45853 = ( n16649 & ~n34841 ) | ( n16649 & n45852 ) | ( ~n34841 & n45852 ) ;
  assign n45854 = ( n3715 & n18105 ) | ( n3715 & n25369 ) | ( n18105 & n25369 ) ;
  assign n45855 = ~n14149 & n45854 ;
  assign n45856 = n7709 & n45855 ;
  assign n45858 = n14352 ^ n388 ^ 1'b0 ;
  assign n45857 = ~n10666 & n12973 ;
  assign n45859 = n45858 ^ n45857 ^ 1'b0 ;
  assign n45860 = ~n3398 & n41685 ;
  assign n45861 = n42481 & n45860 ;
  assign n45862 = n35683 ^ n31714 ^ n8856 ;
  assign n45863 = n37766 ^ n31678 ^ n18877 ;
  assign n45864 = ( n24116 & n44814 ) | ( n24116 & ~n45863 ) | ( n44814 & ~n45863 ) ;
  assign n45865 = n45864 ^ n10777 ^ n7755 ;
  assign n45866 = n5460 ^ n3887 ^ 1'b0 ;
  assign n45867 = n18148 & n45866 ;
  assign n45868 = ( n11944 & n22221 ) | ( n11944 & ~n45867 ) | ( n22221 & ~n45867 ) ;
  assign n45869 = n45868 ^ n42662 ^ n33676 ;
  assign n45873 = ( ~n8051 & n26958 ) | ( ~n8051 & n42626 ) | ( n26958 & n42626 ) ;
  assign n45870 = ~n23266 & n30148 ;
  assign n45871 = n45870 ^ n11566 ^ 1'b0 ;
  assign n45872 = n22036 | n45871 ;
  assign n45874 = n45873 ^ n45872 ^ n13250 ;
  assign n45875 = n27165 ^ n13906 ^ n9183 ;
  assign n45879 = n474 & ~n13740 ;
  assign n45880 = n45879 ^ n18608 ^ 1'b0 ;
  assign n45876 = n18627 ^ n4570 ^ n4213 ;
  assign n45877 = n45876 ^ n26160 ^ n3971 ;
  assign n45878 = n45877 ^ n28820 ^ 1'b0 ;
  assign n45881 = n45880 ^ n45878 ^ n42907 ;
  assign n45882 = ( n4216 & n9706 ) | ( n4216 & ~n16459 ) | ( n9706 & ~n16459 ) ;
  assign n45883 = ( n3010 & n33165 ) | ( n3010 & n45882 ) | ( n33165 & n45882 ) ;
  assign n45884 = n13084 | n14045 ;
  assign n45885 = n45884 ^ n30562 ^ 1'b0 ;
  assign n45886 = ( n10978 & ~n13150 ) | ( n10978 & n16117 ) | ( ~n13150 & n16117 ) ;
  assign n45887 = ( ~n4344 & n20296 ) | ( ~n4344 & n40239 ) | ( n20296 & n40239 ) ;
  assign n45888 = n31085 & ~n40794 ;
  assign n45889 = ( n23833 & n40009 ) | ( n23833 & ~n45888 ) | ( n40009 & ~n45888 ) ;
  assign n45890 = ( n13946 & ~n45887 ) | ( n13946 & n45889 ) | ( ~n45887 & n45889 ) ;
  assign n45891 = ( n5676 & n24798 ) | ( n5676 & ~n29390 ) | ( n24798 & ~n29390 ) ;
  assign n45892 = n33226 ^ n20887 ^ n11041 ;
  assign n45893 = n45892 ^ n27878 ^ n19811 ;
  assign n45894 = ( n12765 & n18661 ) | ( n12765 & n40078 ) | ( n18661 & n40078 ) ;
  assign n45895 = n20828 & ~n45894 ;
  assign n45896 = n4397 & n37497 ;
  assign n45897 = n45896 ^ n22981 ^ 1'b0 ;
  assign n45898 = n45897 ^ n22604 ^ 1'b0 ;
  assign n45899 = ( n13582 & ~n29964 ) | ( n13582 & n45898 ) | ( ~n29964 & n45898 ) ;
  assign n45900 = ( n5384 & n29882 ) | ( n5384 & ~n37709 ) | ( n29882 & ~n37709 ) ;
  assign n45901 = n23592 ^ n10030 ^ 1'b0 ;
  assign n45902 = n45900 & ~n45901 ;
  assign n45903 = n45902 ^ n2575 ^ 1'b0 ;
  assign n45904 = ~n22094 & n45903 ;
  assign n45905 = ~n2102 & n11467 ;
  assign n45906 = n45905 ^ n29683 ^ 1'b0 ;
  assign n45907 = n39571 ^ n34046 ^ n14262 ;
  assign n45908 = n14081 ^ n7959 ^ n7890 ;
  assign n45909 = ~n5314 & n20642 ;
  assign n45910 = ( n35773 & ~n45908 ) | ( n35773 & n45909 ) | ( ~n45908 & n45909 ) ;
  assign n45911 = ( n33697 & n37749 ) | ( n33697 & ~n45910 ) | ( n37749 & ~n45910 ) ;
  assign n45912 = n45911 ^ n39939 ^ n15433 ;
  assign n45915 = ( n1742 & n8871 ) | ( n1742 & n39486 ) | ( n8871 & n39486 ) ;
  assign n45913 = n3987 | n32379 ;
  assign n45914 = n45913 ^ n2165 ^ 1'b0 ;
  assign n45916 = n45915 ^ n45914 ^ n19514 ;
  assign n45917 = n45916 ^ n15535 ^ 1'b0 ;
  assign n45918 = n7119 | n25798 ;
  assign n45919 = n45918 ^ n4910 ^ n1235 ;
  assign n45920 = ( n13343 & ~n41435 ) | ( n13343 & n45919 ) | ( ~n41435 & n45919 ) ;
  assign n45921 = n15585 & ~n28510 ;
  assign n45922 = n45921 ^ n11007 ^ 1'b0 ;
  assign n45923 = ( n6397 & ~n7577 ) | ( n6397 & n7822 ) | ( ~n7577 & n7822 ) ;
  assign n45924 = n27461 | n45923 ;
  assign n45925 = n18257 ^ n14437 ^ n13345 ;
  assign n45926 = n45925 ^ n5587 ^ n706 ;
  assign n45927 = ( n10205 & n19846 ) | ( n10205 & n40923 ) | ( n19846 & n40923 ) ;
  assign n45928 = n45927 ^ n20210 ^ x156 ;
  assign n45929 = n26811 ^ n3088 ^ 1'b0 ;
  assign n45930 = ( n18029 & n22756 ) | ( n18029 & ~n41334 ) | ( n22756 & ~n41334 ) ;
  assign n45931 = n45930 ^ n11987 ^ 1'b0 ;
  assign n45933 = ( ~n286 & n11017 ) | ( ~n286 & n22498 ) | ( n11017 & n22498 ) ;
  assign n45932 = ( n7613 & n10086 ) | ( n7613 & n21724 ) | ( n10086 & n21724 ) ;
  assign n45934 = n45933 ^ n45932 ^ n6100 ;
  assign n45935 = n45934 ^ n16681 ^ n11470 ;
  assign n45938 = ( n8652 & n8986 ) | ( n8652 & ~n18286 ) | ( n8986 & ~n18286 ) ;
  assign n45936 = n42365 ^ n28808 ^ n12337 ;
  assign n45937 = ~n2024 & n45936 ;
  assign n45939 = n45938 ^ n45937 ^ x39 ;
  assign n45940 = n45863 ^ n11071 ^ n5030 ;
  assign n45941 = ( n13860 & ~n19829 ) | ( n13860 & n45940 ) | ( ~n19829 & n45940 ) ;
  assign n45942 = ( n9011 & n10477 ) | ( n9011 & n37056 ) | ( n10477 & n37056 ) ;
  assign n45943 = n5691 | n6480 ;
  assign n45945 = n36893 ^ n20946 ^ n3568 ;
  assign n45944 = n20955 | n41014 ;
  assign n45946 = n45945 ^ n45944 ^ 1'b0 ;
  assign n45947 = ( n24463 & ~n30747 ) | ( n24463 & n45946 ) | ( ~n30747 & n45946 ) ;
  assign n45948 = ( ~n10028 & n36604 ) | ( ~n10028 & n45947 ) | ( n36604 & n45947 ) ;
  assign n45949 = ( n16558 & n21405 ) | ( n16558 & n41817 ) | ( n21405 & n41817 ) ;
  assign n45951 = n8139 & n36247 ;
  assign n45952 = n45951 ^ n16638 ^ 1'b0 ;
  assign n45950 = ( n2323 & n9787 ) | ( n2323 & n12503 ) | ( n9787 & n12503 ) ;
  assign n45953 = n45952 ^ n45950 ^ n40982 ;
  assign n45954 = n34630 | n45953 ;
  assign n45955 = ( ~n4005 & n9681 ) | ( ~n4005 & n23103 ) | ( n9681 & n23103 ) ;
  assign n45956 = n45955 ^ n30952 ^ n16109 ;
  assign n45957 = n45956 ^ n18859 ^ n3029 ;
  assign n45958 = n32794 ^ n19860 ^ x102 ;
  assign n45959 = ( n21898 & n39738 ) | ( n21898 & n45958 ) | ( n39738 & n45958 ) ;
  assign n45960 = ( n3923 & ~n35981 ) | ( n3923 & n45959 ) | ( ~n35981 & n45959 ) ;
  assign n45961 = ( n12683 & ~n44211 ) | ( n12683 & n45960 ) | ( ~n44211 & n45960 ) ;
  assign n45962 = n13731 & n45961 ;
  assign n45963 = n20245 & n45962 ;
  assign n45964 = ( n2188 & n7470 ) | ( n2188 & ~n34656 ) | ( n7470 & ~n34656 ) ;
  assign n45965 = n31029 ^ n9102 ^ 1'b0 ;
  assign n45966 = n45964 & n45965 ;
  assign n45967 = n26625 ^ n18758 ^ n7048 ;
  assign n45968 = n4920 & n5405 ;
  assign n45969 = ~n45967 & n45968 ;
  assign n45970 = ( ~n28648 & n39016 ) | ( ~n28648 & n41265 ) | ( n39016 & n41265 ) ;
  assign n45971 = n33615 ^ n2632 ^ 1'b0 ;
  assign n45972 = n14651 & n16103 ;
  assign n45973 = n14525 ^ n2982 ^ n1324 ;
  assign n45974 = n45973 ^ n39284 ^ 1'b0 ;
  assign n45976 = n9955 ^ n7265 ^ n5271 ;
  assign n45977 = n45976 ^ n16843 ^ n11906 ;
  assign n45975 = n7795 ^ n3965 ^ n2421 ;
  assign n45978 = n45977 ^ n45975 ^ n32187 ;
  assign n45979 = n45978 ^ n45485 ^ n12201 ;
  assign n45980 = n34640 ^ n24140 ^ n8006 ;
  assign n45981 = n45980 ^ n26339 ^ 1'b0 ;
  assign n45982 = ( n721 & n9091 ) | ( n721 & ~n30278 ) | ( n9091 & ~n30278 ) ;
  assign n45983 = ( n7162 & ~n24228 ) | ( n7162 & n45982 ) | ( ~n24228 & n45982 ) ;
  assign n45984 = n38044 & ~n43199 ;
  assign n45985 = n25827 & n45984 ;
  assign n45988 = n2973 & n19135 ;
  assign n45989 = n45988 ^ n29151 ^ 1'b0 ;
  assign n45986 = n11090 & ~n22010 ;
  assign n45987 = n45986 ^ n3543 ^ 1'b0 ;
  assign n45990 = n45989 ^ n45987 ^ n30378 ;
  assign n45991 = n35413 & ~n45990 ;
  assign n45992 = n45991 ^ n14300 ^ 1'b0 ;
  assign n45993 = n45992 ^ n33940 ^ n18903 ;
  assign n45994 = n39494 & ~n45993 ;
  assign n45995 = ~n14379 & n45994 ;
  assign n45996 = n27303 ^ n6269 ^ 1'b0 ;
  assign n45997 = n18395 | n36074 ;
  assign n45998 = ( ~n5164 & n8333 ) | ( ~n5164 & n14520 ) | ( n8333 & n14520 ) ;
  assign n45999 = n26298 ^ n14723 ^ 1'b0 ;
  assign n46000 = n13203 & ~n45999 ;
  assign n46001 = ( n2302 & ~n40462 ) | ( n2302 & n46000 ) | ( ~n40462 & n46000 ) ;
  assign n46002 = ( n25798 & ~n45998 ) | ( n25798 & n46001 ) | ( ~n45998 & n46001 ) ;
  assign n46003 = n4019 | n41909 ;
  assign n46004 = n46003 ^ n16262 ^ 1'b0 ;
  assign n46005 = n6801 & ~n12471 ;
  assign n46006 = n46005 ^ n27427 ^ 1'b0 ;
  assign n46007 = n46004 & n46006 ;
  assign n46008 = n13480 ^ n4414 ^ 1'b0 ;
  assign n46009 = n2932 & n46008 ;
  assign n46010 = ( n8494 & n13770 ) | ( n8494 & ~n46009 ) | ( n13770 & ~n46009 ) ;
  assign n46011 = n46010 ^ n27762 ^ n11580 ;
  assign n46012 = ( n6909 & n44790 ) | ( n6909 & ~n46011 ) | ( n44790 & ~n46011 ) ;
  assign n46013 = ( n4344 & n7083 ) | ( n4344 & n24239 ) | ( n7083 & n24239 ) ;
  assign n46014 = n46013 ^ n32936 ^ n8951 ;
  assign n46015 = n31741 ^ n14129 ^ n12496 ;
  assign n46016 = ( ~n11443 & n46014 ) | ( ~n11443 & n46015 ) | ( n46014 & n46015 ) ;
  assign n46017 = n32986 ^ n18471 ^ n17341 ;
  assign n46018 = n46017 ^ n15286 ^ 1'b0 ;
  assign n46019 = ( n7515 & ~n12333 ) | ( n7515 & n18136 ) | ( ~n12333 & n18136 ) ;
  assign n46020 = n46019 ^ n40828 ^ 1'b0 ;
  assign n46021 = n46018 | n46020 ;
  assign n46022 = n34498 ^ n24602 ^ 1'b0 ;
  assign n46023 = n43590 & ~n46022 ;
  assign n46024 = n32243 ^ n27867 ^ n727 ;
  assign n46025 = n20055 ^ n4659 ^ 1'b0 ;
  assign n46026 = n32437 ^ n15269 ^ 1'b0 ;
  assign n46027 = ( n18987 & n26216 ) | ( n18987 & n46026 ) | ( n26216 & n46026 ) ;
  assign n46028 = ( ~n26908 & n46025 ) | ( ~n26908 & n46027 ) | ( n46025 & n46027 ) ;
  assign n46029 = n33993 ^ n14267 ^ x29 ;
  assign n46030 = n46029 ^ n45361 ^ n4853 ;
  assign n46033 = ( ~n11020 & n11304 ) | ( ~n11020 & n14596 ) | ( n11304 & n14596 ) ;
  assign n46034 = n46033 ^ n19636 ^ n4743 ;
  assign n46031 = n26074 ^ n15772 ^ n10890 ;
  assign n46032 = n46031 ^ n25811 ^ n22256 ;
  assign n46035 = n46034 ^ n46032 ^ n36689 ;
  assign n46036 = n29521 ^ n15953 ^ n14501 ;
  assign n46038 = n43108 ^ n30792 ^ n16172 ;
  assign n46037 = ( n14888 & n17630 ) | ( n14888 & n42070 ) | ( n17630 & n42070 ) ;
  assign n46039 = n46038 ^ n46037 ^ n19057 ;
  assign n46040 = ~n45335 & n46039 ;
  assign n46041 = n10673 & n11612 ;
  assign n46044 = n10438 | n25868 ;
  assign n46045 = n29197 & ~n46044 ;
  assign n46042 = ( n16974 & ~n22026 ) | ( n16974 & n34296 ) | ( ~n22026 & n34296 ) ;
  assign n46043 = n46042 ^ n31136 ^ 1'b0 ;
  assign n46046 = n46045 ^ n46043 ^ n31806 ;
  assign n46047 = n38705 ^ n30599 ^ n23229 ;
  assign n46048 = ( n9673 & n10382 ) | ( n9673 & ~n16922 ) | ( n10382 & ~n16922 ) ;
  assign n46049 = ( n13462 & n32701 ) | ( n13462 & n46048 ) | ( n32701 & n46048 ) ;
  assign n46050 = ( n9642 & ~n13593 ) | ( n9642 & n46049 ) | ( ~n13593 & n46049 ) ;
  assign n46051 = n22747 ^ n20817 ^ n14306 ;
  assign n46052 = n46051 ^ n21798 ^ n4015 ;
  assign n46053 = ( n46047 & n46050 ) | ( n46047 & ~n46052 ) | ( n46050 & ~n46052 ) ;
  assign n46054 = ~n10118 & n37553 ;
  assign n46055 = n46054 ^ n28050 ^ 1'b0 ;
  assign n46056 = n33073 ^ n24026 ^ n14109 ;
  assign n46057 = ( n18940 & n19203 ) | ( n18940 & ~n46056 ) | ( n19203 & ~n46056 ) ;
  assign n46058 = n38650 ^ n26389 ^ n6575 ;
  assign n46059 = ( n4176 & n27177 ) | ( n4176 & n44410 ) | ( n27177 & n44410 ) ;
  assign n46060 = ( n6164 & n7266 ) | ( n6164 & n32975 ) | ( n7266 & n32975 ) ;
  assign n46061 = ( n25815 & n28428 ) | ( n25815 & n46060 ) | ( n28428 & n46060 ) ;
  assign n46062 = ( ~n9944 & n14187 ) | ( ~n9944 & n33062 ) | ( n14187 & n33062 ) ;
  assign n46063 = n14323 & ~n46062 ;
  assign n46064 = ~n19184 & n46063 ;
  assign n46065 = x185 & ~n3696 ;
  assign n46066 = ~n29924 & n46065 ;
  assign n46067 = ( n11314 & n45666 ) | ( n11314 & ~n46066 ) | ( n45666 & ~n46066 ) ;
  assign n46068 = n6848 ^ n1837 ^ n487 ;
  assign n46069 = n836 & n46068 ;
  assign n46070 = ~n46067 & n46069 ;
  assign n46071 = n42687 ^ n36150 ^ n25384 ;
  assign n46072 = n28890 & ~n46071 ;
  assign n46073 = n46072 ^ n35734 ^ 1'b0 ;
  assign n46074 = n36185 ^ n32036 ^ n13844 ;
  assign n46075 = n15460 | n18185 ;
  assign n46076 = n12290 & ~n46075 ;
  assign n46077 = ( n29291 & n34828 ) | ( n29291 & ~n46076 ) | ( n34828 & ~n46076 ) ;
  assign n46078 = n46077 ^ n18609 ^ n9817 ;
  assign n46079 = n46078 ^ n23587 ^ n16540 ;
  assign n46080 = n42347 ^ n31476 ^ 1'b0 ;
  assign n46081 = n19558 ^ n1731 ^ 1'b0 ;
  assign n46082 = ~n25061 & n46081 ;
  assign n46083 = ( n6747 & n9379 ) | ( n6747 & n39248 ) | ( n9379 & n39248 ) ;
  assign n46084 = n46083 ^ n17519 ^ n445 ;
  assign n46085 = ( n2617 & ~n12221 ) | ( n2617 & n41170 ) | ( ~n12221 & n41170 ) ;
  assign n46086 = n46085 ^ n23903 ^ n13331 ;
  assign n46087 = ( ~n9033 & n27192 ) | ( ~n9033 & n29970 ) | ( n27192 & n29970 ) ;
  assign n46088 = n46087 ^ n9120 ^ n7287 ;
  assign n46089 = n23359 ^ n17849 ^ n15772 ;
  assign n46090 = ( n3695 & ~n19469 ) | ( n3695 & n46089 ) | ( ~n19469 & n46089 ) ;
  assign n46091 = n14368 & ~n36019 ;
  assign n46092 = n46090 & n46091 ;
  assign n46093 = n31596 ^ n19687 ^ 1'b0 ;
  assign n46094 = n30220 ^ n10290 ^ 1'b0 ;
  assign n46095 = n27111 ^ n19971 ^ x85 ;
  assign n46096 = n35588 ^ n32164 ^ n1057 ;
  assign n46097 = n43635 ^ n37616 ^ n12307 ;
  assign n46098 = n46097 ^ n39714 ^ 1'b0 ;
  assign n46099 = n38732 ^ n17936 ^ n14791 ;
  assign n46100 = ( n1667 & n15829 ) | ( n1667 & n45809 ) | ( n15829 & n45809 ) ;
  assign n46102 = ( n11593 & n25214 ) | ( n11593 & n30548 ) | ( n25214 & n30548 ) ;
  assign n46101 = ~n4576 & n17005 ;
  assign n46103 = n46102 ^ n46101 ^ 1'b0 ;
  assign n46104 = n7637 | n46103 ;
  assign n46105 = n18982 & ~n46104 ;
  assign n46106 = ( n6074 & ~n12841 ) | ( n6074 & n15076 ) | ( ~n12841 & n15076 ) ;
  assign n46107 = n46106 ^ n16887 ^ n3749 ;
  assign n46108 = n15048 | n46107 ;
  assign n46109 = n46108 ^ n32457 ^ 1'b0 ;
  assign n46110 = ( ~n1828 & n23210 ) | ( ~n1828 & n28391 ) | ( n23210 & n28391 ) ;
  assign n46111 = ( x39 & ~n38914 ) | ( x39 & n46110 ) | ( ~n38914 & n46110 ) ;
  assign n46112 = n13968 ^ n13782 ^ n2472 ;
  assign n46113 = n46112 ^ n17754 ^ n16849 ;
  assign n46114 = n46113 ^ n21936 ^ 1'b0 ;
  assign n46115 = n14462 ^ n7673 ^ n7315 ;
  assign n46116 = ( n14407 & n19188 ) | ( n14407 & n46115 ) | ( n19188 & n46115 ) ;
  assign n46118 = n20956 ^ n18603 ^ n906 ;
  assign n46117 = n793 | n11210 ;
  assign n46119 = n46118 ^ n46117 ^ x46 ;
  assign n46120 = n14398 ^ n7904 ^ n6285 ;
  assign n46121 = n20079 ^ n8719 ^ 1'b0 ;
  assign n46122 = n3528 & n46121 ;
  assign n46123 = n46122 ^ n33947 ^ n4915 ;
  assign n46124 = n38954 ^ n9512 ^ n8786 ;
  assign n46125 = n26798 ^ n14899 ^ 1'b0 ;
  assign n46126 = n46125 ^ n36469 ^ n6824 ;
  assign n46127 = n25262 ^ n14322 ^ n1212 ;
  assign n46128 = n36350 & n46127 ;
  assign n46129 = n46128 ^ n6573 ^ n1276 ;
  assign n46130 = ( ~n20764 & n22185 ) | ( ~n20764 & n46129 ) | ( n22185 & n46129 ) ;
  assign n46131 = n37880 ^ n36824 ^ 1'b0 ;
  assign n46132 = ( n21030 & ~n44934 ) | ( n21030 & n46131 ) | ( ~n44934 & n46131 ) ;
  assign n46133 = n34175 ^ n22026 ^ n6394 ;
  assign n46134 = n13756 ^ n8269 ^ x168 ;
  assign n46135 = n11128 ^ n8728 ^ n2760 ;
  assign n46136 = ( ~n19008 & n29289 ) | ( ~n19008 & n35600 ) | ( n29289 & n35600 ) ;
  assign n46137 = ( n4843 & ~n46135 ) | ( n4843 & n46136 ) | ( ~n46135 & n46136 ) ;
  assign n46138 = n380 | n21300 ;
  assign n46139 = n46137 | n46138 ;
  assign n46140 = n12920 & n13203 ;
  assign n46141 = ~n15710 & n46140 ;
  assign n46142 = ( ~x103 & n1084 ) | ( ~x103 & n3517 ) | ( n1084 & n3517 ) ;
  assign n46143 = n46142 ^ n30505 ^ n19181 ;
  assign n46144 = n46143 ^ n11504 ^ n3454 ;
  assign n46145 = ( n1614 & ~n6423 ) | ( n1614 & n13735 ) | ( ~n6423 & n13735 ) ;
  assign n46146 = ( n1879 & ~n16101 ) | ( n1879 & n17715 ) | ( ~n16101 & n17715 ) ;
  assign n46147 = n25093 ^ n18255 ^ n5807 ;
  assign n46148 = n45833 ^ n40406 ^ n33273 ;
  assign n46149 = ( n13101 & n14772 ) | ( n13101 & ~n26751 ) | ( n14772 & ~n26751 ) ;
  assign n46150 = n20591 ^ n17847 ^ n15976 ;
  assign n46151 = ( n530 & n16626 ) | ( n530 & n22875 ) | ( n16626 & n22875 ) ;
  assign n46152 = n14605 | n19824 ;
  assign n46153 = n24956 ^ n11163 ^ n1233 ;
  assign n46154 = ~n19754 & n46153 ;
  assign n46155 = ~n46152 & n46154 ;
  assign n46156 = n12444 | n43734 ;
  assign n46157 = n7396 & ~n46156 ;
  assign n46158 = ~n2743 & n11791 ;
  assign n46159 = n1460 & n46158 ;
  assign n46160 = n46159 ^ n43090 ^ n27980 ;
  assign n46161 = n12848 ^ n12184 ^ n5568 ;
  assign n46162 = ( n16847 & ~n17734 ) | ( n16847 & n46161 ) | ( ~n17734 & n46161 ) ;
  assign n46163 = n14987 & ~n37143 ;
  assign n46164 = ( ~n18539 & n44605 ) | ( ~n18539 & n46163 ) | ( n44605 & n46163 ) ;
  assign n46165 = ( n44051 & n46162 ) | ( n44051 & n46164 ) | ( n46162 & n46164 ) ;
  assign n46166 = n36413 ^ n19551 ^ n1324 ;
  assign n46167 = n35600 ^ n19232 ^ n14228 ;
  assign n46168 = n46167 ^ n13105 ^ n11918 ;
  assign n46169 = n46168 ^ n25672 ^ n922 ;
  assign n46170 = ( ~n9583 & n15512 ) | ( ~n9583 & n46169 ) | ( n15512 & n46169 ) ;
  assign n46171 = n44637 ^ n23383 ^ n16375 ;
  assign n46172 = n45771 ^ n44603 ^ n1744 ;
  assign n46173 = n21863 ^ n21161 ^ n6675 ;
  assign n46174 = ~n4283 & n15023 ;
  assign n46175 = n46174 ^ n25366 ^ 1'b0 ;
  assign n46176 = ~n1216 & n46175 ;
  assign n46177 = n46176 ^ n8383 ^ 1'b0 ;
  assign n46178 = ( n2827 & ~n6272 ) | ( n2827 & n17875 ) | ( ~n6272 & n17875 ) ;
  assign n46179 = n46178 ^ n33760 ^ n13985 ;
  assign n46181 = n38111 ^ n26544 ^ n16574 ;
  assign n46180 = ( ~n11988 & n22466 ) | ( ~n11988 & n23397 ) | ( n22466 & n23397 ) ;
  assign n46182 = n46181 ^ n46180 ^ 1'b0 ;
  assign n46183 = ( ~n1987 & n11517 ) | ( ~n1987 & n45152 ) | ( n11517 & n45152 ) ;
  assign n46184 = n46183 ^ n36500 ^ n36184 ;
  assign n46185 = ( n841 & ~n4712 ) | ( n841 & n10242 ) | ( ~n4712 & n10242 ) ;
  assign n46186 = ( n14650 & n22468 ) | ( n14650 & n46185 ) | ( n22468 & n46185 ) ;
  assign n46187 = ( n430 & n9036 ) | ( n430 & ~n20405 ) | ( n9036 & ~n20405 ) ;
  assign n46188 = ( n21694 & ~n34651 ) | ( n21694 & n46187 ) | ( ~n34651 & n46187 ) ;
  assign n46189 = n46188 ^ n33440 ^ n6848 ;
  assign n46190 = n40551 ^ n4689 ^ 1'b0 ;
  assign n46191 = n11830 & ~n46190 ;
  assign n46192 = ~n14122 & n22230 ;
  assign n46193 = ~n18845 & n46192 ;
  assign n46194 = n15774 ^ n8048 ^ 1'b0 ;
  assign n46195 = ~n3484 & n46194 ;
  assign n46196 = n39910 ^ n36095 ^ n3250 ;
  assign n46197 = ( n9922 & ~n10681 ) | ( n9922 & n30595 ) | ( ~n10681 & n30595 ) ;
  assign n46198 = ( x112 & n36537 ) | ( x112 & n46197 ) | ( n36537 & n46197 ) ;
  assign n46199 = n46198 ^ n44463 ^ n13393 ;
  assign n46200 = n29310 ^ n18156 ^ n6349 ;
  assign n46201 = n19325 ^ n10694 ^ n10067 ;
  assign n46202 = n28930 ^ n24896 ^ n10886 ;
  assign n46203 = ( ~n2551 & n36644 ) | ( ~n2551 & n46202 ) | ( n36644 & n46202 ) ;
  assign n46204 = n42953 ^ n18162 ^ 1'b0 ;
  assign n46205 = n21286 | n46204 ;
  assign n46206 = ( x47 & n5679 ) | ( x47 & ~n10812 ) | ( n5679 & ~n10812 ) ;
  assign n46207 = n46206 ^ n21208 ^ 1'b0 ;
  assign n46208 = n3957 & n46207 ;
  assign n46209 = n1111 & ~n17750 ;
  assign n46210 = n37924 ^ n14050 ^ 1'b0 ;
  assign n46211 = ( n18352 & n19251 ) | ( n18352 & n23744 ) | ( n19251 & n23744 ) ;
  assign n46212 = ( n46209 & n46210 ) | ( n46209 & ~n46211 ) | ( n46210 & ~n46211 ) ;
  assign n46213 = n6274 & n11504 ;
  assign n46214 = n46213 ^ n35355 ^ n1008 ;
  assign n46215 = n14835 ^ n9567 ^ n4791 ;
  assign n46216 = n46215 ^ n33949 ^ n2091 ;
  assign n46217 = ( n34107 & n45372 ) | ( n34107 & ~n46216 ) | ( n45372 & ~n46216 ) ;
  assign n46218 = n38046 ^ n33849 ^ n31444 ;
  assign n46219 = ( ~n9013 & n25966 ) | ( ~n9013 & n46218 ) | ( n25966 & n46218 ) ;
  assign n46220 = ( n2272 & n24112 ) | ( n2272 & ~n34766 ) | ( n24112 & ~n34766 ) ;
  assign n46221 = ( ~n28079 & n28475 ) | ( ~n28079 & n46220 ) | ( n28475 & n46220 ) ;
  assign n46222 = n9241 & ~n46221 ;
  assign n46223 = n46222 ^ n7830 ^ 1'b0 ;
  assign n46225 = ( n18844 & ~n39356 ) | ( n18844 & n43073 ) | ( ~n39356 & n43073 ) ;
  assign n46224 = n7501 & n9041 ;
  assign n46226 = n46225 ^ n46224 ^ 1'b0 ;
  assign n46227 = n46226 ^ n41138 ^ n36196 ;
  assign n46228 = ( n7281 & n46223 ) | ( n7281 & n46227 ) | ( n46223 & n46227 ) ;
  assign n46229 = n5098 ^ n1152 ^ 1'b0 ;
  assign n46230 = n46229 ^ n39819 ^ n20081 ;
  assign n46231 = n32138 ^ n11271 ^ n2998 ;
  assign n46232 = n46231 ^ n36230 ^ n31101 ;
  assign n46233 = n27473 & n33422 ;
  assign n46234 = ~n2677 & n46233 ;
  assign n46235 = n37899 ^ n7016 ^ 1'b0 ;
  assign n46236 = n3005 & ~n46235 ;
  assign n46237 = ~n31239 & n46236 ;
  assign n46238 = n20957 & n46237 ;
  assign n46240 = n23628 ^ n9611 ^ n7039 ;
  assign n46239 = ~n12354 & n29540 ;
  assign n46241 = n46240 ^ n46239 ^ n22846 ;
  assign n46244 = n34426 ^ n14967 ^ n12112 ;
  assign n46242 = n38307 ^ n22443 ^ n13409 ;
  assign n46243 = n46242 ^ n22267 ^ n12871 ;
  assign n46245 = n46244 ^ n46243 ^ n20055 ;
  assign n46246 = n43261 ^ n31730 ^ 1'b0 ;
  assign n46247 = n18241 ^ n15025 ^ 1'b0 ;
  assign n46248 = ~n20868 & n46247 ;
  assign n46249 = ( n899 & n12238 ) | ( n899 & n16203 ) | ( n12238 & n16203 ) ;
  assign n46250 = ( ~n46246 & n46248 ) | ( ~n46246 & n46249 ) | ( n46248 & n46249 ) ;
  assign n46251 = ( ~n13110 & n23854 ) | ( ~n13110 & n39716 ) | ( n23854 & n39716 ) ;
  assign n46252 = n45024 ^ n14813 ^ n5274 ;
  assign n46253 = n18648 & n43221 ;
  assign n46254 = ~n40647 & n46253 ;
  assign n46255 = n46161 ^ n27136 ^ n6577 ;
  assign n46256 = n36945 ^ n35990 ^ n9264 ;
  assign n46257 = n16755 & n37847 ;
  assign n46258 = ~n3672 & n46257 ;
  assign n46259 = ( ~n7477 & n12506 ) | ( ~n7477 & n46258 ) | ( n12506 & n46258 ) ;
  assign n46260 = n26566 & ~n46259 ;
  assign n46261 = n17764 & ~n46260 ;
  assign n46262 = n37004 ^ n20337 ^ n8532 ;
  assign n46263 = ( n10134 & ~n12283 ) | ( n10134 & n42665 ) | ( ~n12283 & n42665 ) ;
  assign n46264 = n37528 ^ n21081 ^ n4466 ;
  assign n46265 = ( ~n1612 & n10882 ) | ( ~n1612 & n31930 ) | ( n10882 & n31930 ) ;
  assign n46266 = ( n9140 & ~n28285 ) | ( n9140 & n46265 ) | ( ~n28285 & n46265 ) ;
  assign n46267 = n46266 ^ n7063 ^ 1'b0 ;
  assign n46268 = ( n5264 & ~n46264 ) | ( n5264 & n46267 ) | ( ~n46264 & n46267 ) ;
  assign n46269 = ( ~n21851 & n23740 ) | ( ~n21851 & n46268 ) | ( n23740 & n46268 ) ;
  assign n46270 = n46269 ^ n26267 ^ n1530 ;
  assign n46271 = n36467 ^ n4099 ^ n2628 ;
  assign n46272 = n40647 ^ n27989 ^ 1'b0 ;
  assign n46273 = n13133 ^ n12245 ^ 1'b0 ;
  assign n46274 = ~n45673 & n46273 ;
  assign n46275 = ~n38711 & n46274 ;
  assign n46276 = ~n11277 & n46275 ;
  assign n46277 = ( ~n26785 & n27858 ) | ( ~n26785 & n41442 ) | ( n27858 & n41442 ) ;
  assign n46278 = n19498 & n38599 ;
  assign n46279 = n19182 | n28803 ;
  assign n46280 = n46279 ^ n37707 ^ 1'b0 ;
  assign n46281 = ( n12077 & n45410 ) | ( n12077 & ~n46280 ) | ( n45410 & ~n46280 ) ;
  assign n46282 = ( n34003 & n46278 ) | ( n34003 & ~n46281 ) | ( n46278 & ~n46281 ) ;
  assign n46283 = n9262 ^ n5512 ^ x139 ;
  assign n46284 = n22935 ^ n17827 ^ n748 ;
  assign n46285 = ( n23992 & n31823 ) | ( n23992 & ~n46284 ) | ( n31823 & ~n46284 ) ;
  assign n46286 = n13681 ^ n2432 ^ n2212 ;
  assign n46287 = ( n1717 & n8473 ) | ( n1717 & n46286 ) | ( n8473 & n46286 ) ;
  assign n46288 = n46287 ^ n12044 ^ n6899 ;
  assign n46289 = ( n3185 & n17183 ) | ( n3185 & n24122 ) | ( n17183 & n24122 ) ;
  assign n46290 = n20959 & ~n46289 ;
  assign n46291 = n46290 ^ n36644 ^ n7415 ;
  assign n46292 = n26351 ^ n11711 ^ 1'b0 ;
  assign n46293 = n46292 ^ n44399 ^ n11448 ;
  assign n46294 = n4575 & ~n33957 ;
  assign n46295 = n46294 ^ n8839 ^ 1'b0 ;
  assign n46296 = n11440 ^ n10820 ^ n2937 ;
  assign n46297 = ( ~n20105 & n22056 ) | ( ~n20105 & n46296 ) | ( n22056 & n46296 ) ;
  assign n46298 = n9783 | n16187 ;
  assign n46299 = ( ~n6684 & n44202 ) | ( ~n6684 & n46298 ) | ( n44202 & n46298 ) ;
  assign n46300 = n46299 ^ n9964 ^ n9494 ;
  assign n46301 = n44055 ^ n10651 ^ 1'b0 ;
  assign n46302 = n10824 | n41509 ;
  assign n46303 = n46302 ^ n2570 ^ 1'b0 ;
  assign n46304 = ( n12845 & n40197 ) | ( n12845 & ~n46303 ) | ( n40197 & ~n46303 ) ;
  assign n46305 = n29214 ^ n14306 ^ n9114 ;
  assign n46306 = n44943 ^ n30654 ^ n8127 ;
  assign n46307 = n6018 & ~n24360 ;
  assign n46308 = ~n3599 & n46307 ;
  assign n46309 = n19726 & n46308 ;
  assign n46310 = ( n29282 & n46306 ) | ( n29282 & ~n46309 ) | ( n46306 & ~n46309 ) ;
  assign n46311 = n46310 ^ n7682 ^ n5061 ;
  assign n46312 = ( n19216 & ~n46305 ) | ( n19216 & n46311 ) | ( ~n46305 & n46311 ) ;
  assign n46313 = n42556 ^ n39632 ^ n26828 ;
  assign n46314 = n29078 ^ n11164 ^ n2315 ;
  assign n46315 = n46314 ^ n21556 ^ 1'b0 ;
  assign n46316 = n17545 & n38689 ;
  assign n46318 = n27679 ^ n17248 ^ n6703 ;
  assign n46317 = n11166 & n11218 ;
  assign n46319 = n46318 ^ n46317 ^ n5942 ;
  assign n46320 = n11520 ^ n8551 ^ 1'b0 ;
  assign n46321 = n5894 | n46320 ;
  assign n46322 = n2005 & ~n46321 ;
  assign n46323 = ( n2598 & n5603 ) | ( n2598 & n16120 ) | ( n5603 & n16120 ) ;
  assign n46324 = ( n23431 & ~n34521 ) | ( n23431 & n46323 ) | ( ~n34521 & n46323 ) ;
  assign n46325 = n25425 ^ n16774 ^ 1'b0 ;
  assign n46326 = n27040 | n46071 ;
  assign n46327 = ( n5132 & ~n46325 ) | ( n5132 & n46326 ) | ( ~n46325 & n46326 ) ;
  assign n46328 = ~n623 & n25604 ;
  assign n46329 = n20875 ^ n19415 ^ 1'b0 ;
  assign n46330 = ( n11347 & ~n12716 ) | ( n11347 & n46329 ) | ( ~n12716 & n46329 ) ;
  assign n46331 = n12882 & ~n22877 ;
  assign n46332 = n46331 ^ n39377 ^ 1'b0 ;
  assign n46333 = ( n446 & ~n4340 ) | ( n446 & n23682 ) | ( ~n4340 & n23682 ) ;
  assign n46334 = n46333 ^ n18083 ^ n10122 ;
  assign n46335 = n10924 & ~n24268 ;
  assign n46336 = n46335 ^ n34258 ^ 1'b0 ;
  assign n46337 = n37425 & ~n46336 ;
  assign n46338 = n13724 ^ n11132 ^ n10801 ;
  assign n46339 = n46338 ^ n22457 ^ n11061 ;
  assign n46340 = n33673 ^ n18536 ^ n11814 ;
  assign n46341 = ( n6148 & ~n19591 ) | ( n6148 & n26607 ) | ( ~n19591 & n26607 ) ;
  assign n46342 = ~n25737 & n46341 ;
  assign n46343 = n37504 & n39891 ;
  assign n46344 = ( n1830 & ~n23355 ) | ( n1830 & n46343 ) | ( ~n23355 & n46343 ) ;
  assign n46345 = n23417 ^ n15642 ^ n15314 ;
  assign n46346 = ( ~n24579 & n25235 ) | ( ~n24579 & n46345 ) | ( n25235 & n46345 ) ;
  assign n46347 = n24029 ^ n22597 ^ n8692 ;
  assign n46348 = n1955 & n32349 ;
  assign n46349 = n17794 & n23408 ;
  assign n46350 = n7700 & n14339 ;
  assign n46351 = n46350 ^ n18943 ^ n2799 ;
  assign n46352 = n11340 & ~n28434 ;
  assign n46353 = ( n14738 & ~n46351 ) | ( n14738 & n46352 ) | ( ~n46351 & n46352 ) ;
  assign n46354 = ( n7627 & ~n14698 ) | ( n7627 & n36562 ) | ( ~n14698 & n36562 ) ;
  assign n46355 = n34591 | n39117 ;
  assign n46356 = n35137 & ~n46355 ;
  assign n46357 = ( ~n12341 & n39356 ) | ( ~n12341 & n46356 ) | ( n39356 & n46356 ) ;
  assign n46358 = ( n26626 & n38597 ) | ( n26626 & n46357 ) | ( n38597 & n46357 ) ;
  assign n46359 = ( n6014 & n15581 ) | ( n6014 & ~n40167 ) | ( n15581 & ~n40167 ) ;
  assign n46360 = n24372 ^ n15767 ^ n2076 ;
  assign n46361 = ( n1790 & n28434 ) | ( n1790 & n36640 ) | ( n28434 & n36640 ) ;
  assign n46362 = ( ~n11014 & n33715 ) | ( ~n11014 & n46361 ) | ( n33715 & n46361 ) ;
  assign n46363 = n13819 & ~n27497 ;
  assign n46364 = n46363 ^ n4156 ^ 1'b0 ;
  assign n46365 = n19594 ^ n13687 ^ n6196 ;
  assign n46366 = ( n498 & ~n7821 ) | ( n498 & n23325 ) | ( ~n7821 & n23325 ) ;
  assign n46367 = n46366 ^ n35754 ^ n18379 ;
  assign n46368 = ( n12770 & ~n22095 ) | ( n12770 & n33111 ) | ( ~n22095 & n33111 ) ;
  assign n46369 = n46368 ^ n38370 ^ n35930 ;
  assign n46370 = n28120 ^ n26063 ^ n25939 ;
  assign n46371 = n23584 ^ n2710 ^ n312 ;
  assign n46372 = n46371 ^ n17834 ^ 1'b0 ;
  assign n46373 = n41915 ^ n35587 ^ n2315 ;
  assign n46374 = n32425 ^ n11088 ^ n716 ;
  assign n46375 = n46374 ^ n42218 ^ n12620 ;
  assign n46376 = n9770 & n21377 ;
  assign n46377 = n9260 ^ n6290 ^ 1'b0 ;
  assign n46379 = ( n9896 & ~n19711 ) | ( n9896 & n36497 ) | ( ~n19711 & n36497 ) ;
  assign n46380 = ( n25043 & ~n42529 ) | ( n25043 & n46379 ) | ( ~n42529 & n46379 ) ;
  assign n46381 = n46380 ^ n28830 ^ n22767 ;
  assign n46378 = n36123 ^ n20764 ^ n11528 ;
  assign n46382 = n46381 ^ n46378 ^ n12247 ;
  assign n46383 = ( n12885 & n21353 ) | ( n12885 & n30942 ) | ( n21353 & n30942 ) ;
  assign n46384 = ( n25232 & ~n38908 ) | ( n25232 & n46383 ) | ( ~n38908 & n46383 ) ;
  assign n46385 = n13173 ^ n5267 ^ n3019 ;
  assign n46386 = n1751 | n9027 ;
  assign n46387 = n46386 ^ n4835 ^ 1'b0 ;
  assign n46388 = n46387 ^ n12811 ^ n12531 ;
  assign n46389 = ~n1440 & n12107 ;
  assign n46390 = ~n28312 & n46389 ;
  assign n46391 = n14614 | n46390 ;
  assign n46392 = n35876 ^ n29288 ^ n8710 ;
  assign n46393 = n28771 ^ n19424 ^ n1512 ;
  assign n46397 = n4072 & ~n7062 ;
  assign n46398 = n46397 ^ n37900 ^ n34487 ;
  assign n46394 = n43412 ^ n20399 ^ n2161 ;
  assign n46395 = ~n7685 & n46394 ;
  assign n46396 = n34759 & n46395 ;
  assign n46399 = n46398 ^ n46396 ^ n45424 ;
  assign n46400 = n38092 ^ n21658 ^ n8858 ;
  assign n46401 = ( ~n12039 & n14088 ) | ( ~n12039 & n46400 ) | ( n14088 & n46400 ) ;
  assign n46402 = n2159 | n2437 ;
  assign n46403 = n7368 | n46402 ;
  assign n46404 = n40015 & n46403 ;
  assign n46405 = n32261 ^ n30004 ^ n12370 ;
  assign n46406 = n38213 | n46405 ;
  assign n46407 = n38678 ^ n7687 ^ n1898 ;
  assign n46408 = ( n7495 & n28101 ) | ( n7495 & ~n46407 ) | ( n28101 & ~n46407 ) ;
  assign n46409 = n43611 ^ n35582 ^ n4408 ;
  assign n46410 = ( ~n17736 & n38344 ) | ( ~n17736 & n46409 ) | ( n38344 & n46409 ) ;
  assign n46411 = ( n42800 & n46408 ) | ( n42800 & n46410 ) | ( n46408 & n46410 ) ;
  assign n46412 = n2008 ^ n832 ^ n830 ;
  assign n46413 = n22510 ^ n13965 ^ n12046 ;
  assign n46414 = n17801 ^ n3995 ^ 1'b0 ;
  assign n46415 = n46413 | n46414 ;
  assign n46416 = n3487 | n46415 ;
  assign n46417 = n46416 ^ n4017 ^ 1'b0 ;
  assign n46418 = n43904 ^ n20857 ^ n16799 ;
  assign n46419 = n4500 & ~n46418 ;
  assign n46420 = ~n1197 & n21461 ;
  assign n46421 = ( n9135 & ~n25472 ) | ( n9135 & n46420 ) | ( ~n25472 & n46420 ) ;
  assign n46422 = n40653 ^ n31311 ^ n9683 ;
  assign n46423 = n46422 ^ n38636 ^ n34682 ;
  assign n46424 = n46318 ^ n33836 ^ 1'b0 ;
  assign n46425 = n46424 ^ n7762 ^ n4476 ;
  assign n46426 = n42303 ^ n35341 ^ n13940 ;
  assign n46427 = ~n19064 & n43835 ;
  assign n46428 = ( x97 & ~n46426 ) | ( x97 & n46427 ) | ( ~n46426 & n46427 ) ;
  assign n46429 = n13781 & ~n38591 ;
  assign n46430 = n16047 ^ n11399 ^ n2080 ;
  assign n46431 = ( n23181 & ~n27634 ) | ( n23181 & n46430 ) | ( ~n27634 & n46430 ) ;
  assign n46432 = n44168 ^ n23707 ^ n11608 ;
  assign n46433 = ( n17275 & ~n46431 ) | ( n17275 & n46432 ) | ( ~n46431 & n46432 ) ;
  assign n46434 = n13237 | n18608 ;
  assign n46435 = n46434 ^ n33976 ^ 1'b0 ;
  assign n46436 = n5777 | n13738 ;
  assign n46437 = n46435 & ~n46436 ;
  assign n46438 = n28983 ^ n10165 ^ 1'b0 ;
  assign n46439 = n25205 | n46438 ;
  assign n46440 = ( n14839 & ~n17703 ) | ( n14839 & n18664 ) | ( ~n17703 & n18664 ) ;
  assign n46441 = ( n11530 & n37243 ) | ( n11530 & n46440 ) | ( n37243 & n46440 ) ;
  assign n46442 = ( n713 & n7062 ) | ( n713 & ~n22336 ) | ( n7062 & ~n22336 ) ;
  assign n46443 = ( n15331 & n22108 ) | ( n15331 & ~n24508 ) | ( n22108 & ~n24508 ) ;
  assign n46447 = ( ~n9418 & n20299 ) | ( ~n9418 & n36452 ) | ( n20299 & n36452 ) ;
  assign n46444 = ~n2364 & n30727 ;
  assign n46445 = n43470 ^ n43136 ^ 1'b0 ;
  assign n46446 = n46444 | n46445 ;
  assign n46448 = n46447 ^ n46446 ^ n1601 ;
  assign n46449 = n21925 ^ n14343 ^ n10111 ;
  assign n46450 = n16733 & n46449 ;
  assign n46451 = n20002 | n46450 ;
  assign n46452 = n21591 ^ n20086 ^ n7530 ;
  assign n46453 = ( n11214 & n13799 ) | ( n11214 & n18860 ) | ( n13799 & n18860 ) ;
  assign n46454 = n46453 ^ n25761 ^ n6707 ;
  assign n46455 = n43103 ^ n28345 ^ n6096 ;
  assign n46456 = n32439 ^ n17966 ^ n8884 ;
  assign n46457 = n11731 & n46456 ;
  assign n46458 = n46457 ^ n13847 ^ 1'b0 ;
  assign n46463 = n42777 ^ n525 ^ 1'b0 ;
  assign n46464 = n20109 | n46463 ;
  assign n46465 = n46464 ^ n1785 ^ 1'b0 ;
  assign n46459 = n498 & n7834 ;
  assign n46460 = n46459 ^ n30046 ^ 1'b0 ;
  assign n46461 = ( ~n1726 & n13905 ) | ( ~n1726 & n46460 ) | ( n13905 & n46460 ) ;
  assign n46462 = ( n25498 & ~n28663 ) | ( n25498 & n46461 ) | ( ~n28663 & n46461 ) ;
  assign n46466 = n46465 ^ n46462 ^ n36339 ;
  assign n46467 = n25181 & n26445 ;
  assign n46468 = ( ~n835 & n2933 ) | ( ~n835 & n30115 ) | ( n2933 & n30115 ) ;
  assign n46469 = n46468 ^ n12833 ^ n7048 ;
  assign n46470 = ( n2794 & n10154 ) | ( n2794 & n10642 ) | ( n10154 & n10642 ) ;
  assign n46471 = x132 & n31495 ;
  assign n46472 = ( ~n7125 & n9861 ) | ( ~n7125 & n46471 ) | ( n9861 & n46471 ) ;
  assign n46473 = n46472 ^ n45288 ^ n2703 ;
  assign n46474 = n23927 ^ n20871 ^ n11114 ;
  assign n46475 = ( n6620 & n31326 ) | ( n6620 & n46474 ) | ( n31326 & n46474 ) ;
  assign n46482 = ( ~n1561 & n1588 ) | ( ~n1561 & n21529 ) | ( n1588 & n21529 ) ;
  assign n46483 = n46482 ^ n18738 ^ 1'b0 ;
  assign n46484 = n7297 & ~n46483 ;
  assign n46485 = n46484 ^ n7217 ^ n5289 ;
  assign n46486 = ( ~n15598 & n18136 ) | ( ~n15598 & n46485 ) | ( n18136 & n46485 ) ;
  assign n46478 = n15677 | n19757 ;
  assign n46479 = n41699 | n46478 ;
  assign n46480 = n46479 ^ n46266 ^ n20713 ;
  assign n46481 = ( n17856 & n33976 ) | ( n17856 & ~n46480 ) | ( n33976 & ~n46480 ) ;
  assign n46487 = n46486 ^ n46481 ^ n36557 ;
  assign n46476 = n15027 ^ n10643 ^ n7562 ;
  assign n46477 = n8530 & n46476 ;
  assign n46488 = n46487 ^ n46477 ^ 1'b0 ;
  assign n46490 = n8035 ^ n2704 ^ x25 ;
  assign n46489 = n25080 ^ n10444 ^ 1'b0 ;
  assign n46491 = n46490 ^ n46489 ^ 1'b0 ;
  assign n46498 = n33158 ^ n26387 ^ 1'b0 ;
  assign n46492 = n21829 ^ n4454 ^ 1'b0 ;
  assign n46493 = n12343 | n46492 ;
  assign n46494 = n46493 ^ n22747 ^ 1'b0 ;
  assign n46495 = ( n9683 & ~n14677 ) | ( n9683 & n46494 ) | ( ~n14677 & n46494 ) ;
  assign n46496 = n44037 & ~n46495 ;
  assign n46497 = n46496 ^ n46468 ^ 1'b0 ;
  assign n46499 = n46498 ^ n46497 ^ n7426 ;
  assign n46502 = n39016 ^ n12281 ^ n7272 ;
  assign n46503 = n46502 ^ n21439 ^ n13625 ;
  assign n46500 = n33521 & n44605 ;
  assign n46501 = ~n43592 & n46500 ;
  assign n46504 = n46503 ^ n46501 ^ n43065 ;
  assign n46505 = n29884 ^ n16696 ^ 1'b0 ;
  assign n46506 = n20509 & n37153 ;
  assign n46507 = n46506 ^ n18389 ^ 1'b0 ;
  assign n46508 = ~n46505 & n46507 ;
  assign n46509 = n46508 ^ n1822 ^ 1'b0 ;
  assign n46510 = n31317 ^ n10671 ^ n9868 ;
  assign n46511 = n46510 ^ n5558 ^ 1'b0 ;
  assign n46512 = n2920 & n46511 ;
  assign n46513 = n46512 ^ n21698 ^ n2593 ;
  assign n46514 = ( n33253 & ~n33510 ) | ( n33253 & n42551 ) | ( ~n33510 & n42551 ) ;
  assign n46515 = ( n5056 & n45546 ) | ( n5056 & ~n46514 ) | ( n45546 & ~n46514 ) ;
  assign n46516 = n46515 ^ n43718 ^ 1'b0 ;
  assign n46517 = n46516 ^ n7672 ^ n600 ;
  assign n46523 = ( n7137 & n15929 ) | ( n7137 & ~n16276 ) | ( n15929 & ~n16276 ) ;
  assign n46524 = ( ~n2708 & n12555 ) | ( ~n2708 & n46523 ) | ( n12555 & n46523 ) ;
  assign n46520 = n14069 ^ n7034 ^ n2325 ;
  assign n46521 = n46520 ^ n2280 ^ 1'b0 ;
  assign n46518 = ( n6336 & n9588 ) | ( n6336 & ~n41213 ) | ( n9588 & ~n41213 ) ;
  assign n46519 = n46518 ^ n7738 ^ 1'b0 ;
  assign n46522 = n46521 ^ n46519 ^ n24922 ;
  assign n46525 = n46524 ^ n46522 ^ n42422 ;
  assign n46526 = n12710 | n27685 ;
  assign n46527 = n33615 & ~n46526 ;
  assign n46528 = n6550 & n9968 ;
  assign n46529 = n1352 & n46528 ;
  assign n46530 = n28988 ^ n6069 ^ 1'b0 ;
  assign n46531 = n38264 & ~n46530 ;
  assign n46532 = ~n25314 & n34498 ;
  assign n46533 = ~n28124 & n46532 ;
  assign n46534 = ( n23012 & n35330 ) | ( n23012 & ~n46533 ) | ( n35330 & ~n46533 ) ;
  assign n46535 = n22198 & n29064 ;
  assign n46536 = ~n798 & n46535 ;
  assign n46537 = n46536 ^ n2477 ^ 1'b0 ;
  assign n46538 = n46018 ^ n38778 ^ n9132 ;
  assign n46539 = n46537 & n46538 ;
  assign n46540 = n42509 ^ n18937 ^ n18212 ;
  assign n46541 = n36134 ^ n18997 ^ n503 ;
  assign n46548 = ( n835 & n6549 ) | ( n835 & n7478 ) | ( n6549 & n7478 ) ;
  assign n46545 = n46440 ^ n29036 ^ n19581 ;
  assign n46546 = ( n28196 & n39665 ) | ( n28196 & n46545 ) | ( n39665 & n46545 ) ;
  assign n46544 = n41509 ^ n27506 ^ n18206 ;
  assign n46542 = ( n7204 & n10712 ) | ( n7204 & n14118 ) | ( n10712 & n14118 ) ;
  assign n46543 = ( n19496 & ~n34117 ) | ( n19496 & n46542 ) | ( ~n34117 & n46542 ) ;
  assign n46547 = n46546 ^ n46544 ^ n46543 ;
  assign n46549 = n46548 ^ n46547 ^ n22002 ;
  assign n46550 = n38632 ^ n21937 ^ 1'b0 ;
  assign n46551 = n46550 ^ n29411 ^ n2268 ;
  assign n46552 = ( n5004 & ~n17743 ) | ( n5004 & n18265 ) | ( ~n17743 & n18265 ) ;
  assign n46553 = ( n37982 & n45910 ) | ( n37982 & ~n46552 ) | ( n45910 & ~n46552 ) ;
  assign n46554 = n28142 ^ n19236 ^ n3733 ;
  assign n46555 = ~n4208 & n23611 ;
  assign n46556 = ~n46554 & n46555 ;
  assign n46557 = n46553 & n46556 ;
  assign n46558 = n5953 & ~n9749 ;
  assign n46559 = n46558 ^ n19112 ^ 1'b0 ;
  assign n46560 = ( n20923 & ~n24164 ) | ( n20923 & n40915 ) | ( ~n24164 & n40915 ) ;
  assign n46561 = n32841 & n46560 ;
  assign n46568 = ( n5549 & ~n10318 ) | ( n5549 & n23471 ) | ( ~n10318 & n23471 ) ;
  assign n46569 = ~n6067 & n46568 ;
  assign n46567 = ( n3360 & n12733 ) | ( n3360 & n28706 ) | ( n12733 & n28706 ) ;
  assign n46570 = n46569 ^ n46567 ^ n3546 ;
  assign n46564 = n30350 ^ n29151 ^ n19113 ;
  assign n46565 = ( ~n4713 & n30265 ) | ( ~n4713 & n46564 ) | ( n30265 & n46564 ) ;
  assign n46562 = ~n19031 & n21071 ;
  assign n46563 = n9714 & n46562 ;
  assign n46566 = n46565 ^ n46563 ^ n9067 ;
  assign n46571 = n46570 ^ n46566 ^ 1'b0 ;
  assign n46572 = n13370 & ~n34413 ;
  assign n46573 = n46572 ^ n5829 ^ 1'b0 ;
  assign n46574 = ( n26131 & n42277 ) | ( n26131 & ~n46573 ) | ( n42277 & ~n46573 ) ;
  assign n46575 = ( n1246 & n22701 ) | ( n1246 & n39082 ) | ( n22701 & n39082 ) ;
  assign n46576 = n32368 ^ n6374 ^ n2219 ;
  assign n46577 = ( n18357 & n35736 ) | ( n18357 & ~n46576 ) | ( n35736 & ~n46576 ) ;
  assign n46578 = ( n397 & n11541 ) | ( n397 & n43128 ) | ( n11541 & n43128 ) ;
  assign n46579 = n31112 ^ n18583 ^ n16461 ;
  assign n46580 = ( ~n9177 & n24256 ) | ( ~n9177 & n46579 ) | ( n24256 & n46579 ) ;
  assign n46581 = n28123 | n36840 ;
  assign n46582 = n27781 ^ n21258 ^ 1'b0 ;
  assign n46583 = n46582 ^ n19829 ^ n7385 ;
  assign n46584 = n23273 ^ n19042 ^ 1'b0 ;
  assign n46585 = ~n15844 & n46584 ;
  assign n46586 = n8348 ^ n5546 ^ n2016 ;
  assign n46587 = n17824 & n23552 ;
  assign n46588 = n46586 & n46587 ;
  assign n46589 = n19039 & n19817 ;
  assign n46590 = n46589 ^ n34511 ^ n29922 ;
  assign n46591 = ( n6773 & n16597 ) | ( n6773 & n17717 ) | ( n16597 & n17717 ) ;
  assign n46592 = n6036 | n18690 ;
  assign n46593 = n46592 ^ n15930 ^ 1'b0 ;
  assign n46594 = ( n2066 & n46591 ) | ( n2066 & ~n46593 ) | ( n46591 & ~n46593 ) ;
  assign n46595 = n46594 ^ n40655 ^ 1'b0 ;
  assign n46596 = n46590 & ~n46595 ;
  assign n46597 = ~n11715 & n35213 ;
  assign n46598 = n46597 ^ n4034 ^ 1'b0 ;
  assign n46599 = ( ~n6158 & n16728 ) | ( ~n6158 & n46598 ) | ( n16728 & n46598 ) ;
  assign n46600 = ( n3084 & n4695 ) | ( n3084 & ~n12620 ) | ( n4695 & ~n12620 ) ;
  assign n46601 = n46600 ^ x246 ^ 1'b0 ;
  assign n46602 = n46599 & n46601 ;
  assign n46603 = ( n42070 & ~n45026 ) | ( n42070 & n46602 ) | ( ~n45026 & n46602 ) ;
  assign n46604 = n28184 & ~n30655 ;
  assign n46605 = ( n11243 & n45349 ) | ( n11243 & n46604 ) | ( n45349 & n46604 ) ;
  assign n46606 = n43199 ^ n35392 ^ n26403 ;
  assign n46607 = n35223 ^ n22735 ^ n3383 ;
  assign n46609 = n24896 & ~n41023 ;
  assign n46610 = n46609 ^ n10376 ^ 1'b0 ;
  assign n46608 = ( ~n8082 & n8419 ) | ( ~n8082 & n43652 ) | ( n8419 & n43652 ) ;
  assign n46611 = n46610 ^ n46608 ^ n6856 ;
  assign n46612 = ( x151 & n8100 ) | ( x151 & ~n12795 ) | ( n8100 & ~n12795 ) ;
  assign n46613 = n28433 ^ n23566 ^ n10212 ;
  assign n46614 = ( n27824 & n30813 ) | ( n27824 & ~n46613 ) | ( n30813 & ~n46613 ) ;
  assign n46615 = n39643 ^ n8233 ^ n6208 ;
  assign n46616 = n46615 ^ n36891 ^ n28355 ;
  assign n46617 = ( x55 & ~n5661 ) | ( x55 & n10447 ) | ( ~n5661 & n10447 ) ;
  assign n46618 = n46617 ^ n16943 ^ n11392 ;
  assign n46619 = n46618 ^ n10277 ^ 1'b0 ;
  assign n46620 = ~n46616 & n46619 ;
  assign n46621 = n46620 ^ n487 ^ 1'b0 ;
  assign n46622 = n27257 ^ n21921 ^ n1122 ;
  assign n46626 = ( ~n5734 & n7274 ) | ( ~n5734 & n15015 ) | ( n7274 & n15015 ) ;
  assign n46624 = n24136 ^ n8729 ^ 1'b0 ;
  assign n46625 = n46624 ^ n35483 ^ n31964 ;
  assign n46623 = n40876 ^ n30340 ^ n7331 ;
  assign n46627 = n46626 ^ n46625 ^ n46623 ;
  assign n46628 = n25259 ^ n17594 ^ 1'b0 ;
  assign n46629 = n17886 & n46628 ;
  assign n46630 = n19625 ^ n16091 ^ n7799 ;
  assign n46631 = ( n13022 & n46629 ) | ( n13022 & n46630 ) | ( n46629 & n46630 ) ;
  assign n46632 = ~n15697 & n29209 ;
  assign n46633 = n8245 & ~n46632 ;
  assign n46634 = n318 | n30197 ;
  assign n46635 = n28935 | n46634 ;
  assign n46636 = n30180 ^ n7703 ^ 1'b0 ;
  assign n46637 = n18424 | n46636 ;
  assign n46639 = n11766 & ~n22575 ;
  assign n46638 = n46206 ^ n18969 ^ 1'b0 ;
  assign n46640 = n46639 ^ n46638 ^ n32663 ;
  assign n46641 = ( n3820 & n4314 ) | ( n3820 & ~n15535 ) | ( n4314 & ~n15535 ) ;
  assign n46642 = n607 & n1353 ;
  assign n46643 = n46642 ^ n43256 ^ 1'b0 ;
  assign n46644 = ( ~n19431 & n35602 ) | ( ~n19431 & n46643 ) | ( n35602 & n46643 ) ;
  assign n46645 = n46644 ^ n14393 ^ n12798 ;
  assign n46646 = n21637 ^ n14206 ^ n14153 ;
  assign n46647 = n46646 ^ n40802 ^ n16532 ;
  assign n46648 = n5650 & ~n46647 ;
  assign n46649 = n46648 ^ n12947 ^ n546 ;
  assign n46650 = n23112 ^ n16433 ^ 1'b0 ;
  assign n46651 = n46650 ^ n30720 ^ n12437 ;
  assign n46652 = ~n2979 & n6313 ;
  assign n46653 = n46652 ^ n12235 ^ n6417 ;
  assign n46654 = n46653 ^ n45115 ^ n24586 ;
  assign n46656 = n11425 ^ n8846 ^ n571 ;
  assign n46655 = n26576 ^ n7593 ^ n4758 ;
  assign n46657 = n46656 ^ n46655 ^ n30024 ;
  assign n46658 = n9890 ^ n1430 ^ 1'b0 ;
  assign n46659 = ~n19902 & n46658 ;
  assign n46660 = n31733 & n38384 ;
  assign n46661 = ~n46659 & n46660 ;
  assign n46662 = ~n11044 & n14016 ;
  assign n46663 = ~n22761 & n46662 ;
  assign n46664 = n35355 ^ n9059 ^ 1'b0 ;
  assign n46665 = ( n682 & n46663 ) | ( n682 & ~n46664 ) | ( n46663 & ~n46664 ) ;
  assign n46666 = n33091 ^ n11907 ^ n4037 ;
  assign n46667 = ( n2797 & n12340 ) | ( n2797 & n46666 ) | ( n12340 & n46666 ) ;
  assign n46669 = ( ~n3630 & n17056 ) | ( ~n3630 & n18697 ) | ( n17056 & n18697 ) ;
  assign n46668 = n18912 ^ n15646 ^ n2909 ;
  assign n46670 = n46669 ^ n46668 ^ n22829 ;
  assign n46671 = ( n24604 & n46403 ) | ( n24604 & ~n46670 ) | ( n46403 & ~n46670 ) ;
  assign n46672 = ( ~n16884 & n23308 ) | ( ~n16884 & n25960 ) | ( n23308 & n25960 ) ;
  assign n46673 = n46672 ^ n23802 ^ n8448 ;
  assign n46674 = n45339 ^ n1404 ^ n1402 ;
  assign n46675 = n26051 ^ n1106 ^ 1'b0 ;
  assign n46676 = ( n6047 & n23537 ) | ( n6047 & n46675 ) | ( n23537 & n46675 ) ;
  assign n46677 = ( n2758 & n23105 ) | ( n2758 & n38032 ) | ( n23105 & n38032 ) ;
  assign n46678 = ~n10270 & n46677 ;
  assign n46679 = ~n33836 & n46678 ;
  assign n46680 = n6816 | n44988 ;
  assign n46681 = n46680 ^ n9437 ^ 1'b0 ;
  assign n46682 = n14339 ^ n8629 ^ x175 ;
  assign n46683 = n46682 ^ n44650 ^ 1'b0 ;
  assign n46684 = n9203 | n11577 ;
  assign n46685 = n46684 ^ n6445 ^ n1501 ;
  assign n46686 = n26203 ^ n10320 ^ n4799 ;
  assign n46687 = n46686 ^ n41911 ^ n20224 ;
  assign n46688 = n46687 ^ n25771 ^ 1'b0 ;
  assign n46689 = n11046 ^ n7746 ^ 1'b0 ;
  assign n46690 = ( n15631 & n38753 ) | ( n15631 & ~n46689 ) | ( n38753 & ~n46689 ) ;
  assign n46691 = n36211 ^ n20315 ^ n1504 ;
  assign n46692 = n46691 ^ n19491 ^ n18818 ;
  assign n46693 = ( n7606 & n17278 ) | ( n7606 & n46692 ) | ( n17278 & n46692 ) ;
  assign n46694 = n28128 ^ n15742 ^ 1'b0 ;
  assign n46695 = n16982 & ~n33669 ;
  assign n46696 = n46695 ^ n42751 ^ 1'b0 ;
  assign n46697 = n6143 & n13020 ;
  assign n46698 = ( n11335 & n11826 ) | ( n11335 & n29464 ) | ( n11826 & n29464 ) ;
  assign n46699 = ( n669 & ~n7562 ) | ( n669 & n10236 ) | ( ~n7562 & n10236 ) ;
  assign n46700 = n46699 ^ n9928 ^ 1'b0 ;
  assign n46701 = n46698 | n46700 ;
  assign n46702 = n3035 & ~n46701 ;
  assign n46703 = ~n46697 & n46702 ;
  assign n46704 = n32334 ^ n20031 ^ n5264 ;
  assign n46705 = n25716 ^ n12856 ^ n10692 ;
  assign n46706 = ( n36696 & ~n46704 ) | ( n36696 & n46705 ) | ( ~n46704 & n46705 ) ;
  assign n46707 = n9284 ^ n7695 ^ n4162 ;
  assign n46708 = ~n42560 & n46707 ;
  assign n46709 = n16745 ^ n14153 ^ n2883 ;
  assign n46710 = ( n2703 & ~n14295 ) | ( n2703 & n32862 ) | ( ~n14295 & n32862 ) ;
  assign n46711 = n26087 & ~n40845 ;
  assign n46712 = ( n340 & n11702 ) | ( n340 & ~n46711 ) | ( n11702 & ~n46711 ) ;
  assign n46713 = n20540 ^ n16088 ^ 1'b0 ;
  assign n46714 = n25412 ^ n10380 ^ 1'b0 ;
  assign n46722 = n6443 ^ n4511 ^ n3317 ;
  assign n46723 = n46722 ^ n32703 ^ n11769 ;
  assign n46724 = n20230 ^ n7384 ^ 1'b0 ;
  assign n46725 = n46723 & ~n46724 ;
  assign n46717 = n33188 | n43457 ;
  assign n46718 = n21811 & ~n46717 ;
  assign n46719 = n2891 | n46718 ;
  assign n46720 = n42792 | n46719 ;
  assign n46715 = ~n4269 & n9916 ;
  assign n46716 = n46715 ^ n44476 ^ 1'b0 ;
  assign n46721 = n46720 ^ n46716 ^ n6366 ;
  assign n46726 = n46725 ^ n46721 ^ n31594 ;
  assign n46727 = ( n5123 & n31901 ) | ( n5123 & n41291 ) | ( n31901 & n41291 ) ;
  assign n46728 = ( n1514 & n20181 ) | ( n1514 & ~n31608 ) | ( n20181 & ~n31608 ) ;
  assign n46729 = n33256 ^ n31574 ^ n17500 ;
  assign n46730 = n11332 ^ n5350 ^ 1'b0 ;
  assign n46731 = n21265 & ~n46730 ;
  assign n46732 = ( n1157 & n19952 ) | ( n1157 & n46731 ) | ( n19952 & n46731 ) ;
  assign n46733 = ( n15465 & n20750 ) | ( n15465 & ~n33701 ) | ( n20750 & ~n33701 ) ;
  assign n46734 = ~n11492 & n36561 ;
  assign n46735 = ~n19910 & n46734 ;
  assign n46736 = n36254 ^ n512 ^ 1'b0 ;
  assign n46737 = n41883 | n46736 ;
  assign n46738 = ( n3262 & n5522 ) | ( n3262 & n9858 ) | ( n5522 & n9858 ) ;
  assign n46739 = ( n6164 & n16333 ) | ( n6164 & n46738 ) | ( n16333 & n46738 ) ;
  assign n46740 = n5671 & ~n46739 ;
  assign n46741 = n29948 ^ n6167 ^ n753 ;
  assign n46742 = ( n2497 & ~n23412 ) | ( n2497 & n39166 ) | ( ~n23412 & n39166 ) ;
  assign n46743 = n16495 ^ n1112 ^ 1'b0 ;
  assign n46744 = ( n46741 & ~n46742 ) | ( n46741 & n46743 ) | ( ~n46742 & n46743 ) ;
  assign n46746 = n9044 ^ n4677 ^ n926 ;
  assign n46747 = n2307 ^ n1741 ^ x124 ;
  assign n46748 = ( n9913 & n46746 ) | ( n9913 & n46747 ) | ( n46746 & n46747 ) ;
  assign n46745 = ( n5331 & n20850 ) | ( n5331 & n23967 ) | ( n20850 & n23967 ) ;
  assign n46749 = n46748 ^ n46745 ^ n30333 ;
  assign n46750 = ( n2170 & n5506 ) | ( n2170 & ~n18725 ) | ( n5506 & ~n18725 ) ;
  assign n46751 = ~n7331 & n46750 ;
  assign n46752 = n44454 ^ n21801 ^ n21563 ;
  assign n46753 = n11402 & n46752 ;
  assign n46754 = n46751 & n46753 ;
  assign n46755 = n31222 & ~n46754 ;
  assign n46756 = ( n1457 & n17070 ) | ( n1457 & ~n46755 ) | ( n17070 & ~n46755 ) ;
  assign n46760 = n19490 ^ n15419 ^ n5482 ;
  assign n46759 = ~n23430 & n32631 ;
  assign n46757 = n32933 ^ n15608 ^ n11345 ;
  assign n46758 = n46757 ^ n23559 ^ n11386 ;
  assign n46761 = n46760 ^ n46759 ^ n46758 ;
  assign n46762 = ( n33654 & n43916 ) | ( n33654 & n46013 ) | ( n43916 & n46013 ) ;
  assign n46763 = ( ~n9811 & n20375 ) | ( ~n9811 & n44324 ) | ( n20375 & n44324 ) ;
  assign n46764 = ~n13360 & n29201 ;
  assign n46765 = ~n19706 & n46764 ;
  assign n46766 = n41355 ^ n19718 ^ n9749 ;
  assign n46767 = n46766 ^ n46183 ^ n1846 ;
  assign n46768 = n46767 ^ n21998 ^ n14154 ;
  assign n46769 = ( n9193 & n32337 ) | ( n9193 & ~n37511 ) | ( n32337 & ~n37511 ) ;
  assign n46770 = ( ~n3514 & n6897 ) | ( ~n3514 & n46769 ) | ( n6897 & n46769 ) ;
  assign n46771 = ( n11179 & n19150 ) | ( n11179 & ~n22169 ) | ( n19150 & ~n22169 ) ;
  assign n46772 = ( n10650 & n23503 ) | ( n10650 & n46771 ) | ( n23503 & n46771 ) ;
  assign n46773 = n35657 ^ n34588 ^ n26047 ;
  assign n46774 = ( ~n17338 & n46772 ) | ( ~n17338 & n46773 ) | ( n46772 & n46773 ) ;
  assign n46775 = n3416 | n4192 ;
  assign n46776 = n46775 ^ n16357 ^ 1'b0 ;
  assign n46777 = n26936 ^ n23483 ^ n13496 ;
  assign n46778 = ( n44298 & n46776 ) | ( n44298 & ~n46777 ) | ( n46776 & ~n46777 ) ;
  assign n46779 = ( n1878 & ~n39287 ) | ( n1878 & n40556 ) | ( ~n39287 & n40556 ) ;
  assign n46780 = n21612 & ~n46779 ;
  assign n46781 = n46780 ^ n38350 ^ n26257 ;
  assign n46782 = n27181 ^ n15445 ^ n8732 ;
  assign n46783 = n46782 ^ n20890 ^ n3203 ;
  assign n46784 = n44064 ^ n34828 ^ n23427 ;
  assign n46785 = n18166 ^ x221 ^ 1'b0 ;
  assign n46786 = n21587 | n46785 ;
  assign n46787 = n21870 ^ n15539 ^ 1'b0 ;
  assign n46788 = n38350 | n46787 ;
  assign n46791 = ( n1559 & n11894 ) | ( n1559 & ~n19857 ) | ( n11894 & ~n19857 ) ;
  assign n46792 = n46791 ^ n24825 ^ n20505 ;
  assign n46789 = ( n1474 & n16926 ) | ( n1474 & ~n22393 ) | ( n16926 & ~n22393 ) ;
  assign n46790 = x13 & n46789 ;
  assign n46793 = n46792 ^ n46790 ^ n28781 ;
  assign n46794 = n46617 ^ n6773 ^ 1'b0 ;
  assign n46795 = n22404 & ~n46794 ;
  assign n46796 = n36246 ^ n13636 ^ 1'b0 ;
  assign n46797 = n46795 & ~n46796 ;
  assign n46798 = n5353 | n23991 ;
  assign n46799 = n46798 ^ n12490 ^ 1'b0 ;
  assign n46800 = n46799 ^ n42209 ^ n16427 ;
  assign n46801 = ( n15522 & ~n46797 ) | ( n15522 & n46800 ) | ( ~n46797 & n46800 ) ;
  assign n46802 = n15418 & ~n40700 ;
  assign n46803 = n46802 ^ n46722 ^ n9249 ;
  assign n46804 = n46803 ^ n30058 ^ 1'b0 ;
  assign n46805 = ( ~n8081 & n32855 ) | ( ~n8081 & n36095 ) | ( n32855 & n36095 ) ;
  assign n46806 = n40703 ^ n13687 ^ 1'b0 ;
  assign n46807 = n12230 & n46806 ;
  assign n46808 = ( n1008 & n46805 ) | ( n1008 & ~n46807 ) | ( n46805 & ~n46807 ) ;
  assign n46809 = n15800 ^ n14573 ^ n13861 ;
  assign n46810 = ( n2439 & n4244 ) | ( n2439 & ~n4739 ) | ( n4244 & ~n4739 ) ;
  assign n46813 = n15122 ^ n9020 ^ 1'b0 ;
  assign n46811 = n46017 ^ n25798 ^ n2733 ;
  assign n46812 = n46811 ^ n21306 ^ n16137 ;
  assign n46814 = n46813 ^ n46812 ^ n23470 ;
  assign n46815 = ( n22095 & n46810 ) | ( n22095 & n46814 ) | ( n46810 & n46814 ) ;
  assign n46816 = n1094 & n27368 ;
  assign n46817 = ( ~n4850 & n17473 ) | ( ~n4850 & n19174 ) | ( n17473 & n19174 ) ;
  assign n46818 = n46817 ^ n8891 ^ 1'b0 ;
  assign n46819 = n46816 | n46818 ;
  assign n46820 = n41126 ^ n2911 ^ 1'b0 ;
  assign n46821 = n3476 | n46820 ;
  assign n46822 = n26380 ^ n14484 ^ n3743 ;
  assign n46823 = n25323 ^ n2258 ^ 1'b0 ;
  assign n46824 = n46823 ^ n38341 ^ n32425 ;
  assign n46825 = n46824 ^ n25965 ^ 1'b0 ;
  assign n46826 = n46014 ^ n19039 ^ n15332 ;
  assign n46827 = n46826 ^ n21021 ^ n7979 ;
  assign n46828 = n46827 ^ n43662 ^ n8784 ;
  assign n46829 = n23388 ^ n17440 ^ 1'b0 ;
  assign n46830 = n27924 & ~n46829 ;
  assign n46831 = n46830 ^ n25698 ^ n20850 ;
  assign n46832 = ( n633 & ~n29136 ) | ( n633 & n32545 ) | ( ~n29136 & n32545 ) ;
  assign n46833 = ( n30057 & ~n31689 ) | ( n30057 & n46832 ) | ( ~n31689 & n46832 ) ;
  assign n46834 = n22647 ^ n14886 ^ n12975 ;
  assign n46835 = n2459 & n29204 ;
  assign n46836 = n46835 ^ n8561 ^ 1'b0 ;
  assign n46837 = n5200 ^ n3041 ^ 1'b0 ;
  assign n46838 = n6465 & n46837 ;
  assign n46839 = ( n19188 & ~n31004 ) | ( n19188 & n31876 ) | ( ~n31004 & n31876 ) ;
  assign n46840 = ( n8479 & n38651 ) | ( n8479 & ~n46839 ) | ( n38651 & ~n46839 ) ;
  assign n46841 = n26197 ^ n10783 ^ 1'b0 ;
  assign n46842 = ( n6157 & n11312 ) | ( n6157 & ~n12755 ) | ( n11312 & ~n12755 ) ;
  assign n46843 = ~n11152 & n46842 ;
  assign n46844 = ( n40255 & ~n46841 ) | ( n40255 & n46843 ) | ( ~n46841 & n46843 ) ;
  assign n46845 = n10663 ^ n9840 ^ n3303 ;
  assign n46846 = n46845 ^ n15286 ^ n6745 ;
  assign n46847 = n46846 ^ n8860 ^ n1414 ;
  assign n46848 = n46278 ^ n5489 ^ 1'b0 ;
  assign n46849 = n8482 & ~n46848 ;
  assign n46850 = n18433 & n46849 ;
  assign n46851 = n46850 ^ n5101 ^ 1'b0 ;
  assign n46852 = n46851 ^ n22563 ^ n19515 ;
  assign n46856 = ( n3267 & n16335 ) | ( n3267 & n27854 ) | ( n16335 & n27854 ) ;
  assign n46853 = n7750 & n14982 ;
  assign n46854 = n46853 ^ n34503 ^ 1'b0 ;
  assign n46855 = n46854 ^ n21155 ^ n12661 ;
  assign n46857 = n46856 ^ n46855 ^ n31311 ;
  assign n46858 = n37089 ^ n13856 ^ n1733 ;
  assign n46859 = ~n3108 & n29989 ;
  assign n46860 = n46859 ^ n29871 ^ 1'b0 ;
  assign n46861 = n40137 & ~n40745 ;
  assign n46862 = n46861 ^ n2064 ^ 1'b0 ;
  assign n46863 = n27383 ^ n27017 ^ n7679 ;
  assign n46864 = n46863 ^ n29344 ^ n1731 ;
  assign n46867 = ( n13071 & n14233 ) | ( n13071 & ~n45998 ) | ( n14233 & ~n45998 ) ;
  assign n46865 = n7474 ^ n6167 ^ n5976 ;
  assign n46866 = ( ~n8024 & n15113 ) | ( ~n8024 & n46865 ) | ( n15113 & n46865 ) ;
  assign n46868 = n46867 ^ n46866 ^ n33692 ;
  assign n46869 = ( ~n8573 & n14588 ) | ( ~n8573 & n21292 ) | ( n14588 & n21292 ) ;
  assign n46870 = ( ~n4372 & n39081 ) | ( ~n4372 & n41368 ) | ( n39081 & n41368 ) ;
  assign n46871 = n25995 ^ n20981 ^ n9192 ;
  assign n46872 = ( ~n46869 & n46870 ) | ( ~n46869 & n46871 ) | ( n46870 & n46871 ) ;
  assign n46873 = n21005 ^ n9226 ^ x181 ;
  assign n46874 = n46873 ^ n34004 ^ n9905 ;
  assign n46875 = ~n18320 & n46874 ;
  assign n46876 = n46875 ^ n7582 ^ n5056 ;
  assign n46877 = n17002 ^ n12251 ^ 1'b0 ;
  assign n46878 = n6630 & ~n9636 ;
  assign n46879 = n46878 ^ n22426 ^ 1'b0 ;
  assign n46880 = n15315 & ~n46879 ;
  assign n46881 = n46880 ^ n2151 ^ 1'b0 ;
  assign n46882 = n46881 ^ n39210 ^ n4074 ;
  assign n46883 = n34296 ^ n32118 ^ n711 ;
  assign n46884 = n28717 ^ n1659 ^ 1'b0 ;
  assign n46885 = n46883 & ~n46884 ;
  assign n46887 = n39920 ^ n7182 ^ n2520 ;
  assign n46886 = ~n10188 & n17566 ;
  assign n46888 = n46887 ^ n46886 ^ 1'b0 ;
  assign n46889 = n27814 ^ n17802 ^ 1'b0 ;
  assign n46890 = ~n29651 & n46889 ;
  assign n46891 = ( ~n941 & n13683 ) | ( ~n941 & n37499 ) | ( n13683 & n37499 ) ;
  assign n46892 = ( n4314 & ~n15192 ) | ( n4314 & n46891 ) | ( ~n15192 & n46891 ) ;
  assign n46893 = n46892 ^ n40820 ^ n5308 ;
  assign n46894 = n46893 ^ n32060 ^ n8550 ;
  assign n46895 = ( n9173 & n39841 ) | ( n9173 & n45751 ) | ( n39841 & n45751 ) ;
  assign n46896 = n27978 ^ n11697 ^ n5135 ;
  assign n46898 = n8175 ^ n7757 ^ n6886 ;
  assign n46897 = n2760 | n3878 ;
  assign n46899 = n46898 ^ n46897 ^ n783 ;
  assign n46901 = ( n7364 & n24028 ) | ( n7364 & ~n33911 ) | ( n24028 & ~n33911 ) ;
  assign n46900 = ( n10444 & ~n18251 ) | ( n10444 & n34234 ) | ( ~n18251 & n34234 ) ;
  assign n46902 = n46901 ^ n46900 ^ n29357 ;
  assign n46903 = ( n22367 & ~n25310 ) | ( n22367 & n46902 ) | ( ~n25310 & n46902 ) ;
  assign n46904 = ( n6204 & n7984 ) | ( n6204 & n44084 ) | ( n7984 & n44084 ) ;
  assign n46905 = n27617 ^ n14417 ^ 1'b0 ;
  assign n46906 = n30337 ^ n14308 ^ 1'b0 ;
  assign n46907 = n39615 & n46906 ;
  assign n46910 = ( n1911 & n30007 ) | ( n1911 & n40654 ) | ( n30007 & n40654 ) ;
  assign n46908 = n34207 ^ n16974 ^ n16580 ;
  assign n46909 = n5782 & ~n46908 ;
  assign n46911 = n46910 ^ n46909 ^ 1'b0 ;
  assign n46912 = n3110 | n42376 ;
  assign n46913 = n46912 ^ n2765 ^ 1'b0 ;
  assign n46914 = n18415 ^ n7106 ^ 1'b0 ;
  assign n46915 = n46914 ^ n26365 ^ 1'b0 ;
  assign n46916 = n46915 ^ n39676 ^ n4503 ;
  assign n46917 = n46916 ^ n36644 ^ n9524 ;
  assign n46918 = n1866 & ~n41390 ;
  assign n46919 = n46918 ^ n21065 ^ 1'b0 ;
  assign n46920 = ( n7010 & n9064 ) | ( n7010 & ~n46919 ) | ( n9064 & ~n46919 ) ;
  assign n46923 = n15408 & ~n25091 ;
  assign n46921 = ~n11401 & n39673 ;
  assign n46922 = ( ~n33645 & n37050 ) | ( ~n33645 & n46921 ) | ( n37050 & n46921 ) ;
  assign n46924 = n46923 ^ n46922 ^ n9288 ;
  assign n46926 = n38267 ^ n34469 ^ n15034 ;
  assign n46925 = n37665 ^ n29854 ^ 1'b0 ;
  assign n46927 = n46926 ^ n46925 ^ n36165 ;
  assign n46928 = n39620 ^ n39488 ^ n25561 ;
  assign n46929 = n11267 & ~n38947 ;
  assign n46930 = ~n42351 & n46929 ;
  assign n46931 = n42669 ^ n38067 ^ n37201 ;
  assign n46932 = ( n10538 & n22609 ) | ( n10538 & ~n28847 ) | ( n22609 & ~n28847 ) ;
  assign n46933 = ~n8634 & n34031 ;
  assign n46934 = n46933 ^ n36846 ^ n15134 ;
  assign n46935 = n42530 ^ n2150 ^ n1747 ;
  assign n46936 = n3097 | n10938 ;
  assign n46937 = n41071 & ~n46936 ;
  assign n46938 = n757 & ~n26216 ;
  assign n46939 = n46938 ^ n41912 ^ 1'b0 ;
  assign n46940 = ( n32897 & n46937 ) | ( n32897 & n46939 ) | ( n46937 & n46939 ) ;
  assign n46941 = ( n16442 & n19856 ) | ( n16442 & ~n44988 ) | ( n19856 & ~n44988 ) ;
  assign n46942 = n46941 ^ n7481 ^ 1'b0 ;
  assign n46943 = ~n5134 & n46942 ;
  assign n46944 = n11493 ^ n6156 ^ 1'b0 ;
  assign n46945 = n46944 ^ n34263 ^ 1'b0 ;
  assign n46946 = n43120 & ~n46945 ;
  assign n46947 = ( ~n9075 & n24215 ) | ( ~n9075 & n33436 ) | ( n24215 & n33436 ) ;
  assign n46948 = n46947 ^ n19099 ^ n13880 ;
  assign n46949 = n46948 ^ n21240 ^ 1'b0 ;
  assign n46950 = ( n19783 & n42075 ) | ( n19783 & ~n46949 ) | ( n42075 & ~n46949 ) ;
  assign n46951 = ~n20512 & n39673 ;
  assign n46952 = ( n8094 & n24359 ) | ( n8094 & ~n46951 ) | ( n24359 & ~n46951 ) ;
  assign n46953 = ( ~n2629 & n32000 ) | ( ~n2629 & n44992 ) | ( n32000 & n44992 ) ;
  assign n46954 = ( ~x32 & n31422 ) | ( ~x32 & n34193 ) | ( n31422 & n34193 ) ;
  assign n46958 = ~n1476 & n22226 ;
  assign n46956 = n18547 ^ n11324 ^ 1'b0 ;
  assign n46955 = ~n487 & n25979 ;
  assign n46957 = n46956 ^ n46955 ^ 1'b0 ;
  assign n46959 = n46958 ^ n46957 ^ n41948 ;
  assign n46960 = ( ~n2682 & n18618 ) | ( ~n2682 & n40982 ) | ( n18618 & n40982 ) ;
  assign n46961 = n13973 | n44943 ;
  assign n46962 = ( n24851 & n44014 ) | ( n24851 & ~n46961 ) | ( n44014 & ~n46961 ) ;
  assign n46963 = n46962 ^ n14756 ^ n12465 ;
  assign n46964 = ( n17897 & n42067 ) | ( n17897 & n46963 ) | ( n42067 & n46963 ) ;
  assign n46965 = n26719 ^ n26174 ^ 1'b0 ;
  assign n46966 = n8482 & ~n46965 ;
  assign n46967 = ( n1674 & ~n28554 ) | ( n1674 & n33049 ) | ( ~n28554 & n33049 ) ;
  assign n46968 = n23624 ^ n12240 ^ 1'b0 ;
  assign n46969 = n46865 | n46968 ;
  assign n46970 = n14357 ^ n10465 ^ n1692 ;
  assign n46971 = ( n39778 & n46969 ) | ( n39778 & ~n46970 ) | ( n46969 & ~n46970 ) ;
  assign n46972 = n7644 & ~n14555 ;
  assign n46973 = n46972 ^ n8295 ^ 1'b0 ;
  assign n46974 = ( ~n3229 & n19020 ) | ( ~n3229 & n46973 ) | ( n19020 & n46973 ) ;
  assign n46975 = n30081 ^ n19922 ^ n2500 ;
  assign n46976 = n46975 ^ n12737 ^ 1'b0 ;
  assign n46977 = n43077 ^ n31245 ^ n2916 ;
  assign n46978 = ( n24604 & ~n43150 ) | ( n24604 & n46977 ) | ( ~n43150 & n46977 ) ;
  assign n46979 = n46978 ^ n39050 ^ n27479 ;
  assign n46980 = n35061 ^ n24173 ^ n2035 ;
  assign n46981 = n46980 ^ n10619 ^ n5331 ;
  assign n46982 = ( ~n15616 & n29195 ) | ( ~n15616 & n46981 ) | ( n29195 & n46981 ) ;
  assign n46983 = ( n5950 & n10324 ) | ( n5950 & ~n12995 ) | ( n10324 & ~n12995 ) ;
  assign n46984 = ~n46131 & n46983 ;
  assign n46985 = n8752 & ~n46984 ;
  assign n46986 = ~n22363 & n46985 ;
  assign n46987 = ( ~n17160 & n23296 ) | ( ~n17160 & n46986 ) | ( n23296 & n46986 ) ;
  assign n46988 = n1991 | n12000 ;
  assign n46989 = n46988 ^ n5971 ^ 1'b0 ;
  assign n46990 = ( n14281 & n14635 ) | ( n14281 & n46989 ) | ( n14635 & n46989 ) ;
  assign n46991 = n18496 ^ n15019 ^ 1'b0 ;
  assign n46992 = x78 & n46991 ;
  assign n46993 = n33297 ^ n6519 ^ 1'b0 ;
  assign n46994 = n25821 & ~n46993 ;
  assign n46995 = n42888 ^ n40671 ^ n34651 ;
  assign n46996 = n27473 ^ n22774 ^ n10086 ;
  assign n46997 = n21495 | n46996 ;
  assign n46998 = n41223 ^ n1344 ^ 1'b0 ;
  assign n46999 = ( n10824 & n25614 ) | ( n10824 & n46998 ) | ( n25614 & n46998 ) ;
  assign n47000 = ( n16155 & n24798 ) | ( n16155 & ~n28883 ) | ( n24798 & ~n28883 ) ;
  assign n47001 = n15862 ^ n6797 ^ n5610 ;
  assign n47002 = ( n18013 & n18770 ) | ( n18013 & n47001 ) | ( n18770 & n47001 ) ;
  assign n47003 = ~n2467 & n26499 ;
  assign n47004 = n28888 ^ n26643 ^ 1'b0 ;
  assign n47005 = ( ~n25784 & n28278 ) | ( ~n25784 & n47004 ) | ( n28278 & n47004 ) ;
  assign n47006 = ( n21658 & ~n24818 ) | ( n21658 & n47005 ) | ( ~n24818 & n47005 ) ;
  assign n47007 = ( ~n5978 & n9000 ) | ( ~n5978 & n25161 ) | ( n9000 & n25161 ) ;
  assign n47008 = n47007 ^ n17862 ^ n7297 ;
  assign n47009 = ~n1274 & n10720 ;
  assign n47010 = ~n17939 & n47009 ;
  assign n47012 = ( n7273 & ~n9853 ) | ( n7273 & n32522 ) | ( ~n9853 & n32522 ) ;
  assign n47011 = n7337 & ~n34151 ;
  assign n47013 = n47012 ^ n47011 ^ n28123 ;
  assign n47014 = n32898 ^ n21242 ^ n4755 ;
  assign n47015 = n47014 ^ n14594 ^ n10121 ;
  assign n47016 = ( n9341 & n11478 ) | ( n9341 & n11647 ) | ( n11478 & n11647 ) ;
  assign n47017 = ( n20458 & n32248 ) | ( n20458 & ~n47016 ) | ( n32248 & ~n47016 ) ;
  assign n47018 = ( n6399 & n9405 ) | ( n6399 & n12076 ) | ( n9405 & n12076 ) ;
  assign n47019 = ( ~n40215 & n45651 ) | ( ~n40215 & n47018 ) | ( n45651 & n47018 ) ;
  assign n47020 = ( n22052 & ~n47017 ) | ( n22052 & n47019 ) | ( ~n47017 & n47019 ) ;
  assign n47021 = n22744 ^ n20004 ^ n5673 ;
  assign n47022 = n47021 ^ n30355 ^ n9418 ;
  assign n47023 = n18776 ^ n9363 ^ 1'b0 ;
  assign n47024 = n15469 & ~n47023 ;
  assign n47025 = ( ~n1404 & n13154 ) | ( ~n1404 & n31497 ) | ( n13154 & n31497 ) ;
  assign n47029 = n24370 ^ n10185 ^ n4963 ;
  assign n47030 = ( n34517 & n45909 ) | ( n34517 & ~n47029 ) | ( n45909 & ~n47029 ) ;
  assign n47026 = x147 & ~n33904 ;
  assign n47027 = n47026 ^ n27339 ^ 1'b0 ;
  assign n47028 = n47027 ^ n34845 ^ n22358 ;
  assign n47031 = n47030 ^ n47028 ^ n4264 ;
  assign n47032 = ( ~n47024 & n47025 ) | ( ~n47024 & n47031 ) | ( n47025 & n47031 ) ;
  assign n47033 = n37565 ^ n32724 ^ 1'b0 ;
  assign n47034 = n11696 | n47033 ;
  assign n47035 = n3229 | n47034 ;
  assign n47036 = n24372 & ~n47035 ;
  assign n47037 = n47036 ^ n24207 ^ n14122 ;
  assign n47038 = n43296 ^ n40034 ^ 1'b0 ;
  assign n47039 = n26031 ^ n8046 ^ n4509 ;
  assign n47040 = n24391 ^ n13102 ^ n3461 ;
  assign n47041 = ( ~n4787 & n23293 ) | ( ~n4787 & n47040 ) | ( n23293 & n47040 ) ;
  assign n47042 = ( x166 & n6110 ) | ( x166 & ~n47041 ) | ( n6110 & ~n47041 ) ;
  assign n47043 = n319 & n10532 ;
  assign n47044 = n47043 ^ n14352 ^ n12382 ;
  assign n47045 = n27472 ^ n22366 ^ n16901 ;
  assign n47046 = ( ~n445 & n13740 ) | ( ~n445 & n47045 ) | ( n13740 & n47045 ) ;
  assign n47047 = ( ~n1508 & n30513 ) | ( ~n1508 & n36791 ) | ( n30513 & n36791 ) ;
  assign n47048 = ( ~n12797 & n18377 ) | ( ~n12797 & n47047 ) | ( n18377 & n47047 ) ;
  assign n47049 = n4540 & ~n31296 ;
  assign n47050 = n47049 ^ n14718 ^ 1'b0 ;
  assign n47051 = ( n24638 & n47048 ) | ( n24638 & n47050 ) | ( n47048 & n47050 ) ;
  assign n47055 = n41769 ^ n38929 ^ n27207 ;
  assign n47052 = n3462 | n19539 ;
  assign n47053 = n11332 | n47052 ;
  assign n47054 = ~n20804 & n47053 ;
  assign n47056 = n47055 ^ n47054 ^ 1'b0 ;
  assign n47057 = n4441 & ~n25940 ;
  assign n47058 = ~n42534 & n47057 ;
  assign n47059 = ( n5895 & ~n47056 ) | ( n5895 & n47058 ) | ( ~n47056 & n47058 ) ;
  assign n47060 = n15889 ^ n10334 ^ 1'b0 ;
  assign n47061 = n47060 ^ n41463 ^ n30444 ;
  assign n47062 = n47061 ^ n45640 ^ n31485 ;
  assign n47063 = n16786 & n46551 ;
  assign n47064 = n2905 & ~n4812 ;
  assign n47065 = ~n6945 & n47064 ;
  assign n47066 = n47065 ^ n10023 ^ 1'b0 ;
  assign n47067 = n24101 & ~n47066 ;
  assign n47068 = n47067 ^ n21381 ^ 1'b0 ;
  assign n47069 = n3376 & ~n47068 ;
  assign n47070 = ( n8382 & n17566 ) | ( n8382 & n29057 ) | ( n17566 & n29057 ) ;
  assign n47071 = ( n1792 & ~n37360 ) | ( n1792 & n47070 ) | ( ~n37360 & n47070 ) ;
  assign n47072 = n47071 ^ n43604 ^ n1639 ;
  assign n47073 = n31857 ^ n21476 ^ n9641 ;
  assign n47074 = n47073 ^ n37107 ^ n33286 ;
  assign n47075 = n15720 ^ n10444 ^ n6485 ;
  assign n47076 = n900 | n2052 ;
  assign n47077 = ( n26429 & n44970 ) | ( n26429 & ~n47076 ) | ( n44970 & ~n47076 ) ;
  assign n47078 = n16327 ^ n14196 ^ 1'b0 ;
  assign n47079 = n33736 & ~n42426 ;
  assign n47080 = ( ~n8819 & n29200 ) | ( ~n8819 & n47079 ) | ( n29200 & n47079 ) ;
  assign n47081 = n14673 ^ n1188 ^ 1'b0 ;
  assign n47082 = ( n19211 & n24805 ) | ( n19211 & n26092 ) | ( n24805 & n26092 ) ;
  assign n47083 = n47082 ^ n8068 ^ n3007 ;
  assign n47084 = n11749 ^ n8835 ^ n8780 ;
  assign n47085 = n47084 ^ x74 ^ 1'b0 ;
  assign n47086 = ~n47083 & n47085 ;
  assign n47087 = ~n13605 & n24551 ;
  assign n47088 = n31913 & n47087 ;
  assign n47089 = n18446 | n33027 ;
  assign n47090 = n47089 ^ n36487 ^ 1'b0 ;
  assign n47092 = ( ~x53 & n9798 ) | ( ~x53 & n36169 ) | ( n9798 & n36169 ) ;
  assign n47091 = ( n5471 & n17081 ) | ( n5471 & n17443 ) | ( n17081 & n17443 ) ;
  assign n47093 = n47092 ^ n47091 ^ n41515 ;
  assign n47094 = n34676 ^ n29070 ^ n2024 ;
  assign n47095 = n47094 ^ n45347 ^ 1'b0 ;
  assign n47096 = n12610 ^ n12369 ^ n1989 ;
  assign n47097 = ( ~n6249 & n20153 ) | ( ~n6249 & n47096 ) | ( n20153 & n47096 ) ;
  assign n47098 = n47097 ^ n28910 ^ n28422 ;
  assign n47099 = ( n8668 & ~n47095 ) | ( n8668 & n47098 ) | ( ~n47095 & n47098 ) ;
  assign n47100 = n47099 ^ n9239 ^ 1'b0 ;
  assign n47104 = ( n12235 & ~n26000 ) | ( n12235 & n28150 ) | ( ~n26000 & n28150 ) ;
  assign n47103 = ( n4576 & n6048 ) | ( n4576 & ~n16147 ) | ( n6048 & ~n16147 ) ;
  assign n47101 = ( n2633 & n3445 ) | ( n2633 & n4651 ) | ( n3445 & n4651 ) ;
  assign n47102 = ( n4227 & ~n41333 ) | ( n4227 & n47101 ) | ( ~n41333 & n47101 ) ;
  assign n47105 = n47104 ^ n47103 ^ n47102 ;
  assign n47106 = ( n1292 & ~n10067 ) | ( n1292 & n14041 ) | ( ~n10067 & n14041 ) ;
  assign n47107 = ( ~n20845 & n24497 ) | ( ~n20845 & n27229 ) | ( n24497 & n27229 ) ;
  assign n47108 = ( n18715 & n39487 ) | ( n18715 & n47107 ) | ( n39487 & n47107 ) ;
  assign n47109 = ( n12218 & n47106 ) | ( n12218 & ~n47108 ) | ( n47106 & ~n47108 ) ;
  assign n47110 = n22392 & n35436 ;
  assign n47111 = n40858 ^ n34604 ^ 1'b0 ;
  assign n47112 = ( n46424 & n47110 ) | ( n46424 & n47111 ) | ( n47110 & n47111 ) ;
  assign n47113 = n12836 | n36370 ;
  assign n47114 = n47113 ^ n42526 ^ 1'b0 ;
  assign n47115 = n47114 ^ n21442 ^ n3519 ;
  assign n47116 = ~n12807 & n47115 ;
  assign n47117 = n11574 & n47116 ;
  assign n47118 = n10706 ^ n3679 ^ 1'b0 ;
  assign n47119 = n45932 & ~n47118 ;
  assign n47120 = n47119 ^ n39853 ^ n15934 ;
  assign n47121 = ( n4677 & ~n16338 ) | ( n4677 & n19574 ) | ( ~n16338 & n19574 ) ;
  assign n47122 = n47121 ^ n39234 ^ n15376 ;
  assign n47124 = n7185 ^ n5916 ^ x128 ;
  assign n47125 = n47124 ^ n16454 ^ n16271 ;
  assign n47123 = ( n5954 & n16210 ) | ( n5954 & n34115 ) | ( n16210 & n34115 ) ;
  assign n47126 = n47125 ^ n47123 ^ 1'b0 ;
  assign n47127 = ~n47122 & n47126 ;
  assign n47128 = ~n40127 & n47127 ;
  assign n47129 = ~n47120 & n47128 ;
  assign n47130 = ( ~n2199 & n9808 ) | ( ~n2199 & n13192 ) | ( n9808 & n13192 ) ;
  assign n47131 = n47130 ^ n40732 ^ n23221 ;
  assign n47132 = n47131 ^ n14307 ^ 1'b0 ;
  assign n47133 = n28189 & n47132 ;
  assign n47134 = n32167 & n47133 ;
  assign n47135 = ~n35250 & n47134 ;
  assign n47136 = n30366 ^ n10840 ^ n9081 ;
  assign n47138 = ( n2111 & ~n10121 ) | ( n2111 & n23166 ) | ( ~n10121 & n23166 ) ;
  assign n47137 = n7406 ^ n6634 ^ n4827 ;
  assign n47139 = n47138 ^ n47137 ^ n40836 ;
  assign n47144 = n5448 & n28923 ;
  assign n47145 = ~n32169 & n47144 ;
  assign n47146 = ~n19694 & n47145 ;
  assign n47140 = n24419 ^ n21259 ^ n9226 ;
  assign n47141 = n40808 & ~n47140 ;
  assign n47142 = n24788 & n47141 ;
  assign n47143 = n47142 ^ n22472 ^ n20905 ;
  assign n47147 = n47146 ^ n47143 ^ n2938 ;
  assign n47148 = n623 & ~n7988 ;
  assign n47149 = ~n35211 & n47148 ;
  assign n47150 = ~n38214 & n39094 ;
  assign n47151 = n14632 & ~n42620 ;
  assign n47152 = n47150 & n47151 ;
  assign n47153 = n16366 ^ n5528 ^ 1'b0 ;
  assign n47154 = n5812 & n47153 ;
  assign n47155 = ( n22187 & ~n25877 ) | ( n22187 & n47154 ) | ( ~n25877 & n47154 ) ;
  assign n47156 = n7756 ^ n2783 ^ 1'b0 ;
  assign n47157 = n47155 & n47156 ;
  assign n47158 = ( n10229 & ~n22879 ) | ( n10229 & n35112 ) | ( ~n22879 & n35112 ) ;
  assign n47159 = n47158 ^ n46085 ^ n18516 ;
  assign n47160 = n47159 ^ n31038 ^ n25772 ;
  assign n47161 = ( ~n3875 & n20434 ) | ( ~n3875 & n35876 ) | ( n20434 & n35876 ) ;
  assign n47162 = n36208 ^ n33010 ^ 1'b0 ;
  assign n47163 = n28433 & n47162 ;
  assign n47164 = n44366 ^ n27237 ^ n20793 ;
  assign n47165 = n47164 ^ n1837 ^ 1'b0 ;
  assign n47166 = n21585 ^ n8180 ^ n666 ;
  assign n47167 = ( n16466 & n46867 ) | ( n16466 & n47166 ) | ( n46867 & n47166 ) ;
  assign n47168 = ( n25049 & ~n47165 ) | ( n25049 & n47167 ) | ( ~n47165 & n47167 ) ;
  assign n47169 = n2097 & n47168 ;
  assign n47170 = ~n47163 & n47169 ;
  assign n47171 = n38206 ^ n25908 ^ n20484 ;
  assign n47172 = n47171 ^ n40149 ^ n19960 ;
  assign n47173 = ( x187 & n47170 ) | ( x187 & ~n47172 ) | ( n47170 & ~n47172 ) ;
  assign n47174 = n39716 ^ n14170 ^ 1'b0 ;
  assign n47175 = ( n16082 & n18356 ) | ( n16082 & ~n47174 ) | ( n18356 & ~n47174 ) ;
  assign n47176 = ~n18650 & n43050 ;
  assign n47177 = n47176 ^ n27720 ^ 1'b0 ;
  assign n47180 = ( ~n9609 & n11782 ) | ( ~n9609 & n16534 ) | ( n11782 & n16534 ) ;
  assign n47178 = n30007 | n31531 ;
  assign n47179 = n47178 ^ n2447 ^ 1'b0 ;
  assign n47181 = n47180 ^ n47179 ^ n24089 ;
  assign n47182 = n30162 ^ n26758 ^ 1'b0 ;
  assign n47183 = n32667 & ~n47030 ;
  assign n47184 = n32888 & n47183 ;
  assign n47185 = n30324 ^ n16230 ^ n12649 ;
  assign n47186 = n27939 | n46231 ;
  assign n47187 = n47185 & ~n47186 ;
  assign n47188 = n31017 ^ n29311 ^ 1'b0 ;
  assign n47189 = n23356 & ~n47188 ;
  assign n47190 = n15248 ^ n9493 ^ n3336 ;
  assign n47191 = n35544 ^ n6869 ^ 1'b0 ;
  assign n47192 = ( n7599 & n8819 ) | ( n7599 & n21362 ) | ( n8819 & n21362 ) ;
  assign n47193 = ~n40344 & n47192 ;
  assign n47194 = ~n3294 & n47193 ;
  assign n47195 = ( n3463 & n5696 ) | ( n3463 & ~n47194 ) | ( n5696 & ~n47194 ) ;
  assign n47196 = ( n21819 & n33637 ) | ( n21819 & ~n47195 ) | ( n33637 & ~n47195 ) ;
  assign n47197 = ( n15701 & n31112 ) | ( n15701 & n47196 ) | ( n31112 & n47196 ) ;
  assign n47198 = n26749 ^ n3204 ^ 1'b0 ;
  assign n47199 = n28036 ^ n18915 ^ n8326 ;
  assign n47200 = n26087 ^ n11167 ^ n9038 ;
  assign n47201 = n47200 ^ n15535 ^ n6696 ;
  assign n47202 = ( n13000 & n25101 ) | ( n13000 & ~n40350 ) | ( n25101 & ~n40350 ) ;
  assign n47203 = ( n699 & n3431 ) | ( n699 & n47202 ) | ( n3431 & n47202 ) ;
  assign n47204 = n25657 ^ n269 ^ 1'b0 ;
  assign n47205 = n33672 & n47204 ;
  assign n47206 = ~n814 & n9129 ;
  assign n47207 = n41345 & n47206 ;
  assign n47208 = n13013 & n42683 ;
  assign n47209 = n43988 & n47208 ;
  assign n47210 = n47209 ^ n32797 ^ n11949 ;
  assign n47211 = n25970 ^ n11260 ^ n1780 ;
  assign n47212 = n8442 & ~n47211 ;
  assign n47213 = n28203 ^ n17900 ^ n16644 ;
  assign n47214 = ( n3213 & n27837 ) | ( n3213 & n44915 ) | ( n27837 & n44915 ) ;
  assign n47215 = ( n19952 & n47213 ) | ( n19952 & n47214 ) | ( n47213 & n47214 ) ;
  assign n47216 = n21213 ^ n20965 ^ 1'b0 ;
  assign n47218 = n33698 ^ n6447 ^ 1'b0 ;
  assign n47217 = n17781 ^ n16778 ^ n12800 ;
  assign n47219 = n47218 ^ n47217 ^ 1'b0 ;
  assign n47220 = n47219 ^ n45027 ^ n28885 ;
  assign n47221 = n14821 | n26826 ;
  assign n47222 = n11564 | n47221 ;
  assign n47223 = n34951 ^ n31692 ^ n16336 ;
  assign n47224 = ~n15935 & n21477 ;
  assign n47225 = ( ~n8007 & n29099 ) | ( ~n8007 & n47224 ) | ( n29099 & n47224 ) ;
  assign n47226 = n47225 ^ n23925 ^ n19020 ;
  assign n47227 = ( n5034 & ~n8020 ) | ( n5034 & n47226 ) | ( ~n8020 & n47226 ) ;
  assign n47228 = n354 & ~n47227 ;
  assign n47229 = ~n47223 & n47228 ;
  assign n47230 = n27710 ^ n8976 ^ 1'b0 ;
  assign n47231 = ~n44686 & n47230 ;
  assign n47232 = ( n4732 & n43051 ) | ( n4732 & n47231 ) | ( n43051 & n47231 ) ;
  assign n47237 = n21905 ^ n17541 ^ n5665 ;
  assign n47233 = n19127 ^ n1028 ^ 1'b0 ;
  assign n47234 = ( ~n3898 & n4277 ) | ( ~n3898 & n6886 ) | ( n4277 & n6886 ) ;
  assign n47235 = n30950 & n47234 ;
  assign n47236 = ~n47233 & n47235 ;
  assign n47238 = n47237 ^ n47236 ^ n41154 ;
  assign n47239 = ( ~n5616 & n9681 ) | ( ~n5616 & n28844 ) | ( n9681 & n28844 ) ;
  assign n47240 = n47239 ^ n10614 ^ n5566 ;
  assign n47241 = ( ~n34074 & n34186 ) | ( ~n34074 & n36553 ) | ( n34186 & n36553 ) ;
  assign n47242 = ( ~n45013 & n47240 ) | ( ~n45013 & n47241 ) | ( n47240 & n47241 ) ;
  assign n47243 = n19348 ^ n11576 ^ n9796 ;
  assign n47251 = ~n13356 & n29254 ;
  assign n47245 = n10844 ^ n7209 ^ n1673 ;
  assign n47246 = ( ~n16455 & n19921 ) | ( ~n16455 & n33724 ) | ( n19921 & n33724 ) ;
  assign n47247 = ( ~n13755 & n18958 ) | ( ~n13755 & n47246 ) | ( n18958 & n47246 ) ;
  assign n47248 = ~n3027 & n8573 ;
  assign n47249 = n20768 & n47248 ;
  assign n47250 = ( n47245 & n47247 ) | ( n47245 & n47249 ) | ( n47247 & n47249 ) ;
  assign n47244 = ( n305 & n20687 ) | ( n305 & n44560 ) | ( n20687 & n44560 ) ;
  assign n47252 = n47251 ^ n47250 ^ n47244 ;
  assign n47253 = n38199 ^ n5941 ^ n4686 ;
  assign n47254 = n39192 ^ n28541 ^ n11602 ;
  assign n47255 = n44090 ^ n18422 ^ 1'b0 ;
  assign n47256 = n39273 & ~n47255 ;
  assign n47257 = n5839 ^ n1382 ^ 1'b0 ;
  assign n47258 = n43844 & ~n47257 ;
  assign n47259 = ~n1063 & n29504 ;
  assign n47260 = n47259 ^ n9328 ^ 1'b0 ;
  assign n47261 = n18161 ^ n10478 ^ n6030 ;
  assign n47262 = n47261 ^ n44463 ^ n12897 ;
  assign n47263 = n29790 ^ x227 ^ 1'b0 ;
  assign n47264 = ( ~n20232 & n27751 ) | ( ~n20232 & n34934 ) | ( n27751 & n34934 ) ;
  assign n47265 = n46181 ^ n22711 ^ n8052 ;
  assign n47266 = ( ~n15803 & n24271 ) | ( ~n15803 & n44455 ) | ( n24271 & n44455 ) ;
  assign n47267 = n44532 ^ n9958 ^ n7922 ;
  assign n47268 = ( n7395 & n14506 ) | ( n7395 & n38361 ) | ( n14506 & n38361 ) ;
  assign n47269 = n43295 ^ n40234 ^ n7185 ;
  assign n47270 = ( n9482 & ~n19609 ) | ( n9482 & n27645 ) | ( ~n19609 & n27645 ) ;
  assign n47271 = ~n47269 & n47270 ;
  assign n47272 = ~n5791 & n5846 ;
  assign n47273 = ( ~n1013 & n6431 ) | ( ~n1013 & n14092 ) | ( n6431 & n14092 ) ;
  assign n47274 = ~n34435 & n47273 ;
  assign n47275 = ~n47272 & n47274 ;
  assign n47278 = ( ~n2703 & n7149 ) | ( ~n2703 & n21479 ) | ( n7149 & n21479 ) ;
  assign n47277 = ( n15567 & n29278 ) | ( n15567 & ~n33076 ) | ( n29278 & ~n33076 ) ;
  assign n47276 = n16450 ^ n9217 ^ n5101 ;
  assign n47279 = n47278 ^ n47277 ^ n47276 ;
  assign n47280 = ( n9969 & n33724 ) | ( n9969 & ~n39094 ) | ( n33724 & ~n39094 ) ;
  assign n47281 = n11681 & ~n26043 ;
  assign n47282 = n47281 ^ n16863 ^ 1'b0 ;
  assign n47283 = ( ~n680 & n19177 ) | ( ~n680 & n47282 ) | ( n19177 & n47282 ) ;
  assign n47284 = n42077 ^ n32840 ^ n2283 ;
  assign n47285 = n47284 ^ n44988 ^ n24397 ;
  assign n47286 = ( n31719 & ~n34010 ) | ( n31719 & n47285 ) | ( ~n34010 & n47285 ) ;
  assign n47287 = n19546 & ~n24884 ;
  assign n47288 = n11630 & ~n43710 ;
  assign n47289 = ~n41685 & n47288 ;
  assign n47290 = n36548 ^ n28392 ^ n10749 ;
  assign n47291 = n34417 ^ n20986 ^ 1'b0 ;
  assign n47292 = n38253 ^ n28585 ^ n3384 ;
  assign n47293 = n47292 ^ n35523 ^ 1'b0 ;
  assign n47294 = n47293 ^ n15827 ^ 1'b0 ;
  assign n47295 = n39144 ^ n28764 ^ n1460 ;
  assign n47296 = ( n21960 & n31047 ) | ( n21960 & n47295 ) | ( n31047 & n47295 ) ;
  assign n47297 = ( ~x232 & n730 ) | ( ~x232 & n25755 ) | ( n730 & n25755 ) ;
  assign n47298 = n47297 ^ n38669 ^ n6393 ;
  assign n47299 = n8367 ^ n1445 ^ 1'b0 ;
  assign n47300 = n47299 ^ n30316 ^ n28534 ;
  assign n47301 = ( ~n4042 & n29489 ) | ( ~n4042 & n44127 ) | ( n29489 & n44127 ) ;
  assign n47302 = ( n12432 & n31096 ) | ( n12432 & n31977 ) | ( n31096 & n31977 ) ;
  assign n47306 = n15772 ^ n5057 ^ n1723 ;
  assign n47307 = ( ~n18148 & n39170 ) | ( ~n18148 & n47306 ) | ( n39170 & n47306 ) ;
  assign n47303 = n21030 ^ n14908 ^ n9006 ;
  assign n47304 = n42152 ^ n9261 ^ 1'b0 ;
  assign n47305 = ~n47303 & n47304 ;
  assign n47308 = n47307 ^ n47305 ^ n30350 ;
  assign n47309 = n27444 ^ n19020 ^ n4716 ;
  assign n47310 = n47309 ^ n5296 ^ n4306 ;
  assign n47311 = n31773 ^ n13376 ^ n7832 ;
  assign n47312 = ( n1229 & ~n5600 ) | ( n1229 & n27046 ) | ( ~n5600 & n27046 ) ;
  assign n47313 = n47312 ^ n18065 ^ n11111 ;
  assign n47314 = ( n44578 & n47311 ) | ( n44578 & ~n47313 ) | ( n47311 & ~n47313 ) ;
  assign n47315 = n47314 ^ n42160 ^ n10040 ;
  assign n47319 = n35938 ^ n30478 ^ n18256 ;
  assign n47317 = n11619 ^ n854 ^ x225 ;
  assign n47318 = n9058 & ~n47317 ;
  assign n47320 = n47319 ^ n47318 ^ n7638 ;
  assign n47316 = ( n8142 & n32337 ) | ( n8142 & n35390 ) | ( n32337 & n35390 ) ;
  assign n47321 = n47320 ^ n47316 ^ n3097 ;
  assign n47322 = n19710 & ~n28343 ;
  assign n47323 = ( ~n2780 & n15602 ) | ( ~n2780 & n47322 ) | ( n15602 & n47322 ) ;
  assign n47324 = ( n2699 & n4217 ) | ( n2699 & ~n47323 ) | ( n4217 & ~n47323 ) ;
  assign n47325 = ( n29763 & n43674 ) | ( n29763 & n47324 ) | ( n43674 & n47324 ) ;
  assign n47326 = n27590 ^ n11494 ^ n4781 ;
  assign n47327 = n47326 ^ n27339 ^ 1'b0 ;
  assign n47328 = n14900 & n47327 ;
  assign n47329 = n47328 ^ n18389 ^ 1'b0 ;
  assign n47330 = n2362 & n19746 ;
  assign n47331 = n10228 & ~n30731 ;
  assign n47332 = n47331 ^ n3085 ^ 1'b0 ;
  assign n47333 = ~n47330 & n47332 ;
  assign n47334 = ( n11409 & n30093 ) | ( n11409 & ~n46051 ) | ( n30093 & ~n46051 ) ;
  assign n47335 = n3209 & ~n12392 ;
  assign n47336 = n26520 | n47335 ;
  assign n47337 = n47334 & ~n47336 ;
  assign n47338 = ( n8027 & ~n20940 ) | ( n8027 & n45911 ) | ( ~n20940 & n45911 ) ;
  assign n47339 = n45575 ^ n32311 ^ n947 ;
  assign n47341 = n21005 & ~n31887 ;
  assign n47340 = n29919 ^ n19887 ^ n2744 ;
  assign n47342 = n47341 ^ n47340 ^ n36952 ;
  assign n47343 = n33464 ^ n22917 ^ n4399 ;
  assign n47344 = n33384 ^ n11079 ^ 1'b0 ;
  assign n47345 = ( n2374 & n33896 ) | ( n2374 & ~n47344 ) | ( n33896 & ~n47344 ) ;
  assign n47346 = n32609 ^ n26979 ^ n10062 ;
  assign n47347 = n9975 ^ n9240 ^ n5670 ;
  assign n47348 = n46221 | n47347 ;
  assign n47349 = n44070 ^ n3086 ^ n2764 ;
  assign n47350 = n16105 ^ n4466 ^ 1'b0 ;
  assign n47351 = n11260 & n47350 ;
  assign n47353 = n15379 ^ x132 ^ 1'b0 ;
  assign n47354 = n47353 ^ n9884 ^ n5267 ;
  assign n47352 = n4035 | n7592 ;
  assign n47355 = n47354 ^ n47352 ^ 1'b0 ;
  assign n47356 = n40971 ^ n5859 ^ n3985 ;
  assign n47357 = ( ~n19531 & n29122 ) | ( ~n19531 & n47356 ) | ( n29122 & n47356 ) ;
  assign n47358 = ~n28637 & n47357 ;
  assign n47359 = ( n4166 & n9144 ) | ( n4166 & ~n41987 ) | ( n9144 & ~n41987 ) ;
  assign n47360 = ( n5731 & n8865 ) | ( n5731 & ~n47359 ) | ( n8865 & ~n47359 ) ;
  assign n47361 = n22033 ^ n8933 ^ n1569 ;
  assign n47362 = n1794 & ~n29313 ;
  assign n47363 = n47362 ^ n47138 ^ n23578 ;
  assign n47364 = n8942 & n47363 ;
  assign n47365 = x176 & n20299 ;
  assign n47366 = ~n14150 & n47365 ;
  assign n47367 = ( ~n1724 & n3678 ) | ( ~n1724 & n37854 ) | ( n3678 & n37854 ) ;
  assign n47368 = ( n13894 & n20841 ) | ( n13894 & n26223 ) | ( n20841 & n26223 ) ;
  assign n47369 = n47368 ^ n11281 ^ n5240 ;
  assign n47370 = n47369 ^ n5988 ^ n5869 ;
  assign n47371 = n10895 & ~n47370 ;
  assign n47372 = ~n20445 & n47031 ;
  assign n47373 = n19185 ^ n15163 ^ n10567 ;
  assign n47374 = n47373 ^ n15867 ^ 1'b0 ;
  assign n47375 = n46383 | n47374 ;
  assign n47376 = ( n10514 & n24139 ) | ( n10514 & ~n47375 ) | ( n24139 & ~n47375 ) ;
  assign n47377 = n42391 ^ n17316 ^ n3302 ;
  assign n47378 = n47377 ^ n27551 ^ n1709 ;
  assign n47379 = ( n23190 & ~n28902 ) | ( n23190 & n30791 ) | ( ~n28902 & n30791 ) ;
  assign n47380 = ( ~n26118 & n26308 ) | ( ~n26118 & n31685 ) | ( n26308 & n31685 ) ;
  assign n47381 = ( x106 & ~n13147 ) | ( x106 & n17784 ) | ( ~n13147 & n17784 ) ;
  assign n47382 = n3194 & n47381 ;
  assign n47383 = ~n8967 & n47382 ;
  assign n47384 = ( n8573 & n22911 ) | ( n8573 & ~n33911 ) | ( n22911 & ~n33911 ) ;
  assign n47385 = n23265 ^ n21732 ^ n13701 ;
  assign n47386 = n45957 & ~n47385 ;
  assign n47387 = n47384 & n47386 ;
  assign n47388 = ( n23246 & n33001 ) | ( n23246 & n39473 ) | ( n33001 & n39473 ) ;
  assign n47389 = ( n8299 & ~n14461 ) | ( n8299 & n22609 ) | ( ~n14461 & n22609 ) ;
  assign n47390 = ( n4471 & ~n5878 ) | ( n4471 & n47389 ) | ( ~n5878 & n47389 ) ;
  assign n47391 = ( n20887 & ~n24661 ) | ( n20887 & n47390 ) | ( ~n24661 & n47390 ) ;
  assign n47392 = n38738 ^ n7522 ^ 1'b0 ;
  assign n47393 = n18982 ^ n14532 ^ 1'b0 ;
  assign n47394 = ( n4382 & ~n4963 ) | ( n4382 & n47393 ) | ( ~n4963 & n47393 ) ;
  assign n47395 = n17681 & ~n47394 ;
  assign n47396 = n7511 & n21282 ;
  assign n47397 = n2110 & n47396 ;
  assign n47398 = n24602 ^ n14748 ^ n9318 ;
  assign n47399 = ( n463 & ~n1996 ) | ( n463 & n47398 ) | ( ~n1996 & n47398 ) ;
  assign n47400 = ( n6218 & n6484 ) | ( n6218 & ~n41384 ) | ( n6484 & ~n41384 ) ;
  assign n47401 = n3577 | n34222 ;
  assign n47402 = ( n1145 & n9881 ) | ( n1145 & ~n20420 ) | ( n9881 & ~n20420 ) ;
  assign n47403 = ( n13528 & n18784 ) | ( n13528 & n46643 ) | ( n18784 & n46643 ) ;
  assign n47404 = n31482 ^ n21438 ^ n9156 ;
  assign n47405 = ( n7732 & n47403 ) | ( n7732 & ~n47404 ) | ( n47403 & ~n47404 ) ;
  assign n47406 = n1032 & ~n16444 ;
  assign n47407 = ( ~n10496 & n15848 ) | ( ~n10496 & n18103 ) | ( n15848 & n18103 ) ;
  assign n47408 = ( n3275 & ~n38224 ) | ( n3275 & n47407 ) | ( ~n38224 & n47407 ) ;
  assign n47409 = ( ~n686 & n1021 ) | ( ~n686 & n27031 ) | ( n1021 & n27031 ) ;
  assign n47410 = ( n2225 & n20976 ) | ( n2225 & n31120 ) | ( n20976 & n31120 ) ;
  assign n47411 = ( n28990 & n47409 ) | ( n28990 & n47410 ) | ( n47409 & n47410 ) ;
  assign n47412 = n8702 ^ n1329 ^ 1'b0 ;
  assign n47413 = ( ~n12932 & n41456 ) | ( ~n12932 & n47412 ) | ( n41456 & n47412 ) ;
  assign n47419 = n3223 & ~n4318 ;
  assign n47420 = n19215 & n47419 ;
  assign n47414 = n24011 | n30012 ;
  assign n47415 = n37267 | n47414 ;
  assign n47416 = n1983 & n4544 ;
  assign n47417 = n47416 ^ n20232 ^ 1'b0 ;
  assign n47418 = ( n39285 & n47415 ) | ( n39285 & n47417 ) | ( n47415 & n47417 ) ;
  assign n47421 = n47420 ^ n47418 ^ n4694 ;
  assign n47425 = n5088 & n9601 ;
  assign n47422 = n16001 | n19869 ;
  assign n47423 = n47422 ^ n24016 ^ 1'b0 ;
  assign n47424 = ~n8246 & n47423 ;
  assign n47426 = n47425 ^ n47424 ^ 1'b0 ;
  assign n47427 = n44106 ^ n12069 ^ 1'b0 ;
  assign n47428 = ~n12665 & n19592 ;
  assign n47429 = n40311 ^ n6055 ^ n5247 ;
  assign n47430 = n8826 & ~n47429 ;
  assign n47431 = n15443 ^ n11889 ^ 1'b0 ;
  assign n47432 = n47431 ^ n14573 ^ n14308 ;
  assign n47433 = n47432 ^ n30378 ^ n8204 ;
  assign n47434 = n47433 ^ n13490 ^ n2880 ;
  assign n47441 = n11352 ^ n11034 ^ n2996 ;
  assign n47442 = n1148 & ~n47441 ;
  assign n47443 = ~n16513 & n47442 ;
  assign n47439 = n23435 ^ n13992 ^ n8810 ;
  assign n47435 = n2219 & n25242 ;
  assign n47436 = ~n38624 & n47435 ;
  assign n47437 = n36889 ^ n22590 ^ n10171 ;
  assign n47438 = ( n41641 & ~n47436 ) | ( n41641 & n47437 ) | ( ~n47436 & n47437 ) ;
  assign n47440 = n47439 ^ n47438 ^ n43259 ;
  assign n47444 = n47443 ^ n47440 ^ n5899 ;
  assign n47445 = n37782 ^ n19815 ^ n11433 ;
  assign n47446 = ( x102 & ~n15558 ) | ( x102 & n47445 ) | ( ~n15558 & n47445 ) ;
  assign n47447 = ( n12547 & n17993 ) | ( n12547 & ~n47446 ) | ( n17993 & ~n47446 ) ;
  assign n47448 = ( ~n10908 & n35704 ) | ( ~n10908 & n37811 ) | ( n35704 & n37811 ) ;
  assign n47450 = ~n6562 & n9832 ;
  assign n47451 = n47450 ^ n5754 ^ 1'b0 ;
  assign n47449 = n5514 & n13313 ;
  assign n47452 = n47451 ^ n47449 ^ n39261 ;
  assign n47453 = n1757 | n7096 ;
  assign n47454 = n39418 | n47453 ;
  assign n47455 = n13792 ^ n582 ^ 1'b0 ;
  assign n47456 = n14145 | n47455 ;
  assign n47457 = n47456 ^ n19305 ^ n4043 ;
  assign n47458 = n47457 ^ n2401 ^ 1'b0 ;
  assign n47459 = n7230 ^ n747 ^ 1'b0 ;
  assign n47460 = n15894 ^ n1481 ^ 1'b0 ;
  assign n47461 = n17456 & n47460 ;
  assign n47462 = n7513 | n22176 ;
  assign n47463 = n5379 & ~n47462 ;
  assign n47464 = ( ~n13826 & n13898 ) | ( ~n13826 & n47463 ) | ( n13898 & n47463 ) ;
  assign n47465 = ( n8958 & n47461 ) | ( n8958 & n47464 ) | ( n47461 & n47464 ) ;
  assign n47466 = ( n36169 & n47459 ) | ( n36169 & n47465 ) | ( n47459 & n47465 ) ;
  assign n47467 = ( n4039 & n6854 ) | ( n4039 & n7607 ) | ( n6854 & n7607 ) ;
  assign n47468 = n47467 ^ n23843 ^ n10000 ;
  assign n47469 = ( n32660 & ~n44173 ) | ( n32660 & n47468 ) | ( ~n44173 & n47468 ) ;
  assign n47470 = n31340 ^ n27204 ^ 1'b0 ;
  assign n47471 = n33303 ^ n4515 ^ 1'b0 ;
  assign n47472 = n47471 ^ n7082 ^ n6213 ;
  assign n47473 = ( ~n5326 & n46169 ) | ( ~n5326 & n47472 ) | ( n46169 & n47472 ) ;
  assign n47474 = n44984 ^ n15353 ^ n15133 ;
  assign n47475 = ( n4094 & ~n8569 ) | ( n4094 & n47474 ) | ( ~n8569 & n47474 ) ;
  assign n47476 = n32842 ^ n11966 ^ n3069 ;
  assign n47477 = ~n24008 & n38214 ;
  assign n47478 = ( n3855 & ~n47476 ) | ( n3855 & n47477 ) | ( ~n47476 & n47477 ) ;
  assign n47479 = ( ~n22750 & n31554 ) | ( ~n22750 & n47478 ) | ( n31554 & n47478 ) ;
  assign n47480 = ( ~n13037 & n28307 ) | ( ~n13037 & n43116 ) | ( n28307 & n43116 ) ;
  assign n47481 = n31248 ^ n25330 ^ n4562 ;
  assign n47482 = n45450 ^ n8233 ^ n3361 ;
  assign n47483 = n47482 ^ n19511 ^ 1'b0 ;
  assign n47484 = n39111 ^ n27697 ^ x51 ;
  assign n47485 = ( ~n7515 & n27778 ) | ( ~n7515 & n47484 ) | ( n27778 & n47484 ) ;
  assign n47486 = ( n11012 & n11111 ) | ( n11012 & n41140 ) | ( n11111 & n41140 ) ;
  assign n47487 = ~n45841 & n47486 ;
  assign n47488 = n33884 & n47487 ;
  assign n47489 = n34369 ^ n32273 ^ n24694 ;
  assign n47490 = n25759 ^ n6929 ^ 1'b0 ;
  assign n47491 = ( n32914 & n33576 ) | ( n32914 & ~n37588 ) | ( n33576 & ~n37588 ) ;
  assign n47492 = ( n8191 & ~n12643 ) | ( n8191 & n47129 ) | ( ~n12643 & n47129 ) ;
  assign n47493 = n6861 ^ n4676 ^ 1'b0 ;
  assign n47494 = ( n2443 & n16953 ) | ( n2443 & ~n30794 ) | ( n16953 & ~n30794 ) ;
  assign n47495 = n45383 ^ n26752 ^ n5902 ;
  assign n47496 = ( ~n12368 & n47494 ) | ( ~n12368 & n47495 ) | ( n47494 & n47495 ) ;
  assign n47497 = n9210 & n18041 ;
  assign n47498 = ~n6355 & n16034 ;
  assign n47499 = ~n47497 & n47498 ;
  assign n47500 = n36101 | n47499 ;
  assign n47501 = n46048 | n47500 ;
  assign n47503 = n16789 | n26998 ;
  assign n47504 = n11582 | n47503 ;
  assign n47502 = n11388 & ~n33130 ;
  assign n47505 = n47504 ^ n47502 ^ 1'b0 ;
  assign n47506 = ( ~n6435 & n26651 ) | ( ~n6435 & n31723 ) | ( n26651 & n31723 ) ;
  assign n47507 = ( x68 & n2107 ) | ( x68 & ~n26795 ) | ( n2107 & ~n26795 ) ;
  assign n47508 = n23779 ^ n9530 ^ n7474 ;
  assign n47509 = n29294 ^ n19455 ^ n3284 ;
  assign n47510 = n8709 & ~n30919 ;
  assign n47511 = n41995 ^ n30322 ^ n13305 ;
  assign n47512 = n45763 ^ n19431 ^ 1'b0 ;
  assign n47513 = n7990 & ~n47512 ;
  assign n47514 = n47513 ^ n13081 ^ 1'b0 ;
  assign n47515 = ( n23207 & n34258 ) | ( n23207 & ~n47514 ) | ( n34258 & ~n47514 ) ;
  assign n47516 = ~n4120 & n15759 ;
  assign n47517 = n42431 ^ n7478 ^ 1'b0 ;
  assign n47518 = n47516 & ~n47517 ;
  assign n47519 = ~n14684 & n37386 ;
  assign n47520 = n47519 ^ n24435 ^ 1'b0 ;
  assign n47532 = ( n7275 & ~n12419 ) | ( n7275 & n15518 ) | ( ~n12419 & n15518 ) ;
  assign n47533 = n47532 ^ n2598 ^ 1'b0 ;
  assign n47530 = ( n18000 & n36237 ) | ( n18000 & n42221 ) | ( n36237 & n42221 ) ;
  assign n47531 = ( n3887 & n34304 ) | ( n3887 & n47530 ) | ( n34304 & n47530 ) ;
  assign n47522 = ~n4738 & n33668 ;
  assign n47523 = ~n6119 & n47522 ;
  assign n47521 = ( n1560 & n2426 ) | ( n1560 & ~n43018 ) | ( n2426 & ~n43018 ) ;
  assign n47524 = n47523 ^ n47521 ^ n4874 ;
  assign n47525 = ~n8256 & n12721 ;
  assign n47526 = n31344 ^ n8070 ^ 1'b0 ;
  assign n47527 = ( n47524 & n47525 ) | ( n47524 & n47526 ) | ( n47525 & n47526 ) ;
  assign n47528 = n12518 & ~n47527 ;
  assign n47529 = ~n23071 & n47528 ;
  assign n47534 = n47533 ^ n47531 ^ n47529 ;
  assign n47535 = ( n7515 & ~n24430 ) | ( n7515 & n35969 ) | ( ~n24430 & n35969 ) ;
  assign n47536 = ( n15034 & n23967 ) | ( n15034 & n37814 ) | ( n23967 & n37814 ) ;
  assign n47537 = ( ~n17701 & n20390 ) | ( ~n17701 & n38789 ) | ( n20390 & n38789 ) ;
  assign n47538 = ( n43927 & n47536 ) | ( n43927 & ~n47537 ) | ( n47536 & ~n47537 ) ;
  assign n47541 = ( ~n1262 & n1862 ) | ( ~n1262 & n25336 ) | ( n1862 & n25336 ) ;
  assign n47539 = n10245 & n18720 ;
  assign n47540 = ~n20491 & n47539 ;
  assign n47542 = n47541 ^ n47540 ^ n12204 ;
  assign n47543 = n37427 ^ n34319 ^ 1'b0 ;
  assign n47544 = ~n2215 & n47543 ;
  assign n47545 = n18592 ^ n15541 ^ 1'b0 ;
  assign n47546 = ( n6464 & n10485 ) | ( n6464 & n30188 ) | ( n10485 & n30188 ) ;
  assign n47547 = ~n13566 & n45810 ;
  assign n47548 = n26362 ^ n5271 ^ n4576 ;
  assign n47549 = ( n6993 & ~n23120 ) | ( n6993 & n32007 ) | ( ~n23120 & n32007 ) ;
  assign n47550 = n22300 & ~n35704 ;
  assign n47551 = n47550 ^ n16813 ^ n13017 ;
  assign n47552 = n47551 ^ n34160 ^ n15430 ;
  assign n47554 = n29283 ^ n6687 ^ n2465 ;
  assign n47555 = ~n23815 & n47554 ;
  assign n47556 = n47555 ^ n44512 ^ 1'b0 ;
  assign n47553 = n29432 ^ n486 ^ 1'b0 ;
  assign n47557 = n47556 ^ n47553 ^ n33877 ;
  assign n47558 = n40775 & n45068 ;
  assign n47559 = ~n4458 & n47558 ;
  assign n47560 = n40362 ^ n20660 ^ 1'b0 ;
  assign n47561 = ( n3326 & ~n22468 ) | ( n3326 & n28592 ) | ( ~n22468 & n28592 ) ;
  assign n47562 = ( n1137 & ~n20946 ) | ( n1137 & n45894 ) | ( ~n20946 & n45894 ) ;
  assign n47563 = n38904 ^ n28239 ^ n13697 ;
  assign n47564 = n47563 ^ n31617 ^ n19017 ;
  assign n47565 = ( n19370 & n42652 ) | ( n19370 & ~n47564 ) | ( n42652 & ~n47564 ) ;
  assign n47566 = ( ~n1667 & n25938 ) | ( ~n1667 & n35051 ) | ( n25938 & n35051 ) ;
  assign n47567 = ( n16205 & n23701 ) | ( n16205 & ~n47566 ) | ( n23701 & ~n47566 ) ;
  assign n47568 = n24778 ^ n9594 ^ 1'b0 ;
  assign n47569 = ~n1973 & n47568 ;
  assign n47570 = n28520 ^ n9284 ^ 1'b0 ;
  assign n47571 = ( n47468 & n47569 ) | ( n47468 & ~n47570 ) | ( n47569 & ~n47570 ) ;
  assign n47572 = n27165 ^ n20901 ^ n2691 ;
  assign n47573 = ( n4481 & n14200 ) | ( n4481 & n25877 ) | ( n14200 & n25877 ) ;
  assign n47574 = n47573 ^ n11524 ^ n6181 ;
  assign n47575 = n38814 ^ n17080 ^ 1'b0 ;
  assign n47576 = n35929 ^ n27461 ^ n11760 ;
  assign n47577 = n16604 ^ n8851 ^ n3315 ;
  assign n47578 = ( n572 & n23746 ) | ( n572 & n47577 ) | ( n23746 & n47577 ) ;
  assign n47579 = n12288 | n47578 ;
  assign n47580 = n18291 ^ n13559 ^ n1663 ;
  assign n47581 = n47580 ^ n5380 ^ 1'b0 ;
  assign n47582 = ( n2537 & n24313 ) | ( n2537 & n26243 ) | ( n24313 & n26243 ) ;
  assign n47583 = ( n19709 & n37998 ) | ( n19709 & n47582 ) | ( n37998 & n47582 ) ;
  assign n47584 = n24439 ^ n20272 ^ 1'b0 ;
  assign n47585 = n47584 ^ n41164 ^ n34115 ;
  assign n47586 = n47585 ^ n26075 ^ n1647 ;
  assign n47587 = n47586 ^ n13777 ^ n12314 ;
  assign n47588 = n10070 ^ n8605 ^ n3773 ;
  assign n47589 = n47588 ^ n18817 ^ n4822 ;
  assign n47590 = n1363 & ~n47589 ;
  assign n47591 = n6564 & n6703 ;
  assign n47592 = n41098 ^ n17138 ^ 1'b0 ;
  assign n47593 = n24094 ^ n11136 ^ n1508 ;
  assign n47594 = n24654 ^ n13582 ^ 1'b0 ;
  assign n47595 = n47594 ^ n14444 ^ 1'b0 ;
  assign n47596 = ~n47593 & n47595 ;
  assign n47597 = ( n1733 & ~n6063 ) | ( n1733 & n46356 ) | ( ~n6063 & n46356 ) ;
  assign n47598 = ~n10098 & n10563 ;
  assign n47599 = n47598 ^ n13328 ^ x4 ;
  assign n47600 = n47599 ^ n42427 ^ n11264 ;
  assign n47601 = n47600 ^ n43335 ^ n23736 ;
  assign n47602 = n388 & ~n35713 ;
  assign n47603 = n47602 ^ n24162 ^ n6766 ;
  assign n47604 = n7632 ^ n1016 ^ 1'b0 ;
  assign n47605 = n39618 ^ n35686 ^ 1'b0 ;
  assign n47606 = n14857 ^ n9606 ^ 1'b0 ;
  assign n47607 = ( n17966 & n29243 ) | ( n17966 & n47606 ) | ( n29243 & n47606 ) ;
  assign n47608 = n1592 & n12480 ;
  assign n47609 = ( n10598 & n34213 ) | ( n10598 & ~n47608 ) | ( n34213 & ~n47608 ) ;
  assign n47610 = ( n47605 & ~n47607 ) | ( n47605 & n47609 ) | ( ~n47607 & n47609 ) ;
  assign n47611 = n12496 ^ n12063 ^ n7738 ;
  assign n47612 = n47611 ^ n29138 ^ n5777 ;
  assign n47613 = ( n10664 & ~n29269 ) | ( n10664 & n37354 ) | ( ~n29269 & n37354 ) ;
  assign n47614 = ~n26172 & n46723 ;
  assign n47615 = ~n17301 & n47614 ;
  assign n47616 = n13102 ^ n321 ^ 1'b0 ;
  assign n47617 = ~n45304 & n47616 ;
  assign n47618 = ( n10301 & n21890 ) | ( n10301 & n24065 ) | ( n21890 & n24065 ) ;
  assign n47619 = n20873 & n33094 ;
  assign n47620 = ~n30880 & n47619 ;
  assign n47621 = n47620 ^ n30846 ^ n4430 ;
  assign n47622 = n47621 ^ n26224 ^ 1'b0 ;
  assign n47623 = n44425 ^ n34220 ^ n4396 ;
  assign n47631 = n38181 ^ n4394 ^ 1'b0 ;
  assign n47629 = n15434 ^ n5359 ^ 1'b0 ;
  assign n47625 = n28599 ^ n23430 ^ n17834 ;
  assign n47624 = n16443 ^ n5088 ^ 1'b0 ;
  assign n47626 = n47625 ^ n47624 ^ n43073 ;
  assign n47627 = n9533 & n47626 ;
  assign n47628 = n47627 ^ n39531 ^ 1'b0 ;
  assign n47630 = n47629 ^ n47628 ^ n9723 ;
  assign n47632 = n47631 ^ n47630 ^ n16519 ;
  assign n47633 = ( n2220 & n28595 ) | ( n2220 & ~n29302 ) | ( n28595 & ~n29302 ) ;
  assign n47634 = n5860 ^ n3350 ^ n468 ;
  assign n47635 = n47634 ^ n2283 ^ 1'b0 ;
  assign n47636 = n47635 ^ n2790 ^ 1'b0 ;
  assign n47637 = n14293 & ~n29925 ;
  assign n47638 = x227 & ~n24129 ;
  assign n47639 = n33550 & n47638 ;
  assign n47640 = ( n9353 & n21326 ) | ( n9353 & n22903 ) | ( n21326 & n22903 ) ;
  assign n47641 = n25992 & ~n47640 ;
  assign n47642 = n17463 & n47641 ;
  assign n47643 = n25737 ^ n14141 ^ n12794 ;
  assign n47646 = n42009 ^ n41481 ^ 1'b0 ;
  assign n47644 = n9535 ^ n5271 ^ 1'b0 ;
  assign n47645 = ( n1439 & ~n10852 ) | ( n1439 & n47644 ) | ( ~n10852 & n47644 ) ;
  assign n47647 = n47646 ^ n47645 ^ n15261 ;
  assign n47648 = ( n1077 & n7371 ) | ( n1077 & ~n17775 ) | ( n7371 & ~n17775 ) ;
  assign n47649 = n47648 ^ n6059 ^ n5531 ;
  assign n47650 = n31562 & n41326 ;
  assign n47651 = ( ~n2844 & n4806 ) | ( ~n2844 & n12666 ) | ( n4806 & n12666 ) ;
  assign n47652 = n47651 ^ n9276 ^ n818 ;
  assign n47653 = ( n47649 & n47650 ) | ( n47649 & ~n47652 ) | ( n47650 & ~n47652 ) ;
  assign n47654 = n47653 ^ n25590 ^ n3020 ;
  assign n47655 = n38865 ^ n4500 ^ 1'b0 ;
  assign n47656 = n47655 ^ n20223 ^ n20210 ;
  assign n47657 = n24891 ^ n12251 ^ n11709 ;
  assign n47658 = ( n6845 & n22702 ) | ( n6845 & ~n30308 ) | ( n22702 & ~n30308 ) ;
  assign n47659 = n47658 ^ n26693 ^ n19370 ;
  assign n47660 = ( n14228 & ~n36222 ) | ( n14228 & n47659 ) | ( ~n36222 & n47659 ) ;
  assign n47661 = ( n6769 & n47657 ) | ( n6769 & ~n47660 ) | ( n47657 & ~n47660 ) ;
  assign n47662 = n40019 ^ n37833 ^ n27740 ;
  assign n47665 = n16486 ^ n11068 ^ n2413 ;
  assign n47666 = n47665 ^ n16332 ^ n15250 ;
  assign n47667 = n6817 | n47666 ;
  assign n47663 = n13757 ^ n6658 ^ n3360 ;
  assign n47664 = ( ~n18973 & n29419 ) | ( ~n18973 & n47663 ) | ( n29419 & n47663 ) ;
  assign n47668 = n47667 ^ n47664 ^ n2294 ;
  assign n47669 = n42150 & ~n45880 ;
  assign n47670 = n47669 ^ n21780 ^ n15086 ;
  assign n47671 = n24337 ^ n18756 ^ n4175 ;
  assign n47672 = n47671 ^ n39112 ^ n19067 ;
  assign n47673 = n47670 & ~n47672 ;
  assign n47674 = ~n22309 & n47673 ;
  assign n47675 = ( ~n3728 & n14843 ) | ( ~n3728 & n15170 ) | ( n14843 & n15170 ) ;
  assign n47676 = n10361 ^ n7423 ^ 1'b0 ;
  assign n47677 = n47675 | n47676 ;
  assign n47678 = ( n15274 & ~n15640 ) | ( n15274 & n26930 ) | ( ~n15640 & n26930 ) ;
  assign n47679 = n37867 ^ n24192 ^ n17384 ;
  assign n47680 = ( n3968 & ~n9305 ) | ( n3968 & n42393 ) | ( ~n9305 & n42393 ) ;
  assign n47681 = n1088 & n38236 ;
  assign n47682 = n47681 ^ n2115 ^ 1'b0 ;
  assign n47683 = n22498 ^ n22137 ^ n17121 ;
  assign n47684 = ( n33211 & n47682 ) | ( n33211 & ~n47683 ) | ( n47682 & ~n47683 ) ;
  assign n47685 = ( n7554 & ~n16250 ) | ( n7554 & n36231 ) | ( ~n16250 & n36231 ) ;
  assign n47687 = ( n25661 & ~n27313 ) | ( n25661 & n35426 ) | ( ~n27313 & n35426 ) ;
  assign n47688 = n47687 ^ n25391 ^ n12853 ;
  assign n47686 = n3447 & n5929 ;
  assign n47689 = n47688 ^ n47686 ^ 1'b0 ;
  assign n47690 = n9200 | n36998 ;
  assign n47691 = n22782 | n47690 ;
  assign n47692 = n34339 ^ n29777 ^ n4553 ;
  assign n47693 = n28820 ^ x248 ^ 1'b0 ;
  assign n47694 = ( n8713 & n19671 ) | ( n8713 & ~n21485 ) | ( n19671 & ~n21485 ) ;
  assign n47695 = n412 | n47694 ;
  assign n47696 = n47695 ^ n35896 ^ 1'b0 ;
  assign n47697 = n47696 ^ n29468 ^ n22576 ;
  assign n47698 = n10416 ^ n7053 ^ n6080 ;
  assign n47699 = ( n5750 & ~n6232 ) | ( n5750 & n24089 ) | ( ~n6232 & n24089 ) ;
  assign n47700 = n47699 ^ n19576 ^ n11793 ;
  assign n47701 = n40833 ^ n26958 ^ 1'b0 ;
  assign n47702 = ~n3820 & n47701 ;
  assign n47703 = n47702 ^ n19357 ^ n8140 ;
  assign n47704 = n43245 ^ n17803 ^ 1'b0 ;
  assign n47705 = ~n1450 & n47704 ;
  assign n47706 = ( ~n4247 & n13605 ) | ( ~n4247 & n47705 ) | ( n13605 & n47705 ) ;
  assign n47707 = n46209 ^ n12080 ^ n6456 ;
  assign n47708 = ~n13123 & n47707 ;
  assign n47709 = n47708 ^ n18530 ^ 1'b0 ;
  assign n47710 = ( n3501 & ~n15704 ) | ( n3501 & n24701 ) | ( ~n15704 & n24701 ) ;
  assign n47711 = n5679 & ~n17331 ;
  assign n47712 = ( n7222 & n43486 ) | ( n7222 & ~n47711 ) | ( n43486 & ~n47711 ) ;
  assign n47713 = ( n12178 & n47710 ) | ( n12178 & ~n47712 ) | ( n47710 & ~n47712 ) ;
  assign n47714 = n31829 ^ n13088 ^ 1'b0 ;
  assign n47715 = n47714 ^ n37293 ^ n32829 ;
  assign n47716 = n47715 ^ n13173 ^ 1'b0 ;
  assign n47717 = ( n7526 & n32421 ) | ( n7526 & ~n47716 ) | ( n32421 & ~n47716 ) ;
  assign n47718 = n24472 ^ n23945 ^ n17003 ;
  assign n47719 = ( n4588 & ~n16271 ) | ( n4588 & n22666 ) | ( ~n16271 & n22666 ) ;
  assign n47720 = ( n2150 & n26731 ) | ( n2150 & ~n47719 ) | ( n26731 & ~n47719 ) ;
  assign n47721 = ( n2485 & n10490 ) | ( n2485 & ~n22880 ) | ( n10490 & ~n22880 ) ;
  assign n47722 = n47721 ^ n39519 ^ n5536 ;
  assign n47723 = n45987 & n47722 ;
  assign n47724 = n36455 ^ n19955 ^ n979 ;
  assign n47725 = ( n13719 & n44747 ) | ( n13719 & ~n45009 ) | ( n44747 & ~n45009 ) ;
  assign n47726 = ( n5448 & ~n22041 ) | ( n5448 & n47725 ) | ( ~n22041 & n47725 ) ;
  assign n47727 = n13684 ^ n2107 ^ 1'b0 ;
  assign n47728 = n31146 & n47727 ;
  assign n47729 = n6599 & n34444 ;
  assign n47730 = ~n47728 & n47729 ;
  assign n47731 = n47730 ^ n13074 ^ n12490 ;
  assign n47732 = n31532 ^ n11173 ^ 1'b0 ;
  assign n47733 = n36021 ^ n12797 ^ n7211 ;
  assign n47734 = n47733 ^ n35291 ^ 1'b0 ;
  assign n47735 = n47734 ^ n38872 ^ 1'b0 ;
  assign n47736 = n28726 ^ n22517 ^ n20161 ;
  assign n47737 = n31642 ^ n30403 ^ 1'b0 ;
  assign n47743 = n26315 ^ n8387 ^ 1'b0 ;
  assign n47741 = n18894 | n28943 ;
  assign n47742 = n47741 ^ n34490 ^ 1'b0 ;
  assign n47738 = n31003 ^ n12506 ^ n9611 ;
  assign n47739 = ~n9353 & n47738 ;
  assign n47740 = ~n35369 & n47739 ;
  assign n47744 = n47743 ^ n47742 ^ n47740 ;
  assign n47745 = ~n25663 & n43430 ;
  assign n47746 = n46202 & n47745 ;
  assign n47747 = n16744 & ~n47746 ;
  assign n47748 = n18637 & n47747 ;
  assign n47749 = n41849 ^ n40456 ^ 1'b0 ;
  assign n47750 = n32902 & ~n47749 ;
  assign n47751 = n22196 ^ n10523 ^ n6716 ;
  assign n47752 = n47751 ^ n45113 ^ n34987 ;
  assign n47753 = n46424 ^ n46050 ^ n10664 ;
  assign n47754 = n23573 ^ n14762 ^ 1'b0 ;
  assign n47755 = ~n16843 & n47754 ;
  assign n47756 = ( n3075 & ~n21503 ) | ( n3075 & n40724 ) | ( ~n21503 & n40724 ) ;
  assign n47757 = ( n34425 & n47755 ) | ( n34425 & n47756 ) | ( n47755 & n47756 ) ;
  assign n47758 = ( n7521 & n15111 ) | ( n7521 & n28729 ) | ( n15111 & n28729 ) ;
  assign n47759 = n47758 ^ n22480 ^ n6593 ;
  assign n47760 = n10296 | n20295 ;
  assign n47761 = n1367 & ~n47760 ;
  assign n47762 = ( ~n25493 & n27814 ) | ( ~n25493 & n47761 ) | ( n27814 & n47761 ) ;
  assign n47763 = n28310 ^ n4526 ^ n3960 ;
  assign n47764 = n9042 ^ n8124 ^ n6602 ;
  assign n47765 = ( ~n12303 & n38450 ) | ( ~n12303 & n47764 ) | ( n38450 & n47764 ) ;
  assign n47766 = n47765 ^ n41127 ^ n16669 ;
  assign n47768 = n13775 ^ n6057 ^ n3469 ;
  assign n47769 = n35857 ^ n17863 ^ n11664 ;
  assign n47770 = n47769 ^ n10463 ^ 1'b0 ;
  assign n47771 = n4238 & n47770 ;
  assign n47772 = n47768 & n47771 ;
  assign n47767 = ( n10282 & ~n11822 ) | ( n10282 & n25475 ) | ( ~n11822 & n25475 ) ;
  assign n47773 = n47772 ^ n47767 ^ n38639 ;
  assign n47774 = ( n6136 & n17144 ) | ( n6136 & ~n17389 ) | ( n17144 & ~n17389 ) ;
  assign n47775 = n12572 & ~n47774 ;
  assign n47776 = n47775 ^ n946 ^ 1'b0 ;
  assign n47778 = n5457 ^ n3497 ^ n3437 ;
  assign n47779 = ( ~n7912 & n18829 ) | ( ~n7912 & n47778 ) | ( n18829 & n47778 ) ;
  assign n47777 = n44718 ^ n17434 ^ 1'b0 ;
  assign n47780 = n47779 ^ n47777 ^ n41944 ;
  assign n47781 = n18516 ^ n16793 ^ n9824 ;
  assign n47782 = n26083 & ~n47781 ;
  assign n47783 = n47780 & n47782 ;
  assign n47784 = n11398 ^ n1318 ^ n431 ;
  assign n47785 = n27105 & n47784 ;
  assign n47789 = ( n18717 & n19747 ) | ( n18717 & n24933 ) | ( n19747 & n24933 ) ;
  assign n47786 = n25442 ^ n11416 ^ 1'b0 ;
  assign n47787 = ~n35970 & n47786 ;
  assign n47788 = n47787 ^ n34010 ^ n14252 ;
  assign n47790 = n47789 ^ n47788 ^ 1'b0 ;
  assign n47791 = n9923 ^ n9044 ^ n3260 ;
  assign n47792 = n47791 ^ n19786 ^ n3796 ;
  assign n47793 = ( n4665 & ~n13301 ) | ( n4665 & n21831 ) | ( ~n13301 & n21831 ) ;
  assign n47794 = n47793 ^ n44329 ^ n1856 ;
  assign n47795 = ( ~n4628 & n11949 ) | ( ~n4628 & n43901 ) | ( n11949 & n43901 ) ;
  assign n47796 = n47795 ^ n28465 ^ n23112 ;
  assign n47797 = n37811 | n47796 ;
  assign n47798 = n26063 & ~n47797 ;
  assign n47799 = n29952 ^ n23482 ^ n20170 ;
  assign n47800 = n47799 ^ n39091 ^ n3570 ;
  assign n47801 = ( n12174 & n22356 ) | ( n12174 & ~n47800 ) | ( n22356 & ~n47800 ) ;
  assign n47802 = ~n9351 & n47801 ;
  assign n47803 = ~n14876 & n47802 ;
  assign n47804 = n1405 & n11742 ;
  assign n47805 = ~n7413 & n47804 ;
  assign n47806 = ( n2615 & n14941 ) | ( n2615 & n20032 ) | ( n14941 & n20032 ) ;
  assign n47807 = ( n3335 & n26216 ) | ( n3335 & ~n47806 ) | ( n26216 & ~n47806 ) ;
  assign n47808 = ( ~n28876 & n45142 ) | ( ~n28876 & n47807 ) | ( n45142 & n47807 ) ;
  assign n47809 = n30033 ^ n6819 ^ n4094 ;
  assign n47810 = n29699 ^ n4813 ^ n1736 ;
  assign n47811 = ~n46131 & n46795 ;
  assign n47812 = n47811 ^ n45616 ^ n23628 ;
  assign n47813 = n6294 ^ n3532 ^ n927 ;
  assign n47814 = n42547 ^ n33449 ^ n5777 ;
  assign n47815 = ( n26220 & ~n47813 ) | ( n26220 & n47814 ) | ( ~n47813 & n47814 ) ;
  assign n47816 = ( n18873 & ~n31370 ) | ( n18873 & n33592 ) | ( ~n31370 & n33592 ) ;
  assign n47817 = ( n22007 & ~n23709 ) | ( n22007 & n46566 ) | ( ~n23709 & n46566 ) ;
  assign n47818 = n42547 ^ n35976 ^ n32760 ;
  assign n47819 = ( n3572 & n14331 ) | ( n3572 & ~n24740 ) | ( n14331 & ~n24740 ) ;
  assign n47820 = n29018 & ~n47819 ;
  assign n47821 = ~n20462 & n47820 ;
  assign n47822 = n3745 & ~n14140 ;
  assign n47823 = n47822 ^ n10780 ^ 1'b0 ;
  assign n47824 = n34111 & n44446 ;
  assign n47825 = n47824 ^ n46850 ^ n12519 ;
  assign n47826 = ( ~n4770 & n7927 ) | ( ~n4770 & n14635 ) | ( n7927 & n14635 ) ;
  assign n47827 = n47826 ^ n35694 ^ n5246 ;
  assign n47828 = ( n5175 & n35003 ) | ( n5175 & n47827 ) | ( n35003 & n47827 ) ;
  assign n47829 = n4078 & ~n12127 ;
  assign n47830 = n47829 ^ n11841 ^ 1'b0 ;
  assign n47831 = ( n2766 & n23074 ) | ( n2766 & ~n47830 ) | ( n23074 & ~n47830 ) ;
  assign n47832 = n41641 ^ n31528 ^ n5390 ;
  assign n47833 = n25369 ^ n21007 ^ n11434 ;
  assign n47834 = ( n14488 & n47780 ) | ( n14488 & ~n47833 ) | ( n47780 & ~n47833 ) ;
  assign n47835 = n12180 ^ n9072 ^ n7557 ;
  assign n47836 = n2883 ^ n1770 ^ 1'b0 ;
  assign n47837 = n35532 ^ n17870 ^ n6128 ;
  assign n47838 = n47837 ^ n15208 ^ 1'b0 ;
  assign n47840 = n38872 ^ n817 ^ 1'b0 ;
  assign n47839 = n2349 | n29739 ;
  assign n47841 = n47840 ^ n47839 ^ 1'b0 ;
  assign n47842 = n508 & ~n2006 ;
  assign n47843 = n47842 ^ n3989 ^ 1'b0 ;
  assign n47844 = n47843 ^ n16744 ^ n2750 ;
  assign n47845 = n47844 ^ n1770 ^ 1'b0 ;
  assign n47846 = n19207 ^ n12525 ^ n2753 ;
  assign n47847 = x135 | n47846 ;
  assign n47848 = ( ~x39 & n5264 ) | ( ~x39 & n34192 ) | ( n5264 & n34192 ) ;
  assign n47849 = n47848 ^ n21276 ^ 1'b0 ;
  assign n47850 = ( n23901 & n27214 ) | ( n23901 & ~n35734 ) | ( n27214 & ~n35734 ) ;
  assign n47851 = ( n5142 & n34317 ) | ( n5142 & ~n38901 ) | ( n34317 & ~n38901 ) ;
  assign n47852 = ( n14555 & n47850 ) | ( n14555 & ~n47851 ) | ( n47850 & ~n47851 ) ;
  assign n47853 = ( n9678 & n13417 ) | ( n9678 & n47852 ) | ( n13417 & n47852 ) ;
  assign n47854 = n12413 ^ n8515 ^ n1809 ;
  assign n47855 = n12947 & n47854 ;
  assign n47856 = ( n1902 & ~n7339 ) | ( n1902 & n27778 ) | ( ~n7339 & n27778 ) ;
  assign n47857 = ( n3096 & n14680 ) | ( n3096 & n47856 ) | ( n14680 & n47856 ) ;
  assign n47858 = n24390 ^ n4190 ^ n356 ;
  assign n47859 = n47858 ^ n42478 ^ 1'b0 ;
  assign n47860 = n47859 ^ n43617 ^ n7330 ;
  assign n47864 = n23867 ^ n15724 ^ n2802 ;
  assign n47861 = ( n19057 & n22478 ) | ( n19057 & ~n47778 ) | ( n22478 & ~n47778 ) ;
  assign n47862 = n29231 | n47861 ;
  assign n47863 = n47862 ^ n41993 ^ 1'b0 ;
  assign n47865 = n47864 ^ n47863 ^ 1'b0 ;
  assign n47866 = n47865 ^ n46666 ^ n15436 ;
  assign n47867 = n7241 ^ n4525 ^ n2900 ;
  assign n47868 = n709 & n47867 ;
  assign n47869 = n15435 & n47868 ;
  assign n47870 = n1165 | n47869 ;
  assign n47871 = n47870 ^ n6059 ^ 1'b0 ;
  assign n47872 = ( ~n35195 & n41039 ) | ( ~n35195 & n43238 ) | ( n41039 & n43238 ) ;
  assign n47873 = n47872 ^ n4265 ^ 1'b0 ;
  assign n47874 = n17991 ^ n12957 ^ n6465 ;
  assign n47875 = ( n22462 & ~n35967 ) | ( n22462 & n47874 ) | ( ~n35967 & n47874 ) ;
  assign n47876 = n1061 | n37952 ;
  assign n47877 = n27232 ^ n17520 ^ n5365 ;
  assign n47878 = n47877 ^ n27075 ^ 1'b0 ;
  assign n47879 = n20991 ^ n16723 ^ 1'b0 ;
  assign n47880 = n47879 ^ n38239 ^ n16746 ;
  assign n47881 = n21037 ^ n15129 ^ n662 ;
  assign n47882 = ( n9989 & n38978 ) | ( n9989 & ~n47881 ) | ( n38978 & ~n47881 ) ;
  assign n47883 = ( n30478 & n47880 ) | ( n30478 & ~n47882 ) | ( n47880 & ~n47882 ) ;
  assign n47884 = ( n5923 & ~n26044 ) | ( n5923 & n29340 ) | ( ~n26044 & n29340 ) ;
  assign n47885 = ( n4184 & n38557 ) | ( n4184 & ~n47696 ) | ( n38557 & ~n47696 ) ;
  assign n47886 = ( n8848 & n16524 ) | ( n8848 & n47885 ) | ( n16524 & n47885 ) ;
  assign n47887 = n3942 | n20223 ;
  assign n47888 = n22163 & ~n47887 ;
  assign n47889 = ( n8389 & n21084 ) | ( n8389 & ~n31370 ) | ( n21084 & ~n31370 ) ;
  assign n47890 = ( ~n23815 & n47888 ) | ( ~n23815 & n47889 ) | ( n47888 & n47889 ) ;
  assign n47891 = n13538 | n47524 ;
  assign n47892 = n30543 & n47891 ;
  assign n47893 = ~n37780 & n47892 ;
  assign n47894 = n47893 ^ n1541 ^ n345 ;
  assign n47895 = n19983 | n34099 ;
  assign n47896 = n8757 & n41946 ;
  assign n47897 = n9712 & n47896 ;
  assign n47898 = n35244 & ~n47897 ;
  assign n47899 = n14323 ^ n5100 ^ n4094 ;
  assign n47900 = n47541 ^ n18705 ^ n17134 ;
  assign n47901 = ( n2041 & ~n14353 ) | ( n2041 & n47900 ) | ( ~n14353 & n47900 ) ;
  assign n47902 = n29493 ^ n17899 ^ n5828 ;
  assign n47903 = n41333 ^ n14037 ^ 1'b0 ;
  assign n47904 = n33757 & n47903 ;
  assign n47905 = ~n35315 & n47904 ;
  assign n47906 = n47902 & n47905 ;
  assign n47907 = n35395 ^ n5417 ^ n4410 ;
  assign n47908 = ( n13519 & n19382 ) | ( n13519 & n35815 ) | ( n19382 & n35815 ) ;
  assign n47909 = ( n6324 & n44511 ) | ( n6324 & n47908 ) | ( n44511 & n47908 ) ;
  assign n47910 = n31234 ^ n19971 ^ 1'b0 ;
  assign n47911 = ~n8723 & n29396 ;
  assign n47912 = ( n20721 & ~n45767 ) | ( n20721 & n47911 ) | ( ~n45767 & n47911 ) ;
  assign n47913 = n47846 ^ n6161 ^ x122 ;
  assign n47914 = n47913 ^ n35026 ^ n23771 ;
  assign n47915 = ~n6907 & n42526 ;
  assign n47916 = ( n6607 & n10558 ) | ( n6607 & ~n47915 ) | ( n10558 & ~n47915 ) ;
  assign n47917 = n34548 & n47916 ;
  assign n47918 = n24939 | n42058 ;
  assign n47919 = n19296 ^ n19256 ^ n5627 ;
  assign n47920 = n9624 & ~n42922 ;
  assign n47921 = n46718 ^ n19951 ^ n7352 ;
  assign n47922 = n44755 ^ n34175 ^ n13428 ;
  assign n47923 = n47922 ^ n3623 ^ n2556 ;
  assign n47924 = ( n7165 & n47921 ) | ( n7165 & ~n47923 ) | ( n47921 & ~n47923 ) ;
  assign n47925 = ( ~n1412 & n9745 ) | ( ~n1412 & n12712 ) | ( n9745 & n12712 ) ;
  assign n47926 = n47925 ^ n26053 ^ n16105 ;
  assign n47927 = ( n12775 & ~n40333 ) | ( n12775 & n47926 ) | ( ~n40333 & n47926 ) ;
  assign n47928 = n17674 ^ n5661 ^ 1'b0 ;
  assign n47929 = ( n18389 & n33949 ) | ( n18389 & ~n47928 ) | ( n33949 & ~n47928 ) ;
  assign n47930 = n5670 ^ n5193 ^ 1'b0 ;
  assign n47931 = n35051 ^ n16142 ^ n555 ;
  assign n47932 = n47930 & n47931 ;
  assign n47933 = n42243 ^ n2342 ^ 1'b0 ;
  assign n47934 = n32687 & ~n45220 ;
  assign n47935 = n32886 ^ n12073 ^ x22 ;
  assign n47936 = n47935 ^ n18128 ^ n346 ;
  assign n47937 = ~n37420 & n47936 ;
  assign n47938 = n47937 ^ n22380 ^ n19535 ;
  assign n47939 = n40985 ^ n28199 ^ n3008 ;
  assign n47940 = n47939 ^ n43699 ^ n39654 ;
  assign n47941 = n39934 ^ n29691 ^ 1'b0 ;
  assign n47942 = n47648 ^ n25793 ^ n6436 ;
  assign n47943 = n4014 ^ n1279 ^ 1'b0 ;
  assign n47944 = n24285 ^ n8826 ^ n1321 ;
  assign n47945 = n10873 & n47944 ;
  assign n47946 = n26084 | n46350 ;
  assign n47947 = n47946 ^ n21984 ^ 1'b0 ;
  assign n47948 = ( n5784 & n7644 ) | ( n5784 & ~n10533 ) | ( n7644 & ~n10533 ) ;
  assign n47949 = n47948 ^ n47239 ^ n25563 ;
  assign n47950 = ( n17955 & ~n38857 ) | ( n17955 & n47949 ) | ( ~n38857 & n47949 ) ;
  assign n47951 = n20940 ^ n4354 ^ n2227 ;
  assign n47952 = n9455 ^ n4026 ^ 1'b0 ;
  assign n47953 = n47952 ^ n32004 ^ n1676 ;
  assign n47954 = n47953 ^ n35688 ^ n1557 ;
  assign n47955 = n15406 ^ n9057 ^ n9009 ;
  assign n47956 = n45082 ^ n34629 ^ n31139 ;
  assign n47957 = n26347 & ~n32211 ;
  assign n47958 = n47957 ^ n47611 ^ 1'b0 ;
  assign n47959 = ( ~n28254 & n31686 ) | ( ~n28254 & n41481 ) | ( n31686 & n41481 ) ;
  assign n47960 = n10308 & n11690 ;
  assign n47961 = n47960 ^ n16869 ^ 1'b0 ;
  assign n47962 = n5964 & ~n47961 ;
  assign n47963 = n47959 & n47962 ;
  assign n47964 = ( n5950 & ~n8360 ) | ( n5950 & n8692 ) | ( ~n8360 & n8692 ) ;
  assign n47965 = n47964 ^ n28070 ^ n22168 ;
  assign n47966 = n43213 ^ n21698 ^ n7368 ;
  assign n47967 = n6062 & ~n16194 ;
  assign n47968 = ~n1801 & n47967 ;
  assign n47969 = n47968 ^ n42008 ^ n21831 ;
  assign n47970 = n36643 ^ n17642 ^ n5229 ;
  assign n47971 = n47970 ^ n41886 ^ n19917 ;
  assign n47972 = n12654 ^ n3635 ^ 1'b0 ;
  assign n47974 = ( n36394 & n42948 ) | ( n36394 & ~n47955 ) | ( n42948 & ~n47955 ) ;
  assign n47973 = n3996 ^ n1447 ^ 1'b0 ;
  assign n47975 = n47974 ^ n47973 ^ 1'b0 ;
  assign n47976 = n10860 ^ n8454 ^ 1'b0 ;
  assign n47977 = n47976 ^ n17041 ^ n3865 ;
  assign n47978 = n1103 & n47977 ;
  assign n47979 = n47978 ^ n38874 ^ n24317 ;
  assign n47980 = ( n21073 & n30775 ) | ( n21073 & ~n47979 ) | ( n30775 & ~n47979 ) ;
  assign n47981 = n5840 & ~n47980 ;
  assign n47982 = n47981 ^ n20772 ^ 1'b0 ;
  assign n47983 = n3001 & n26244 ;
  assign n47984 = n47983 ^ n44511 ^ 1'b0 ;
  assign n47985 = n31749 ^ n22411 ^ n5921 ;
  assign n47986 = n47985 ^ n27165 ^ n25599 ;
  assign n47987 = n28624 ^ n21682 ^ 1'b0 ;
  assign n47988 = ~n5178 & n7385 ;
  assign n47989 = n47988 ^ n3993 ^ 1'b0 ;
  assign n47990 = ( n12045 & ~n14203 ) | ( n12045 & n47989 ) | ( ~n14203 & n47989 ) ;
  assign n47991 = n962 & ~n10852 ;
  assign n47992 = n16271 & n47991 ;
  assign n47993 = n47992 ^ n15614 ^ n13201 ;
  assign n47994 = n22363 ^ n15346 ^ n14569 ;
  assign n47995 = n44917 ^ n14865 ^ 1'b0 ;
  assign n47996 = ( n2361 & n11310 ) | ( n2361 & ~n14772 ) | ( n11310 & ~n14772 ) ;
  assign n47997 = ~n10548 & n22769 ;
  assign n47998 = n47996 & n47997 ;
  assign n47999 = ( n5853 & ~n7274 ) | ( n5853 & n22107 ) | ( ~n7274 & n22107 ) ;
  assign n48000 = n47999 ^ n45326 ^ n1317 ;
  assign n48001 = n48000 ^ n7875 ^ 1'b0 ;
  assign n48002 = ~n20374 & n48001 ;
  assign n48003 = n6743 | n21294 ;
  assign n48004 = ( ~n4603 & n13117 ) | ( ~n4603 & n14331 ) | ( n13117 & n14331 ) ;
  assign n48005 = ( ~n10302 & n26597 ) | ( ~n10302 & n48004 ) | ( n26597 & n48004 ) ;
  assign n48006 = ( n23992 & ~n37491 ) | ( n23992 & n48005 ) | ( ~n37491 & n48005 ) ;
  assign n48007 = ( n27560 & n39307 ) | ( n27560 & n42003 ) | ( n39307 & n42003 ) ;
  assign n48008 = ( ~n3831 & n7574 ) | ( ~n3831 & n7909 ) | ( n7574 & n7909 ) ;
  assign n48009 = n48008 ^ n7019 ^ 1'b0 ;
  assign n48010 = ( ~n6290 & n12646 ) | ( ~n6290 & n13747 ) | ( n12646 & n13747 ) ;
  assign n48011 = n33359 ^ n29357 ^ 1'b0 ;
  assign n48012 = ( n36486 & n48010 ) | ( n36486 & ~n48011 ) | ( n48010 & ~n48011 ) ;
  assign n48013 = n20012 ^ n19311 ^ 1'b0 ;
  assign n48015 = n29759 ^ n8946 ^ n2981 ;
  assign n48014 = ~n13070 & n45517 ;
  assign n48016 = n48015 ^ n48014 ^ 1'b0 ;
  assign n48017 = n6760 & ~n42892 ;
  assign n48018 = n48017 ^ n17951 ^ 1'b0 ;
  assign n48019 = n26472 & ~n28320 ;
  assign n48020 = n7116 | n48019 ;
  assign n48021 = n48020 ^ n2150 ^ 1'b0 ;
  assign n48022 = n15160 | n16493 ;
  assign n48023 = ( n1597 & ~n34394 ) | ( n1597 & n40268 ) | ( ~n34394 & n40268 ) ;
  assign n48026 = n46264 ^ n12556 ^ n2674 ;
  assign n48024 = n13861 & ~n36662 ;
  assign n48025 = n48024 ^ n25009 ^ 1'b0 ;
  assign n48027 = n48026 ^ n48025 ^ n19933 ;
  assign n48030 = n8314 ^ n5255 ^ n3622 ;
  assign n48028 = ~n14640 & n27791 ;
  assign n48029 = n1467 & n48028 ;
  assign n48031 = n48030 ^ n48029 ^ 1'b0 ;
  assign n48032 = n41260 ^ n12191 ^ n7085 ;
  assign n48033 = n46307 ^ n26738 ^ 1'b0 ;
  assign n48034 = ~n48032 & n48033 ;
  assign n48035 = n10137 & n48034 ;
  assign n48036 = n47179 ^ n32004 ^ 1'b0 ;
  assign n48037 = ( n19659 & n30250 ) | ( n19659 & ~n36636 ) | ( n30250 & ~n36636 ) ;
  assign n48038 = ( n1015 & n19334 ) | ( n1015 & n48037 ) | ( n19334 & n48037 ) ;
  assign n48039 = n48038 ^ n8067 ^ 1'b0 ;
  assign n48040 = ( n2550 & n5858 ) | ( n2550 & ~n10412 ) | ( n5858 & ~n10412 ) ;
  assign n48041 = ~n7148 & n47409 ;
  assign n48042 = n48040 & n48041 ;
  assign n48043 = n32612 ^ n32265 ^ 1'b0 ;
  assign n48044 = x193 & n48043 ;
  assign n48045 = ( n19218 & n32064 ) | ( n19218 & ~n37382 ) | ( n32064 & ~n37382 ) ;
  assign n48046 = ( n12838 & n29990 ) | ( n12838 & ~n41418 ) | ( n29990 & ~n41418 ) ;
  assign n48047 = n25428 ^ n8101 ^ n5159 ;
  assign n48048 = ( n6407 & n20918 ) | ( n6407 & n39569 ) | ( n20918 & n39569 ) ;
  assign n48049 = ( ~n20257 & n27727 ) | ( ~n20257 & n48048 ) | ( n27727 & n48048 ) ;
  assign n48050 = n17149 ^ n10135 ^ n4177 ;
  assign n48051 = n48050 ^ n42181 ^ n5363 ;
  assign n48052 = n13809 | n37594 ;
  assign n48053 = n1047 | n48052 ;
  assign n48054 = n36987 & n48053 ;
  assign n48055 = n48054 ^ n25038 ^ 1'b0 ;
  assign n48056 = n48055 ^ n32232 ^ n13142 ;
  assign n48057 = n25191 & ~n48056 ;
  assign n48058 = n28807 ^ n26383 ^ n16603 ;
  assign n48060 = ~n27573 & n43862 ;
  assign n48059 = ( x206 & ~n12493 ) | ( x206 & n29051 ) | ( ~n12493 & n29051 ) ;
  assign n48061 = n48060 ^ n48059 ^ n23517 ;
  assign n48062 = n13744 ^ n3107 ^ 1'b0 ;
  assign n48063 = n23724 | n48062 ;
  assign n48064 = ~n14506 & n34160 ;
  assign n48065 = ~n44511 & n48064 ;
  assign n48066 = ~n17555 & n20365 ;
  assign n48067 = n48065 & n48066 ;
  assign n48068 = n16436 | n45841 ;
  assign n48069 = n48067 & ~n48068 ;
  assign n48070 = n26344 ^ n12980 ^ n3353 ;
  assign n48071 = n48070 ^ n42868 ^ n2973 ;
  assign n48072 = n333 & n26251 ;
  assign n48073 = n48072 ^ n33693 ^ 1'b0 ;
  assign n48074 = ( ~n4650 & n33016 ) | ( ~n4650 & n48073 ) | ( n33016 & n48073 ) ;
  assign n48075 = n36198 ^ n8452 ^ 1'b0 ;
  assign n48076 = n17611 & n48075 ;
  assign n48077 = n48076 ^ n18544 ^ n5123 ;
  assign n48078 = ( n3673 & ~n23101 ) | ( n3673 & n34383 ) | ( ~n23101 & n34383 ) ;
  assign n48079 = n48078 ^ n28339 ^ n3110 ;
  assign n48080 = n48079 ^ n36603 ^ n24746 ;
  assign n48081 = n30471 ^ n25404 ^ n4859 ;
  assign n48082 = n34964 ^ n32974 ^ n8314 ;
  assign n48083 = n5905 ^ n5736 ^ n795 ;
  assign n48084 = n48083 ^ n9811 ^ n1684 ;
  assign n48085 = n48084 ^ n11760 ^ 1'b0 ;
  assign n48086 = ( n8337 & n19641 ) | ( n8337 & n35444 ) | ( n19641 & n35444 ) ;
  assign n48087 = n19471 ^ n18006 ^ n15915 ;
  assign n48088 = ( ~n40348 & n48086 ) | ( ~n40348 & n48087 ) | ( n48086 & n48087 ) ;
  assign n48089 = n22303 & ~n27015 ;
  assign n48090 = n10989 & n48089 ;
  assign n48091 = n1954 & ~n2041 ;
  assign n48092 = n48091 ^ n1223 ^ 1'b0 ;
  assign n48093 = n5891 & ~n48092 ;
  assign n48094 = n48093 ^ n10111 ^ 1'b0 ;
  assign n48095 = n9445 | n12556 ;
  assign n48096 = n44888 ^ n3232 ^ 1'b0 ;
  assign n48097 = ~n41995 & n48096 ;
  assign n48098 = n48097 ^ n8690 ^ 1'b0 ;
  assign n48099 = n37714 ^ n5376 ^ 1'b0 ;
  assign n48100 = n23592 & n48099 ;
  assign n48101 = n48100 ^ n47778 ^ 1'b0 ;
  assign n48102 = n48101 ^ n25329 ^ 1'b0 ;
  assign n48103 = ( ~n8784 & n48098 ) | ( ~n8784 & n48102 ) | ( n48098 & n48102 ) ;
  assign n48104 = n22063 ^ n10549 ^ n8559 ;
  assign n48105 = n33032 ^ n17756 ^ n3469 ;
  assign n48106 = ( n14452 & ~n17155 ) | ( n14452 & n34134 ) | ( ~n17155 & n34134 ) ;
  assign n48107 = n48106 ^ n28226 ^ n23074 ;
  assign n48108 = n48107 ^ n17862 ^ n10111 ;
  assign n48109 = ( n660 & ~n15015 ) | ( n660 & n21546 ) | ( ~n15015 & n21546 ) ;
  assign n48110 = ( n9884 & n26549 ) | ( n9884 & n48109 ) | ( n26549 & n48109 ) ;
  assign n48111 = n19488 ^ n1703 ^ 1'b0 ;
  assign n48112 = ( n3981 & ~n17464 ) | ( n3981 & n47895 ) | ( ~n17464 & n47895 ) ;
  assign n48114 = n43507 ^ n13009 ^ n1315 ;
  assign n48113 = ( n16434 & n17178 ) | ( n16434 & ~n32362 ) | ( n17178 & ~n32362 ) ;
  assign n48115 = n48114 ^ n48113 ^ n7515 ;
  assign n48117 = ( n16030 & ~n20957 ) | ( n16030 & n41082 ) | ( ~n20957 & n41082 ) ;
  assign n48116 = ( n24905 & n26279 ) | ( n24905 & n27697 ) | ( n26279 & n27697 ) ;
  assign n48118 = n48117 ^ n48116 ^ n1791 ;
  assign n48119 = ( n30596 & n45215 ) | ( n30596 & n48118 ) | ( n45215 & n48118 ) ;
  assign n48120 = n39423 ^ n36649 ^ n27573 ;
  assign n48121 = n2759 ^ n1175 ^ 1'b0 ;
  assign n48125 = n9578 & n27553 ;
  assign n48124 = n14051 ^ n5522 ^ 1'b0 ;
  assign n48122 = n1565 & ~n2910 ;
  assign n48123 = n48122 ^ n11594 ^ 1'b0 ;
  assign n48126 = n48125 ^ n48124 ^ n48123 ;
  assign n48127 = ( n5964 & ~n17485 ) | ( n5964 & n23785 ) | ( ~n17485 & n23785 ) ;
  assign n48128 = n37662 ^ n17003 ^ n10855 ;
  assign n48129 = n12267 & ~n25130 ;
  assign n48130 = n16870 & n25005 ;
  assign n48131 = n48130 ^ n22488 ^ 1'b0 ;
  assign n48132 = n29327 & n39546 ;
  assign n48133 = ~n13559 & n48132 ;
  assign n48137 = ( n5453 & n12511 ) | ( n5453 & n21879 ) | ( n12511 & n21879 ) ;
  assign n48138 = ( n2727 & ~n22833 ) | ( n2727 & n48137 ) | ( ~n22833 & n48137 ) ;
  assign n48134 = n14894 ^ n2911 ^ 1'b0 ;
  assign n48135 = n2397 & n48134 ;
  assign n48136 = ( n10123 & n10928 ) | ( n10123 & ~n48135 ) | ( n10928 & ~n48135 ) ;
  assign n48139 = n48138 ^ n48136 ^ n5014 ;
  assign n48140 = n28293 ^ n7197 ^ n3206 ;
  assign n48141 = ( n17359 & n18744 ) | ( n17359 & n33027 ) | ( n18744 & n33027 ) ;
  assign n48142 = ( n21834 & n34736 ) | ( n21834 & n37660 ) | ( n34736 & n37660 ) ;
  assign n48143 = n48142 ^ n20515 ^ 1'b0 ;
  assign n48144 = n12246 & ~n21681 ;
  assign n48145 = n48144 ^ n25940 ^ n22933 ;
  assign n48146 = n14605 | n23595 ;
  assign n48147 = ( n2474 & ~n5260 ) | ( n2474 & n42992 ) | ( ~n5260 & n42992 ) ;
  assign n48148 = ( n2156 & n35724 ) | ( n2156 & ~n48147 ) | ( n35724 & ~n48147 ) ;
  assign n48149 = ~n25228 & n46415 ;
  assign n48150 = ( ~n9572 & n24733 ) | ( ~n9572 & n48078 ) | ( n24733 & n48078 ) ;
  assign n48151 = n453 & n31626 ;
  assign n48152 = ~n48150 & n48151 ;
  assign n48153 = n29057 ^ n23936 ^ 1'b0 ;
  assign n48154 = n42369 & n48153 ;
  assign n48155 = n48154 ^ n35910 ^ n4824 ;
  assign n48156 = ( n6057 & n37034 ) | ( n6057 & ~n47320 ) | ( n37034 & ~n47320 ) ;
  assign n48157 = n48156 ^ n39676 ^ n30398 ;
  assign n48158 = n48155 & ~n48157 ;
  assign n48159 = ~n8734 & n19544 ;
  assign n48160 = ( ~n10892 & n41786 ) | ( ~n10892 & n48159 ) | ( n41786 & n48159 ) ;
  assign n48161 = ( ~n2775 & n32161 ) | ( ~n2775 & n39506 ) | ( n32161 & n39506 ) ;
  assign n48162 = n29320 ^ n21172 ^ n7929 ;
  assign n48163 = n19558 ^ n12269 ^ 1'b0 ;
  assign n48164 = ~n32050 & n48163 ;
  assign n48165 = n48164 ^ n46742 ^ n16006 ;
  assign n48166 = ( n34053 & n44459 ) | ( n34053 & n48165 ) | ( n44459 & n48165 ) ;
  assign n48167 = n42692 ^ n24127 ^ n16778 ;
  assign n48168 = ( n28339 & n45082 ) | ( n28339 & ~n48167 ) | ( n45082 & ~n48167 ) ;
  assign n48170 = n27101 ^ n18370 ^ n559 ;
  assign n48169 = n41288 ^ n19219 ^ n3326 ;
  assign n48171 = n48170 ^ n48169 ^ n45648 ;
  assign n48172 = ~n3203 & n48171 ;
  assign n48175 = n16184 ^ n15445 ^ n5006 ;
  assign n48174 = ~n28341 & n38779 ;
  assign n48176 = n48175 ^ n48174 ^ n39588 ;
  assign n48173 = n3086 & ~n33004 ;
  assign n48177 = n48176 ^ n48173 ^ 1'b0 ;
  assign n48178 = n36677 ^ n23020 ^ n14597 ;
  assign n48179 = n13324 & ~n48178 ;
  assign n48181 = ( n7446 & n22866 ) | ( n7446 & n33825 ) | ( n22866 & n33825 ) ;
  assign n48180 = n19918 ^ n14070 ^ n6807 ;
  assign n48182 = n48181 ^ n48180 ^ 1'b0 ;
  assign n48183 = n48179 & ~n48182 ;
  assign n48184 = n45533 ^ n28691 ^ 1'b0 ;
  assign n48185 = n21870 | n48184 ;
  assign n48186 = n27633 & n46479 ;
  assign n48187 = n48186 ^ n3370 ^ 1'b0 ;
  assign n48188 = ( n8897 & n13969 ) | ( n8897 & ~n39458 ) | ( n13969 & ~n39458 ) ;
  assign n48189 = ( ~n5889 & n26264 ) | ( ~n5889 & n44642 ) | ( n26264 & n44642 ) ;
  assign n48190 = n18171 | n48189 ;
  assign n48191 = n29817 & n48190 ;
  assign n48192 = n48191 ^ n36327 ^ 1'b0 ;
  assign n48193 = n15717 ^ n12556 ^ 1'b0 ;
  assign n48194 = n48192 & n48193 ;
  assign n48195 = n48194 ^ n34500 ^ n8896 ;
  assign n48196 = ( n15309 & n21684 ) | ( n15309 & n22481 ) | ( n21684 & n22481 ) ;
  assign n48197 = ( n23091 & n23710 ) | ( n23091 & n48196 ) | ( n23710 & n48196 ) ;
  assign n48198 = n27269 ^ n24895 ^ n4128 ;
  assign n48199 = ( ~n13753 & n29940 ) | ( ~n13753 & n33273 ) | ( n29940 & n33273 ) ;
  assign n48200 = n1775 & ~n10368 ;
  assign n48201 = n48199 & n48200 ;
  assign n48202 = n23329 ^ n14223 ^ n8652 ;
  assign n48203 = n48202 ^ n21216 ^ n1462 ;
  assign n48204 = n41137 ^ n15010 ^ 1'b0 ;
  assign n48205 = ( n18132 & n25844 ) | ( n18132 & n27538 ) | ( n25844 & n27538 ) ;
  assign n48206 = n48205 ^ n46622 ^ 1'b0 ;
  assign n48207 = n22147 ^ n21614 ^ n7583 ;
  assign n48208 = n48207 ^ n42258 ^ n13638 ;
  assign n48209 = n37066 ^ n36143 ^ n6662 ;
  assign n48213 = n27571 ^ n26394 ^ n20390 ;
  assign n48210 = ( n272 & ~n3480 ) | ( n272 & n24370 ) | ( ~n3480 & n24370 ) ;
  assign n48211 = ( n27449 & n35066 ) | ( n27449 & n48210 ) | ( n35066 & n48210 ) ;
  assign n48212 = n48211 ^ n25950 ^ n4187 ;
  assign n48214 = n48213 ^ n48212 ^ n8792 ;
  assign n48215 = n19590 ^ n6434 ^ 1'b0 ;
  assign n48216 = ~n1652 & n48215 ;
  assign n48217 = n7803 ^ n6472 ^ n3025 ;
  assign n48218 = n46208 ^ n37204 ^ 1'b0 ;
  assign n48219 = ~n48217 & n48218 ;
  assign n48220 = ( ~n21006 & n22126 ) | ( ~n21006 & n35929 ) | ( n22126 & n35929 ) ;
  assign n48221 = ( n11848 & n41291 ) | ( n11848 & n48220 ) | ( n41291 & n48220 ) ;
  assign n48222 = n31982 ^ n17620 ^ n16352 ;
  assign n48223 = n18109 & ~n48222 ;
  assign n48224 = ( n950 & n32487 ) | ( n950 & n42202 ) | ( n32487 & n42202 ) ;
  assign n48225 = n48224 ^ n44410 ^ n11970 ;
  assign n48226 = n45216 ^ n34409 ^ n13146 ;
  assign n48227 = n46089 ^ n31054 ^ n4547 ;
  assign n48228 = n34467 ^ n8382 ^ 1'b0 ;
  assign n48229 = n44996 ^ n40769 ^ 1'b0 ;
  assign n48230 = n13324 & n47832 ;
  assign n48231 = n48230 ^ n32041 ^ 1'b0 ;
  assign n48232 = n15757 & ~n32385 ;
  assign n48237 = ( n3174 & ~n23371 ) | ( n3174 & n26372 ) | ( ~n23371 & n26372 ) ;
  assign n48238 = ( ~n5368 & n12995 ) | ( ~n5368 & n48237 ) | ( n12995 & n48237 ) ;
  assign n48239 = n29692 ^ n14315 ^ n4176 ;
  assign n48240 = ( ~n46629 & n48238 ) | ( ~n46629 & n48239 ) | ( n48238 & n48239 ) ;
  assign n48233 = ~n5299 & n12005 ;
  assign n48234 = n24917 & n48233 ;
  assign n48235 = ( n12721 & ~n24938 ) | ( n12721 & n48234 ) | ( ~n24938 & n48234 ) ;
  assign n48236 = n48235 ^ n23762 ^ n20925 ;
  assign n48241 = n48240 ^ n48236 ^ n45854 ;
  assign n48242 = ( n13574 & ~n16024 ) | ( n13574 & n26279 ) | ( ~n16024 & n26279 ) ;
  assign n48243 = ( n25330 & ~n30524 ) | ( n25330 & n48242 ) | ( ~n30524 & n48242 ) ;
  assign n48244 = n18843 ^ n10908 ^ n914 ;
  assign n48245 = ( n31168 & n38245 ) | ( n31168 & ~n38839 ) | ( n38245 & ~n38839 ) ;
  assign n48246 = n12359 & n48245 ;
  assign n48247 = n48244 & n48246 ;
  assign n48248 = ( n22615 & n36845 ) | ( n22615 & n48247 ) | ( n36845 & n48247 ) ;
  assign n48249 = n7450 & n14233 ;
  assign n48250 = n9416 ^ n7358 ^ 1'b0 ;
  assign n48251 = ( ~n21451 & n23196 ) | ( ~n21451 & n48250 ) | ( n23196 & n48250 ) ;
  assign n48252 = ( n5228 & n48249 ) | ( n5228 & ~n48251 ) | ( n48249 & ~n48251 ) ;
  assign n48253 = ( n16168 & n22499 ) | ( n16168 & n34348 ) | ( n22499 & n34348 ) ;
  assign n48254 = ( n8336 & n15663 ) | ( n8336 & ~n26931 ) | ( n15663 & ~n26931 ) ;
  assign n48255 = n29136 ^ n3913 ^ 1'b0 ;
  assign n48256 = n33429 ^ n25376 ^ n4858 ;
  assign n48257 = ( n14974 & ~n48255 ) | ( n14974 & n48256 ) | ( ~n48255 & n48256 ) ;
  assign n48258 = n15685 ^ n12498 ^ 1'b0 ;
  assign n48259 = n5834 & n48258 ;
  assign n48260 = n37384 ^ n14554 ^ n4729 ;
  assign n48261 = n24904 & ~n48260 ;
  assign n48262 = n13285 & n48261 ;
  assign n48263 = n48259 | n48262 ;
  assign n48264 = n45571 ^ n30615 ^ n2738 ;
  assign n48265 = n48264 ^ n44029 ^ n11611 ;
  assign n48268 = n21383 ^ n14806 ^ n2721 ;
  assign n48267 = ( n6539 & n13544 ) | ( n6539 & n39161 ) | ( n13544 & n39161 ) ;
  assign n48266 = n24492 | n46309 ;
  assign n48269 = n48268 ^ n48267 ^ n48266 ;
  assign n48270 = n43490 ^ n15777 ^ 1'b0 ;
  assign n48271 = ( n16763 & n41631 ) | ( n16763 & n48113 ) | ( n41631 & n48113 ) ;
  assign n48272 = n13493 ^ n9641 ^ n3007 ;
  assign n48273 = n31559 & ~n48272 ;
  assign n48274 = ~n12943 & n27035 ;
  assign n48275 = n46544 ^ n31111 ^ n6563 ;
  assign n48278 = n20624 ^ n14348 ^ 1'b0 ;
  assign n48279 = n48278 ^ n19713 ^ n19008 ;
  assign n48276 = ( ~n24575 & n35164 ) | ( ~n24575 & n47631 ) | ( n35164 & n47631 ) ;
  assign n48277 = ~n29811 & n48276 ;
  assign n48280 = n48279 ^ n48277 ^ 1'b0 ;
  assign n48281 = n19962 ^ n6787 ^ n1894 ;
  assign n48282 = ( n5487 & n22752 ) | ( n5487 & ~n48281 ) | ( n22752 & ~n48281 ) ;
  assign n48283 = n9543 | n29231 ;
  assign n48284 = n48282 | n48283 ;
  assign n48285 = ~n14344 & n17014 ;
  assign n48286 = n24359 & n48285 ;
  assign n48288 = n3277 | n37081 ;
  assign n48289 = n48288 ^ n33498 ^ 1'b0 ;
  assign n48290 = n47683 & ~n48289 ;
  assign n48291 = n48290 ^ n20280 ^ 1'b0 ;
  assign n48287 = n39514 ^ n36112 ^ n653 ;
  assign n48292 = n48291 ^ n48287 ^ n8489 ;
  assign n48293 = n28487 ^ n3298 ^ n2795 ;
  assign n48294 = n48293 ^ n10216 ^ n7727 ;
  assign n48295 = n45429 | n46432 ;
  assign n48296 = n13721 ^ n3352 ^ n464 ;
  assign n48297 = n48296 ^ n47225 ^ n16163 ;
  assign n48298 = ( n6571 & ~n9598 ) | ( n6571 & n13673 ) | ( ~n9598 & n13673 ) ;
  assign n48299 = ( n1339 & n6694 ) | ( n1339 & ~n21593 ) | ( n6694 & ~n21593 ) ;
  assign n48300 = n48299 ^ n2171 ^ 1'b0 ;
  assign n48301 = n29409 ^ n14322 ^ 1'b0 ;
  assign n48302 = ~n48300 & n48301 ;
  assign n48303 = n48302 ^ n2564 ^ 1'b0 ;
  assign n48304 = n23180 ^ n11277 ^ n1549 ;
  assign n48305 = ( n3392 & n10256 ) | ( n3392 & n48304 ) | ( n10256 & n48304 ) ;
  assign n48306 = n30681 ^ n7444 ^ 1'b0 ;
  assign n48307 = n9061 ^ x186 ^ 1'b0 ;
  assign n48308 = n1560 | n48307 ;
  assign n48309 = ( n11785 & n21073 ) | ( n11785 & ~n21250 ) | ( n21073 & ~n21250 ) ;
  assign n48310 = n29992 ^ n19513 ^ n17633 ;
  assign n48311 = n48309 | n48310 ;
  assign n48312 = ( n4335 & n29140 ) | ( n4335 & n39117 ) | ( n29140 & n39117 ) ;
  assign n48313 = n48312 ^ n42640 ^ n8872 ;
  assign n48314 = n44090 ^ n17233 ^ n3443 ;
  assign n48315 = n48314 ^ n45149 ^ n35656 ;
  assign n48316 = ( n25375 & n42077 ) | ( n25375 & n45223 ) | ( n42077 & n45223 ) ;
  assign n48317 = n41189 ^ n33531 ^ n6564 ;
  assign n48318 = n48317 ^ n14371 ^ n4684 ;
  assign n48319 = ( n15313 & ~n30700 ) | ( n15313 & n48224 ) | ( ~n30700 & n48224 ) ;
  assign n48320 = n48319 ^ n38017 ^ n8162 ;
  assign n48321 = n39094 ^ n20508 ^ n3521 ;
  assign n48322 = n29584 & ~n48321 ;
  assign n48323 = n48322 ^ n44301 ^ 1'b0 ;
  assign n48324 = n6809 | n7904 ;
  assign n48325 = n48324 ^ n8997 ^ 1'b0 ;
  assign n48326 = ( n1729 & ~n7297 ) | ( n1729 & n22996 ) | ( ~n7297 & n22996 ) ;
  assign n48327 = ( ~n23251 & n37624 ) | ( ~n23251 & n48326 ) | ( n37624 & n48326 ) ;
  assign n48328 = n48327 ^ n8224 ^ 1'b0 ;
  assign n48329 = n48325 | n48328 ;
  assign n48330 = n39813 ^ n21376 ^ n9302 ;
  assign n48331 = n48330 ^ n6058 ^ 1'b0 ;
  assign n48332 = n32752 | n48331 ;
  assign n48333 = ( ~n6272 & n11050 ) | ( ~n6272 & n22249 ) | ( n11050 & n22249 ) ;
  assign n48334 = ( n9834 & ~n36565 ) | ( n9834 & n48333 ) | ( ~n36565 & n48333 ) ;
  assign n48335 = n48334 ^ n25985 ^ n20006 ;
  assign n48336 = ( n6424 & n11163 ) | ( n6424 & ~n48335 ) | ( n11163 & ~n48335 ) ;
  assign n48337 = n48336 ^ n38052 ^ n8569 ;
  assign n48338 = n22525 ^ n19899 ^ n19539 ;
  assign n48339 = n45632 ^ n32295 ^ n592 ;
  assign n48340 = ( n27982 & ~n48338 ) | ( n27982 & n48339 ) | ( ~n48338 & n48339 ) ;
  assign n48341 = n34351 & n36257 ;
  assign n48342 = n29499 ^ n8121 ^ n7732 ;
  assign n48343 = n48342 ^ n38752 ^ n3433 ;
  assign n48344 = n48343 ^ n46031 ^ n33597 ;
  assign n48345 = ( n45210 & n48341 ) | ( n45210 & ~n48344 ) | ( n48341 & ~n48344 ) ;
  assign n48346 = n38287 ^ n36264 ^ n25537 ;
  assign n48347 = n47621 | n48346 ;
  assign n48348 = n14938 & n48347 ;
  assign n48349 = ( n3825 & n8886 ) | ( n3825 & ~n20284 ) | ( n8886 & ~n20284 ) ;
  assign n48350 = ( n20109 & n38438 ) | ( n20109 & ~n48349 ) | ( n38438 & ~n48349 ) ;
  assign n48351 = ( ~n3094 & n8528 ) | ( ~n3094 & n48350 ) | ( n8528 & n48350 ) ;
  assign n48352 = ~n13145 & n36856 ;
  assign n48353 = ~n1487 & n48352 ;
  assign n48354 = ( ~n9662 & n34647 ) | ( ~n9662 & n48353 ) | ( n34647 & n48353 ) ;
  assign n48355 = ~n5734 & n8040 ;
  assign n48356 = ~n36635 & n38766 ;
  assign n48359 = n37757 ^ n32232 ^ n1924 ;
  assign n48360 = n48359 ^ n16450 ^ n15642 ;
  assign n48357 = ( n6570 & ~n10155 ) | ( n6570 & n10287 ) | ( ~n10155 & n10287 ) ;
  assign n48358 = n48357 ^ n12837 ^ n2589 ;
  assign n48361 = n48360 ^ n48358 ^ n28479 ;
  assign n48362 = n48361 ^ n5000 ^ 1'b0 ;
  assign n48363 = n48362 ^ n18626 ^ 1'b0 ;
  assign n48364 = n48356 | n48363 ;
  assign n48365 = n48364 ^ n22819 ^ n20361 ;
  assign n48366 = n24796 ^ n18652 ^ n4518 ;
  assign n48367 = n15909 ^ n13571 ^ 1'b0 ;
  assign n48368 = n48367 ^ n2727 ^ n2293 ;
  assign n48369 = ( n2182 & ~n48366 ) | ( n2182 & n48368 ) | ( ~n48366 & n48368 ) ;
  assign n48374 = n14618 ^ n10473 ^ n7387 ;
  assign n48370 = n7097 ^ n6137 ^ 1'b0 ;
  assign n48371 = n48370 ^ n22623 ^ n10971 ;
  assign n48372 = ( ~n6503 & n7180 ) | ( ~n6503 & n31685 ) | ( n7180 & n31685 ) ;
  assign n48373 = n48371 & n48372 ;
  assign n48375 = n48374 ^ n48373 ^ n17420 ;
  assign n48376 = n12497 & ~n46113 ;
  assign n48377 = n48376 ^ n11070 ^ 1'b0 ;
  assign n48378 = n12166 & n20373 ;
  assign n48379 = n34441 ^ n11970 ^ n5015 ;
  assign n48380 = n28694 ^ n2014 ^ 1'b0 ;
  assign n48381 = n24770 & ~n48380 ;
  assign n48382 = ( n14275 & ~n31783 ) | ( n14275 & n48381 ) | ( ~n31783 & n48381 ) ;
  assign n48383 = ( ~n4914 & n16565 ) | ( ~n4914 & n48382 ) | ( n16565 & n48382 ) ;
  assign n48384 = n44686 ^ n29181 ^ n331 ;
  assign n48385 = ( ~n34975 & n39278 ) | ( ~n34975 & n48384 ) | ( n39278 & n48384 ) ;
  assign n48386 = n48385 ^ n12951 ^ n1535 ;
  assign n48387 = ~n14768 & n45813 ;
  assign n48388 = n48387 ^ n15351 ^ n4077 ;
  assign n48389 = n48388 ^ n6777 ^ n2947 ;
  assign n48390 = ( n2943 & n5329 ) | ( n2943 & ~n13787 ) | ( n5329 & ~n13787 ) ;
  assign n48391 = n17541 | n28751 ;
  assign n48392 = n48391 ^ n11416 ^ n5899 ;
  assign n48393 = n869 | n8133 ;
  assign n48394 = ~n3862 & n16353 ;
  assign n48395 = n20137 & n48394 ;
  assign n48396 = ( ~n16480 & n32064 ) | ( ~n16480 & n48395 ) | ( n32064 & n48395 ) ;
  assign n48397 = n8567 ^ n4388 ^ 1'b0 ;
  assign n48398 = ~n2244 & n48397 ;
  assign n48399 = n14824 ^ n7666 ^ n1868 ;
  assign n48400 = ( n10037 & n29862 ) | ( n10037 & ~n39284 ) | ( n29862 & ~n39284 ) ;
  assign n48401 = n48399 & ~n48400 ;
  assign n48402 = ~n15088 & n48401 ;
  assign n48403 = n48402 ^ n32665 ^ 1'b0 ;
  assign n48404 = ( n5234 & ~n10697 ) | ( n5234 & n20722 ) | ( ~n10697 & n20722 ) ;
  assign n48405 = n46610 ^ n34054 ^ n8454 ;
  assign n48406 = ( n40664 & n48404 ) | ( n40664 & n48405 ) | ( n48404 & n48405 ) ;
  assign n48408 = ( ~n1224 & n3167 ) | ( ~n1224 & n14845 ) | ( n3167 & n14845 ) ;
  assign n48407 = n2728 & ~n7779 ;
  assign n48409 = n48408 ^ n48407 ^ n17391 ;
  assign n48410 = n13348 & n20200 ;
  assign n48411 = ( ~n4591 & n21289 ) | ( ~n4591 & n24751 ) | ( n21289 & n24751 ) ;
  assign n48412 = n32487 ^ n11004 ^ 1'b0 ;
  assign n48413 = n25230 | n29197 ;
  assign n48414 = n3402 & ~n6194 ;
  assign n48415 = n9222 & n48414 ;
  assign n48416 = n37939 ^ n1944 ^ 1'b0 ;
  assign n48417 = n39552 & n48416 ;
  assign n48418 = ( n9144 & n20742 ) | ( n9144 & ~n22175 ) | ( n20742 & ~n22175 ) ;
  assign n48419 = n48418 ^ n42114 ^ n9962 ;
  assign n48420 = ( n16725 & n40294 ) | ( n16725 & ~n48419 ) | ( n40294 & ~n48419 ) ;
  assign n48421 = n28143 ^ n21012 ^ n3361 ;
  assign n48422 = ~n8960 & n47018 ;
  assign n48426 = ( n13427 & n16926 ) | ( n13427 & ~n43259 ) | ( n16926 & ~n43259 ) ;
  assign n48424 = n20492 ^ n17479 ^ 1'b0 ;
  assign n48423 = n22628 ^ n8825 ^ n6505 ;
  assign n48425 = n48424 ^ n48423 ^ n6342 ;
  assign n48427 = n48426 ^ n48425 ^ n18326 ;
  assign n48428 = n39882 ^ n18292 ^ n1410 ;
  assign n48429 = ( n8803 & ~n12851 ) | ( n8803 & n29456 ) | ( ~n12851 & n29456 ) ;
  assign n48430 = n22084 ^ n11989 ^ 1'b0 ;
  assign n48431 = ( ~n4471 & n8934 ) | ( ~n4471 & n12375 ) | ( n8934 & n12375 ) ;
  assign n48432 = n48431 ^ n19315 ^ 1'b0 ;
  assign n48433 = n28964 | n48432 ;
  assign n48434 = n25694 ^ n19546 ^ n17814 ;
  assign n48435 = ( ~n48430 & n48433 ) | ( ~n48430 & n48434 ) | ( n48433 & n48434 ) ;
  assign n48436 = n48435 ^ n34842 ^ n17802 ;
  assign n48439 = ( n8606 & n25867 ) | ( n8606 & ~n28855 ) | ( n25867 & ~n28855 ) ;
  assign n48437 = n16611 ^ n8856 ^ n3327 ;
  assign n48438 = n27453 & ~n48437 ;
  assign n48440 = n48439 ^ n48438 ^ 1'b0 ;
  assign n48444 = n10770 & ~n22836 ;
  assign n48445 = n48444 ^ n8081 ^ 1'b0 ;
  assign n48441 = n14910 ^ n8157 ^ 1'b0 ;
  assign n48442 = ~n24544 & n48441 ;
  assign n48443 = ~n7312 & n48442 ;
  assign n48446 = n48445 ^ n48443 ^ 1'b0 ;
  assign n48447 = n31362 ^ n8054 ^ n7385 ;
  assign n48448 = n48447 ^ n21609 ^ n11940 ;
  assign n48449 = n48448 ^ n1326 ^ 1'b0 ;
  assign n48450 = n48449 ^ n672 ^ 1'b0 ;
  assign n48451 = ( ~n4551 & n16492 ) | ( ~n4551 & n16532 ) | ( n16492 & n16532 ) ;
  assign n48452 = n22854 & ~n30673 ;
  assign n48453 = ~n48451 & n48452 ;
  assign n48454 = n48453 ^ n33292 ^ n9937 ;
  assign n48455 = ( ~n23978 & n24115 ) | ( ~n23978 & n27552 ) | ( n24115 & n27552 ) ;
  assign n48456 = ( n25176 & n25421 ) | ( n25176 & n39824 ) | ( n25421 & n39824 ) ;
  assign n48457 = n17779 & n32689 ;
  assign n48458 = n48457 ^ n16017 ^ 1'b0 ;
  assign n48459 = ~n23112 & n48458 ;
  assign n48460 = n8893 & n48459 ;
  assign n48461 = n1886 & ~n13306 ;
  assign n48462 = n24653 & n48461 ;
  assign n48463 = n26498 ^ n20125 ^ n12629 ;
  assign n48464 = ( n13316 & n26740 ) | ( n13316 & ~n31353 ) | ( n26740 & ~n31353 ) ;
  assign n48465 = n48464 ^ n43598 ^ n38709 ;
  assign n48466 = n42967 ^ n3245 ^ n798 ;
  assign n48467 = ( n27856 & n33282 ) | ( n27856 & ~n48466 ) | ( n33282 & ~n48466 ) ;
  assign n48468 = n41337 ^ n27292 ^ x87 ;
  assign n48469 = n8223 ^ n7797 ^ 1'b0 ;
  assign n48470 = ~n7448 & n17208 ;
  assign n48471 = n48470 ^ n22271 ^ 1'b0 ;
  assign n48472 = ( n39333 & n48469 ) | ( n39333 & ~n48471 ) | ( n48469 & ~n48471 ) ;
  assign n48473 = n32328 & n40652 ;
  assign n48474 = n48473 ^ n8269 ^ 1'b0 ;
  assign n48475 = n37465 ^ n16977 ^ n6741 ;
  assign n48476 = n48475 ^ n44598 ^ n13637 ;
  assign n48477 = n4333 | n7029 ;
  assign n48478 = n48477 ^ n28496 ^ n17722 ;
  assign n48479 = n41263 ^ n33228 ^ n13587 ;
  assign n48480 = n26508 ^ n20855 ^ n5067 ;
  assign n48481 = ( n3910 & ~n17929 ) | ( n3910 & n48480 ) | ( ~n17929 & n48480 ) ;
  assign n48482 = n25561 ^ n18291 ^ n6295 ;
  assign n48483 = n37438 ^ n11329 ^ n10367 ;
  assign n48484 = n48483 ^ n32125 ^ 1'b0 ;
  assign n48486 = n44795 ^ n26130 ^ n10811 ;
  assign n48485 = n7301 | n26887 ;
  assign n48487 = n48486 ^ n48485 ^ 1'b0 ;
  assign n48488 = n37315 ^ n1846 ^ 1'b0 ;
  assign n48489 = n7401 & n48488 ;
  assign n48490 = n28585 ^ n5090 ^ 1'b0 ;
  assign n48491 = n48490 ^ n36559 ^ n32779 ;
  assign n48492 = n28920 ^ n5285 ^ n2290 ;
  assign n48493 = ( ~n3021 & n30352 ) | ( ~n3021 & n48492 ) | ( n30352 & n48492 ) ;
  assign n48494 = n35201 ^ n20437 ^ n12623 ;
  assign n48495 = ( ~n4637 & n29825 ) | ( ~n4637 & n43881 ) | ( n29825 & n43881 ) ;
  assign n48496 = n44554 ^ n1090 ^ 1'b0 ;
  assign n48499 = n26717 ^ n20735 ^ n11924 ;
  assign n48497 = n5420 & ~n5822 ;
  assign n48498 = n48497 ^ n26047 ^ n6998 ;
  assign n48500 = n48499 ^ n48498 ^ n19371 ;
  assign n48501 = ( n10562 & n26441 ) | ( n10562 & ~n40017 ) | ( n26441 & ~n40017 ) ;
  assign n48502 = n10541 ^ n6028 ^ 1'b0 ;
  assign n48503 = ( n11876 & n42431 ) | ( n11876 & n48502 ) | ( n42431 & n48502 ) ;
  assign n48504 = n2442 | n21699 ;
  assign n48505 = ~n7339 & n42750 ;
  assign n48506 = n27101 ^ n25404 ^ n6601 ;
  assign n48507 = ( n14716 & n21883 ) | ( n14716 & n25060 ) | ( n21883 & n25060 ) ;
  assign n48508 = ~n29760 & n48507 ;
  assign n48509 = n48506 & n48508 ;
  assign n48510 = n46303 ^ n37178 ^ n15879 ;
  assign n48511 = ( n4170 & n23157 ) | ( n4170 & ~n47041 ) | ( n23157 & ~n47041 ) ;
  assign n48512 = ( n469 & n4652 ) | ( n469 & ~n46944 ) | ( n4652 & ~n46944 ) ;
  assign n48513 = n48512 ^ n22399 ^ 1'b0 ;
  assign n48514 = n19404 & ~n20016 ;
  assign n48515 = n15168 ^ n10742 ^ x238 ;
  assign n48516 = n22772 | n48515 ;
  assign n48517 = n48516 ^ n1408 ^ 1'b0 ;
  assign n48518 = ( n34086 & n48514 ) | ( n34086 & ~n48517 ) | ( n48514 & ~n48517 ) ;
  assign n48519 = n48518 ^ n28666 ^ n27026 ;
  assign n48520 = n22506 ^ n15703 ^ n5285 ;
  assign n48521 = n5507 ^ x26 ^ 1'b0 ;
  assign n48522 = n48521 ^ n25326 ^ n17406 ;
  assign n48523 = n40482 & ~n48522 ;
  assign n48524 = ~n39478 & n48523 ;
  assign n48525 = ( n27144 & n48520 ) | ( n27144 & n48524 ) | ( n48520 & n48524 ) ;
  assign n48526 = n38672 ^ n6690 ^ 1'b0 ;
  assign n48527 = ~n12712 & n25260 ;
  assign n48528 = n265 | n41538 ;
  assign n48529 = n6998 ^ n6099 ^ n2834 ;
  assign n48530 = ( n24941 & n36453 ) | ( n24941 & n48529 ) | ( n36453 & n48529 ) ;
  assign n48531 = n5008 & n46131 ;
  assign n48532 = n48531 ^ n39421 ^ 1'b0 ;
  assign n48533 = n48532 ^ n33327 ^ n4856 ;
  assign n48534 = n41353 ^ n20920 ^ n13863 ;
  assign n48535 = ( ~n3849 & n12266 ) | ( ~n3849 & n13807 ) | ( n12266 & n13807 ) ;
  assign n48536 = ( n20101 & n26743 ) | ( n20101 & n48535 ) | ( n26743 & n48535 ) ;
  assign n48537 = ~n38758 & n47566 ;
  assign n48538 = n46314 & n48537 ;
  assign n48539 = n48538 ^ n33911 ^ 1'b0 ;
  assign n48540 = ( n27145 & ~n48536 ) | ( n27145 & n48539 ) | ( ~n48536 & n48539 ) ;
  assign n48541 = n20146 ^ n15155 ^ x239 ;
  assign n48542 = n48541 ^ n12565 ^ n1378 ;
  assign n48543 = ( n5084 & n23239 ) | ( n5084 & n47671 ) | ( n23239 & n47671 ) ;
  assign n48544 = ( n5021 & ~n13730 ) | ( n5021 & n37581 ) | ( ~n13730 & n37581 ) ;
  assign n48545 = n48544 ^ n40694 ^ n27636 ;
  assign n48546 = n44544 ^ n38979 ^ n9801 ;
  assign n48547 = n47499 | n48546 ;
  assign n48548 = n48547 ^ n40794 ^ 1'b0 ;
  assign n48549 = n9375 | n48548 ;
  assign n48550 = n48545 | n48549 ;
  assign n48551 = n48550 ^ n10392 ^ n10073 ;
  assign n48552 = n48551 ^ n14636 ^ 1'b0 ;
  assign n48553 = n39017 & ~n48552 ;
  assign n48554 = ~n6210 & n7514 ;
  assign n48555 = ~n31820 & n48554 ;
  assign n48556 = n44955 ^ n43743 ^ n28583 ;
  assign n48557 = n48556 ^ n34371 ^ n32474 ;
  assign n48558 = n48557 ^ n30329 ^ n6575 ;
  assign n48559 = n17028 | n18823 ;
  assign n48560 = n21210 | n48559 ;
  assign n48561 = n48560 ^ n44005 ^ n9392 ;
  assign n48562 = n48561 ^ n36284 ^ n2818 ;
  assign n48563 = ( n18856 & n24094 ) | ( n18856 & ~n28031 ) | ( n24094 & ~n28031 ) ;
  assign n48564 = n48563 ^ n43076 ^ n1705 ;
  assign n48565 = n9537 | n27345 ;
  assign n48566 = n48565 ^ n7798 ^ 1'b0 ;
  assign n48567 = n48566 ^ n15311 ^ 1'b0 ;
  assign n48568 = n24078 ^ n21373 ^ n18474 ;
  assign n48569 = ( n1431 & n7390 ) | ( n1431 & ~n40421 ) | ( n7390 & ~n40421 ) ;
  assign n48570 = n40092 ^ n17361 ^ n8464 ;
  assign n48571 = n6472 & n11794 ;
  assign n48572 = ( n40562 & n48570 ) | ( n40562 & n48571 ) | ( n48570 & n48571 ) ;
  assign n48573 = ( n29078 & ~n48569 ) | ( n29078 & n48572 ) | ( ~n48569 & n48572 ) ;
  assign n48574 = n48573 ^ n2564 ^ 1'b0 ;
  assign n48575 = n46524 ^ n19226 ^ 1'b0 ;
  assign n48576 = n48575 ^ n43271 ^ n10592 ;
  assign n48577 = n48576 ^ n42675 ^ n18250 ;
  assign n48578 = ~n12102 & n23543 ;
  assign n48579 = n38461 & n48578 ;
  assign n48580 = ( n2743 & ~n13460 ) | ( n2743 & n24834 ) | ( ~n13460 & n24834 ) ;
  assign n48581 = n48580 ^ n11019 ^ 1'b0 ;
  assign n48582 = ( n26951 & ~n39645 ) | ( n26951 & n47594 ) | ( ~n39645 & n47594 ) ;
  assign n48583 = n48582 ^ n7292 ^ 1'b0 ;
  assign n48584 = ( n11129 & ~n20893 ) | ( n11129 & n37390 ) | ( ~n20893 & n37390 ) ;
  assign n48585 = ( x199 & n3875 ) | ( x199 & n7062 ) | ( n3875 & n7062 ) ;
  assign n48586 = n10336 & ~n22271 ;
  assign n48587 = n48586 ^ n16268 ^ 1'b0 ;
  assign n48588 = ( n1511 & n12913 ) | ( n1511 & n48587 ) | ( n12913 & n48587 ) ;
  assign n48589 = ( ~n3306 & n8404 ) | ( ~n3306 & n9782 ) | ( n8404 & n9782 ) ;
  assign n48593 = n31792 ^ n23872 ^ 1'b0 ;
  assign n48590 = n27167 ^ n3029 ^ n1023 ;
  assign n48591 = n439 | n25680 ;
  assign n48592 = n48590 | n48591 ;
  assign n48594 = n48593 ^ n48592 ^ n28344 ;
  assign n48595 = n33207 | n45543 ;
  assign n48596 = ( n11592 & ~n12737 ) | ( n11592 & n20981 ) | ( ~n12737 & n20981 ) ;
  assign n48597 = n48596 ^ n22218 ^ 1'b0 ;
  assign n48598 = ~n31246 & n48597 ;
  assign n48605 = n39871 ^ n14616 ^ n8072 ;
  assign n48599 = n34910 ^ n13634 ^ 1'b0 ;
  assign n48600 = ~n6549 & n48599 ;
  assign n48601 = ~n12104 & n48600 ;
  assign n48602 = n48601 ^ n20175 ^ 1'b0 ;
  assign n48603 = ( n1146 & ~n15592 ) | ( n1146 & n48602 ) | ( ~n15592 & n48602 ) ;
  assign n48604 = ( n29130 & n34864 ) | ( n29130 & ~n48603 ) | ( n34864 & ~n48603 ) ;
  assign n48606 = n48605 ^ n48604 ^ n15405 ;
  assign n48607 = n36421 ^ n31997 ^ n7921 ;
  assign n48608 = n48607 ^ n33833 ^ n11435 ;
  assign n48614 = n37814 & n41326 ;
  assign n48609 = n16302 ^ n14295 ^ n372 ;
  assign n48610 = n48609 ^ n19907 ^ 1'b0 ;
  assign n48611 = n8352 & ~n48610 ;
  assign n48612 = n48611 ^ n16813 ^ 1'b0 ;
  assign n48613 = ~n15935 & n48612 ;
  assign n48615 = n48614 ^ n48613 ^ n30385 ;
  assign n48616 = ( ~n10998 & n15597 ) | ( ~n10998 & n47320 ) | ( n15597 & n47320 ) ;
  assign n48617 = ( ~n15378 & n23908 ) | ( ~n15378 & n31044 ) | ( n23908 & n31044 ) ;
  assign n48618 = ( n21176 & n44969 ) | ( n21176 & n48617 ) | ( n44969 & n48617 ) ;
  assign n48619 = ~n11453 & n20860 ;
  assign n48620 = n48619 ^ n14130 ^ 1'b0 ;
  assign n48621 = n31147 ^ n30358 ^ n19191 ;
  assign n48622 = n23874 & ~n48621 ;
  assign n48623 = n48622 ^ n11493 ^ 1'b0 ;
  assign n48624 = n7257 | n23813 ;
  assign n48625 = n48623 | n48624 ;
  assign n48626 = n18952 ^ n6718 ^ 1'b0 ;
  assign n48627 = n48626 ^ n28999 ^ n905 ;
  assign n48628 = n24934 ^ n19356 ^ 1'b0 ;
  assign n48629 = ~n5219 & n48628 ;
  assign n48630 = n48629 ^ n35256 ^ 1'b0 ;
  assign n48631 = ~n8796 & n11850 ;
  assign n48632 = ~n37589 & n48631 ;
  assign n48633 = ( ~n27693 & n46548 ) | ( ~n27693 & n48632 ) | ( n46548 & n48632 ) ;
  assign n48634 = n24664 ^ n18486 ^ n582 ;
  assign n48635 = n13612 ^ n10094 ^ n4064 ;
  assign n48636 = n48635 ^ n34822 ^ n30048 ;
  assign n48637 = n32177 ^ n28798 ^ n19881 ;
  assign n48638 = n35328 ^ n6106 ^ 1'b0 ;
  assign n48639 = n48638 ^ n19149 ^ n6606 ;
  assign n48640 = n48639 ^ n10170 ^ n4601 ;
  assign n48641 = n22356 ^ n628 ^ 1'b0 ;
  assign n48642 = ~n23840 & n48641 ;
  assign n48643 = n48642 ^ n15005 ^ n8258 ;
  assign n48644 = n48643 ^ n42857 ^ n18842 ;
  assign n48645 = n12315 & n36422 ;
  assign n48646 = n48645 ^ n20075 ^ 1'b0 ;
  assign n48647 = ( n22415 & n28568 ) | ( n22415 & n29419 ) | ( n28568 & n29419 ) ;
  assign n48648 = n29022 & ~n48647 ;
  assign n48649 = ( n565 & n2818 ) | ( n565 & ~n45772 ) | ( n2818 & ~n45772 ) ;
  assign n48650 = n17137 & ~n48649 ;
  assign n48651 = ( ~n13940 & n20491 ) | ( ~n13940 & n45575 ) | ( n20491 & n45575 ) ;
  assign n48652 = n46019 ^ n22513 ^ n17947 ;
  assign n48653 = n13387 | n19193 ;
  assign n48654 = ( ~n4807 & n36409 ) | ( ~n4807 & n48653 ) | ( n36409 & n48653 ) ;
  assign n48655 = n44063 ^ n40481 ^ 1'b0 ;
  assign n48656 = n19317 | n48655 ;
  assign n48657 = n25265 ^ n18746 ^ n8822 ;
  assign n48658 = ~n8307 & n38734 ;
  assign n48659 = ~n48657 & n48658 ;
  assign n48660 = n30796 ^ n307 ^ 1'b0 ;
  assign n48661 = n14557 & n48660 ;
  assign n48662 = ( n4277 & n17070 ) | ( n4277 & ~n39432 ) | ( n17070 & ~n39432 ) ;
  assign n48663 = n38499 ^ n17280 ^ n2717 ;
  assign n48664 = n48663 ^ n39685 ^ n27281 ;
  assign n48665 = ( n1844 & n2905 ) | ( n1844 & ~n33305 ) | ( n2905 & ~n33305 ) ;
  assign n48666 = n8004 ^ n7881 ^ 1'b0 ;
  assign n48667 = n48666 ^ n8990 ^ n3016 ;
  assign n48668 = n48667 ^ n18608 ^ n17080 ;
  assign n48669 = n48668 ^ n29597 ^ n4014 ;
  assign n48670 = ( n14922 & ~n29663 ) | ( n14922 & n38263 ) | ( ~n29663 & n38263 ) ;
  assign n48671 = ( n15646 & n40519 ) | ( n15646 & n48670 ) | ( n40519 & n48670 ) ;
  assign n48672 = n31684 ^ n25115 ^ n3835 ;
  assign n48673 = ( n23298 & n24024 ) | ( n23298 & n37937 ) | ( n24024 & n37937 ) ;
  assign n48674 = n18379 ^ n8632 ^ n1695 ;
  assign n48675 = n19555 & ~n48674 ;
  assign n48676 = ( n28401 & n48673 ) | ( n28401 & n48675 ) | ( n48673 & n48675 ) ;
  assign n48677 = ( ~n8905 & n18856 ) | ( ~n8905 & n24791 ) | ( n18856 & n24791 ) ;
  assign n48678 = n1523 & n48677 ;
  assign n48679 = n48678 ^ n25344 ^ 1'b0 ;
  assign n48680 = ~n15951 & n48679 ;
  assign n48683 = n18207 ^ n17368 ^ n9473 ;
  assign n48681 = n11261 ^ n6485 ^ n5094 ;
  assign n48682 = ( ~n27753 & n46210 ) | ( ~n27753 & n48681 ) | ( n46210 & n48681 ) ;
  assign n48684 = n48683 ^ n48682 ^ n28308 ;
  assign n48685 = n38530 ^ n36705 ^ n1453 ;
  assign n48686 = n13364 ^ n1432 ^ 1'b0 ;
  assign n48687 = n40036 ^ n7548 ^ n3798 ;
  assign n48688 = ( n10019 & n23773 ) | ( n10019 & n25705 ) | ( n23773 & n25705 ) ;
  assign n48689 = ( ~n38386 & n43453 ) | ( ~n38386 & n48688 ) | ( n43453 & n48688 ) ;
  assign n48690 = n16683 ^ n7573 ^ n1844 ;
  assign n48691 = ( n33483 & n42427 ) | ( n33483 & ~n48690 ) | ( n42427 & ~n48690 ) ;
  assign n48692 = ( n8933 & n11516 ) | ( n8933 & ~n21665 ) | ( n11516 & ~n21665 ) ;
  assign n48693 = ( n936 & ~n20635 ) | ( n936 & n48692 ) | ( ~n20635 & n48692 ) ;
  assign n48694 = ~n8685 & n48693 ;
  assign n48695 = n48694 ^ n10975 ^ 1'b0 ;
  assign n48696 = ( n13460 & n48691 ) | ( n13460 & n48695 ) | ( n48691 & n48695 ) ;
  assign n48697 = n29251 ^ n3186 ^ n2951 ;
  assign n48698 = n11411 ^ n6438 ^ 1'b0 ;
  assign n48699 = n48698 ^ n43627 ^ 1'b0 ;
  assign n48700 = ( n7732 & ~n48697 ) | ( n7732 & n48699 ) | ( ~n48697 & n48699 ) ;
  assign n48701 = ( ~n4233 & n7934 ) | ( ~n4233 & n20204 ) | ( n7934 & n20204 ) ;
  assign n48702 = n48701 ^ n42319 ^ 1'b0 ;
  assign n48703 = n9976 | n48702 ;
  assign n48704 = n15428 | n26818 ;
  assign n48705 = n40654 & ~n48704 ;
  assign n48706 = n37619 ^ n4646 ^ 1'b0 ;
  assign n48707 = ~n5080 & n48706 ;
  assign n48708 = n27989 ^ n3831 ^ x223 ;
  assign n48709 = ( n10115 & n42520 ) | ( n10115 & ~n48708 ) | ( n42520 & ~n48708 ) ;
  assign n48710 = n48709 ^ n47621 ^ n7563 ;
  assign n48711 = n48710 ^ n43563 ^ n19596 ;
  assign n48712 = ( n4990 & n12159 ) | ( n4990 & ~n16587 ) | ( n12159 & ~n16587 ) ;
  assign n48713 = n23864 ^ n15475 ^ 1'b0 ;
  assign n48714 = n31732 ^ n15895 ^ n12062 ;
  assign n48715 = n25404 & ~n29929 ;
  assign n48716 = n48715 ^ n11928 ^ 1'b0 ;
  assign n48718 = n45196 ^ n5210 ^ n842 ;
  assign n48717 = n8936 & n16117 ;
  assign n48719 = n48718 ^ n48717 ^ 1'b0 ;
  assign n48720 = n38972 ^ n24498 ^ n23473 ;
  assign n48721 = n41294 ^ n38036 ^ n8422 ;
  assign n48722 = n31338 & n33181 ;
  assign n48723 = n34821 & n48722 ;
  assign n48724 = ( n1979 & n23431 ) | ( n1979 & ~n48723 ) | ( n23431 & ~n48723 ) ;
  assign n48725 = ( n6074 & n16981 ) | ( n6074 & n22110 ) | ( n16981 & n22110 ) ;
  assign n48726 = ~n12934 & n16609 ;
  assign n48727 = n48726 ^ n35848 ^ 1'b0 ;
  assign n48728 = n20619 ^ n15563 ^ 1'b0 ;
  assign n48729 = n31484 | n48728 ;
  assign n48730 = n48729 ^ n7009 ^ n4300 ;
  assign n48731 = ( ~x215 & n5059 ) | ( ~x215 & n14351 ) | ( n5059 & n14351 ) ;
  assign n48732 = n32672 | n48731 ;
  assign n48733 = n48732 ^ n45354 ^ 1'b0 ;
  assign n48734 = n19231 & n38678 ;
  assign n48735 = ( n3431 & n28785 ) | ( n3431 & n47237 ) | ( n28785 & n47237 ) ;
  assign n48736 = ( ~n14385 & n14721 ) | ( ~n14385 & n39185 ) | ( n14721 & n39185 ) ;
  assign n48737 = n43595 ^ n10317 ^ n7319 ;
  assign n48738 = n48737 ^ n16613 ^ 1'b0 ;
  assign n48739 = n35128 ^ n11293 ^ n7458 ;
  assign n48740 = n48739 ^ n15463 ^ n7053 ;
  assign n48741 = n48740 ^ n37972 ^ n13367 ;
  assign n48742 = ( n893 & n3146 ) | ( n893 & n5215 ) | ( n3146 & n5215 ) ;
  assign n48743 = ( n12382 & n28871 ) | ( n12382 & ~n48742 ) | ( n28871 & ~n48742 ) ;
  assign n48744 = ( n31912 & n38632 ) | ( n31912 & n48743 ) | ( n38632 & n48743 ) ;
  assign n48745 = ~n5302 & n23925 ;
  assign n48746 = n48745 ^ n31704 ^ n15133 ;
  assign n48747 = n40447 ^ n7099 ^ n466 ;
  assign n48748 = n19490 & n48747 ;
  assign n48749 = ( n1315 & n7512 ) | ( n1315 & ~n48748 ) | ( n7512 & ~n48748 ) ;
  assign n48750 = n34413 ^ n2087 ^ 1'b0 ;
  assign n48751 = n27928 ^ n10559 ^ n10285 ;
  assign n48752 = n48751 ^ n32015 ^ n19922 ;
  assign n48753 = ( ~n689 & n15789 ) | ( ~n689 & n48752 ) | ( n15789 & n48752 ) ;
  assign n48754 = ~n31135 & n48753 ;
  assign n48755 = n48754 ^ n14628 ^ 1'b0 ;
  assign n48756 = n16778 ^ n4858 ^ 1'b0 ;
  assign n48757 = n48756 ^ n1352 ^ n654 ;
  assign n48758 = n36887 ^ n23473 ^ 1'b0 ;
  assign n48759 = ( ~n21377 & n48757 ) | ( ~n21377 & n48758 ) | ( n48757 & n48758 ) ;
  assign n48760 = n25208 ^ n18779 ^ n16269 ;
  assign n48761 = ( ~n25901 & n40916 ) | ( ~n25901 & n48760 ) | ( n40916 & n48760 ) ;
  assign n48762 = n12594 | n36943 ;
  assign n48763 = ( n14186 & ~n33918 ) | ( n14186 & n47774 ) | ( ~n33918 & n47774 ) ;
  assign n48764 = n48763 ^ n44583 ^ 1'b0 ;
  assign n48765 = ( n11349 & ~n19095 ) | ( n11349 & n48764 ) | ( ~n19095 & n48764 ) ;
  assign n48766 = n46343 ^ n31628 ^ 1'b0 ;
  assign n48767 = n9104 | n48766 ;
  assign n48768 = ~n48765 & n48767 ;
  assign n48769 = n38173 ^ n18037 ^ n9498 ;
  assign n48770 = n46058 ^ n8017 ^ 1'b0 ;
  assign n48771 = n12795 | n48770 ;
  assign n48772 = n23442 ^ n15550 ^ n868 ;
  assign n48773 = n48772 ^ n39992 ^ n27878 ;
  assign n48774 = n13630 ^ n1013 ^ 1'b0 ;
  assign n48775 = n30490 | n48774 ;
  assign n48776 = ( n22009 & n26094 ) | ( n22009 & n48775 ) | ( n26094 & n48775 ) ;
  assign n48777 = n13516 ^ n3417 ^ 1'b0 ;
  assign n48778 = n23503 & n48777 ;
  assign n48779 = ~n16809 & n48778 ;
  assign n48780 = n48779 ^ n44762 ^ 1'b0 ;
  assign n48781 = n48780 ^ n38208 ^ n16445 ;
  assign n48782 = n28752 ^ n17354 ^ 1'b0 ;
  assign n48783 = n39343 ^ n13241 ^ n2316 ;
  assign n48784 = ( n4581 & n27145 ) | ( n4581 & ~n36192 ) | ( n27145 & ~n36192 ) ;
  assign n48785 = n12909 | n16480 ;
  assign n48786 = n48785 ^ n27209 ^ 1'b0 ;
  assign n48787 = n7632 & ~n44928 ;
  assign n48788 = ~n17863 & n48787 ;
  assign n48789 = n48171 ^ n21124 ^ n5059 ;
  assign n48790 = ( n10461 & n25691 ) | ( n10461 & ~n48789 ) | ( n25691 & ~n48789 ) ;
  assign n48791 = n13187 | n24361 ;
  assign n48792 = n5215 | n48791 ;
  assign n48793 = n48792 ^ n15155 ^ n7837 ;
  assign n48794 = n31636 ^ n27030 ^ n5595 ;
  assign n48795 = ( n12892 & ~n31484 ) | ( n12892 & n32388 ) | ( ~n31484 & n32388 ) ;
  assign n48796 = n5528 & ~n13019 ;
  assign n48797 = ~n11178 & n48796 ;
  assign n48798 = ( n13916 & ~n27352 ) | ( n13916 & n40439 ) | ( ~n27352 & n40439 ) ;
  assign n48799 = ( n9437 & n48797 ) | ( n9437 & n48798 ) | ( n48797 & n48798 ) ;
  assign n48800 = n3190 ^ n1351 ^ n479 ;
  assign n48801 = n48800 ^ n26391 ^ 1'b0 ;
  assign n48802 = ( n959 & n10761 ) | ( n959 & ~n15938 ) | ( n10761 & ~n15938 ) ;
  assign n48803 = n48802 ^ n43356 ^ n28122 ;
  assign n48804 = ( ~n9475 & n47368 ) | ( ~n9475 & n48803 ) | ( n47368 & n48803 ) ;
  assign n48805 = ( n19855 & n48801 ) | ( n19855 & n48804 ) | ( n48801 & n48804 ) ;
  assign n48806 = n25475 ^ n16638 ^ 1'b0 ;
  assign n48807 = n48806 ^ n36151 ^ n18884 ;
  assign n48808 = n48807 ^ n9527 ^ n4761 ;
  assign n48809 = n9929 & ~n38416 ;
  assign n48810 = n48809 ^ n3236 ^ 1'b0 ;
  assign n48811 = n1953 ^ x246 ^ 1'b0 ;
  assign n48812 = ( n29935 & ~n31325 ) | ( n29935 & n31469 ) | ( ~n31325 & n31469 ) ;
  assign n48813 = n23757 ^ n15031 ^ 1'b0 ;
  assign n48814 = n47970 & ~n48813 ;
  assign n48815 = ( n48811 & n48812 ) | ( n48811 & ~n48814 ) | ( n48812 & ~n48814 ) ;
  assign n48816 = n23643 ^ n4784 ^ 1'b0 ;
  assign n48817 = n48816 ^ n5174 ^ 1'b0 ;
  assign n48818 = n29759 ^ n24089 ^ n14318 ;
  assign n48819 = n17322 ^ n2015 ^ 1'b0 ;
  assign n48820 = n48819 ^ n40680 ^ 1'b0 ;
  assign n48821 = n27655 ^ n14743 ^ n652 ;
  assign n48822 = n48821 ^ n34547 ^ n2962 ;
  assign n48823 = ( ~n12063 & n39394 ) | ( ~n12063 & n48822 ) | ( n39394 & n48822 ) ;
  assign n48824 = n38132 ^ n3400 ^ n2726 ;
  assign n48825 = ~n3064 & n16339 ;
  assign n48826 = n48825 ^ n36013 ^ n8901 ;
  assign n48827 = n16243 & n43621 ;
  assign n48828 = n48827 ^ n28307 ^ 1'b0 ;
  assign n48829 = n34672 ^ n33955 ^ n2923 ;
  assign n48830 = n19365 ^ n5686 ^ 1'b0 ;
  assign n48831 = n38040 & ~n48830 ;
  assign n48832 = n48831 ^ n9993 ^ n4124 ;
  assign n48833 = ~n12101 & n42083 ;
  assign n48834 = n48833 ^ n5323 ^ 1'b0 ;
  assign n48835 = n27043 & ~n48834 ;
  assign n48836 = n48835 ^ n28929 ^ 1'b0 ;
  assign n48837 = ( ~n22083 & n23356 ) | ( ~n22083 & n28197 ) | ( n23356 & n28197 ) ;
  assign n48838 = ( n33942 & n36324 ) | ( n33942 & ~n38150 ) | ( n36324 & ~n38150 ) ;
  assign n48839 = n39848 ^ n2976 ^ 1'b0 ;
  assign n48840 = n12206 & ~n25861 ;
  assign n48841 = ~n514 & n48840 ;
  assign n48842 = n47478 ^ x63 ^ 1'b0 ;
  assign n48843 = n3973 | n48842 ;
  assign n48844 = ( n2537 & ~n8915 ) | ( n2537 & n42878 ) | ( ~n8915 & n42878 ) ;
  assign n48845 = ( n1444 & ~n8896 ) | ( n1444 & n31092 ) | ( ~n8896 & n31092 ) ;
  assign n48846 = n48845 ^ n26806 ^ n18489 ;
  assign n48847 = n48846 ^ n3841 ^ n3259 ;
  assign n48848 = ( ~n2226 & n23737 ) | ( ~n2226 & n36068 ) | ( n23737 & n36068 ) ;
  assign n48849 = n19141 ^ n6845 ^ n1576 ;
  assign n48850 = ( ~n6087 & n33641 ) | ( ~n6087 & n48849 ) | ( n33641 & n48849 ) ;
  assign n48851 = n789 & n24025 ;
  assign n48852 = ~n21617 & n48851 ;
  assign n48853 = ( n41032 & n48850 ) | ( n41032 & ~n48852 ) | ( n48850 & ~n48852 ) ;
  assign n48854 = n36897 ^ n14588 ^ 1'b0 ;
  assign n48855 = n48854 ^ n34282 ^ n9058 ;
  assign n48856 = ( n24115 & n48165 ) | ( n24115 & ~n48855 ) | ( n48165 & ~n48855 ) ;
  assign n48857 = n38945 ^ n19839 ^ n7279 ;
  assign n48858 = ~n8427 & n20963 ;
  assign n48859 = n48858 ^ n38274 ^ n34016 ;
  assign n48860 = ( ~n13324 & n37338 ) | ( ~n13324 & n48859 ) | ( n37338 & n48859 ) ;
  assign n48861 = n19258 & ~n21229 ;
  assign n48862 = n48861 ^ n41945 ^ n18104 ;
  assign n48863 = n46867 ^ n15904 ^ n3433 ;
  assign n48864 = n38130 ^ n20781 ^ n18317 ;
  assign n48869 = n15303 ^ n6159 ^ n2325 ;
  assign n48867 = ( n2941 & ~n8773 ) | ( n2941 & n13501 ) | ( ~n8773 & n13501 ) ;
  assign n48865 = ( n3075 & n17063 ) | ( n3075 & n31260 ) | ( n17063 & n31260 ) ;
  assign n48866 = n48865 ^ n16202 ^ x102 ;
  assign n48868 = n48867 ^ n48866 ^ n1871 ;
  assign n48870 = n48869 ^ n48868 ^ n18602 ;
  assign n48871 = n18239 ^ n17714 ^ n2318 ;
  assign n48872 = ( n12063 & ~n19896 ) | ( n12063 & n48871 ) | ( ~n19896 & n48871 ) ;
  assign n48873 = n48872 ^ n37262 ^ n8652 ;
  assign n48874 = ( ~n19420 & n35490 ) | ( ~n19420 & n48873 ) | ( n35490 & n48873 ) ;
  assign n48875 = n6744 | n35395 ;
  assign n48876 = n32566 ^ n4117 ^ 1'b0 ;
  assign n48877 = ( n4876 & n16318 ) | ( n4876 & ~n30424 ) | ( n16318 & ~n30424 ) ;
  assign n48879 = ( n8808 & n11826 ) | ( n8808 & n20002 ) | ( n11826 & n20002 ) ;
  assign n48878 = n13530 | n26835 ;
  assign n48880 = n48879 ^ n48878 ^ 1'b0 ;
  assign n48881 = ( n14423 & n28120 ) | ( n14423 & ~n48880 ) | ( n28120 & ~n48880 ) ;
  assign n48882 = ( n2735 & n30684 ) | ( n2735 & ~n48881 ) | ( n30684 & ~n48881 ) ;
  assign n48883 = n25896 ^ n20427 ^ n6958 ;
  assign n48884 = n48883 ^ n5117 ^ 1'b0 ;
  assign n48885 = n31702 | n48884 ;
  assign n48886 = n15422 ^ n13663 ^ n4213 ;
  assign n48887 = n48886 ^ n37176 ^ n16285 ;
  assign n48888 = n21888 ^ n10613 ^ 1'b0 ;
  assign n48889 = ~n48887 & n48888 ;
  assign n48890 = n873 & ~n7078 ;
  assign n48891 = n48890 ^ n2248 ^ 1'b0 ;
  assign n48892 = n48891 ^ n27495 ^ n9143 ;
  assign n48893 = ( n14383 & n19078 ) | ( n14383 & ~n48892 ) | ( n19078 & ~n48892 ) ;
  assign n48894 = ( n3813 & n8772 ) | ( n3813 & n27428 ) | ( n8772 & n27428 ) ;
  assign n48895 = n47854 ^ n17345 ^ n946 ;
  assign n48896 = ( n29493 & ~n32722 ) | ( n29493 & n48895 ) | ( ~n32722 & n48895 ) ;
  assign n48897 = ( n14549 & n20731 ) | ( n14549 & n32203 ) | ( n20731 & n32203 ) ;
  assign n48898 = n48897 ^ n48181 ^ n15628 ;
  assign n48899 = ( n14716 & n18041 ) | ( n14716 & ~n41359 ) | ( n18041 & ~n41359 ) ;
  assign n48900 = n13167 ^ n9221 ^ n3545 ;
  assign n48901 = n48900 ^ n24449 ^ n6208 ;
  assign n48902 = ( ~n18704 & n19983 ) | ( ~n18704 & n26274 ) | ( n19983 & n26274 ) ;
  assign n48903 = n48902 ^ n44686 ^ n31665 ;
  assign n48904 = ( ~n11325 & n48901 ) | ( ~n11325 & n48903 ) | ( n48901 & n48903 ) ;
  assign n48905 = n10897 ^ n2824 ^ n1390 ;
  assign n48906 = n8615 ^ n6519 ^ 1'b0 ;
  assign n48907 = ~n6647 & n48906 ;
  assign n48908 = n48907 ^ n38550 ^ n12302 ;
  assign n48909 = ~n7933 & n48742 ;
  assign n48910 = n48909 ^ n1708 ^ 1'b0 ;
  assign n48911 = n24411 ^ n9135 ^ n2580 ;
  assign n48912 = n48911 ^ n44869 ^ 1'b0 ;
  assign n48913 = n48910 & n48912 ;
  assign n48914 = n27703 ^ n26740 ^ n22767 ;
  assign n48915 = n48914 ^ n39036 ^ 1'b0 ;
  assign n48916 = ( n8949 & n18941 ) | ( n8949 & ~n36128 ) | ( n18941 & ~n36128 ) ;
  assign n48917 = n48916 ^ n45133 ^ 1'b0 ;
  assign n48918 = ( n18716 & n22308 ) | ( n18716 & n36247 ) | ( n22308 & n36247 ) ;
  assign n48919 = n19735 ^ n7330 ^ n5022 ;
  assign n48920 = n15341 ^ n1246 ^ 1'b0 ;
  assign n48921 = n20213 ^ n2991 ^ 1'b0 ;
  assign n48922 = n48921 ^ n22224 ^ n20710 ;
  assign n48923 = ( ~n27017 & n48920 ) | ( ~n27017 & n48922 ) | ( n48920 & n48922 ) ;
  assign n48924 = n9199 & n15416 ;
  assign n48925 = n36723 & n48924 ;
  assign n48926 = ( n3405 & n24157 ) | ( n3405 & ~n48925 ) | ( n24157 & ~n48925 ) ;
  assign n48928 = ( n861 & ~n2185 ) | ( n861 & n16644 ) | ( ~n2185 & n16644 ) ;
  assign n48927 = ( n6811 & n14893 ) | ( n6811 & n36513 ) | ( n14893 & n36513 ) ;
  assign n48929 = n48928 ^ n48927 ^ n40561 ;
  assign n48930 = n41883 ^ n4249 ^ 1'b0 ;
  assign n48931 = n1942 & n48930 ;
  assign n48932 = n7577 & n45661 ;
  assign n48933 = ~n48931 & n48932 ;
  assign n48934 = ( n1552 & n1725 ) | ( n1552 & n3315 ) | ( n1725 & n3315 ) ;
  assign n48935 = n9789 | n48934 ;
  assign n48936 = n36996 ^ n6181 ^ 1'b0 ;
  assign n48937 = n12223 | n48936 ;
  assign n48938 = ( ~n19071 & n39851 ) | ( ~n19071 & n47094 ) | ( n39851 & n47094 ) ;
  assign n48939 = ( n9341 & n43104 ) | ( n9341 & n48938 ) | ( n43104 & n48938 ) ;
  assign n48940 = ~n13843 & n17883 ;
  assign n48941 = n48940 ^ n40089 ^ n4747 ;
  assign n48942 = n48521 ^ n21021 ^ n14579 ;
  assign n48943 = ( n1242 & n5997 ) | ( n1242 & ~n15484 ) | ( n5997 & ~n15484 ) ;
  assign n48944 = n48943 ^ n10390 ^ n1695 ;
  assign n48945 = ( n31922 & n45238 ) | ( n31922 & n48944 ) | ( n45238 & n48944 ) ;
  assign n48946 = n48945 ^ n46941 ^ n39303 ;
  assign n48947 = ( ~n8243 & n36425 ) | ( ~n8243 & n39734 ) | ( n36425 & n39734 ) ;
  assign n48948 = n22220 & ~n30351 ;
  assign n48949 = n16830 ^ n2332 ^ 1'b0 ;
  assign n48950 = n882 | n48949 ;
  assign n48951 = n48950 ^ n46675 ^ n15907 ;
  assign n48952 = n19301 & ~n48951 ;
  assign n48953 = ( ~n15325 & n25864 ) | ( ~n15325 & n34244 ) | ( n25864 & n34244 ) ;
  assign n48954 = ~n45910 & n48953 ;
  assign n48955 = n8980 & ~n26287 ;
  assign n48956 = ~n24647 & n48955 ;
  assign n48957 = ( ~n33073 & n40899 ) | ( ~n33073 & n41521 ) | ( n40899 & n41521 ) ;
  assign n48958 = ~n48956 & n48957 ;
  assign n48959 = n36503 ^ n9339 ^ n3837 ;
  assign n48960 = ( n22201 & n28031 ) | ( n22201 & n42861 ) | ( n28031 & n42861 ) ;
  assign n48961 = n420 & n48960 ;
  assign n48962 = n48959 & n48961 ;
  assign n48963 = n23074 ^ n11098 ^ 1'b0 ;
  assign n48964 = n34775 ^ n32125 ^ n6771 ;
  assign n48965 = n4943 ^ n1970 ^ n457 ;
  assign n48966 = n22825 ^ n14209 ^ n5531 ;
  assign n48967 = n48966 ^ n18391 ^ 1'b0 ;
  assign n48968 = n9822 & n48967 ;
  assign n48969 = ( ~n12841 & n22098 ) | ( ~n12841 & n48968 ) | ( n22098 & n48968 ) ;
  assign n48973 = ( n5477 & n5493 ) | ( n5477 & n22031 ) | ( n5493 & n22031 ) ;
  assign n48971 = n31931 & n35976 ;
  assign n48972 = ~n18594 & n48971 ;
  assign n48970 = ( n8900 & n23290 ) | ( n8900 & ~n44885 ) | ( n23290 & ~n44885 ) ;
  assign n48974 = n48973 ^ n48972 ^ n48970 ;
  assign n48975 = n4211 & ~n36963 ;
  assign n48976 = n48975 ^ n44484 ^ 1'b0 ;
  assign n48977 = n16997 ^ n13603 ^ n10311 ;
  assign n48978 = ( n45347 & n48976 ) | ( n45347 & n48977 ) | ( n48976 & n48977 ) ;
  assign n48979 = n48978 ^ n42396 ^ n37555 ;
  assign n48981 = n14765 ^ n3845 ^ n796 ;
  assign n48980 = n30524 & ~n32961 ;
  assign n48982 = n48981 ^ n48980 ^ 1'b0 ;
  assign n48983 = x154 & ~n48982 ;
  assign n48984 = ~n24224 & n48983 ;
  assign n48985 = n15616 ^ n9454 ^ 1'b0 ;
  assign n48986 = n19158 | n48985 ;
  assign n48987 = n31963 ^ n13048 ^ n10245 ;
  assign n48989 = ( n1181 & n14301 ) | ( n1181 & ~n34506 ) | ( n14301 & ~n34506 ) ;
  assign n48990 = ( n10433 & ~n13624 ) | ( n10433 & n48989 ) | ( ~n13624 & n48989 ) ;
  assign n48991 = ( ~n34596 & n35452 ) | ( ~n34596 & n48990 ) | ( n35452 & n48990 ) ;
  assign n48988 = n29949 ^ n18150 ^ n7246 ;
  assign n48992 = n48991 ^ n48988 ^ n45069 ;
  assign n48993 = ( n2707 & n5664 ) | ( n2707 & ~n21061 ) | ( n5664 & ~n21061 ) ;
  assign n48994 = ~n14170 & n30720 ;
  assign n48995 = ~n48993 & n48994 ;
  assign n48996 = n48995 ^ n42092 ^ n4327 ;
  assign n48997 = ~n20510 & n32854 ;
  assign n49000 = n47599 ^ n1850 ^ 1'b0 ;
  assign n49001 = n6954 & ~n20876 ;
  assign n49002 = n20445 & n49001 ;
  assign n49003 = ( n28191 & ~n36862 ) | ( n28191 & n49002 ) | ( ~n36862 & n49002 ) ;
  assign n49004 = ( n6886 & n49000 ) | ( n6886 & n49003 ) | ( n49000 & n49003 ) ;
  assign n48998 = n24645 ^ n20795 ^ n17048 ;
  assign n48999 = ( n24117 & ~n41364 ) | ( n24117 & n48998 ) | ( ~n41364 & n48998 ) ;
  assign n49005 = n49004 ^ n48999 ^ n17398 ;
  assign n49006 = ( n9853 & ~n23655 ) | ( n9853 & n46274 ) | ( ~n23655 & n46274 ) ;
  assign n49007 = n11182 & ~n43860 ;
  assign n49008 = n9303 & n49007 ;
  assign n49010 = ( n7277 & n24795 ) | ( n7277 & ~n30879 ) | ( n24795 & ~n30879 ) ;
  assign n49009 = n21543 & ~n33483 ;
  assign n49011 = n49010 ^ n49009 ^ 1'b0 ;
  assign n49012 = n38324 ^ n19225 ^ n6693 ;
  assign n49013 = ( ~n4894 & n47683 ) | ( ~n4894 & n49012 ) | ( n47683 & n49012 ) ;
  assign n49014 = n5223 | n8776 ;
  assign n49015 = n32394 | n49014 ;
  assign n49016 = n49015 ^ n35465 ^ n1669 ;
  assign n49017 = n47223 ^ n20750 ^ n12143 ;
  assign n49018 = ( n11926 & n12126 ) | ( n11926 & n26318 ) | ( n12126 & n26318 ) ;
  assign n49019 = n49018 ^ n17504 ^ n3004 ;
  assign n49020 = n10740 & n11619 ;
  assign n49021 = n26391 & n49020 ;
  assign n49022 = ( n20062 & n21387 ) | ( n20062 & n34669 ) | ( n21387 & n34669 ) ;
  assign n49023 = ( n24574 & ~n29038 ) | ( n24574 & n31982 ) | ( ~n29038 & n31982 ) ;
  assign n49024 = n49023 ^ n13050 ^ n12798 ;
  assign n49025 = ~n15846 & n48220 ;
  assign n49026 = ~n49024 & n49025 ;
  assign n49027 = ( ~n49021 & n49022 ) | ( ~n49021 & n49026 ) | ( n49022 & n49026 ) ;
  assign n49028 = n44574 ^ n1150 ^ 1'b0 ;
  assign n49029 = n49028 ^ n48178 ^ n8767 ;
  assign n49030 = ~n3309 & n7133 ;
  assign n49031 = ~n2538 & n49030 ;
  assign n49032 = n30188 & ~n40582 ;
  assign n49033 = n11773 & n49032 ;
  assign n49034 = n3944 | n45575 ;
  assign n49035 = n49034 ^ n14184 ^ 1'b0 ;
  assign n49037 = n9085 ^ n4378 ^ 1'b0 ;
  assign n49038 = n11604 ^ n6153 ^ 1'b0 ;
  assign n49039 = n49037 & ~n49038 ;
  assign n49040 = n49039 ^ n38916 ^ n21466 ;
  assign n49036 = ( n7029 & ~n26944 ) | ( n7029 & n40107 ) | ( ~n26944 & n40107 ) ;
  assign n49041 = n49040 ^ n49036 ^ n3004 ;
  assign n49042 = n45714 ^ n44170 ^ n26273 ;
  assign n49043 = n11048 ^ n9485 ^ n5370 ;
  assign n49044 = n12415 | n36024 ;
  assign n49045 = n49044 ^ n8716 ^ 1'b0 ;
  assign n49051 = n10778 ^ n1242 ^ 1'b0 ;
  assign n49052 = n6519 & ~n49051 ;
  assign n49050 = n23928 ^ n5584 ^ n2604 ;
  assign n49049 = ~n17285 & n19428 ;
  assign n49053 = n49052 ^ n49050 ^ n49049 ;
  assign n49046 = n14998 ^ n14398 ^ 1'b0 ;
  assign n49047 = n49046 ^ n19110 ^ 1'b0 ;
  assign n49048 = n48855 & n49047 ;
  assign n49054 = n49053 ^ n49048 ^ n26157 ;
  assign n49055 = ( n49043 & n49045 ) | ( n49043 & n49054 ) | ( n49045 & n49054 ) ;
  assign n49056 = n36400 ^ n33581 ^ n11041 ;
  assign n49057 = ( n3708 & n3754 ) | ( n3708 & n9278 ) | ( n3754 & n9278 ) ;
  assign n49058 = ( ~n7047 & n24330 ) | ( ~n7047 & n49057 ) | ( n24330 & n49057 ) ;
  assign n49059 = ( n27491 & n30487 ) | ( n27491 & n48217 ) | ( n30487 & n48217 ) ;
  assign n49060 = ( n4384 & ~n33658 ) | ( n4384 & n38808 ) | ( ~n33658 & n38808 ) ;
  assign n49062 = ( ~n1052 & n5772 ) | ( ~n1052 & n11906 ) | ( n5772 & n11906 ) ;
  assign n49061 = ( n2506 & ~n15750 ) | ( n2506 & n45298 ) | ( ~n15750 & n45298 ) ;
  assign n49063 = n49062 ^ n49061 ^ n25661 ;
  assign n49064 = ( n47780 & n49060 ) | ( n47780 & n49063 ) | ( n49060 & n49063 ) ;
  assign n49065 = n8419 & ~n31399 ;
  assign n49066 = n49065 ^ n38182 ^ n8517 ;
  assign n49067 = n6454 | n8423 ;
  assign n49068 = n27934 ^ n25761 ^ n10242 ;
  assign n49069 = ~n35179 & n49068 ;
  assign n49070 = ~n23504 & n28529 ;
  assign n49071 = ~n49069 & n49070 ;
  assign n49072 = ( ~n3131 & n8830 ) | ( ~n3131 & n18625 ) | ( n8830 & n18625 ) ;
  assign n49073 = n49072 ^ n44196 ^ n12667 ;
  assign n49074 = n49073 ^ n32323 ^ n1958 ;
  assign n49075 = ( n4371 & n4872 ) | ( n4371 & ~n20337 ) | ( n4872 & ~n20337 ) ;
  assign n49076 = ( n7896 & n16432 ) | ( n7896 & ~n49075 ) | ( n16432 & ~n49075 ) ;
  assign n49077 = ( n13002 & ~n21514 ) | ( n13002 & n47043 ) | ( ~n21514 & n47043 ) ;
  assign n49078 = n48617 ^ n45353 ^ n8834 ;
  assign n49079 = ( ~n1404 & n7187 ) | ( ~n1404 & n13158 ) | ( n7187 & n13158 ) ;
  assign n49080 = n1639 | n2206 ;
  assign n49081 = ( n4394 & n49079 ) | ( n4394 & n49080 ) | ( n49079 & n49080 ) ;
  assign n49082 = n34664 & n36146 ;
  assign n49083 = ~n36882 & n49082 ;
  assign n49084 = ( n20665 & n21610 ) | ( n20665 & ~n49083 ) | ( n21610 & ~n49083 ) ;
  assign n49085 = ( ~n2787 & n4155 ) | ( ~n2787 & n30187 ) | ( n4155 & n30187 ) ;
  assign n49086 = ~n849 & n8500 ;
  assign n49087 = n49086 ^ n17796 ^ 1'b0 ;
  assign n49088 = n5283 & n43831 ;
  assign n49089 = n19995 & n33705 ;
  assign n49090 = n49089 ^ n14535 ^ 1'b0 ;
  assign n49091 = ( n5461 & n7012 ) | ( n5461 & n49090 ) | ( n7012 & n49090 ) ;
  assign n49092 = ( ~n10290 & n16519 ) | ( ~n10290 & n49091 ) | ( n16519 & n49091 ) ;
  assign n49093 = n12334 ^ n6323 ^ n4493 ;
  assign n49095 = ( ~n315 & n26142 ) | ( ~n315 & n27503 ) | ( n26142 & n27503 ) ;
  assign n49094 = ~n16860 & n19877 ;
  assign n49096 = n49095 ^ n49094 ^ n16245 ;
  assign n49097 = n34644 ^ n8317 ^ 1'b0 ;
  assign n49101 = n31964 ^ n11281 ^ n2782 ;
  assign n49098 = n13613 ^ n10200 ^ n9022 ;
  assign n49099 = n49098 ^ n9231 ^ n7176 ;
  assign n49100 = ( ~n16780 & n40818 ) | ( ~n16780 & n49099 ) | ( n40818 & n49099 ) ;
  assign n49102 = n49101 ^ n49100 ^ n24053 ;
  assign n49103 = n49102 ^ n38590 ^ n4845 ;
  assign n49104 = n880 & n15286 ;
  assign n49105 = ~n4448 & n49104 ;
  assign n49106 = ( ~n8591 & n13983 ) | ( ~n8591 & n49105 ) | ( n13983 & n49105 ) ;
  assign n49107 = n31959 ^ n4764 ^ 1'b0 ;
  assign n49108 = n27191 & ~n49107 ;
  assign n49109 = ( n3134 & ~n49106 ) | ( n3134 & n49108 ) | ( ~n49106 & n49108 ) ;
  assign n49110 = n12338 ^ n2366 ^ 1'b0 ;
  assign n49111 = n47334 | n49110 ;
  assign n49112 = n25464 ^ n12452 ^ n5276 ;
  assign n49113 = n49112 ^ n20219 ^ 1'b0 ;
  assign n49114 = ( n9188 & ~n32072 ) | ( n9188 & n38239 ) | ( ~n32072 & n38239 ) ;
  assign n49115 = ( ~n12769 & n24022 ) | ( ~n12769 & n34351 ) | ( n24022 & n34351 ) ;
  assign n49118 = n29094 | n41477 ;
  assign n49116 = n2330 & ~n17954 ;
  assign n49117 = n19762 & n49116 ;
  assign n49119 = n49118 ^ n49117 ^ n9361 ;
  assign n49120 = ( n2052 & n11849 ) | ( n2052 & ~n26991 ) | ( n11849 & ~n26991 ) ;
  assign n49121 = ( n12056 & ~n47944 ) | ( n12056 & n49120 ) | ( ~n47944 & n49120 ) ;
  assign n49124 = n25961 ^ n17678 ^ 1'b0 ;
  assign n49125 = n3483 & ~n49124 ;
  assign n49122 = n37081 ^ n11754 ^ 1'b0 ;
  assign n49123 = n33283 & ~n49122 ;
  assign n49126 = n49125 ^ n49123 ^ n46556 ;
  assign n49127 = ( n7399 & n20373 ) | ( n7399 & ~n44335 ) | ( n20373 & ~n44335 ) ;
  assign n49128 = ( ~n3532 & n47837 ) | ( ~n3532 & n49127 ) | ( n47837 & n49127 ) ;
  assign n49130 = n4360 ^ n3908 ^ n3781 ;
  assign n49131 = ~n2219 & n49130 ;
  assign n49129 = ( n3216 & ~n5073 ) | ( n3216 & n44912 ) | ( ~n5073 & n44912 ) ;
  assign n49132 = n49131 ^ n49129 ^ n20508 ;
  assign n49133 = n49132 ^ n41684 ^ n5056 ;
  assign n49134 = ( n1056 & n7413 ) | ( n1056 & n23253 ) | ( n7413 & n23253 ) ;
  assign n49135 = ( n15724 & n26459 ) | ( n15724 & ~n49134 ) | ( n26459 & ~n49134 ) ;
  assign n49136 = n4143 | n18597 ;
  assign n49137 = n49136 ^ n25915 ^ 1'b0 ;
  assign n49138 = ~n545 & n33317 ;
  assign n49139 = n49137 & n49138 ;
  assign n49140 = n18959 ^ n8775 ^ n2456 ;
  assign n49141 = n11183 ^ n4854 ^ 1'b0 ;
  assign n49142 = ~n49140 & n49141 ;
  assign n49143 = n39960 ^ n17063 ^ n6224 ;
  assign n49144 = ( n9863 & ~n37709 ) | ( n9863 & n40449 ) | ( ~n37709 & n40449 ) ;
  assign n49145 = n49144 ^ n38789 ^ n12515 ;
  assign n49146 = n35011 ^ n32660 ^ n13313 ;
  assign n49147 = ( n4774 & ~n6445 ) | ( n4774 & n8688 ) | ( ~n6445 & n8688 ) ;
  assign n49148 = n49147 ^ n6232 ^ 1'b0 ;
  assign n49149 = ( ~n2931 & n8899 ) | ( ~n2931 & n23566 ) | ( n8899 & n23566 ) ;
  assign n49150 = n49149 ^ n3421 ^ n3296 ;
  assign n49151 = n1660 & n21627 ;
  assign n49152 = ~n24248 & n49151 ;
  assign n49153 = ( n16523 & n22110 ) | ( n16523 & ~n49152 ) | ( n22110 & ~n49152 ) ;
  assign n49154 = n14282 | n33621 ;
  assign n49155 = n49154 ^ n21449 ^ 1'b0 ;
  assign n49156 = n49155 ^ n15646 ^ n12751 ;
  assign n49157 = n42526 & ~n43213 ;
  assign n49158 = n38253 ^ n9881 ^ 1'b0 ;
  assign n49159 = n5056 & n49158 ;
  assign n49160 = n29807 ^ n22560 ^ n932 ;
  assign n49161 = ( n23494 & n32969 ) | ( n23494 & n49160 ) | ( n32969 & n49160 ) ;
  assign n49162 = n49161 ^ n3794 ^ 1'b0 ;
  assign n49163 = n4376 & ~n49162 ;
  assign n49164 = ( n5270 & ~n6098 ) | ( n5270 & n40591 ) | ( ~n6098 & n40591 ) ;
  assign n49168 = n24819 ^ n17426 ^ 1'b0 ;
  assign n49165 = ~n4404 & n4982 ;
  assign n49166 = n49165 ^ n3366 ^ 1'b0 ;
  assign n49167 = n49166 ^ n6155 ^ n3010 ;
  assign n49169 = n49168 ^ n49167 ^ n19362 ;
  assign n49170 = n11688 ^ n8985 ^ 1'b0 ;
  assign n49171 = n44257 & n49170 ;
  assign n49172 = ~n4166 & n49171 ;
  assign n49173 = n41683 ^ n34836 ^ n5840 ;
  assign n49174 = ( n5882 & n44617 ) | ( n5882 & ~n49173 ) | ( n44617 & ~n49173 ) ;
  assign n49175 = ( n41027 & ~n49172 ) | ( n41027 & n49174 ) | ( ~n49172 & n49174 ) ;
  assign n49176 = n15013 & n16488 ;
  assign n49177 = n49176 ^ n28571 ^ 1'b0 ;
  assign n49178 = ( n9604 & n17920 ) | ( n9604 & ~n49177 ) | ( n17920 & ~n49177 ) ;
  assign n49179 = ( ~n35605 & n38757 ) | ( ~n35605 & n45468 ) | ( n38757 & n45468 ) ;
  assign n49180 = n35387 & n46381 ;
  assign n49181 = n13322 & n15339 ;
  assign n49182 = n22725 & n49181 ;
  assign n49183 = ( n23505 & n29392 ) | ( n23505 & ~n49182 ) | ( n29392 & ~n49182 ) ;
  assign n49184 = ( n8724 & n46298 ) | ( n8724 & n49183 ) | ( n46298 & n49183 ) ;
  assign n49185 = n22780 & n27835 ;
  assign n49186 = n49185 ^ n18848 ^ 1'b0 ;
  assign n49188 = n12425 ^ n6485 ^ n3828 ;
  assign n49187 = ( ~n10112 & n10247 ) | ( ~n10112 & n29841 ) | ( n10247 & n29841 ) ;
  assign n49189 = n49188 ^ n49187 ^ n14567 ;
  assign n49190 = n49189 ^ n49173 ^ n20085 ;
  assign n49191 = n7805 & n14039 ;
  assign n49192 = n49191 ^ n18316 ^ 1'b0 ;
  assign n49193 = n1092 & ~n49192 ;
  assign n49194 = ( n5361 & n32945 ) | ( n5361 & n42732 ) | ( n32945 & n42732 ) ;
  assign n49195 = ( ~n9633 & n12825 ) | ( ~n9633 & n20354 ) | ( n12825 & n20354 ) ;
  assign n49196 = n29534 & ~n49195 ;
  assign n49197 = ~n44050 & n49196 ;
  assign n49198 = ( n21748 & ~n49194 ) | ( n21748 & n49197 ) | ( ~n49194 & n49197 ) ;
  assign n49199 = ( ~n8555 & n13685 ) | ( ~n8555 & n31051 ) | ( n13685 & n31051 ) ;
  assign n49200 = n49199 ^ n21431 ^ n12080 ;
  assign n49201 = n28294 ^ n12000 ^ n5317 ;
  assign n49202 = n49201 ^ n20756 ^ 1'b0 ;
  assign n49203 = n25140 & n44319 ;
  assign n49204 = ( ~n14374 & n25203 ) | ( ~n14374 & n47851 ) | ( n25203 & n47851 ) ;
  assign n49209 = ~n764 & n4565 ;
  assign n49210 = n1036 & n49209 ;
  assign n49207 = n19093 ^ n11293 ^ 1'b0 ;
  assign n49208 = n21798 | n49207 ;
  assign n49205 = ~n25615 & n26882 ;
  assign n49206 = n49205 ^ n29306 ^ 1'b0 ;
  assign n49211 = n49210 ^ n49208 ^ n49206 ;
  assign n49213 = n39868 ^ n34115 ^ n624 ;
  assign n49212 = n43662 ^ n39850 ^ n4853 ;
  assign n49214 = n49213 ^ n49212 ^ 1'b0 ;
  assign n49219 = n28154 & ~n35656 ;
  assign n49215 = n19921 ^ n9137 ^ n3181 ;
  assign n49216 = ( ~n13345 & n36872 ) | ( ~n13345 & n49215 ) | ( n36872 & n49215 ) ;
  assign n49217 = n6607 & ~n49216 ;
  assign n49218 = n49217 ^ n28764 ^ 1'b0 ;
  assign n49220 = n49219 ^ n49218 ^ n30451 ;
  assign n49222 = n7973 | n16573 ;
  assign n49223 = n49222 ^ n33620 ^ 1'b0 ;
  assign n49224 = n11374 ^ n2597 ^ 1'b0 ;
  assign n49225 = ( n29272 & n49223 ) | ( n29272 & n49224 ) | ( n49223 & n49224 ) ;
  assign n49221 = ( ~n32264 & n35033 ) | ( ~n32264 & n48858 ) | ( n35033 & n48858 ) ;
  assign n49226 = n49225 ^ n49221 ^ n22950 ;
  assign n49227 = ( ~n28669 & n29995 ) | ( ~n28669 & n32416 ) | ( n29995 & n32416 ) ;
  assign n49228 = n9429 & ~n47944 ;
  assign n49229 = n27223 ^ n5684 ^ 1'b0 ;
  assign n49230 = x138 & n49229 ;
  assign n49231 = n31496 ^ n8910 ^ n6201 ;
  assign n49232 = n49230 & ~n49231 ;
  assign n49233 = n47031 ^ n26767 ^ 1'b0 ;
  assign n49234 = n5591 & n49233 ;
  assign n49235 = n42559 ^ n13997 ^ n11846 ;
  assign n49236 = n32185 ^ n31530 ^ n9958 ;
  assign n49237 = n41127 ^ n29372 ^ n3654 ;
  assign n49238 = n26371 ^ n7789 ^ 1'b0 ;
  assign n49239 = n49238 ^ n33363 ^ n2880 ;
  assign n49240 = n49239 ^ n39287 ^ n36047 ;
  assign n49241 = n31034 ^ n17232 ^ n7408 ;
  assign n49242 = n22050 ^ n19545 ^ n8794 ;
  assign n49243 = ( n11549 & n49241 ) | ( n11549 & ~n49242 ) | ( n49241 & ~n49242 ) ;
  assign n49244 = n49243 ^ n35746 ^ n10397 ;
  assign n49245 = n9500 & ~n17989 ;
  assign n49246 = n49245 ^ n12259 ^ n1669 ;
  assign n49247 = ( n18096 & n23496 ) | ( n18096 & n33147 ) | ( n23496 & n33147 ) ;
  assign n49248 = n22480 | n42778 ;
  assign n49249 = n49248 ^ n45717 ^ 1'b0 ;
  assign n49250 = n6528 | n17640 ;
  assign n49251 = n33436 & ~n49250 ;
  assign n49252 = n16850 & n24463 ;
  assign n49253 = ~n13132 & n49252 ;
  assign n49254 = ( n6361 & n44022 ) | ( n6361 & ~n49253 ) | ( n44022 & ~n49253 ) ;
  assign n49255 = n31771 & n49254 ;
  assign n49256 = n49255 ^ n15115 ^ 1'b0 ;
  assign n49257 = ( n28808 & n37761 ) | ( n28808 & ~n41608 ) | ( n37761 & ~n41608 ) ;
  assign n49258 = n47123 ^ n46225 ^ n3592 ;
  assign n49259 = n23171 ^ n8638 ^ n7749 ;
  assign n49260 = ( n3376 & n6120 ) | ( n3376 & n49259 ) | ( n6120 & n49259 ) ;
  assign n49261 = n43213 ^ n6739 ^ 1'b0 ;
  assign n49262 = n49261 ^ n16287 ^ n952 ;
  assign n49263 = ( n6891 & n6905 ) | ( n6891 & ~n12278 ) | ( n6905 & ~n12278 ) ;
  assign n49264 = ( n621 & ~n770 ) | ( n621 & n49263 ) | ( ~n770 & n49263 ) ;
  assign n49265 = n23265 | n49264 ;
  assign n49266 = n1766 | n49265 ;
  assign n49267 = ( n3464 & n41436 ) | ( n3464 & ~n49266 ) | ( n41436 & ~n49266 ) ;
  assign n49268 = ( n19961 & ~n49262 ) | ( n19961 & n49267 ) | ( ~n49262 & n49267 ) ;
  assign n49269 = n49268 ^ n31181 ^ n17686 ;
  assign n49270 = n43417 ^ n43029 ^ n9086 ;
  assign n49271 = ( ~n18740 & n30777 ) | ( ~n18740 & n49270 ) | ( n30777 & n49270 ) ;
  assign n49272 = n12247 & n19500 ;
  assign n49273 = n49272 ^ n36632 ^ 1'b0 ;
  assign n49274 = ( ~n10515 & n49271 ) | ( ~n10515 & n49273 ) | ( n49271 & n49273 ) ;
  assign n49275 = ( n3541 & n6952 ) | ( n3541 & ~n19235 ) | ( n6952 & ~n19235 ) ;
  assign n49276 = n3146 | n7565 ;
  assign n49277 = n49276 ^ n34056 ^ 1'b0 ;
  assign n49278 = n49277 ^ n33276 ^ 1'b0 ;
  assign n49279 = n49278 ^ n42303 ^ n7026 ;
  assign n49280 = n2857 & ~n34576 ;
  assign n49281 = n49280 ^ n3096 ^ 1'b0 ;
  assign n49282 = n8707 ^ n5752 ^ n2065 ;
  assign n49283 = ( n41094 & ~n49281 ) | ( n41094 & n49282 ) | ( ~n49281 & n49282 ) ;
  assign n49284 = ( n13909 & n21311 ) | ( n13909 & n49283 ) | ( n21311 & n49283 ) ;
  assign n49285 = n49284 ^ n13242 ^ 1'b0 ;
  assign n49286 = n38450 & n49285 ;
  assign n49287 = ( ~n2884 & n13455 ) | ( ~n2884 & n31678 ) | ( n13455 & n31678 ) ;
  assign n49288 = ( n10963 & n20767 ) | ( n10963 & ~n49287 ) | ( n20767 & ~n49287 ) ;
  assign n49289 = ( ~n11458 & n33641 ) | ( ~n11458 & n49288 ) | ( n33641 & n49288 ) ;
  assign n49293 = ( n30478 & ~n31498 ) | ( n30478 & n38213 ) | ( ~n31498 & n38213 ) ;
  assign n49292 = n12776 ^ n6745 ^ n3969 ;
  assign n49294 = n49293 ^ n49292 ^ n9425 ;
  assign n49291 = n21470 ^ n4589 ^ n2531 ;
  assign n49290 = n42366 ^ n27951 ^ n21656 ;
  assign n49295 = n49294 ^ n49291 ^ n49290 ;
  assign n49296 = n5559 ^ n1575 ^ n939 ;
  assign n49297 = n37129 & n42220 ;
  assign n49298 = n36421 ^ n7888 ^ 1'b0 ;
  assign n49299 = ( ~n45101 & n49297 ) | ( ~n45101 & n49298 ) | ( n49297 & n49298 ) ;
  assign n49300 = ( n31489 & n42215 ) | ( n31489 & ~n49299 ) | ( n42215 & ~n49299 ) ;
  assign n49305 = n33291 ^ n25842 ^ n12074 ;
  assign n49301 = n24551 & n28021 ;
  assign n49302 = ~n17501 & n49301 ;
  assign n49303 = n49302 ^ n32897 ^ n10037 ;
  assign n49304 = n49303 ^ n19914 ^ n801 ;
  assign n49306 = n49305 ^ n49304 ^ n12129 ;
  assign n49308 = n26160 ^ n7271 ^ n2877 ;
  assign n49309 = ( n5894 & n12840 ) | ( n5894 & ~n26460 ) | ( n12840 & ~n26460 ) ;
  assign n49310 = ( n16041 & n49308 ) | ( n16041 & ~n49309 ) | ( n49308 & ~n49309 ) ;
  assign n49307 = n4588 & n29203 ;
  assign n49311 = n49310 ^ n49307 ^ 1'b0 ;
  assign n49312 = ( n5497 & n29931 ) | ( n5497 & ~n49311 ) | ( n29931 & ~n49311 ) ;
  assign n49317 = n36352 ^ n11954 ^ n11188 ;
  assign n49313 = n12318 ^ n7044 ^ n4432 ;
  assign n49314 = n15296 & ~n25069 ;
  assign n49315 = ~n49313 & n49314 ;
  assign n49316 = n49315 ^ n16535 ^ 1'b0 ;
  assign n49318 = n49317 ^ n49316 ^ n46747 ;
  assign n49319 = n37698 ^ n31085 ^ n4992 ;
  assign n49320 = n49319 ^ n6092 ^ 1'b0 ;
  assign n49321 = ~n9741 & n49320 ;
  assign n49322 = n19967 ^ n13630 ^ n1831 ;
  assign n49323 = n49322 ^ n2199 ^ 1'b0 ;
  assign n49324 = ~n16311 & n49323 ;
  assign n49325 = ( n6223 & n7659 ) | ( n6223 & ~n21689 ) | ( n7659 & ~n21689 ) ;
  assign n49326 = n5307 & n49325 ;
  assign n49327 = n19067 & n49326 ;
  assign n49328 = n49327 ^ n40000 ^ 1'b0 ;
  assign n49329 = n14324 ^ n7165 ^ 1'b0 ;
  assign n49330 = ( n12611 & n20822 ) | ( n12611 & n49329 ) | ( n20822 & n49329 ) ;
  assign n49331 = n49330 ^ n16321 ^ n15030 ;
  assign n49332 = ( n353 & n15810 ) | ( n353 & n25939 ) | ( n15810 & n25939 ) ;
  assign n49334 = n776 & n6069 ;
  assign n49335 = n49334 ^ n17026 ^ 1'b0 ;
  assign n49333 = n27497 ^ n22615 ^ n318 ;
  assign n49336 = n49335 ^ n49333 ^ n22565 ;
  assign n49337 = n10276 ^ n1599 ^ n639 ;
  assign n49338 = n49337 ^ n45632 ^ n292 ;
  assign n49339 = n31775 ^ n21487 ^ n7474 ;
  assign n49340 = n49339 ^ n48780 ^ 1'b0 ;
  assign n49342 = n13658 ^ n13561 ^ n867 ;
  assign n49341 = n41082 ^ n34887 ^ n21947 ;
  assign n49343 = n49342 ^ n49341 ^ n4283 ;
  assign n49344 = n42375 ^ n41881 ^ n31884 ;
  assign n49345 = n6349 & ~n43319 ;
  assign n49346 = ~n32591 & n49345 ;
  assign n49347 = n19858 ^ n10094 ^ 1'b0 ;
  assign n49348 = n8077 & ~n49347 ;
  assign n49349 = ( n3652 & ~n18984 ) | ( n3652 & n49348 ) | ( ~n18984 & n49348 ) ;
  assign n49350 = ( ~n5904 & n21151 ) | ( ~n5904 & n35092 ) | ( n21151 & n35092 ) ;
  assign n49351 = n7953 | n33806 ;
  assign n49352 = n25110 | n49351 ;
  assign n49353 = ( n7437 & n49350 ) | ( n7437 & ~n49352 ) | ( n49350 & ~n49352 ) ;
  assign n49354 = n20276 ^ n1106 ^ 1'b0 ;
  assign n49355 = n27977 ^ n2063 ^ n297 ;
  assign n49356 = ( ~n7871 & n9713 ) | ( ~n7871 & n29099 ) | ( n9713 & n29099 ) ;
  assign n49357 = n32595 & n49356 ;
  assign n49358 = ( n2605 & n49355 ) | ( n2605 & n49357 ) | ( n49355 & n49357 ) ;
  assign n49359 = n32460 ^ n7898 ^ 1'b0 ;
  assign n49360 = n49359 ^ n26891 ^ n13612 ;
  assign n49361 = n49360 ^ n31890 ^ n15338 ;
  assign n49362 = n37122 ^ n18852 ^ n14650 ;
  assign n49363 = n49362 ^ n45902 ^ n44019 ;
  assign n49364 = ~n11743 & n21526 ;
  assign n49365 = n39282 ^ n29151 ^ 1'b0 ;
  assign n49366 = ( n8251 & ~n43043 ) | ( n8251 & n43051 ) | ( ~n43043 & n43051 ) ;
  assign n49367 = n47537 ^ n5705 ^ 1'b0 ;
  assign n49370 = n14106 ^ n11168 ^ 1'b0 ;
  assign n49371 = n18350 & ~n49370 ;
  assign n49368 = ( n4739 & n5048 ) | ( n4739 & ~n12423 ) | ( n5048 & ~n12423 ) ;
  assign n49369 = n49368 ^ n34588 ^ n25026 ;
  assign n49372 = n49371 ^ n49369 ^ n44969 ;
  assign n49373 = n40578 ^ n37617 ^ n7578 ;
  assign n49374 = n18397 | n21040 ;
  assign n49375 = n49374 ^ n14076 ^ 1'b0 ;
  assign n49376 = n49375 ^ n10613 ^ n8398 ;
  assign n49377 = n49376 ^ n38017 ^ n16881 ;
  assign n49378 = ~n14495 & n49377 ;
  assign n49379 = n40010 ^ n37175 ^ n7248 ;
  assign n49380 = ( n20338 & n47168 ) | ( n20338 & n49379 ) | ( n47168 & n49379 ) ;
  assign n49381 = n49195 ^ n9100 ^ n368 ;
  assign n49382 = ( ~n1665 & n20182 ) | ( ~n1665 & n49381 ) | ( n20182 & n49381 ) ;
  assign n49383 = n11999 & n33189 ;
  assign n49384 = n25117 & n33163 ;
  assign n49385 = n49384 ^ n16839 ^ 1'b0 ;
  assign n49386 = n4503 ^ n264 ^ 1'b0 ;
  assign n49387 = ( n1920 & ~n11935 ) | ( n1920 & n22094 ) | ( ~n11935 & n22094 ) ;
  assign n49388 = n44061 ^ n19009 ^ 1'b0 ;
  assign n49389 = n41063 ^ n25730 ^ 1'b0 ;
  assign n49390 = n10161 & n49389 ;
  assign n49391 = n32656 ^ n12269 ^ n10048 ;
  assign n49392 = ( ~n23246 & n31795 ) | ( ~n23246 & n36333 ) | ( n31795 & n36333 ) ;
  assign n49394 = ( n5722 & ~n12984 ) | ( n5722 & n14347 ) | ( ~n12984 & n14347 ) ;
  assign n49395 = ( n3294 & n13931 ) | ( n3294 & n49394 ) | ( n13931 & n49394 ) ;
  assign n49393 = n7505 | n47984 ;
  assign n49396 = n49395 ^ n49393 ^ 1'b0 ;
  assign n49397 = n28533 ^ n21945 ^ 1'b0 ;
  assign n49398 = n14084 & ~n49397 ;
  assign n49399 = ( n17518 & ~n21232 ) | ( n17518 & n22685 ) | ( ~n21232 & n22685 ) ;
  assign n49400 = ( n9303 & n28847 ) | ( n9303 & ~n49399 ) | ( n28847 & ~n49399 ) ;
  assign n49401 = n49400 ^ n319 ^ 1'b0 ;
  assign n49402 = n38285 ^ n14382 ^ n10259 ;
  assign n49403 = n37203 & ~n49402 ;
  assign n49404 = n37026 ^ n31872 ^ n23893 ;
  assign n49405 = n34119 & n49404 ;
  assign n49406 = ( n25176 & n45487 ) | ( n25176 & ~n49405 ) | ( n45487 & ~n49405 ) ;
  assign n49407 = ( n4404 & n29622 ) | ( n4404 & ~n32206 ) | ( n29622 & ~n32206 ) ;
  assign n49408 = n49407 ^ n22996 ^ 1'b0 ;
  assign n49416 = n22736 ^ n13007 ^ 1'b0 ;
  assign n49413 = ( n6665 & n7478 ) | ( n6665 & ~n9983 ) | ( n7478 & ~n9983 ) ;
  assign n49414 = n49413 ^ n8080 ^ n5409 ;
  assign n49411 = ~n1857 & n23390 ;
  assign n49410 = n2251 & n2945 ;
  assign n49412 = n49411 ^ n49410 ^ n13878 ;
  assign n49415 = n49414 ^ n49412 ^ n15190 ;
  assign n49409 = ( n18574 & ~n42445 ) | ( n18574 & n48434 ) | ( ~n42445 & n48434 ) ;
  assign n49417 = n49416 ^ n49415 ^ n49409 ;
  assign n49418 = ~n8660 & n27046 ;
  assign n49419 = n23162 & n49418 ;
  assign n49420 = ( n17218 & ~n21876 ) | ( n17218 & n27516 ) | ( ~n21876 & n27516 ) ;
  assign n49421 = ( n19098 & n35892 ) | ( n19098 & ~n49420 ) | ( n35892 & ~n49420 ) ;
  assign n49422 = n49421 ^ n39039 ^ n21271 ;
  assign n49423 = n21592 | n38244 ;
  assign n49424 = n49422 & ~n49423 ;
  assign n49425 = n25350 ^ n12516 ^ 1'b0 ;
  assign n49426 = ( n8230 & ~n10589 ) | ( n8230 & n26506 ) | ( ~n10589 & n26506 ) ;
  assign n49427 = ( n2493 & n5649 ) | ( n2493 & ~n49426 ) | ( n5649 & ~n49426 ) ;
  assign n49428 = ( ~n3863 & n12758 ) | ( ~n3863 & n49427 ) | ( n12758 & n49427 ) ;
  assign n49429 = ( n36362 & n41439 ) | ( n36362 & ~n49428 ) | ( n41439 & ~n49428 ) ;
  assign n49430 = ~n34259 & n40394 ;
  assign n49431 = n42580 ^ n11912 ^ n5988 ;
  assign n49432 = n12321 & n44635 ;
  assign n49433 = ( n3132 & ~n6852 ) | ( n3132 & n49432 ) | ( ~n6852 & n49432 ) ;
  assign n49434 = n1816 ^ n1715 ^ 1'b0 ;
  assign n49435 = n12106 & ~n19426 ;
  assign n49436 = n49435 ^ n5672 ^ 1'b0 ;
  assign n49437 = ( ~n13123 & n22795 ) | ( ~n13123 & n49436 ) | ( n22795 & n49436 ) ;
  assign n49438 = n49437 ^ n16467 ^ n12708 ;
  assign n49439 = ( n893 & ~n12372 ) | ( n893 & n16867 ) | ( ~n12372 & n16867 ) ;
  assign n49440 = n49439 ^ n15554 ^ 1'b0 ;
  assign n49441 = n49440 ^ n35881 ^ n761 ;
  assign n49444 = ( ~n24108 & n33481 ) | ( ~n24108 & n40044 ) | ( n33481 & n40044 ) ;
  assign n49445 = n16149 ^ n14296 ^ 1'b0 ;
  assign n49446 = n49444 & n49445 ;
  assign n49442 = ( ~n19255 & n23520 ) | ( ~n19255 & n26374 ) | ( n23520 & n26374 ) ;
  assign n49443 = n42046 & n49442 ;
  assign n49447 = n49446 ^ n49443 ^ 1'b0 ;
  assign n49448 = n13266 | n26150 ;
  assign n49449 = n4866 & ~n49448 ;
  assign n49450 = n4781 & ~n31433 ;
  assign n49451 = n49450 ^ n38418 ^ 1'b0 ;
  assign n49452 = ( n30912 & ~n32765 ) | ( n30912 & n34003 ) | ( ~n32765 & n34003 ) ;
  assign n49458 = ( n8669 & n14459 ) | ( n8669 & n38932 ) | ( n14459 & n38932 ) ;
  assign n49453 = ( n2440 & n36324 ) | ( n2440 & ~n48522 ) | ( n36324 & ~n48522 ) ;
  assign n49454 = n16712 ^ x44 ^ 1'b0 ;
  assign n49455 = n49453 & ~n49454 ;
  assign n49456 = ( n30830 & ~n32517 ) | ( n30830 & n49455 ) | ( ~n32517 & n49455 ) ;
  assign n49457 = n49456 ^ n19571 ^ n17477 ;
  assign n49459 = n49458 ^ n49457 ^ 1'b0 ;
  assign n49460 = n37666 ^ n28388 ^ n9235 ;
  assign n49461 = n49460 ^ n37215 ^ n2828 ;
  assign n49462 = n49461 ^ n23988 ^ n5340 ;
  assign n49463 = ( n18185 & n26659 ) | ( n18185 & ~n39736 ) | ( n26659 & ~n39736 ) ;
  assign n49464 = n25105 ^ n24559 ^ n19966 ;
  assign n49465 = n35194 ^ n4487 ^ 1'b0 ;
  assign n49466 = n23054 | n45296 ;
  assign n49467 = n49466 ^ n8429 ^ 1'b0 ;
  assign n49468 = n308 & n26370 ;
  assign n49469 = n49468 ^ n12797 ^ 1'b0 ;
  assign n49470 = n7190 & n31588 ;
  assign n49471 = n17028 ^ n5910 ^ 1'b0 ;
  assign n49472 = ( n5980 & ~n8179 ) | ( n5980 & n9057 ) | ( ~n8179 & n9057 ) ;
  assign n49473 = n49472 ^ n12288 ^ n3925 ;
  assign n49474 = n14685 ^ n7992 ^ n642 ;
  assign n49475 = n49474 ^ n13189 ^ n3941 ;
  assign n49476 = n22904 ^ n17808 ^ n11743 ;
  assign n49477 = ( ~n8740 & n49475 ) | ( ~n8740 & n49476 ) | ( n49475 & n49476 ) ;
  assign n49478 = n18066 | n46644 ;
  assign n49479 = n43795 & n49478 ;
  assign n49480 = n48342 ^ n34810 ^ n1165 ;
  assign n49481 = ( n13259 & n17191 ) | ( n13259 & ~n49480 ) | ( n17191 & ~n49480 ) ;
  assign n49482 = n33986 ^ n20292 ^ n4757 ;
  assign n49483 = n25552 & n49482 ;
  assign n49484 = n49483 ^ n28084 ^ 1'b0 ;
  assign n49485 = n38757 ^ n7637 ^ 1'b0 ;
  assign n49486 = n7638 | n10540 ;
  assign n49487 = x97 | n49486 ;
  assign n49488 = ( ~n10304 & n23397 ) | ( ~n10304 & n49487 ) | ( n23397 & n49487 ) ;
  assign n49489 = ( ~n9642 & n14888 ) | ( ~n9642 & n19784 ) | ( n14888 & n19784 ) ;
  assign n49490 = ( n1266 & ~n5244 ) | ( n1266 & n12020 ) | ( ~n5244 & n12020 ) ;
  assign n49491 = ( ~x207 & n30400 ) | ( ~x207 & n30670 ) | ( n30400 & n30670 ) ;
  assign n49492 = n3860 & ~n4051 ;
  assign n49493 = n7316 & ~n49492 ;
  assign n49494 = n49493 ^ n21319 ^ n1355 ;
  assign n49495 = n5341 ^ n3316 ^ 1'b0 ;
  assign n49496 = n14523 | n49495 ;
  assign n49497 = n49496 ^ n49192 ^ n16726 ;
  assign n49498 = n1034 ^ x204 ^ 1'b0 ;
  assign n49499 = n2881 | n49498 ;
  assign n49500 = ( n3176 & n44993 ) | ( n3176 & ~n49499 ) | ( n44993 & ~n49499 ) ;
  assign n49501 = ( n35496 & n47660 ) | ( n35496 & n49500 ) | ( n47660 & n49500 ) ;
  assign n49502 = ( ~n13630 & n14269 ) | ( ~n13630 & n23134 ) | ( n14269 & n23134 ) ;
  assign n49503 = n49502 ^ n23374 ^ n5341 ;
  assign n49504 = n49503 ^ n20556 ^ n15773 ;
  assign n49505 = n44755 ^ n26051 ^ n3376 ;
  assign n49506 = ( ~n8117 & n45816 ) | ( ~n8117 & n49505 ) | ( n45816 & n49505 ) ;
  assign n49507 = ( n2162 & ~n8293 ) | ( n2162 & n19046 ) | ( ~n8293 & n19046 ) ;
  assign n49508 = ( n3049 & ~n12867 ) | ( n3049 & n39866 ) | ( ~n12867 & n39866 ) ;
  assign n49509 = ( n25249 & n49507 ) | ( n25249 & ~n49508 ) | ( n49507 & ~n49508 ) ;
  assign n49510 = ( n12749 & n12839 ) | ( n12749 & n36700 ) | ( n12839 & n36700 ) ;
  assign n49511 = n7063 & ~n15992 ;
  assign n49512 = ( n20764 & ~n35455 ) | ( n20764 & n49511 ) | ( ~n35455 & n49511 ) ;
  assign n49513 = n39043 ^ n34652 ^ 1'b0 ;
  assign n49514 = ~n11827 & n25253 ;
  assign n49515 = n49514 ^ n26028 ^ 1'b0 ;
  assign n49516 = n34662 ^ n15994 ^ 1'b0 ;
  assign n49517 = n47471 ^ n23098 ^ 1'b0 ;
  assign n49518 = n10582 & n49517 ;
  assign n49519 = ( ~n1710 & n42573 ) | ( ~n1710 & n49518 ) | ( n42573 & n49518 ) ;
  assign n49520 = ( n29698 & n30340 ) | ( n29698 & ~n36326 ) | ( n30340 & ~n36326 ) ;
  assign n49521 = n6130 & ~n49520 ;
  assign n49522 = n15301 | n31020 ;
  assign n49523 = n49522 ^ n25294 ^ 1'b0 ;
  assign n49524 = n6216 ^ n5394 ^ n339 ;
  assign n49525 = n49524 ^ n5527 ^ 1'b0 ;
  assign n49526 = n31743 ^ n15310 ^ n8785 ;
  assign n49527 = n9758 ^ n7742 ^ n473 ;
  assign n49528 = n28292 ^ n20374 ^ n7729 ;
  assign n49529 = ( ~n3039 & n37356 ) | ( ~n3039 & n49528 ) | ( n37356 & n49528 ) ;
  assign n49530 = ( n2851 & n9897 ) | ( n2851 & n11466 ) | ( n9897 & n11466 ) ;
  assign n49531 = n49530 ^ n5717 ^ n1623 ;
  assign n49532 = ( n6589 & n15891 ) | ( n6589 & n29724 ) | ( n15891 & n29724 ) ;
  assign n49533 = n49532 ^ n34350 ^ n32162 ;
  assign n49534 = ( n5034 & ~n14673 ) | ( n5034 & n44422 ) | ( ~n14673 & n44422 ) ;
  assign n49535 = ( n8305 & n49533 ) | ( n8305 & ~n49534 ) | ( n49533 & ~n49534 ) ;
  assign n49536 = n39820 ^ n25798 ^ n14070 ;
  assign n49537 = ~n29441 & n37031 ;
  assign n49538 = n49537 ^ n25841 ^ n11699 ;
  assign n49539 = n44917 ^ n22468 ^ n9923 ;
  assign n49540 = n33086 ^ n7455 ^ n1956 ;
  assign n49541 = n42336 ^ n41060 ^ n32125 ;
  assign n49542 = n4488 | n48718 ;
  assign n49543 = n49542 ^ n13481 ^ 1'b0 ;
  assign n49544 = n49543 ^ n15387 ^ 1'b0 ;
  assign n49545 = ~n10693 & n49544 ;
  assign n49546 = n21037 & n49545 ;
  assign n49548 = n35370 ^ n12095 ^ n5918 ;
  assign n49547 = n3128 & n3951 ;
  assign n49549 = n49548 ^ n49547 ^ 1'b0 ;
  assign n49550 = n5745 & n8704 ;
  assign n49551 = ~n17834 & n49550 ;
  assign n49552 = n49551 ^ n35426 ^ n29939 ;
  assign n49553 = n38563 ^ n24579 ^ n5974 ;
  assign n49555 = n39648 ^ n7950 ^ 1'b0 ;
  assign n49556 = n39589 & n49555 ;
  assign n49554 = n8977 | n40775 ;
  assign n49557 = n49556 ^ n49554 ^ n30917 ;
  assign n49558 = ( ~n11448 & n12273 ) | ( ~n11448 & n22849 ) | ( n12273 & n22849 ) ;
  assign n49559 = n49558 ^ n23190 ^ n3879 ;
  assign n49561 = n41408 ^ n9685 ^ n8543 ;
  assign n49562 = n49561 ^ n25057 ^ n14942 ;
  assign n49560 = n27662 ^ n27186 ^ n8422 ;
  assign n49563 = n49562 ^ n49560 ^ n14980 ;
  assign n49564 = n9984 ^ n299 ^ 1'b0 ;
  assign n49565 = n28804 & n49564 ;
  assign n49566 = ( n5339 & ~n37027 ) | ( n5339 & n49565 ) | ( ~n37027 & n49565 ) ;
  assign n49567 = ( n4571 & ~n21419 ) | ( n4571 & n29472 ) | ( ~n21419 & n29472 ) ;
  assign n49568 = ( n1405 & n13210 ) | ( n1405 & ~n44700 ) | ( n13210 & ~n44700 ) ;
  assign n49569 = n290 & ~n41109 ;
  assign n49570 = n40365 ^ n35061 ^ n9094 ;
  assign n49571 = ( n2562 & n14557 ) | ( n2562 & ~n49570 ) | ( n14557 & ~n49570 ) ;
  assign n49572 = n49571 ^ n43565 ^ 1'b0 ;
  assign n49573 = n18349 & n49572 ;
  assign n49574 = n14401 & ~n23741 ;
  assign n49575 = ( ~n17384 & n17639 ) | ( ~n17384 & n47170 ) | ( n17639 & n47170 ) ;
  assign n49576 = n41041 ^ n33315 ^ 1'b0 ;
  assign n49577 = n18902 ^ n15444 ^ 1'b0 ;
  assign n49578 = ~n30724 & n33711 ;
  assign n49579 = ( n12309 & n46733 ) | ( n12309 & n49578 ) | ( n46733 & n49578 ) ;
  assign n49580 = n7794 & ~n31469 ;
  assign n49581 = n49580 ^ n5860 ^ 1'b0 ;
  assign n49582 = ( n4941 & n17863 ) | ( n4941 & n42345 ) | ( n17863 & n42345 ) ;
  assign n49583 = n49582 ^ n18537 ^ n18182 ;
  assign n49584 = ( n8586 & ~n18837 ) | ( n8586 & n49040 ) | ( ~n18837 & n49040 ) ;
  assign n49585 = n26046 ^ n10801 ^ n1991 ;
  assign n49586 = ( n12623 & n15849 ) | ( n12623 & n49585 ) | ( n15849 & n49585 ) ;
  assign n49587 = ( n6034 & ~n13316 ) | ( n6034 & n49586 ) | ( ~n13316 & n49586 ) ;
  assign n49588 = ~n8145 & n11829 ;
  assign n49589 = ~n29140 & n49588 ;
  assign n49590 = n2795 & ~n14267 ;
  assign n49591 = ( n26525 & n49589 ) | ( n26525 & n49590 ) | ( n49589 & n49590 ) ;
  assign n49592 = n47885 ^ n27218 ^ n17404 ;
  assign n49593 = n46143 ^ n6209 ^ n1522 ;
  assign n49594 = ( ~n1736 & n36897 ) | ( ~n1736 & n49593 ) | ( n36897 & n49593 ) ;
  assign n49595 = ( ~n851 & n10620 ) | ( ~n851 & n17307 ) | ( n10620 & n17307 ) ;
  assign n49596 = n25913 ^ n12101 ^ 1'b0 ;
  assign n49597 = n49595 | n49596 ;
  assign n49598 = n11811 & n39967 ;
  assign n49599 = ( n2343 & n4693 ) | ( n2343 & ~n36635 ) | ( n4693 & ~n36635 ) ;
  assign n49602 = n20051 ^ n13098 ^ 1'b0 ;
  assign n49600 = x63 & n1899 ;
  assign n49601 = ( n1948 & n2388 ) | ( n1948 & ~n49600 ) | ( n2388 & ~n49600 ) ;
  assign n49603 = n49602 ^ n49601 ^ n2348 ;
  assign n49605 = n6274 & ~n21225 ;
  assign n49604 = n11734 & n15167 ;
  assign n49606 = n49605 ^ n49604 ^ 1'b0 ;
  assign n49607 = n49606 ^ n44735 ^ n38048 ;
  assign n49608 = n49607 ^ n36092 ^ x209 ;
  assign n49609 = n22246 ^ n14848 ^ n5521 ;
  assign n49610 = ( n17693 & ~n41027 ) | ( n17693 & n49609 ) | ( ~n41027 & n49609 ) ;
  assign n49611 = ( n1670 & n1815 ) | ( n1670 & n49610 ) | ( n1815 & n49610 ) ;
  assign n49612 = n15677 ^ n2339 ^ n1864 ;
  assign n49613 = n26130 ^ n22616 ^ n21496 ;
  assign n49614 = ( ~n21261 & n49612 ) | ( ~n21261 & n49613 ) | ( n49612 & n49613 ) ;
  assign n49615 = n45919 ^ n35156 ^ n22874 ;
  assign n49616 = n33737 ^ n14545 ^ n6986 ;
  assign n49617 = n49616 ^ n37993 ^ n37040 ;
  assign n49618 = ( n2854 & ~n6730 ) | ( n2854 & n20915 ) | ( ~n6730 & n20915 ) ;
  assign n49619 = ( n11857 & ~n49617 ) | ( n11857 & n49618 ) | ( ~n49617 & n49618 ) ;
  assign n49620 = n2178 & ~n22389 ;
  assign n49621 = n49620 ^ n33737 ^ 1'b0 ;
  assign n49622 = n49621 ^ n21566 ^ n11108 ;
  assign n49623 = n3131 & n48368 ;
  assign n49624 = n27427 ^ n10624 ^ n472 ;
  assign n49625 = ( n2533 & ~n12247 ) | ( n2533 & n49624 ) | ( ~n12247 & n49624 ) ;
  assign n49626 = ( n49622 & ~n49623 ) | ( n49622 & n49625 ) | ( ~n49623 & n49625 ) ;
  assign n49627 = ~n323 & n30825 ;
  assign n49628 = ~n4981 & n49627 ;
  assign n49629 = ~n9358 & n31299 ;
  assign n49630 = n49629 ^ n19911 ^ 1'b0 ;
  assign n49631 = n14716 | n49630 ;
  assign n49632 = ( n8573 & n14853 ) | ( n8573 & n20731 ) | ( n14853 & n20731 ) ;
  assign n49633 = ~n14896 & n37089 ;
  assign n49634 = ( n23962 & ~n36567 ) | ( n23962 & n43074 ) | ( ~n36567 & n43074 ) ;
  assign n49635 = n49634 ^ n21791 ^ n594 ;
  assign n49636 = ( n9808 & n20321 ) | ( n9808 & n45277 ) | ( n20321 & n45277 ) ;
  assign n49637 = n49636 ^ n34904 ^ n13358 ;
  assign n49638 = n30236 ^ n12259 ^ n2234 ;
  assign n49640 = ( n14140 & n20670 ) | ( n14140 & n34014 ) | ( n20670 & n34014 ) ;
  assign n49641 = ( n1199 & ~n4910 ) | ( n1199 & n49640 ) | ( ~n4910 & n49640 ) ;
  assign n49639 = ( n16823 & n22211 ) | ( n16823 & n43624 ) | ( n22211 & n43624 ) ;
  assign n49642 = n49641 ^ n49639 ^ n24310 ;
  assign n49643 = ( n6864 & n24211 ) | ( n6864 & ~n38211 ) | ( n24211 & ~n38211 ) ;
  assign n49644 = n33833 ^ n21599 ^ 1'b0 ;
  assign n49645 = ( ~n6004 & n49643 ) | ( ~n6004 & n49644 ) | ( n49643 & n49644 ) ;
  assign n49646 = ( n3961 & ~n36677 ) | ( n3961 & n39886 ) | ( ~n36677 & n39886 ) ;
  assign n49647 = ( n7674 & n9623 ) | ( n7674 & ~n13237 ) | ( n9623 & ~n13237 ) ;
  assign n49648 = ( n21299 & n49646 ) | ( n21299 & ~n49647 ) | ( n49646 & ~n49647 ) ;
  assign n49649 = ( ~n6793 & n37836 ) | ( ~n6793 & n47477 ) | ( n37836 & n47477 ) ;
  assign n49650 = n49649 ^ n34240 ^ n6196 ;
  assign n49651 = n35341 ^ n21288 ^ n15819 ;
  assign n49652 = n4792 ^ n1067 ^ 1'b0 ;
  assign n49653 = n5677 & ~n49652 ;
  assign n49654 = ( ~n44230 & n49651 ) | ( ~n44230 & n49653 ) | ( n49651 & n49653 ) ;
  assign n49655 = n27648 ^ n13202 ^ x105 ;
  assign n49656 = n31593 ^ n18874 ^ n1926 ;
  assign n49657 = ( n10381 & n33969 ) | ( n10381 & n49656 ) | ( n33969 & n49656 ) ;
  assign n49658 = n18401 | n49657 ;
  assign n49659 = ( n1113 & ~n16008 ) | ( n1113 & n30556 ) | ( ~n16008 & n30556 ) ;
  assign n49660 = ( n1712 & n3889 ) | ( n1712 & ~n19213 ) | ( n3889 & ~n19213 ) ;
  assign n49661 = n1567 & n49660 ;
  assign n49662 = n8867 ^ n3786 ^ x111 ;
  assign n49663 = n36167 & n49662 ;
  assign n49664 = n49663 ^ n15057 ^ n5776 ;
  assign n49665 = n49664 ^ n21277 ^ 1'b0 ;
  assign n49666 = n2593 & ~n49665 ;
  assign n49667 = n962 & ~n6929 ;
  assign n49668 = ~n27835 & n49667 ;
  assign n49669 = n22914 ^ n20277 ^ n17257 ;
  assign n49670 = n49669 ^ n32438 ^ n5864 ;
  assign n49671 = n49670 ^ n40582 ^ n13688 ;
  assign n49672 = ~n29737 & n49671 ;
  assign n49673 = ~n19855 & n49672 ;
  assign n49674 = n14656 ^ n13800 ^ x29 ;
  assign n49675 = ( n21061 & ~n30794 ) | ( n21061 & n49674 ) | ( ~n30794 & n49674 ) ;
  assign n49676 = n15602 & n49675 ;
  assign n49677 = n49676 ^ n41069 ^ n37354 ;
  assign n49678 = n10582 ^ n2005 ^ n988 ;
  assign n49679 = n10632 | n30329 ;
  assign n49680 = n6237 & n49679 ;
  assign n49681 = n49680 ^ n40274 ^ 1'b0 ;
  assign n49682 = ( n3341 & ~n11393 ) | ( n3341 & n49681 ) | ( ~n11393 & n49681 ) ;
  assign n49683 = n25274 | n49682 ;
  assign n49684 = n49678 | n49683 ;
  assign n49685 = ( n11395 & n48015 ) | ( n11395 & ~n49684 ) | ( n48015 & ~n49684 ) ;
  assign n49686 = ( ~n13948 & n32305 ) | ( ~n13948 & n49022 ) | ( n32305 & n49022 ) ;
  assign n49687 = n9451 ^ n9333 ^ n4599 ;
  assign n49688 = n49687 ^ n11871 ^ n9729 ;
  assign n49689 = ( n11961 & n30868 ) | ( n11961 & n49688 ) | ( n30868 & n49688 ) ;
  assign n49690 = ( n11383 & ~n22277 ) | ( n11383 & n49689 ) | ( ~n22277 & n49689 ) ;
  assign n49691 = n32543 ^ n21682 ^ n5812 ;
  assign n49692 = n49691 ^ n35020 ^ n4719 ;
  assign n49693 = n29233 ^ n28272 ^ 1'b0 ;
  assign n49699 = n22388 ^ n14203 ^ n6839 ;
  assign n49700 = n49699 ^ n18863 ^ n8431 ;
  assign n49694 = n47644 ^ n20251 ^ n12317 ;
  assign n49695 = n49694 ^ n15955 ^ n2976 ;
  assign n49696 = n49695 ^ n31665 ^ 1'b0 ;
  assign n49697 = ~n13657 & n49696 ;
  assign n49698 = n17754 & n49697 ;
  assign n49701 = n49700 ^ n49698 ^ n21039 ;
  assign n49702 = ~n11223 & n12804 ;
  assign n49703 = n49702 ^ n18886 ^ 1'b0 ;
  assign n49704 = n24214 ^ n23071 ^ n5993 ;
  assign n49705 = n9133 & n49704 ;
  assign n49706 = ~n45668 & n49705 ;
  assign n49707 = n49230 ^ n34285 ^ 1'b0 ;
  assign n49708 = ~n1459 & n4389 ;
  assign n49709 = ~n49707 & n49708 ;
  assign n49710 = n49709 ^ n36135 ^ 1'b0 ;
  assign n49711 = n26539 ^ n22635 ^ n13147 ;
  assign n49712 = ( n26174 & n36292 ) | ( n26174 & ~n49711 ) | ( n36292 & ~n49711 ) ;
  assign n49713 = n49712 ^ n16276 ^ n9426 ;
  assign n49715 = n16242 ^ n15095 ^ n14994 ;
  assign n49714 = n49182 ^ n11786 ^ n2618 ;
  assign n49716 = n49715 ^ n49714 ^ n43862 ;
  assign n49717 = n22145 ^ n10976 ^ n7389 ;
  assign n49718 = ( ~n1157 & n27564 ) | ( ~n1157 & n49717 ) | ( n27564 & n49717 ) ;
  assign n49719 = ( ~n19555 & n28844 ) | ( ~n19555 & n44934 ) | ( n28844 & n44934 ) ;
  assign n49720 = ~n11493 & n27192 ;
  assign n49721 = ~n6952 & n39491 ;
  assign n49722 = n33091 & ~n49721 ;
  assign n49723 = n7798 & ~n13009 ;
  assign n49724 = n49723 ^ n17596 ^ 1'b0 ;
  assign n49725 = n39059 ^ n28039 ^ n22291 ;
  assign n49726 = ~n14213 & n49725 ;
  assign n49727 = n3617 & n43113 ;
  assign n49728 = n49727 ^ n19690 ^ 1'b0 ;
  assign n49729 = ~n5673 & n37131 ;
  assign n49730 = ( ~n3724 & n9900 ) | ( ~n3724 & n23738 ) | ( n9900 & n23738 ) ;
  assign n49731 = ( x28 & n40322 ) | ( x28 & n49730 ) | ( n40322 & n49730 ) ;
  assign n49732 = ( n22061 & n23746 ) | ( n22061 & ~n40888 ) | ( n23746 & ~n40888 ) ;
  assign n49733 = n18822 ^ n3008 ^ 1'b0 ;
  assign n49734 = n48259 ^ n34371 ^ 1'b0 ;
  assign n49735 = n13148 | n49734 ;
  assign n49736 = ( n7118 & n29018 ) | ( n7118 & n49735 ) | ( n29018 & n49735 ) ;
  assign n49737 = ( n32975 & n49733 ) | ( n32975 & n49736 ) | ( n49733 & n49736 ) ;
  assign n49738 = n28639 ^ n15734 ^ 1'b0 ;
  assign n49739 = ~n9720 & n49738 ;
  assign n49740 = ( n9533 & n28840 ) | ( n9533 & n49739 ) | ( n28840 & n49739 ) ;
  assign n49741 = n11256 & n46110 ;
  assign n49742 = n6521 & n27405 ;
  assign n49743 = n29360 & n49742 ;
  assign n49744 = n16065 ^ n379 ^ 1'b0 ;
  assign n49745 = ( n7510 & n15195 ) | ( n7510 & ~n18907 ) | ( n15195 & ~n18907 ) ;
  assign n49746 = ( ~n1407 & n28316 ) | ( ~n1407 & n29891 ) | ( n28316 & n29891 ) ;
  assign n49747 = n49746 ^ n38844 ^ n33116 ;
  assign n49748 = n21030 ^ n17470 ^ 1'b0 ;
  assign n49749 = ~n14331 & n49748 ;
  assign n49750 = n23882 & n36420 ;
  assign n49751 = ( n2008 & ~n49749 ) | ( n2008 & n49750 ) | ( ~n49749 & n49750 ) ;
  assign n49752 = n19786 ^ n1866 ^ 1'b0 ;
  assign n49753 = n49752 ^ n17734 ^ n3706 ;
  assign n49754 = n3660 | n3752 ;
  assign n49755 = ( n21552 & n43430 ) | ( n21552 & n49754 ) | ( n43430 & n49754 ) ;
  assign n49756 = x168 & ~n49195 ;
  assign n49757 = n13727 & ~n16838 ;
  assign n49758 = n49757 ^ n7820 ^ n7696 ;
  assign n49759 = n49756 & n49758 ;
  assign n49760 = ~n3507 & n35408 ;
  assign n49761 = ~n26137 & n49760 ;
  assign n49762 = n20142 ^ n12218 ^ n5736 ;
  assign n49763 = ( n2456 & n13818 ) | ( n2456 & n42645 ) | ( n13818 & n42645 ) ;
  assign n49764 = n40461 ^ n27619 ^ n9254 ;
  assign n49765 = n40015 | n49764 ;
  assign n49766 = n49765 ^ n37271 ^ n15949 ;
  assign n49767 = n26941 & ~n28238 ;
  assign n49768 = n49767 ^ n10570 ^ 1'b0 ;
  assign n49769 = n49768 ^ n47755 ^ n14604 ;
  assign n49770 = n49769 ^ n6739 ^ 1'b0 ;
  assign n49771 = ( n1767 & ~n5158 ) | ( n1767 & n47629 ) | ( ~n5158 & n47629 ) ;
  assign n49772 = ~n26539 & n49771 ;
  assign n49773 = n49772 ^ n7348 ^ 1'b0 ;
  assign n49774 = n41156 ^ n32887 ^ n28313 ;
  assign n49775 = n8409 | n10985 ;
  assign n49776 = n48010 | n49775 ;
  assign n49777 = ~n6117 & n37390 ;
  assign n49778 = n38957 ^ n15710 ^ n13460 ;
  assign n49779 = n42805 ^ n31659 ^ n6357 ;
  assign n49780 = n48326 ^ n21381 ^ n1509 ;
  assign n49781 = ( ~n15817 & n30115 ) | ( ~n15817 & n38513 ) | ( n30115 & n38513 ) ;
  assign n49782 = n49781 ^ n37356 ^ n20413 ;
  assign n49783 = ( n2779 & ~n29231 ) | ( n2779 & n37175 ) | ( ~n29231 & n37175 ) ;
  assign n49784 = n49783 ^ n44813 ^ n29290 ;
  assign n49785 = n13735 ^ n3697 ^ 1'b0 ;
  assign n49786 = n21092 | n49785 ;
  assign n49787 = n27928 ^ n19446 ^ n14948 ;
  assign n49788 = ( n18505 & ~n21377 ) | ( n18505 & n49787 ) | ( ~n21377 & n49787 ) ;
  assign n49789 = n32521 & n49788 ;
  assign n49790 = n9140 & n49789 ;
  assign n49791 = n18041 ^ n17989 ^ 1'b0 ;
  assign n49792 = n33822 & n49791 ;
  assign n49803 = ( n7634 & n12245 ) | ( n7634 & ~n28136 ) | ( n12245 & ~n28136 ) ;
  assign n49804 = ( ~n10876 & n24125 ) | ( ~n10876 & n49803 ) | ( n24125 & n49803 ) ;
  assign n49798 = n28551 ^ n17903 ^ 1'b0 ;
  assign n49799 = n5803 | n49798 ;
  assign n49800 = n49799 ^ n6199 ^ 1'b0 ;
  assign n49801 = ( n22132 & n41576 ) | ( n22132 & n49800 ) | ( n41576 & n49800 ) ;
  assign n49797 = n35718 ^ n34481 ^ n16511 ;
  assign n49795 = n37211 ^ n36867 ^ n19209 ;
  assign n49796 = ( n20752 & ~n46615 ) | ( n20752 & n49795 ) | ( ~n46615 & n49795 ) ;
  assign n49802 = n49801 ^ n49797 ^ n49796 ;
  assign n49793 = n5222 & ~n15692 ;
  assign n49794 = ~n23205 & n49793 ;
  assign n49805 = n49804 ^ n49802 ^ n49794 ;
  assign n49806 = ( n14999 & n17504 ) | ( n14999 & ~n25193 ) | ( n17504 & ~n25193 ) ;
  assign n49807 = n41777 ^ n34072 ^ n3380 ;
  assign n49808 = n49807 ^ n21209 ^ n19418 ;
  assign n49810 = n8532 ^ n3616 ^ 1'b0 ;
  assign n49809 = n4720 & n9808 ;
  assign n49811 = n49810 ^ n49809 ^ n19758 ;
  assign n49812 = ( ~n31164 & n38993 ) | ( ~n31164 & n45660 ) | ( n38993 & n45660 ) ;
  assign n49813 = n19809 ^ n10211 ^ n8671 ;
  assign n49814 = n42830 ^ n26021 ^ 1'b0 ;
  assign n49815 = n43561 ^ n11436 ^ n8701 ;
  assign n49816 = ( n11018 & n49814 ) | ( n11018 & ~n49815 ) | ( n49814 & ~n49815 ) ;
  assign n49817 = n40790 ^ n38274 ^ 1'b0 ;
  assign n49818 = n37304 ^ n15534 ^ 1'b0 ;
  assign n49819 = n49817 | n49818 ;
  assign n49820 = n15637 & ~n44986 ;
  assign n49821 = ( n3102 & n9670 ) | ( n3102 & n36576 ) | ( n9670 & n36576 ) ;
  assign n49822 = ~n15215 & n31089 ;
  assign n49823 = ( n22323 & ~n48302 ) | ( n22323 & n49822 ) | ( ~n48302 & n49822 ) ;
  assign n49824 = ( n10068 & n30016 ) | ( n10068 & n32268 ) | ( n30016 & n32268 ) ;
  assign n49825 = n35768 ^ n25244 ^ 1'b0 ;
  assign n49826 = n49593 ^ n16285 ^ n8526 ;
  assign n49827 = n9668 ^ n7415 ^ n346 ;
  assign n49828 = ( n26059 & ~n49826 ) | ( n26059 & n49827 ) | ( ~n49826 & n49827 ) ;
  assign n49829 = n12472 ^ n9413 ^ n1308 ;
  assign n49830 = n49829 ^ n43436 ^ n6587 ;
  assign n49835 = n366 | n15927 ;
  assign n49831 = n27509 ^ n15288 ^ n1229 ;
  assign n49832 = ( n6665 & n14470 ) | ( n6665 & ~n16753 ) | ( n14470 & ~n16753 ) ;
  assign n49833 = ( n34674 & ~n49831 ) | ( n34674 & n49832 ) | ( ~n49831 & n49832 ) ;
  assign n49834 = n49833 ^ n30868 ^ n23013 ;
  assign n49836 = n49835 ^ n49834 ^ n33286 ;
  assign n49837 = n49836 ^ n9131 ^ n6052 ;
  assign n49838 = n23506 ^ n16195 ^ n708 ;
  assign n49839 = ( n755 & n6926 ) | ( n755 & n19518 ) | ( n6926 & n19518 ) ;
  assign n49840 = ( n379 & n28206 ) | ( n379 & n32721 ) | ( n28206 & n32721 ) ;
  assign n49841 = n4011 | n10856 ;
  assign n49842 = n49841 ^ n660 ^ 1'b0 ;
  assign n49843 = n49842 ^ n11349 ^ n2910 ;
  assign n49844 = n1970 ^ n1808 ^ 1'b0 ;
  assign n49845 = n49843 & n49844 ;
  assign n49846 = n49845 ^ n34862 ^ n14845 ;
  assign n49847 = n12425 ^ n11996 ^ n3173 ;
  assign n49848 = n49847 ^ n25416 ^ 1'b0 ;
  assign n49849 = n49848 ^ n44306 ^ n41464 ;
  assign n49850 = ( n680 & n3777 ) | ( n680 & ~n23890 ) | ( n3777 & ~n23890 ) ;
  assign n49851 = n49850 ^ n11182 ^ n1024 ;
  assign n49852 = ( n24939 & n29387 ) | ( n24939 & n49851 ) | ( n29387 & n49851 ) ;
  assign n49853 = n28039 & ~n47850 ;
  assign n49854 = n16300 & n49853 ;
  assign n49855 = ( n16867 & ~n29922 ) | ( n16867 & n34299 ) | ( ~n29922 & n34299 ) ;
  assign n49856 = ( n3589 & n30097 ) | ( n3589 & ~n49855 ) | ( n30097 & ~n49855 ) ;
  assign n49857 = n49411 ^ n9882 ^ n2729 ;
  assign n49858 = n16432 ^ n16028 ^ n2772 ;
  assign n49859 = ( n18978 & n41718 ) | ( n18978 & ~n49858 ) | ( n41718 & ~n49858 ) ;
  assign n49860 = ( n2875 & n16988 ) | ( n2875 & ~n20084 ) | ( n16988 & ~n20084 ) ;
  assign n49861 = n49860 ^ n12869 ^ 1'b0 ;
  assign n49862 = n44031 ^ n26591 ^ n21308 ;
  assign n49863 = ( n1193 & n8720 ) | ( n1193 & ~n49862 ) | ( n8720 & ~n49862 ) ;
  assign n49864 = ~n1903 & n15347 ;
  assign n49865 = n39824 ^ n6461 ^ 1'b0 ;
  assign n49866 = n14498 | n49865 ;
  assign n49867 = n2618 & ~n49866 ;
  assign n49868 = ( n9029 & n18753 ) | ( n9029 & ~n37403 ) | ( n18753 & ~n37403 ) ;
  assign n49869 = ( n10866 & ~n14318 ) | ( n10866 & n19112 ) | ( ~n14318 & n19112 ) ;
  assign n49870 = n40567 ^ n36228 ^ n22086 ;
  assign n49871 = n41777 ^ n11321 ^ n8043 ;
  assign n49872 = n23555 ^ n12604 ^ 1'b0 ;
  assign n49873 = n49872 ^ n45122 ^ n29682 ;
  assign n49874 = n49873 ^ n33407 ^ n11018 ;
  assign n49875 = n15001 | n15457 ;
  assign n49876 = n49875 ^ n27733 ^ n24723 ;
  assign n49877 = ( ~n11085 & n11312 ) | ( ~n11085 & n31671 ) | ( n11312 & n31671 ) ;
  assign n49878 = n17096 ^ n8977 ^ 1'b0 ;
  assign n49879 = ( n6833 & n33811 ) | ( n6833 & n49878 ) | ( n33811 & n49878 ) ;
  assign n49880 = ~n39257 & n41673 ;
  assign n49881 = n29824 ^ n24555 ^ 1'b0 ;
  assign n49882 = n49881 ^ n47774 ^ n31181 ;
  assign n49883 = n28942 ^ n13928 ^ n7582 ;
  assign n49884 = n11360 | n16245 ;
  assign n49885 = n19183 | n49884 ;
  assign n49886 = n35540 ^ n11539 ^ n8899 ;
  assign n49887 = ( n35107 & n49885 ) | ( n35107 & ~n49886 ) | ( n49885 & ~n49886 ) ;
  assign n49888 = ( n26941 & n28272 ) | ( n26941 & ~n41101 ) | ( n28272 & ~n41101 ) ;
  assign n49889 = n49888 ^ n16795 ^ n8301 ;
  assign n49890 = n49889 ^ n37497 ^ n20955 ;
  assign n49893 = n45499 ^ n44707 ^ n35551 ;
  assign n49891 = ( n6448 & ~n10111 ) | ( n6448 & n45901 ) | ( ~n10111 & n45901 ) ;
  assign n49892 = ( ~n27719 & n30388 ) | ( ~n27719 & n49891 ) | ( n30388 & n49891 ) ;
  assign n49894 = n49893 ^ n49892 ^ n926 ;
  assign n49895 = n24772 ^ n10646 ^ n6579 ;
  assign n49896 = n10705 ^ n9040 ^ n882 ;
  assign n49897 = ( n19978 & n24074 ) | ( n19978 & n49896 ) | ( n24074 & n49896 ) ;
  assign n49898 = n23958 ^ n10888 ^ n2928 ;
  assign n49899 = ( n6201 & ~n11835 ) | ( n6201 & n28350 ) | ( ~n11835 & n28350 ) ;
  assign n49900 = n49899 ^ n35680 ^ 1'b0 ;
  assign n49901 = n4706 & ~n49900 ;
  assign n49902 = n49901 ^ n1862 ^ 1'b0 ;
  assign n49903 = n19098 | n49902 ;
  assign n49904 = ( n1790 & n5904 ) | ( n1790 & n8834 ) | ( n5904 & n8834 ) ;
  assign n49905 = n28121 & n49904 ;
  assign n49906 = ~n45069 & n49905 ;
  assign n49907 = n46197 ^ n13113 ^ n11440 ;
  assign n49908 = n40220 ^ n12184 ^ 1'b0 ;
  assign n49909 = n40180 & n49908 ;
  assign n49910 = ( n46746 & n49907 ) | ( n46746 & n49909 ) | ( n49907 & n49909 ) ;
  assign n49911 = ~n23582 & n33422 ;
  assign n49912 = n49911 ^ n23524 ^ 1'b0 ;
  assign n49913 = ( ~n6890 & n47780 ) | ( ~n6890 & n49912 ) | ( n47780 & n49912 ) ;
  assign n49914 = ( ~n5477 & n10169 ) | ( ~n5477 & n27037 ) | ( n10169 & n27037 ) ;
  assign n49915 = n27794 ^ n27754 ^ 1'b0 ;
  assign n49916 = ( n26361 & n36657 ) | ( n26361 & n49915 ) | ( n36657 & n49915 ) ;
  assign n49917 = ( n20967 & ~n32169 ) | ( n20967 & n33634 ) | ( ~n32169 & n33634 ) ;
  assign n49920 = ( n16509 & n36709 ) | ( n16509 & n44060 ) | ( n36709 & n44060 ) ;
  assign n49918 = n6688 | n38019 ;
  assign n49919 = n49918 ^ n13403 ^ 1'b0 ;
  assign n49921 = n49920 ^ n49919 ^ n5724 ;
  assign n49922 = n33159 ^ n2345 ^ n1486 ;
  assign n49923 = ( n22255 & n35243 ) | ( n22255 & ~n49922 ) | ( n35243 & ~n49922 ) ;
  assign n49924 = ( n14702 & ~n28959 ) | ( n14702 & n34614 ) | ( ~n28959 & n34614 ) ;
  assign n49925 = ( n20115 & n45597 ) | ( n20115 & ~n49924 ) | ( n45597 & ~n49924 ) ;
  assign n49926 = n9791 & ~n32390 ;
  assign n49927 = n49925 & n49926 ;
  assign n49928 = n16037 ^ n9986 ^ n427 ;
  assign n49929 = n49928 ^ n1751 ^ 1'b0 ;
  assign n49930 = n19590 & n49929 ;
  assign n49931 = n49930 ^ n28015 ^ n3789 ;
  assign n49932 = n39240 ^ n6238 ^ 1'b0 ;
  assign n49933 = ( n24212 & n34467 ) | ( n24212 & ~n49932 ) | ( n34467 & ~n49932 ) ;
  assign n49934 = n18474 ^ n1030 ^ 1'b0 ;
  assign n49935 = n36256 ^ n23012 ^ 1'b0 ;
  assign n49936 = n17092 ^ n10259 ^ 1'b0 ;
  assign n49937 = n3952 | n49936 ;
  assign n49938 = n49937 ^ n18120 ^ n3765 ;
  assign n49939 = n7744 & n20936 ;
  assign n49940 = n49939 ^ n11827 ^ 1'b0 ;
  assign n49941 = n49940 ^ n26394 ^ n12738 ;
  assign n49942 = ( n35537 & ~n49938 ) | ( n35537 & n49941 ) | ( ~n49938 & n49941 ) ;
  assign n49943 = n30811 ^ n11084 ^ n9353 ;
  assign n49944 = n10893 | n36204 ;
  assign n49945 = ( n2700 & ~n42962 ) | ( n2700 & n49944 ) | ( ~n42962 & n49944 ) ;
  assign n49946 = ( n17681 & n32093 ) | ( n17681 & n41051 ) | ( n32093 & n41051 ) ;
  assign n49947 = n33001 & n46081 ;
  assign n49949 = ( n4894 & n7083 ) | ( n4894 & n48742 ) | ( n7083 & n48742 ) ;
  assign n49948 = n31321 ^ n27574 ^ n3361 ;
  assign n49950 = n49949 ^ n49948 ^ n14554 ;
  assign n49951 = ( n24513 & n28630 ) | ( n24513 & ~n49950 ) | ( n28630 & ~n49950 ) ;
  assign n49952 = ( n7544 & ~n29685 ) | ( n7544 & n40976 ) | ( ~n29685 & n40976 ) ;
  assign n49953 = n49952 ^ n4213 ^ 1'b0 ;
  assign n49954 = ( n16253 & n39784 ) | ( n16253 & ~n49953 ) | ( n39784 & ~n49953 ) ;
  assign n49955 = n35361 ^ n23819 ^ n20719 ;
  assign n49956 = n49955 ^ n5759 ^ 1'b0 ;
  assign n49957 = ~n16069 & n49956 ;
  assign n49958 = n49957 ^ n15072 ^ n1555 ;
  assign n49959 = n5571 & n32985 ;
  assign n49960 = n49959 ^ n29255 ^ n25299 ;
  assign n49961 = n49960 ^ n32758 ^ n29698 ;
  assign n49962 = n2132 | n10437 ;
  assign n49963 = n25344 ^ n18503 ^ n13887 ;
  assign n49964 = n49963 ^ n44627 ^ 1'b0 ;
  assign n49965 = ( n434 & ~n49962 ) | ( n434 & n49964 ) | ( ~n49962 & n49964 ) ;
  assign n49966 = ( n19591 & n35481 ) | ( n19591 & ~n49965 ) | ( n35481 & ~n49965 ) ;
  assign n49967 = ( n19606 & ~n36101 ) | ( n19606 & n47163 ) | ( ~n36101 & n47163 ) ;
  assign n49968 = n4659 | n10163 ;
  assign n49969 = n49968 ^ n45243 ^ 1'b0 ;
  assign n49970 = n45106 ^ n25181 ^ 1'b0 ;
  assign n49971 = n22385 ^ n14032 ^ 1'b0 ;
  assign n49972 = n2201 & n49971 ;
  assign n49973 = n22560 ^ n13119 ^ n3114 ;
  assign n49974 = n35243 ^ n17261 ^ n2832 ;
  assign n49975 = ( n4156 & n45161 ) | ( n4156 & n49974 ) | ( n45161 & n49974 ) ;
  assign n49976 = n22125 & ~n35332 ;
  assign n49977 = n49976 ^ n16159 ^ 1'b0 ;
  assign n49978 = n20812 ^ n9292 ^ n4589 ;
  assign n49979 = n49978 ^ n42092 ^ n3255 ;
  assign n49980 = n49977 & n49979 ;
  assign n49981 = n45656 ^ n40282 ^ n18338 ;
  assign n49982 = n44018 ^ n34902 ^ n2455 ;
  assign n49983 = n49982 ^ n38663 ^ n29561 ;
  assign n49984 = n24782 ^ n21984 ^ n2428 ;
  assign n49985 = n49984 ^ n15878 ^ n5641 ;
  assign n49986 = n49985 ^ n28527 ^ n23910 ;
  assign n49987 = n39688 ^ n34939 ^ 1'b0 ;
  assign n49988 = ~n7561 & n30467 ;
  assign n49989 = ~n49646 & n49988 ;
  assign n49990 = n19046 ^ n11907 ^ n8298 ;
  assign n49991 = n3845 & n49990 ;
  assign n49992 = n15017 & n49991 ;
  assign n49993 = n36703 ^ n6483 ^ n2867 ;
  assign n49994 = ( ~n788 & n29014 ) | ( ~n788 & n49098 ) | ( n29014 & n49098 ) ;
  assign n49995 = ( n8804 & n29052 ) | ( n8804 & ~n49994 ) | ( n29052 & ~n49994 ) ;
  assign n49996 = ( n42026 & ~n49993 ) | ( n42026 & n49995 ) | ( ~n49993 & n49995 ) ;
  assign n49997 = n14210 ^ n12184 ^ n4361 ;
  assign n49998 = n24110 ^ n14675 ^ n3585 ;
  assign n49999 = n7722 | n49998 ;
  assign n50000 = ( n2155 & ~n46198 ) | ( n2155 & n49999 ) | ( ~n46198 & n49999 ) ;
  assign n50001 = n4545 & n49695 ;
  assign n50002 = n41410 ^ n6151 ^ 1'b0 ;
  assign n50003 = n2115 & n14426 ;
  assign n50004 = ( n2187 & ~n16546 ) | ( n2187 & n28272 ) | ( ~n16546 & n28272 ) ;
  assign n50005 = n9484 & n14061 ;
  assign n50006 = n14978 ^ n14808 ^ n7818 ;
  assign n50007 = ( n9186 & n12809 ) | ( n9186 & ~n20613 ) | ( n12809 & ~n20613 ) ;
  assign n50008 = n50007 ^ n8262 ^ n501 ;
  assign n50009 = n3182 ^ n2133 ^ 1'b0 ;
  assign n50010 = ( n9993 & n18328 ) | ( n9993 & n50009 ) | ( n18328 & n50009 ) ;
  assign n50011 = n50010 ^ n29532 ^ n16194 ;
  assign n50012 = ( ~n10433 & n16778 ) | ( ~n10433 & n44894 ) | ( n16778 & n44894 ) ;
  assign n50015 = n3412 | n24048 ;
  assign n50016 = n50015 ^ n9865 ^ n6421 ;
  assign n50013 = n19656 ^ n18496 ^ 1'b0 ;
  assign n50014 = ~n19843 & n50013 ;
  assign n50017 = n50016 ^ n50014 ^ n23027 ;
  assign n50018 = ( ~n8258 & n17045 ) | ( ~n8258 & n29825 ) | ( n17045 & n29825 ) ;
  assign n50019 = n50018 ^ n22804 ^ 1'b0 ;
  assign n50020 = ( n13200 & n50017 ) | ( n13200 & n50019 ) | ( n50017 & n50019 ) ;
  assign n50021 = n10531 & n19526 ;
  assign n50022 = ~n50020 & n50021 ;
  assign n50023 = ( n5196 & n24811 ) | ( n5196 & ~n50022 ) | ( n24811 & ~n50022 ) ;
  assign n50024 = n21820 ^ n11524 ^ n372 ;
  assign n50025 = n11963 ^ n2832 ^ n1478 ;
  assign n50026 = ( ~n800 & n50024 ) | ( ~n800 & n50025 ) | ( n50024 & n50025 ) ;
  assign n50031 = ( n3093 & n4177 ) | ( n3093 & ~n19232 ) | ( n4177 & ~n19232 ) ;
  assign n50032 = n50031 ^ n5354 ^ 1'b0 ;
  assign n50033 = n13462 | n50032 ;
  assign n50029 = n22395 | n25929 ;
  assign n50027 = ( n5699 & ~n15407 ) | ( n5699 & n34944 ) | ( ~n15407 & n34944 ) ;
  assign n50028 = n50027 ^ n24808 ^ n17193 ;
  assign n50030 = n50029 ^ n50028 ^ n49771 ;
  assign n50034 = n50033 ^ n50030 ^ n18812 ;
  assign n50035 = n44430 ^ n6368 ^ n5931 ;
  assign n50039 = n11569 & ~n46107 ;
  assign n50040 = n2441 & n50039 ;
  assign n50036 = ( n10341 & n23482 ) | ( n10341 & n31070 ) | ( n23482 & n31070 ) ;
  assign n50037 = n50036 ^ n19652 ^ n7269 ;
  assign n50038 = n18478 & ~n50037 ;
  assign n50041 = n50040 ^ n50038 ^ 1'b0 ;
  assign n50042 = n19924 | n27627 ;
  assign n50043 = ~n4356 & n49404 ;
  assign n50044 = n7124 & ~n50043 ;
  assign n50045 = n50044 ^ n36246 ^ 1'b0 ;
  assign n50046 = n15780 ^ n6423 ^ 1'b0 ;
  assign n50047 = ( n6910 & ~n24038 ) | ( n6910 & n43425 ) | ( ~n24038 & n43425 ) ;
  assign n50048 = n5474 & n45105 ;
  assign n50049 = ~n50047 & n50048 ;
  assign n50050 = n50049 ^ n17179 ^ n3522 ;
  assign n50051 = ( n1274 & n11872 ) | ( n1274 & n50050 ) | ( n11872 & n50050 ) ;
  assign n50052 = n48894 ^ n42543 ^ n14081 ;
  assign n50053 = n30211 ^ n22647 ^ n15136 ;
  assign n50054 = n9069 ^ n7242 ^ n3474 ;
  assign n50055 = n50054 ^ n30171 ^ n20617 ;
  assign n50056 = n50055 ^ n34415 ^ n8678 ;
  assign n50058 = n32375 ^ n10956 ^ 1'b0 ;
  assign n50059 = n28505 ^ n5088 ^ 1'b0 ;
  assign n50060 = n50058 | n50059 ;
  assign n50057 = x22 & ~n23165 ;
  assign n50061 = n50060 ^ n50057 ^ 1'b0 ;
  assign n50062 = n2174 & n31536 ;
  assign n50063 = n50062 ^ n28782 ^ 1'b0 ;
  assign n50064 = n50063 ^ n11662 ^ 1'b0 ;
  assign n50065 = n30838 ^ n18330 ^ n2744 ;
  assign n50066 = ( ~n8115 & n46863 ) | ( ~n8115 & n50065 ) | ( n46863 & n50065 ) ;
  assign n50067 = n40321 ^ n33666 ^ 1'b0 ;
  assign n50068 = n49356 ^ n21593 ^ n19420 ;
  assign n50069 = ( n8087 & n50067 ) | ( n8087 & ~n50068 ) | ( n50067 & ~n50068 ) ;
  assign n50070 = n50069 ^ n15809 ^ n1872 ;
  assign n50071 = ( ~n33494 & n39120 ) | ( ~n33494 & n50070 ) | ( n39120 & n50070 ) ;
  assign n50072 = n21091 ^ n13770 ^ n13681 ;
  assign n50073 = ( n9165 & n31017 ) | ( n9165 & n50072 ) | ( n31017 & n50072 ) ;
  assign n50074 = n25376 ^ n17171 ^ n2569 ;
  assign n50075 = n28391 ^ n12705 ^ n10814 ;
  assign n50076 = n50075 ^ n37757 ^ n27571 ;
  assign n50077 = ( n49187 & ~n50074 ) | ( n49187 & n50076 ) | ( ~n50074 & n50076 ) ;
  assign n50078 = n4752 & n5978 ;
  assign n50079 = n50078 ^ n11812 ^ n989 ;
  assign n50080 = n1796 | n44106 ;
  assign n50081 = n28269 ^ n15938 ^ 1'b0 ;
  assign n50082 = ~n15450 & n50081 ;
  assign n50083 = ( n9131 & ~n15708 ) | ( n9131 & n44020 ) | ( ~n15708 & n44020 ) ;
  assign n50084 = n35896 ^ n6177 ^ 1'b0 ;
  assign n50085 = ( ~n8430 & n12337 ) | ( ~n8430 & n50084 ) | ( n12337 & n50084 ) ;
  assign n50086 = n44675 ^ n22630 ^ n8103 ;
  assign n50087 = n11020 | n50086 ;
  assign n50088 = n25247 & ~n50087 ;
  assign n50089 = ( n17428 & n41278 ) | ( n17428 & n50088 ) | ( n41278 & n50088 ) ;
  assign n50090 = ( n7749 & ~n8835 ) | ( n7749 & n11750 ) | ( ~n8835 & n11750 ) ;
  assign n50091 = n50090 ^ n27723 ^ n26460 ;
  assign n50092 = n50091 ^ n38333 ^ n2024 ;
  assign n50093 = ( n13063 & ~n13178 ) | ( n13063 & n37833 ) | ( ~n13178 & n37833 ) ;
  assign n50094 = n11583 ^ n8047 ^ 1'b0 ;
  assign n50095 = n50093 | n50094 ;
  assign n50096 = n50095 ^ n17875 ^ n15792 ;
  assign n50097 = ( ~n41913 & n50092 ) | ( ~n41913 & n50096 ) | ( n50092 & n50096 ) ;
  assign n50098 = n15689 ^ n9873 ^ n1329 ;
  assign n50099 = n19149 ^ n10207 ^ n540 ;
  assign n50100 = ( n10274 & ~n21412 ) | ( n10274 & n50099 ) | ( ~n21412 & n50099 ) ;
  assign n50101 = n29105 ^ n26716 ^ n10390 ;
  assign n50102 = ( n473 & n5510 ) | ( n473 & n50101 ) | ( n5510 & n50101 ) ;
  assign n50103 = ( n17045 & n18143 ) | ( n17045 & n25506 ) | ( n18143 & n25506 ) ;
  assign n50104 = ( n21811 & ~n27985 ) | ( n21811 & n50103 ) | ( ~n27985 & n50103 ) ;
  assign n50105 = n50104 ^ n27856 ^ 1'b0 ;
  assign n50106 = n27940 ^ n6984 ^ n4759 ;
  assign n50109 = ( n2937 & n15432 ) | ( n2937 & ~n18155 ) | ( n15432 & ~n18155 ) ;
  assign n50107 = n35729 ^ n14719 ^ 1'b0 ;
  assign n50108 = n39502 & ~n50107 ;
  assign n50110 = n50109 ^ n50108 ^ n30412 ;
  assign n50111 = n46153 ^ n23621 ^ n4247 ;
  assign n50112 = n28271 ^ n5471 ^ n1699 ;
  assign n50113 = n24076 ^ n16157 ^ n2743 ;
  assign n50114 = n17560 ^ n7817 ^ 1'b0 ;
  assign n50115 = n8604 & n50114 ;
  assign n50116 = ( n8343 & ~n45722 ) | ( n8343 & n50115 ) | ( ~n45722 & n50115 ) ;
  assign n50117 = n4032 & ~n50116 ;
  assign n50118 = ( ~n8160 & n17875 ) | ( ~n8160 & n34278 ) | ( n17875 & n34278 ) ;
  assign n50119 = ( n503 & n9803 ) | ( n503 & n13629 ) | ( n9803 & n13629 ) ;
  assign n50120 = n50119 ^ n12682 ^ n3214 ;
  assign n50121 = ( n13234 & ~n48693 ) | ( n13234 & n50120 ) | ( ~n48693 & n50120 ) ;
  assign n50122 = n4357 & n10498 ;
  assign n50123 = ~n5966 & n15176 ;
  assign n50124 = n7602 & n50123 ;
  assign n50125 = n3374 | n50124 ;
  assign n50126 = n50122 & ~n50125 ;
  assign n50127 = n34213 ^ n30434 ^ n4559 ;
  assign n50128 = n19579 & n50127 ;
  assign n50129 = n44872 ^ n13299 ^ 1'b0 ;
  assign n50130 = n24303 & ~n50129 ;
  assign n50134 = n37249 ^ n16263 ^ n12424 ;
  assign n50133 = n35666 ^ n30303 ^ n4378 ;
  assign n50131 = n14549 ^ n10023 ^ n5132 ;
  assign n50132 = n20434 & n50131 ;
  assign n50135 = n50134 ^ n50133 ^ n50132 ;
  assign n50136 = ( n42475 & n50130 ) | ( n42475 & n50135 ) | ( n50130 & n50135 ) ;
  assign n50137 = n25814 ^ n19255 ^ 1'b0 ;
  assign n50138 = ( n13569 & ~n24088 ) | ( n13569 & n50137 ) | ( ~n24088 & n50137 ) ;
  assign n50139 = n37473 ^ n18391 ^ n12343 ;
  assign n50140 = ( n7370 & ~n24525 ) | ( n7370 & n30717 ) | ( ~n24525 & n30717 ) ;
  assign n50141 = ( ~n25546 & n48092 ) | ( ~n25546 & n50140 ) | ( n48092 & n50140 ) ;
  assign n50142 = n42405 ^ n30835 ^ n6845 ;
  assign n50143 = ( ~n12607 & n34263 ) | ( ~n12607 & n38814 ) | ( n34263 & n38814 ) ;
  assign n50144 = ( ~n1114 & n31746 ) | ( ~n1114 & n39540 ) | ( n31746 & n39540 ) ;
  assign n50145 = n41951 ^ n12071 ^ 1'b0 ;
  assign n50146 = n1921 | n19917 ;
  assign n50147 = n28106 ^ n8314 ^ 1'b0 ;
  assign n50148 = ~n50146 & n50147 ;
  assign n50149 = ~n3098 & n28029 ;
  assign n50150 = n50149 ^ n18515 ^ 1'b0 ;
  assign n50152 = ( ~n16376 & n37732 ) | ( ~n16376 & n45763 ) | ( n37732 & n45763 ) ;
  assign n50153 = n50152 ^ n29042 ^ n26702 ;
  assign n50151 = n48458 ^ n16589 ^ n8377 ;
  assign n50154 = n50153 ^ n50151 ^ n20965 ;
  assign n50155 = n4792 & ~n50154 ;
  assign n50156 = n5903 ^ n2416 ^ n2391 ;
  assign n50157 = n50156 ^ n30058 ^ n27084 ;
  assign n50158 = ( n21504 & n23244 ) | ( n21504 & n43356 ) | ( n23244 & n43356 ) ;
  assign n50159 = ( n2454 & n7898 ) | ( n2454 & ~n50158 ) | ( n7898 & ~n50158 ) ;
  assign n50160 = ( n431 & ~n7081 ) | ( n431 & n16211 ) | ( ~n7081 & n16211 ) ;
  assign n50161 = n50160 ^ n30045 ^ n1815 ;
  assign n50162 = n29924 ^ n7648 ^ n884 ;
  assign n50163 = n50162 ^ n38905 ^ n7991 ;
  assign n50164 = ( n15530 & n22227 ) | ( n15530 & n34347 ) | ( n22227 & n34347 ) ;
  assign n50165 = ( n22089 & n50163 ) | ( n22089 & n50164 ) | ( n50163 & n50164 ) ;
  assign n50166 = ( ~n5401 & n38758 ) | ( ~n5401 & n48800 ) | ( n38758 & n48800 ) ;
  assign n50167 = n12544 ^ n5311 ^ 1'b0 ;
  assign n50168 = n27978 | n50167 ;
  assign n50169 = ( n24950 & ~n39198 ) | ( n24950 & n40016 ) | ( ~n39198 & n40016 ) ;
  assign n50170 = n313 & n50169 ;
  assign n50171 = n50170 ^ x139 ^ 1'b0 ;
  assign n50172 = n25937 ^ n2797 ^ n1036 ;
  assign n50173 = ( n10875 & ~n19029 ) | ( n10875 & n50172 ) | ( ~n19029 & n50172 ) ;
  assign n50174 = n7511 & n50173 ;
  assign n50175 = ~n15444 & n50174 ;
  assign n50176 = n35742 & ~n50175 ;
  assign n50177 = n12769 | n19828 ;
  assign n50178 = ( ~n10277 & n15456 ) | ( ~n10277 & n50177 ) | ( n15456 & n50177 ) ;
  assign n50179 = n50178 ^ n19576 ^ n7944 ;
  assign n50180 = n28827 ^ n11360 ^ n3530 ;
  assign n50181 = n43016 ^ n37562 ^ n26464 ;
  assign n50182 = ( ~n8794 & n33207 ) | ( ~n8794 & n50181 ) | ( n33207 & n50181 ) ;
  assign n50183 = n5543 ^ n4770 ^ 1'b0 ;
  assign n50184 = n15286 ^ n14793 ^ n10961 ;
  assign n50185 = ( n8920 & n23197 ) | ( n8920 & ~n30700 ) | ( n23197 & ~n30700 ) ;
  assign n50186 = n8571 ^ n7731 ^ 1'b0 ;
  assign n50187 = ( n25759 & n50185 ) | ( n25759 & n50186 ) | ( n50185 & n50186 ) ;
  assign n50188 = ( ~n50183 & n50184 ) | ( ~n50183 & n50187 ) | ( n50184 & n50187 ) ;
  assign n50189 = n19776 ^ n16970 ^ n16204 ;
  assign n50190 = n11334 & ~n50189 ;
  assign n50191 = ( n33356 & n45720 ) | ( n33356 & n50190 ) | ( n45720 & n50190 ) ;
  assign n50192 = n32595 ^ n7358 ^ n3109 ;
  assign n50194 = n7009 | n18010 ;
  assign n50195 = n10140 & ~n50194 ;
  assign n50193 = n40879 ^ n2700 ^ 1'b0 ;
  assign n50196 = n50195 ^ n50193 ^ n16635 ;
  assign n50197 = n45933 ^ n17621 ^ n5683 ;
  assign n50198 = n50197 ^ n31914 ^ n8746 ;
  assign n50199 = n19783 & n50198 ;
  assign n50200 = n8056 ^ n7515 ^ 1'b0 ;
  assign n50201 = n37705 & n50200 ;
  assign n50202 = n28774 ^ n22957 ^ 1'b0 ;
  assign n50203 = ~n3837 & n50202 ;
  assign n50204 = ( n28133 & n31004 ) | ( n28133 & n50203 ) | ( n31004 & n50203 ) ;
  assign n50205 = n50204 ^ n42111 ^ n27951 ;
  assign n50206 = n13644 ^ n12494 ^ 1'b0 ;
  assign n50207 = n5681 & n50206 ;
  assign n50208 = n30727 & n50207 ;
  assign n50209 = ( n26798 & n49170 ) | ( n26798 & ~n50208 ) | ( n49170 & ~n50208 ) ;
  assign n50210 = n6961 & n34350 ;
  assign n50211 = ( n800 & ~n6957 ) | ( n800 & n50210 ) | ( ~n6957 & n50210 ) ;
  assign n50212 = n50211 ^ n36246 ^ n21463 ;
  assign n50216 = n37781 ^ n27595 ^ 1'b0 ;
  assign n50213 = n20398 ^ n3532 ^ 1'b0 ;
  assign n50214 = n49293 ^ n22376 ^ 1'b0 ;
  assign n50215 = n50213 & n50214 ;
  assign n50217 = n50216 ^ n50215 ^ n43413 ;
  assign n50218 = ( ~n8242 & n40044 ) | ( ~n8242 & n50217 ) | ( n40044 & n50217 ) ;
  assign n50219 = ( ~n5333 & n24351 ) | ( ~n5333 & n38263 ) | ( n24351 & n38263 ) ;
  assign n50220 = ( n2206 & n15889 ) | ( n2206 & n16950 ) | ( n15889 & n16950 ) ;
  assign n50221 = n27720 & ~n50220 ;
  assign n50222 = ( n30986 & ~n50219 ) | ( n30986 & n50221 ) | ( ~n50219 & n50221 ) ;
  assign n50223 = n37423 ^ n27904 ^ n8860 ;
  assign n50224 = ~n12794 & n44526 ;
  assign n50225 = n50224 ^ n29948 ^ 1'b0 ;
  assign n50226 = n43592 ^ n24161 ^ 1'b0 ;
  assign n50227 = n12685 & ~n50226 ;
  assign n50228 = ~n2200 & n30570 ;
  assign n50229 = n50228 ^ n46410 ^ 1'b0 ;
  assign n50230 = ( n6969 & n33409 ) | ( n6969 & n40836 ) | ( n33409 & n40836 ) ;
  assign n50231 = n50230 ^ n15434 ^ 1'b0 ;
  assign n50232 = n50231 ^ n35654 ^ n2854 ;
  assign n50233 = ( n2363 & n18498 ) | ( n2363 & n50232 ) | ( n18498 & n50232 ) ;
  assign n50234 = n39005 ^ n17827 ^ 1'b0 ;
  assign n50235 = n16615 & ~n50234 ;
  assign n50236 = n50235 ^ n31161 ^ n30655 ;
  assign n50237 = ( n34401 & ~n38933 ) | ( n34401 & n50236 ) | ( ~n38933 & n50236 ) ;
  assign n50238 = n44642 ^ n43998 ^ n20793 ;
  assign n50239 = n20900 ^ n5987 ^ 1'b0 ;
  assign n50241 = ( x164 & n6619 ) | ( x164 & ~n17301 ) | ( n6619 & ~n17301 ) ;
  assign n50240 = n9251 | n49963 ;
  assign n50242 = n50241 ^ n50240 ^ 1'b0 ;
  assign n50243 = n33897 ^ n22875 ^ n17290 ;
  assign n50244 = n22767 ^ n13841 ^ n6401 ;
  assign n50245 = ~n50243 & n50244 ;
  assign n50246 = n50245 ^ n25805 ^ 1'b0 ;
  assign n50247 = n25129 & n28330 ;
  assign n50248 = n27370 & n50247 ;
  assign n50249 = n36908 ^ n20590 ^ n8442 ;
  assign n50250 = n46432 ^ n3495 ^ 1'b0 ;
  assign n50251 = n19752 | n27158 ;
  assign n50256 = n6118 & n16885 ;
  assign n50257 = ~n19817 & n50256 ;
  assign n50252 = n16794 & n24887 ;
  assign n50253 = n1323 & n50252 ;
  assign n50254 = ( n1854 & ~n17185 ) | ( n1854 & n23513 ) | ( ~n17185 & n23513 ) ;
  assign n50255 = ( n39801 & n50253 ) | ( n39801 & ~n50254 ) | ( n50253 & ~n50254 ) ;
  assign n50258 = n50257 ^ n50255 ^ 1'b0 ;
  assign n50261 = ( n13069 & n16381 ) | ( n13069 & n18871 ) | ( n16381 & n18871 ) ;
  assign n50259 = n9527 ^ n3629 ^ n3106 ;
  assign n50260 = ~n682 & n50259 ;
  assign n50262 = n50261 ^ n50260 ^ 1'b0 ;
  assign n50263 = n50262 ^ n14130 ^ 1'b0 ;
  assign n50264 = ( n1131 & ~n5310 ) | ( n1131 & n10761 ) | ( ~n5310 & n10761 ) ;
  assign n50265 = n16035 & ~n42424 ;
  assign n50266 = n50264 & n50265 ;
  assign n50267 = ( n6044 & n12798 ) | ( n6044 & n50266 ) | ( n12798 & n50266 ) ;
  assign n50268 = n7030 & ~n47541 ;
  assign n50269 = n44282 & n50268 ;
  assign n50270 = ( n30046 & ~n37333 ) | ( n30046 & n38968 ) | ( ~n37333 & n38968 ) ;
  assign n50271 = n50270 ^ n45534 ^ n28293 ;
  assign n50275 = ( n480 & n7034 ) | ( n480 & ~n12988 ) | ( n7034 & ~n12988 ) ;
  assign n50273 = n30718 ^ n4340 ^ 1'b0 ;
  assign n50272 = ( ~n13099 & n21856 ) | ( ~n13099 & n24480 ) | ( n21856 & n24480 ) ;
  assign n50274 = n50273 ^ n50272 ^ n3275 ;
  assign n50276 = n50275 ^ n50274 ^ n10962 ;
  assign n50277 = n20915 ^ n15623 ^ n9729 ;
  assign n50278 = n50277 ^ n42154 ^ n20810 ;
  assign n50280 = n6660 ^ n1544 ^ n849 ;
  assign n50279 = n10799 | n24778 ;
  assign n50281 = n50280 ^ n50279 ^ n18299 ;
  assign n50282 = n47014 ^ n10459 ^ n6160 ;
  assign n50283 = ( n11977 & n17110 ) | ( n11977 & n25845 ) | ( n17110 & n25845 ) ;
  assign n50285 = n21285 ^ n9542 ^ 1'b0 ;
  assign n50284 = ~n19310 & n37705 ;
  assign n50286 = n50285 ^ n50284 ^ n19714 ;
  assign n50287 = n10777 & ~n16359 ;
  assign n50288 = ~n44706 & n50287 ;
  assign n50289 = n48260 ^ n32566 ^ n3702 ;
  assign n50290 = n5081 & ~n50289 ;
  assign n50291 = n44295 & n50290 ;
  assign n50292 = n1231 & n5195 ;
  assign n50293 = n957 & n50292 ;
  assign n50294 = ( n23043 & n26564 ) | ( n23043 & n50293 ) | ( n26564 & n50293 ) ;
  assign n50295 = ( n2516 & n2919 ) | ( n2516 & n26877 ) | ( n2919 & n26877 ) ;
  assign n50296 = ( n24879 & ~n26651 ) | ( n24879 & n37736 ) | ( ~n26651 & n37736 ) ;
  assign n50297 = ( n3249 & n50295 ) | ( n3249 & n50296 ) | ( n50295 & n50296 ) ;
  assign n50298 = ( ~n17039 & n35329 ) | ( ~n17039 & n42618 ) | ( n35329 & n42618 ) ;
  assign n50299 = ( n10459 & n12746 ) | ( n10459 & ~n14910 ) | ( n12746 & ~n14910 ) ;
  assign n50300 = n50299 ^ n12605 ^ n5448 ;
  assign n50301 = ( n10393 & n32512 ) | ( n10393 & n50300 ) | ( n32512 & n50300 ) ;
  assign n50302 = ~n19239 & n43388 ;
  assign n50303 = n23651 ^ n11866 ^ n11055 ;
  assign n50304 = n46383 | n50303 ;
  assign n50305 = n10659 | n50304 ;
  assign n50306 = n50305 ^ n47952 ^ n11105 ;
  assign n50307 = ( ~n28594 & n36286 ) | ( ~n28594 & n40086 ) | ( n36286 & n40086 ) ;
  assign n50309 = n13514 | n16768 ;
  assign n50310 = n50309 ^ n16491 ^ 1'b0 ;
  assign n50308 = n16975 & ~n44569 ;
  assign n50311 = n50310 ^ n50308 ^ 1'b0 ;
  assign n50312 = n22321 ^ n14861 ^ n9738 ;
  assign n50313 = ( ~n6330 & n11922 ) | ( ~n6330 & n50312 ) | ( n11922 & n50312 ) ;
  assign n50314 = n50313 ^ x219 ^ 1'b0 ;
  assign n50315 = n24846 ^ n12173 ^ n1981 ;
  assign n50316 = ( n7386 & n32169 ) | ( n7386 & n50315 ) | ( n32169 & n50315 ) ;
  assign n50317 = n50316 ^ n36752 ^ 1'b0 ;
  assign n50318 = n1850 | n50317 ;
  assign n50319 = n47384 ^ n9333 ^ 1'b0 ;
  assign n50320 = n44792 ^ n43981 ^ n43078 ;
  assign n50321 = ( n7107 & n16344 ) | ( n7107 & ~n34295 ) | ( n16344 & ~n34295 ) ;
  assign n50322 = ( n5566 & ~n23302 ) | ( n5566 & n50321 ) | ( ~n23302 & n50321 ) ;
  assign n50324 = n42291 ^ n8760 ^ n2711 ;
  assign n50323 = ( n980 & n18136 ) | ( n980 & n41915 ) | ( n18136 & n41915 ) ;
  assign n50325 = n50324 ^ n50323 ^ n23509 ;
  assign n50326 = ( n34767 & n41222 ) | ( n34767 & ~n45993 ) | ( n41222 & ~n45993 ) ;
  assign n50327 = n41652 ^ n32718 ^ n30557 ;
  assign n50328 = ( n9790 & ~n10599 ) | ( n9790 & n29664 ) | ( ~n10599 & n29664 ) ;
  assign n50329 = ( n26748 & ~n50327 ) | ( n26748 & n50328 ) | ( ~n50327 & n50328 ) ;
  assign n50332 = n23979 ^ n5368 ^ n3076 ;
  assign n50330 = n20175 ^ n11666 ^ 1'b0 ;
  assign n50331 = n11607 & n50330 ;
  assign n50333 = n50332 ^ n50331 ^ 1'b0 ;
  assign n50334 = n5029 & n18536 ;
  assign n50335 = n50334 ^ n18947 ^ 1'b0 ;
  assign n50336 = n13142 | n41682 ;
  assign n50337 = n2747 | n13019 ;
  assign n50338 = n50337 ^ n50152 ^ 1'b0 ;
  assign n50339 = ~n8730 & n50338 ;
  assign n50340 = n39168 & n50339 ;
  assign n50341 = n17295 & ~n27928 ;
  assign n50342 = n50341 ^ n9305 ^ 1'b0 ;
  assign n50343 = ( ~n13637 & n36357 ) | ( ~n13637 & n50342 ) | ( n36357 & n50342 ) ;
  assign n50347 = n11545 ^ n6467 ^ n1436 ;
  assign n50346 = ( n1968 & n11262 ) | ( n1968 & ~n41412 ) | ( n11262 & ~n41412 ) ;
  assign n50344 = ~n41843 & n48458 ;
  assign n50345 = ~n3894 & n50344 ;
  assign n50348 = n50347 ^ n50346 ^ n50345 ;
  assign n50349 = n37113 ^ n2554 ^ 1'b0 ;
  assign n50350 = n6199 & n50349 ;
  assign n50351 = n21987 ^ n9926 ^ n7691 ;
  assign n50354 = n3991 | n21016 ;
  assign n50355 = ( n14078 & n16210 ) | ( n14078 & ~n50354 ) | ( n16210 & ~n50354 ) ;
  assign n50352 = n32235 ^ n1771 ^ 1'b0 ;
  assign n50353 = ( ~n18175 & n27788 ) | ( ~n18175 & n50352 ) | ( n27788 & n50352 ) ;
  assign n50356 = n50355 ^ n50353 ^ n6326 ;
  assign n50357 = ( n10765 & n14008 ) | ( n10765 & n31893 ) | ( n14008 & n31893 ) ;
  assign n50358 = n49912 ^ n6546 ^ 1'b0 ;
  assign n50359 = n1317 & ~n42452 ;
  assign n50360 = n50359 ^ n35110 ^ 1'b0 ;
  assign n50361 = n9486 & n13267 ;
  assign n50362 = ~n3848 & n50361 ;
  assign n50363 = n23422 ^ n21051 ^ 1'b0 ;
  assign n50364 = n50362 | n50363 ;
  assign n50365 = ( n11949 & n17108 ) | ( n11949 & ~n28445 ) | ( n17108 & ~n28445 ) ;
  assign n50366 = ( n13117 & ~n35229 ) | ( n13117 & n50365 ) | ( ~n35229 & n50365 ) ;
  assign n50367 = ( ~n15388 & n28828 ) | ( ~n15388 & n43676 ) | ( n28828 & n43676 ) ;
  assign n50368 = n47846 ^ n9221 ^ n6262 ;
  assign n50369 = n50368 ^ n34299 ^ n9129 ;
  assign n50370 = ( ~n15602 & n26480 ) | ( ~n15602 & n30792 ) | ( n26480 & n30792 ) ;
  assign n50371 = n42500 ^ n31914 ^ n355 ;
  assign n50372 = ( n8918 & n25761 ) | ( n8918 & n32123 ) | ( n25761 & n32123 ) ;
  assign n50373 = n25349 & n50372 ;
  assign n50374 = n50373 ^ n39070 ^ n31895 ;
  assign n50375 = n42601 ^ n38767 ^ n35301 ;
  assign n50376 = n27189 ^ n22429 ^ n15847 ;
  assign n50377 = n5948 & n17835 ;
  assign n50378 = n50377 ^ n12580 ^ 1'b0 ;
  assign n50379 = n24341 & n45889 ;
  assign n50380 = ~n8748 & n50379 ;
  assign n50388 = n45533 ^ n29739 ^ n17742 ;
  assign n50384 = n5370 ^ n4066 ^ n2706 ;
  assign n50381 = n9927 ^ n8472 ^ 1'b0 ;
  assign n50382 = n28310 | n50381 ;
  assign n50383 = ( n21543 & n28438 ) | ( n21543 & n50382 ) | ( n28438 & n50382 ) ;
  assign n50385 = n50384 ^ n50383 ^ n3086 ;
  assign n50386 = n50385 ^ n1157 ^ 1'b0 ;
  assign n50387 = ~n19703 & n50386 ;
  assign n50389 = n50388 ^ n50387 ^ 1'b0 ;
  assign n50390 = n24884 ^ n10704 ^ n5733 ;
  assign n50394 = ( ~x160 & n23189 ) | ( ~x160 & n27898 ) | ( n23189 & n27898 ) ;
  assign n50391 = n28470 ^ n10395 ^ n10320 ;
  assign n50392 = ( ~n2825 & n31865 ) | ( ~n2825 & n50391 ) | ( n31865 & n50391 ) ;
  assign n50393 = ~n5624 & n50392 ;
  assign n50395 = n50394 ^ n50393 ^ 1'b0 ;
  assign n50396 = n50395 ^ n26896 ^ n3367 ;
  assign n50397 = ~n13918 & n50396 ;
  assign n50398 = ( ~n21026 & n21824 ) | ( ~n21026 & n45404 ) | ( n21824 & n45404 ) ;
  assign n50399 = n50398 ^ n21904 ^ 1'b0 ;
  assign n50400 = n13023 ^ n5912 ^ n337 ;
  assign n50401 = ( ~n17151 & n34878 ) | ( ~n17151 & n50400 ) | ( n34878 & n50400 ) ;
  assign n50402 = n25459 ^ n12953 ^ n7854 ;
  assign n50403 = n26282 ^ n15235 ^ n3942 ;
  assign n50404 = ( n30385 & n36551 ) | ( n30385 & n44506 ) | ( n36551 & n44506 ) ;
  assign n50405 = n50404 ^ n14500 ^ n13853 ;
  assign n50406 = ( n40186 & n50403 ) | ( n40186 & ~n50405 ) | ( n50403 & ~n50405 ) ;
  assign n50408 = ( n3880 & n21819 ) | ( n3880 & n26368 ) | ( n21819 & n26368 ) ;
  assign n50407 = n32218 ^ n16334 ^ n8343 ;
  assign n50409 = n50408 ^ n50407 ^ n9940 ;
  assign n50410 = n31117 ^ n6741 ^ 1'b0 ;
  assign n50411 = n32353 ^ n2551 ^ 1'b0 ;
  assign n50412 = ~n50410 & n50411 ;
  assign n50413 = n23190 & ~n39918 ;
  assign n50414 = ~n50412 & n50413 ;
  assign n50415 = ( n17550 & ~n31287 ) | ( n17550 & n36630 ) | ( ~n31287 & n36630 ) ;
  assign n50416 = n50415 ^ n3980 ^ 1'b0 ;
  assign n50417 = n6781 & n50416 ;
  assign n50420 = n20539 ^ n1434 ^ n970 ;
  assign n50418 = n4472 & n33778 ;
  assign n50419 = ~n29726 & n50418 ;
  assign n50421 = n50420 ^ n50419 ^ n2930 ;
  assign n50422 = n28061 ^ n16244 ^ 1'b0 ;
  assign n50423 = ( n1594 & n4440 ) | ( n1594 & n26684 ) | ( n4440 & n26684 ) ;
  assign n50424 = ( ~n16709 & n47658 ) | ( ~n16709 & n50423 ) | ( n47658 & n50423 ) ;
  assign n50427 = ( ~n766 & n9251 ) | ( ~n766 & n34054 ) | ( n9251 & n34054 ) ;
  assign n50425 = n4245 & n41115 ;
  assign n50426 = n7374 & ~n50425 ;
  assign n50428 = n50427 ^ n50426 ^ 1'b0 ;
  assign n50429 = ( n22196 & n35009 ) | ( n22196 & n36339 ) | ( n35009 & n36339 ) ;
  assign n50430 = ( ~n33134 & n50428 ) | ( ~n33134 & n50429 ) | ( n50428 & n50429 ) ;
  assign n50431 = n15757 ^ n7212 ^ 1'b0 ;
  assign n50432 = ( n33458 & n43835 ) | ( n33458 & n50431 ) | ( n43835 & n50431 ) ;
  assign n50433 = n50432 ^ n31912 ^ n13123 ;
  assign n50434 = n37955 ^ n9309 ^ n3824 ;
  assign n50435 = n50434 ^ n6512 ^ 1'b0 ;
  assign n50436 = ~n21779 & n50435 ;
  assign n50437 = ( ~n13006 & n17092 ) | ( ~n13006 & n50436 ) | ( n17092 & n50436 ) ;
  assign n50438 = n18664 ^ n14210 ^ n14072 ;
  assign n50439 = ( ~n7083 & n7235 ) | ( ~n7083 & n36918 ) | ( n7235 & n36918 ) ;
  assign n50440 = ( n8366 & n50438 ) | ( n8366 & n50439 ) | ( n50438 & n50439 ) ;
  assign n50441 = n19343 ^ n13176 ^ 1'b0 ;
  assign n50442 = n50441 ^ n47041 ^ n23632 ;
  assign n50443 = n50442 ^ n29843 ^ n7258 ;
  assign n50444 = n26579 ^ n2150 ^ 1'b0 ;
  assign n50445 = n8549 | n48928 ;
  assign n50446 = n26384 | n50445 ;
  assign n50447 = n2686 & ~n35952 ;
  assign n50448 = n29718 & n41056 ;
  assign n50451 = n15604 ^ n7048 ^ 1'b0 ;
  assign n50452 = n50451 ^ n2586 ^ n2516 ;
  assign n50449 = n23671 ^ n19247 ^ 1'b0 ;
  assign n50450 = n39846 | n50449 ;
  assign n50453 = n50452 ^ n50450 ^ n21257 ;
  assign n50454 = ( n24243 & n50448 ) | ( n24243 & n50453 ) | ( n50448 & n50453 ) ;
  assign n50455 = n45710 ^ n9476 ^ n8258 ;
  assign n50456 = n36083 ^ n30429 ^ n12733 ;
  assign n50457 = n28595 ^ n3918 ^ 1'b0 ;
  assign n50458 = n7699 & n50457 ;
  assign n50459 = ( n3756 & ~n5665 ) | ( n3756 & n10882 ) | ( ~n5665 & n10882 ) ;
  assign n50460 = ( n13142 & n43987 ) | ( n13142 & n50459 ) | ( n43987 & n50459 ) ;
  assign n50461 = n4905 & n16222 ;
  assign n50462 = ~n16968 & n50461 ;
  assign n50463 = n38972 & ~n50462 ;
  assign n50464 = ~n20014 & n50463 ;
  assign n50465 = n21343 ^ n9642 ^ n1255 ;
  assign n50466 = n18536 & ~n50465 ;
  assign n50467 = ~n16746 & n50466 ;
  assign n50468 = n17627 | n25482 ;
  assign n50469 = n8116 | n50468 ;
  assign n50470 = ( n21034 & n26655 ) | ( n21034 & ~n44558 ) | ( n26655 & ~n44558 ) ;
  assign n50471 = ~n13423 & n29905 ;
  assign n50472 = n50471 ^ n28369 ^ n6519 ;
  assign n50473 = n23948 ^ n18974 ^ n8365 ;
  assign n50474 = ( n43104 & ~n47931 ) | ( n43104 & n50473 ) | ( ~n47931 & n50473 ) ;
  assign n50475 = n15017 ^ n11985 ^ 1'b0 ;
  assign n50476 = ( n1314 & n5510 ) | ( n1314 & ~n14610 ) | ( n5510 & ~n14610 ) ;
  assign n50477 = ( n4466 & n26056 ) | ( n4466 & ~n50476 ) | ( n26056 & ~n50476 ) ;
  assign n50478 = ~n12622 & n50477 ;
  assign n50479 = ( n1692 & n18670 ) | ( n1692 & n50478 ) | ( n18670 & n50478 ) ;
  assign n50480 = ( n9557 & n21151 ) | ( n9557 & ~n35806 ) | ( n21151 & ~n35806 ) ;
  assign n50481 = n4405 & n21870 ;
  assign n50482 = n50481 ^ n5338 ^ n4257 ;
  assign n50483 = n50482 ^ n33604 ^ n11374 ;
  assign n50484 = n45786 | n50483 ;
  assign n50485 = n3893 ^ n3468 ^ n2654 ;
  assign n50486 = n50485 ^ n8638 ^ n5875 ;
  assign n50487 = n50486 ^ n14480 ^ n13686 ;
  assign n50488 = ~n19147 & n44970 ;
  assign n50489 = n33450 & n50488 ;
  assign n50490 = n39452 ^ n17890 ^ 1'b0 ;
  assign n50491 = n35426 & ~n50490 ;
  assign n50492 = ~n16555 & n40018 ;
  assign n50493 = n50492 ^ n48629 ^ 1'b0 ;
  assign n50494 = n43002 ^ n21215 ^ 1'b0 ;
  assign n50495 = ( n17493 & ~n19974 ) | ( n17493 & n50494 ) | ( ~n19974 & n50494 ) ;
  assign n50496 = n36984 & ~n50495 ;
  assign n50497 = n50496 ^ n14892 ^ n1382 ;
  assign n50500 = ( n1105 & n15714 ) | ( n1105 & n39762 ) | ( n15714 & n39762 ) ;
  assign n50498 = n41385 ^ n11420 ^ n3521 ;
  assign n50499 = n50498 ^ n24942 ^ n1798 ;
  assign n50501 = n50500 ^ n50499 ^ n11419 ;
  assign n50502 = ( n16592 & n26013 ) | ( n16592 & n50501 ) | ( n26013 & n50501 ) ;
  assign n50503 = ( ~n12802 & n15163 ) | ( ~n12802 & n48900 ) | ( n15163 & n48900 ) ;
  assign n50504 = n9723 & ~n50503 ;
  assign n50505 = n50504 ^ n24921 ^ n16421 ;
  assign n50506 = ( ~n29339 & n37736 ) | ( ~n29339 & n42307 ) | ( n37736 & n42307 ) ;
  assign n50507 = ( n747 & n33615 ) | ( n747 & n50506 ) | ( n33615 & n50506 ) ;
  assign n50508 = n34612 ^ n21957 ^ n5077 ;
  assign n50509 = ( n10262 & n17589 ) | ( n10262 & ~n32252 ) | ( n17589 & ~n32252 ) ;
  assign n50510 = ( n19808 & ~n50508 ) | ( n19808 & n50509 ) | ( ~n50508 & n50509 ) ;
  assign n50511 = n50510 ^ n27820 ^ n24877 ;
  assign n50512 = ( n12287 & n50507 ) | ( n12287 & ~n50511 ) | ( n50507 & ~n50511 ) ;
  assign n50513 = n49402 ^ n24186 ^ n9871 ;
  assign n50514 = n50513 ^ n47658 ^ x71 ;
  assign n50515 = ( ~n13564 & n25038 ) | ( ~n13564 & n50514 ) | ( n25038 & n50514 ) ;
  assign n50516 = n30467 ^ n7577 ^ n6897 ;
  assign n50517 = ( ~n7450 & n19686 ) | ( ~n7450 & n47570 ) | ( n19686 & n47570 ) ;
  assign n50518 = ( n4854 & n30407 ) | ( n4854 & n50009 ) | ( n30407 & n50009 ) ;
  assign n50519 = ( ~n14117 & n15168 ) | ( ~n14117 & n50518 ) | ( n15168 & n50518 ) ;
  assign n50520 = n50519 ^ n37754 ^ n11116 ;
  assign n50521 = n50520 ^ n37005 ^ n905 ;
  assign n50522 = ( n8260 & n22688 ) | ( n8260 & n30476 ) | ( n22688 & n30476 ) ;
  assign n50523 = ~n37663 & n50522 ;
  assign n50524 = ~n26891 & n50523 ;
  assign n50525 = n31729 & ~n39808 ;
  assign n50526 = ~n13802 & n50525 ;
  assign n50527 = n44294 ^ n5911 ^ 1'b0 ;
  assign n50528 = n7779 ^ n4452 ^ n3636 ;
  assign n50529 = n15440 & n19951 ;
  assign n50530 = n50529 ^ n3478 ^ 1'b0 ;
  assign n50531 = ( n8167 & n17869 ) | ( n8167 & ~n50530 ) | ( n17869 & ~n50530 ) ;
  assign n50532 = n50531 ^ n16137 ^ n9595 ;
  assign n50533 = ( ~n9430 & n16295 ) | ( ~n9430 & n50532 ) | ( n16295 & n50532 ) ;
  assign n50534 = ( n22547 & ~n50528 ) | ( n22547 & n50533 ) | ( ~n50528 & n50533 ) ;
  assign n50535 = n15767 ^ n2782 ^ 1'b0 ;
  assign n50536 = n6653 | n50535 ;
  assign n50537 = n50536 ^ n28836 ^ n14308 ;
  assign n50539 = ( n15003 & n15168 ) | ( n15003 & n18742 ) | ( n15168 & n18742 ) ;
  assign n50538 = ( x51 & n1274 ) | ( x51 & n42412 ) | ( n1274 & n42412 ) ;
  assign n50540 = n50539 ^ n50538 ^ n45933 ;
  assign n50541 = n46246 | n47710 ;
  assign n50542 = n14461 & ~n26827 ;
  assign n50543 = ~n50541 & n50542 ;
  assign n50544 = ( n15685 & ~n23126 ) | ( n15685 & n50543 ) | ( ~n23126 & n50543 ) ;
  assign n50545 = n19701 ^ n12244 ^ n6804 ;
  assign n50546 = ( n1569 & n25980 ) | ( n1569 & ~n50545 ) | ( n25980 & ~n50545 ) ;
  assign n50547 = n16615 ^ n7001 ^ 1'b0 ;
  assign n50548 = n20215 & n25266 ;
  assign n50549 = n28235 | n40450 ;
  assign n50550 = n50548 | n50549 ;
  assign n50551 = ( n14099 & ~n50547 ) | ( n14099 & n50550 ) | ( ~n50547 & n50550 ) ;
  assign n50552 = ( ~n14316 & n19651 ) | ( ~n14316 & n23797 ) | ( n19651 & n23797 ) ;
  assign n50553 = n50552 ^ n39210 ^ n27617 ;
  assign n50554 = n46476 ^ n36497 ^ 1'b0 ;
  assign n50555 = ~n20005 & n50554 ;
  assign n50556 = ( n8971 & n9222 ) | ( n8971 & ~n12228 ) | ( n9222 & ~n12228 ) ;
  assign n50557 = n30659 ^ n13738 ^ n7040 ;
  assign n50558 = ~n5769 & n50557 ;
  assign n50559 = n50556 & n50558 ;
  assign n50560 = n9576 ^ n893 ^ 1'b0 ;
  assign n50561 = n24510 & n50560 ;
  assign n50562 = ( n15976 & n20068 ) | ( n15976 & ~n40445 ) | ( n20068 & ~n40445 ) ;
  assign n50563 = ( n2628 & n35338 ) | ( n2628 & ~n50562 ) | ( n35338 & ~n50562 ) ;
  assign n50564 = n48032 ^ n27447 ^ n13496 ;
  assign n50565 = n50564 ^ n43322 ^ n17807 ;
  assign n50566 = n28668 & ~n50565 ;
  assign n50567 = ( n7355 & n15239 ) | ( n7355 & ~n33447 ) | ( n15239 & ~n33447 ) ;
  assign n50568 = ~n3077 & n50567 ;
  assign n50569 = ( n5311 & n7268 ) | ( n5311 & ~n12228 ) | ( n7268 & ~n12228 ) ;
  assign n50570 = n50569 ^ n25079 ^ n15356 ;
  assign n50571 = n49687 ^ n46461 ^ n1202 ;
  assign n50572 = n50571 ^ n37098 ^ n22140 ;
  assign n50573 = n50572 ^ n4901 ^ x239 ;
  assign n50574 = n37262 ^ n30254 ^ n18652 ;
  assign n50575 = ( ~n564 & n16933 ) | ( ~n564 & n50574 ) | ( n16933 & n50574 ) ;
  assign n50576 = n27794 ^ n8417 ^ n3225 ;
  assign n50578 = ~n19117 & n19552 ;
  assign n50579 = n50578 ^ n15916 ^ 1'b0 ;
  assign n50577 = n6456 | n23925 ;
  assign n50580 = n50579 ^ n50577 ^ 1'b0 ;
  assign n50581 = n3105 & ~n6914 ;
  assign n50582 = n50581 ^ n4313 ^ 1'b0 ;
  assign n50587 = ( n2487 & n3129 ) | ( n2487 & ~n11695 ) | ( n3129 & ~n11695 ) ;
  assign n50586 = n37772 ^ n17625 ^ 1'b0 ;
  assign n50583 = n34487 ^ n33412 ^ n24712 ;
  assign n50584 = n50583 ^ n20085 ^ n15839 ;
  assign n50585 = ( ~n17779 & n20704 ) | ( ~n17779 & n50584 ) | ( n20704 & n50584 ) ;
  assign n50588 = n50587 ^ n50586 ^ n50585 ;
  assign n50589 = n50588 ^ n38323 ^ 1'b0 ;
  assign n50590 = n37320 ^ n13728 ^ n7443 ;
  assign n50591 = n50590 ^ n47897 ^ 1'b0 ;
  assign n50592 = n39284 ^ n17451 ^ n13817 ;
  assign n50593 = n50592 ^ n16359 ^ 1'b0 ;
  assign n50594 = n50593 ^ n31226 ^ n12000 ;
  assign n50595 = ( n12363 & n34182 ) | ( n12363 & ~n35420 ) | ( n34182 & ~n35420 ) ;
  assign n50596 = n50595 ^ n36352 ^ 1'b0 ;
  assign n50597 = n50596 ^ n13201 ^ n7515 ;
  assign n50598 = ( n5785 & n6741 ) | ( n5785 & n15282 ) | ( n6741 & n15282 ) ;
  assign n50599 = n50598 ^ n26155 ^ n905 ;
  assign n50600 = ( n3353 & n5237 ) | ( n3353 & ~n10339 ) | ( n5237 & ~n10339 ) ;
  assign n50601 = n7172 ^ n6461 ^ n5010 ;
  assign n50602 = ( n40066 & n50600 ) | ( n40066 & ~n50601 ) | ( n50600 & ~n50601 ) ;
  assign n50605 = n3163 ^ n2802 ^ n1216 ;
  assign n50603 = n11185 & ~n20422 ;
  assign n50604 = n50603 ^ n11486 ^ 1'b0 ;
  assign n50606 = n50605 ^ n50604 ^ n27086 ;
  assign n50607 = n50606 ^ n21775 ^ 1'b0 ;
  assign n50608 = n35257 | n50607 ;
  assign n50609 = n4159 & n12853 ;
  assign n50610 = n50609 ^ n14360 ^ 1'b0 ;
  assign n50611 = n45198 ^ n16685 ^ n6649 ;
  assign n50612 = n24231 ^ n9177 ^ 1'b0 ;
  assign n50613 = ( ~n4686 & n14628 ) | ( ~n4686 & n50612 ) | ( n14628 & n50612 ) ;
  assign n50614 = n25775 | n38483 ;
  assign n50615 = n35065 & ~n50614 ;
  assign n50616 = n50615 ^ n11445 ^ n2440 ;
  assign n50618 = n12520 ^ n9587 ^ x144 ;
  assign n50619 = n612 | n50618 ;
  assign n50620 = n21444 & ~n50619 ;
  assign n50617 = ( n6789 & n26457 ) | ( n6789 & n28935 ) | ( n26457 & n28935 ) ;
  assign n50621 = n50620 ^ n50617 ^ n11040 ;
  assign n50622 = n50621 ^ n33773 ^ n24827 ;
  assign n50626 = ( ~n8839 & n12214 ) | ( ~n8839 & n21701 ) | ( n12214 & n21701 ) ;
  assign n50623 = n6953 & n24583 ;
  assign n50624 = ~n12191 & n50623 ;
  assign n50625 = ( ~n9955 & n16100 ) | ( ~n9955 & n50624 ) | ( n16100 & n50624 ) ;
  assign n50627 = n50626 ^ n50625 ^ n31957 ;
  assign n50630 = ( n6709 & ~n10649 ) | ( n6709 & n17356 ) | ( ~n10649 & n17356 ) ;
  assign n50631 = n50630 ^ n23192 ^ n22788 ;
  assign n50629 = n36009 ^ n17234 ^ 1'b0 ;
  assign n50628 = ( ~n5288 & n42111 ) | ( ~n5288 & n47001 ) | ( n42111 & n47001 ) ;
  assign n50632 = n50631 ^ n50629 ^ n50628 ;
  assign n50633 = n13264 | n38616 ;
  assign n50634 = n4472 | n50633 ;
  assign n50635 = n11006 | n50634 ;
  assign n50636 = n3545 | n36570 ;
  assign n50637 = n50636 ^ n20118 ^ 1'b0 ;
  assign n50638 = n50637 ^ n47433 ^ n12303 ;
  assign n50639 = n21174 ^ x235 ^ 1'b0 ;
  assign n50640 = n33166 | n50138 ;
  assign n50641 = ~n7934 & n18288 ;
  assign n50642 = n50641 ^ n6185 ^ 1'b0 ;
  assign n50643 = n46742 ^ n24340 ^ n1453 ;
  assign n50644 = ( n8067 & ~n15862 ) | ( n8067 & n29059 ) | ( ~n15862 & n29059 ) ;
  assign n50645 = ( n6641 & ~n17559 ) | ( n6641 & n41735 ) | ( ~n17559 & n41735 ) ;
  assign n50646 = n36717 ^ n32014 ^ n31114 ;
  assign n50647 = ( n28668 & n37548 ) | ( n28668 & ~n50646 ) | ( n37548 & ~n50646 ) ;
  assign n50648 = ( ~n3668 & n7139 ) | ( ~n3668 & n32116 ) | ( n7139 & n32116 ) ;
  assign n50649 = n50648 ^ n17639 ^ n9868 ;
  assign n50650 = n8801 ^ n689 ^ 1'b0 ;
  assign n50651 = ~n4877 & n50650 ;
  assign n50652 = n48499 ^ n19519 ^ n18060 ;
  assign n50657 = n21505 ^ n16799 ^ n13627 ;
  assign n50653 = n11156 | n13290 ;
  assign n50654 = n50653 ^ n10954 ^ 1'b0 ;
  assign n50655 = ( n12157 & ~n13754 ) | ( n12157 & n32775 ) | ( ~n13754 & n32775 ) ;
  assign n50656 = ( n14099 & ~n50654 ) | ( n14099 & n50655 ) | ( ~n50654 & n50655 ) ;
  assign n50658 = n50657 ^ n50656 ^ n37553 ;
  assign n50659 = ~n399 & n20711 ;
  assign n50660 = n49923 & n50659 ;
  assign n50661 = ~n12667 & n36752 ;
  assign n50662 = n50661 ^ n49717 ^ n27373 ;
  assign n50663 = ( ~n12715 & n17622 ) | ( ~n12715 & n26898 ) | ( n17622 & n26898 ) ;
  assign n50664 = n24690 ^ n20128 ^ 1'b0 ;
  assign n50665 = ( n24617 & n26097 ) | ( n24617 & ~n41489 ) | ( n26097 & ~n41489 ) ;
  assign n50666 = ~n16786 & n39231 ;
  assign n50667 = n50666 ^ n33921 ^ 1'b0 ;
  assign n50668 = n29628 ^ n15236 ^ 1'b0 ;
  assign n50669 = n50668 ^ n28852 ^ n16106 ;
  assign n50670 = ( n3785 & n6124 ) | ( n3785 & n27791 ) | ( n6124 & n27791 ) ;
  assign n50671 = n49189 ^ n23150 ^ n20079 ;
  assign n50672 = n2451 | n50671 ;
  assign n50673 = n32211 & ~n50672 ;
  assign n50674 = ( ~n24181 & n50670 ) | ( ~n24181 & n50673 ) | ( n50670 & n50673 ) ;
  assign n50675 = ( ~n1987 & n10554 ) | ( ~n1987 & n18486 ) | ( n10554 & n18486 ) ;
  assign n50676 = n50675 ^ n17413 ^ 1'b0 ;
  assign n50677 = n23385 ^ n12254 ^ n2873 ;
  assign n50678 = n50677 ^ n11679 ^ 1'b0 ;
  assign n50680 = n16023 ^ n8129 ^ n5050 ;
  assign n50679 = n50383 ^ n27035 ^ n10558 ;
  assign n50681 = n50680 ^ n50679 ^ n20752 ;
  assign n50682 = n22538 ^ n5156 ^ n4787 ;
  assign n50683 = ( n5035 & n6407 ) | ( n5035 & ~n15195 ) | ( n6407 & ~n15195 ) ;
  assign n50684 = ( n17001 & n27477 ) | ( n17001 & n46842 ) | ( n27477 & n46842 ) ;
  assign n50685 = n50684 ^ n22386 ^ 1'b0 ;
  assign n50686 = ( n15947 & n25700 ) | ( n15947 & n29785 ) | ( n25700 & n29785 ) ;
  assign n50687 = n30343 | n50686 ;
  assign n50688 = n10900 | n50687 ;
  assign n50689 = n18736 ^ n14982 ^ n5162 ;
  assign n50690 = n9649 & ~n19617 ;
  assign n50691 = ~n50689 & n50690 ;
  assign n50692 = n24834 | n26544 ;
  assign n50693 = n50692 ^ n34893 ^ n7379 ;
  assign n50694 = ( n9325 & ~n14980 ) | ( n9325 & n14992 ) | ( ~n14980 & n14992 ) ;
  assign n50695 = n38351 & n50694 ;
  assign n50696 = ( n6975 & n13142 ) | ( n6975 & n24192 ) | ( n13142 & n24192 ) ;
  assign n50697 = n50696 ^ n26162 ^ n8981 ;
  assign n50698 = n50697 ^ n8123 ^ n7439 ;
  assign n50699 = n19826 & ~n28597 ;
  assign n50700 = ( n14013 & n25690 ) | ( n14013 & ~n50699 ) | ( n25690 & ~n50699 ) ;
  assign n50701 = ( ~n3486 & n22615 ) | ( ~n3486 & n50700 ) | ( n22615 & n50700 ) ;
  assign n50702 = n10099 & ~n26421 ;
  assign n50703 = n50702 ^ n31418 ^ n18940 ;
  assign n50704 = ~n9889 & n27934 ;
  assign n50705 = n50704 ^ n50498 ^ n43842 ;
  assign n50706 = ( ~n11202 & n20805 ) | ( ~n11202 & n50705 ) | ( n20805 & n50705 ) ;
  assign n50707 = n4609 | n36981 ;
  assign n50708 = ( n10187 & n28403 ) | ( n10187 & ~n50707 ) | ( n28403 & ~n50707 ) ;
  assign n50709 = ( n10934 & n14193 ) | ( n10934 & n16905 ) | ( n14193 & n16905 ) ;
  assign n50710 = n50709 ^ n8087 ^ n5978 ;
  assign n50711 = n6132 & n19643 ;
  assign n50712 = n25161 | n30947 ;
  assign n50713 = n2755 & ~n50712 ;
  assign n50714 = n18467 ^ n14114 ^ 1'b0 ;
  assign n50715 = ~n17664 & n34671 ;
  assign n50716 = n50715 ^ n2452 ^ 1'b0 ;
  assign n50717 = ( ~n21668 & n25073 ) | ( ~n21668 & n50716 ) | ( n25073 & n50716 ) ;
  assign n50718 = n25698 ^ n24660 ^ n6591 ;
  assign n50719 = ( n13081 & n16522 ) | ( n13081 & ~n36042 ) | ( n16522 & ~n36042 ) ;
  assign n50720 = n2738 & n28509 ;
  assign n50721 = n41408 & n50720 ;
  assign n50722 = ( ~n9911 & n50719 ) | ( ~n9911 & n50721 ) | ( n50719 & n50721 ) ;
  assign n50726 = n48326 ^ n31243 ^ 1'b0 ;
  assign n50727 = n48663 & ~n50726 ;
  assign n50723 = n24895 ^ n10103 ^ 1'b0 ;
  assign n50724 = n22370 ^ n10429 ^ 1'b0 ;
  assign n50725 = n50723 & n50724 ;
  assign n50728 = n50727 ^ n50725 ^ n3163 ;
  assign n50729 = n27945 ^ n26059 ^ 1'b0 ;
  assign n50730 = n14101 | n50729 ;
  assign n50731 = ( n6991 & ~n18749 ) | ( n6991 & n50730 ) | ( ~n18749 & n50730 ) ;
  assign n50732 = n11692 | n24578 ;
  assign n50733 = ( n5940 & n14466 ) | ( n5940 & n19817 ) | ( n14466 & n19817 ) ;
  assign n50734 = ( n38979 & n50732 ) | ( n38979 & n50733 ) | ( n50732 & n50733 ) ;
  assign n50735 = n5921 | n13467 ;
  assign n50736 = ( ~n34088 & n35683 ) | ( ~n34088 & n50735 ) | ( n35683 & n50735 ) ;
  assign n50737 = ( ~n1577 & n4005 ) | ( ~n1577 & n10143 ) | ( n4005 & n10143 ) ;
  assign n50738 = ( n13909 & ~n27511 ) | ( n13909 & n50737 ) | ( ~n27511 & n50737 ) ;
  assign n50739 = n22843 ^ n10961 ^ n7868 ;
  assign n50740 = ( ~n6884 & n16261 ) | ( ~n6884 & n50739 ) | ( n16261 & n50739 ) ;
  assign n50741 = n50740 ^ n48555 ^ 1'b0 ;
  assign n50742 = n50738 | n50741 ;
  assign n50747 = ~n20499 & n31615 ;
  assign n50748 = ~x181 & n50747 ;
  assign n50743 = ( n7263 & n8343 ) | ( n7263 & ~n27084 ) | ( n8343 & ~n27084 ) ;
  assign n50744 = n31241 | n50743 ;
  assign n50745 = n50744 ^ x30 ^ 1'b0 ;
  assign n50746 = ~n572 & n50745 ;
  assign n50749 = n50748 ^ n50746 ^ 1'b0 ;
  assign n50750 = n9288 ^ n4725 ^ n4066 ;
  assign n50751 = n50750 ^ n36258 ^ n5171 ;
  assign n50752 = n50751 ^ n17388 ^ n14388 ;
  assign n50753 = ( n18704 & n43176 ) | ( n18704 & ~n50752 ) | ( n43176 & ~n50752 ) ;
  assign n50754 = n47856 ^ n14255 ^ 1'b0 ;
  assign n50755 = n23076 ^ n20654 ^ n17815 ;
  assign n50756 = ( ~n14935 & n23466 ) | ( ~n14935 & n32076 ) | ( n23466 & n32076 ) ;
  assign n50757 = n50756 ^ n47586 ^ n24548 ;
  assign n50758 = n50755 & n50757 ;
  assign n50759 = n46185 ^ n31083 ^ n29239 ;
  assign n50760 = n5692 & ~n40582 ;
  assign n50761 = n50760 ^ n47516 ^ 1'b0 ;
  assign n50762 = ~n22600 & n36179 ;
  assign n50763 = n50761 & n50762 ;
  assign n50764 = ( n37001 & n47471 ) | ( n37001 & n50763 ) | ( n47471 & n50763 ) ;
  assign n50765 = n2677 & n18698 ;
  assign n50766 = n50765 ^ n3874 ^ 1'b0 ;
  assign n50767 = n9730 & ~n30407 ;
  assign n50768 = n50767 ^ n23319 ^ 1'b0 ;
  assign n50769 = ( n5811 & n6342 ) | ( n5811 & n34432 ) | ( n6342 & n34432 ) ;
  assign n50770 = ~n22251 & n24172 ;
  assign n50771 = n50770 ^ n32328 ^ n17686 ;
  assign n50772 = ( n12179 & ~n47477 ) | ( n12179 & n50771 ) | ( ~n47477 & n50771 ) ;
  assign n50773 = ( ~n44079 & n44286 ) | ( ~n44079 & n47019 ) | ( n44286 & n47019 ) ;
  assign n50774 = n47200 ^ n26765 ^ n5717 ;
  assign n50775 = ( ~n18704 & n28016 ) | ( ~n18704 & n37233 ) | ( n28016 & n37233 ) ;
  assign n50776 = n50775 ^ n49356 ^ 1'b0 ;
  assign n50777 = ( ~n3451 & n33594 ) | ( ~n3451 & n50776 ) | ( n33594 & n50776 ) ;
  assign n50778 = n1270 | n30835 ;
  assign n50779 = ( n15414 & n33801 ) | ( n15414 & ~n50778 ) | ( n33801 & ~n50778 ) ;
  assign n50780 = n26929 ^ n3284 ^ 1'b0 ;
  assign n50783 = n1442 & ~n34119 ;
  assign n50784 = ~n30948 & n50783 ;
  assign n50785 = ( n7806 & n30806 ) | ( n7806 & n50784 ) | ( n30806 & n50784 ) ;
  assign n50781 = ( ~n15465 & n24495 ) | ( ~n15465 & n27516 ) | ( n24495 & n27516 ) ;
  assign n50782 = n50781 ^ n47626 ^ n43105 ;
  assign n50786 = n50785 ^ n50782 ^ n8362 ;
  assign n50787 = n32026 ^ n21139 ^ 1'b0 ;
  assign n50788 = n9222 | n40304 ;
  assign n50789 = n50787 & ~n50788 ;
  assign n50791 = n615 & ~n16940 ;
  assign n50792 = n50791 ^ n33723 ^ 1'b0 ;
  assign n50790 = n18628 & n26829 ;
  assign n50793 = n50792 ^ n50790 ^ 1'b0 ;
  assign n50794 = n27933 ^ n3178 ^ n936 ;
  assign n50795 = n22878 ^ n22583 ^ n20280 ;
  assign n50796 = ( n28318 & n32412 ) | ( n28318 & ~n50055 ) | ( n32412 & ~n50055 ) ;
  assign n50797 = ( n28322 & n50795 ) | ( n28322 & n50796 ) | ( n50795 & n50796 ) ;
  assign n50798 = ( x32 & n21870 ) | ( x32 & ~n33422 ) | ( n21870 & ~n33422 ) ;
  assign n50799 = n6814 | n7819 ;
  assign n50800 = n50799 ^ n42594 ^ 1'b0 ;
  assign n50801 = ( n13017 & n21286 ) | ( n13017 & n50800 ) | ( n21286 & n50800 ) ;
  assign n50802 = ( n3150 & n17446 ) | ( n3150 & ~n26386 ) | ( n17446 & ~n26386 ) ;
  assign n50803 = n50802 ^ n20362 ^ n7165 ;
  assign n50804 = ~n41657 & n45012 ;
  assign n50805 = ( n7804 & ~n16286 ) | ( n7804 & n40512 ) | ( ~n16286 & n40512 ) ;
  assign n50806 = n20695 ^ n6447 ^ n2018 ;
  assign n50807 = n24896 ^ n24653 ^ n22428 ;
  assign n50809 = n26316 ^ n15185 ^ n10435 ;
  assign n50808 = ( n7733 & n8743 ) | ( n7733 & ~n31620 ) | ( n8743 & ~n31620 ) ;
  assign n50810 = n50809 ^ n50808 ^ n8044 ;
  assign n50811 = ( n23495 & n50807 ) | ( n23495 & ~n50810 ) | ( n50807 & ~n50810 ) ;
  assign n50812 = n22593 ^ n19280 ^ 1'b0 ;
  assign n50813 = n7295 & ~n50812 ;
  assign n50814 = ( n50806 & ~n50811 ) | ( n50806 & n50813 ) | ( ~n50811 & n50813 ) ;
  assign n50815 = n29214 ^ n28881 ^ 1'b0 ;
  assign n50816 = ( n697 & n11850 ) | ( n697 & ~n20987 ) | ( n11850 & ~n20987 ) ;
  assign n50817 = n17555 & ~n50816 ;
  assign n50818 = n19033 ^ n14857 ^ 1'b0 ;
  assign n50819 = n17865 & ~n42081 ;
  assign n50820 = ( n30917 & n31175 ) | ( n30917 & ~n37693 ) | ( n31175 & ~n37693 ) ;
  assign n50821 = n17777 & ~n19029 ;
  assign n50822 = n50821 ^ n9834 ^ 1'b0 ;
  assign n50823 = ( n2896 & n4415 ) | ( n2896 & n7518 ) | ( n4415 & n7518 ) ;
  assign n50824 = n6243 & ~n50823 ;
  assign n50825 = n11614 & n50824 ;
  assign n50826 = ( n20997 & ~n50822 ) | ( n20997 & n50825 ) | ( ~n50822 & n50825 ) ;
  assign n50827 = n4625 & ~n20206 ;
  assign n50828 = n50827 ^ n4073 ^ 1'b0 ;
  assign n50829 = n50828 ^ n49558 ^ n24981 ;
  assign n50830 = n2228 & ~n3248 ;
  assign n50831 = n44885 ^ n26827 ^ 1'b0 ;
  assign n50832 = n36253 ^ n11963 ^ n1130 ;
  assign n50833 = n38893 ^ n20733 ^ 1'b0 ;
  assign n50834 = n20826 ^ n8322 ^ n5257 ;
  assign n50835 = n29940 ^ n29273 ^ n13041 ;
  assign n50836 = ( n16852 & n30628 ) | ( n16852 & n37937 ) | ( n30628 & n37937 ) ;
  assign n50837 = ~n4752 & n8303 ;
  assign n50838 = n50837 ^ n21430 ^ n2418 ;
  assign n50839 = n50838 ^ n14441 ^ 1'b0 ;
  assign n50840 = n50836 & ~n50839 ;
  assign n50841 = n50840 ^ n16606 ^ n7736 ;
  assign n50842 = ~n9440 & n32129 ;
  assign n50843 = n50842 ^ n27710 ^ 1'b0 ;
  assign n50846 = n47439 ^ n4597 ^ n377 ;
  assign n50847 = n50846 ^ n19640 ^ 1'b0 ;
  assign n50845 = ( ~n23266 & n25973 ) | ( ~n23266 & n45154 ) | ( n25973 & n45154 ) ;
  assign n50848 = n50847 ^ n50845 ^ n40062 ;
  assign n50844 = n821 & n27892 ;
  assign n50849 = n50848 ^ n50844 ^ 1'b0 ;
  assign n50851 = n23797 & ~n29204 ;
  assign n50850 = n22245 ^ n11006 ^ n8559 ;
  assign n50852 = n50851 ^ n50850 ^ n31904 ;
  assign n50853 = n48710 ^ n40635 ^ n22417 ;
  assign n50855 = n20427 ^ n3976 ^ n2809 ;
  assign n50854 = ( n4596 & n9770 ) | ( n4596 & ~n34418 ) | ( n9770 & ~n34418 ) ;
  assign n50856 = n50855 ^ n50854 ^ n44354 ;
  assign n50857 = n41134 ^ n35097 ^ n2168 ;
  assign n50858 = n49957 ^ n38872 ^ n9545 ;
  assign n50859 = n12680 ^ n2269 ^ n1888 ;
  assign n50860 = n50859 ^ n17633 ^ n12992 ;
  assign n50861 = ( n998 & n1856 ) | ( n998 & ~n23119 ) | ( n1856 & ~n23119 ) ;
  assign n50862 = n9969 ^ n9549 ^ n2305 ;
  assign n50863 = ( ~n11140 & n50684 ) | ( ~n11140 & n50862 ) | ( n50684 & n50862 ) ;
  assign n50867 = n15198 & ~n22429 ;
  assign n50865 = n21378 ^ n10572 ^ n757 ;
  assign n50866 = n7986 & n50865 ;
  assign n50868 = n50867 ^ n50866 ^ n35943 ;
  assign n50864 = ~n5243 & n16357 ;
  assign n50869 = n50868 ^ n50864 ^ 1'b0 ;
  assign n50870 = n19187 & n28384 ;
  assign n50871 = n16942 & n50870 ;
  assign n50875 = ( n5402 & n14985 ) | ( n5402 & ~n22729 ) | ( n14985 & ~n22729 ) ;
  assign n50872 = n37952 ^ n25666 ^ n12586 ;
  assign n50873 = n50872 ^ n24582 ^ n5040 ;
  assign n50874 = ~n33856 & n50873 ;
  assign n50876 = n50875 ^ n50874 ^ 1'b0 ;
  assign n50878 = ( n2114 & n5074 ) | ( n2114 & n15673 ) | ( n5074 & n15673 ) ;
  assign n50879 = n50878 ^ n26072 ^ n8907 ;
  assign n50877 = n19209 | n31048 ;
  assign n50880 = n50879 ^ n50877 ^ 1'b0 ;
  assign n50881 = n20094 & n50880 ;
  assign n50882 = n50881 ^ n11063 ^ n1793 ;
  assign n50883 = ( n3592 & n23230 ) | ( n3592 & n29107 ) | ( n23230 & n29107 ) ;
  assign n50884 = n24411 ^ n21545 ^ n5855 ;
  assign n50885 = ( n17861 & ~n50883 ) | ( n17861 & n50884 ) | ( ~n50883 & n50884 ) ;
  assign n50886 = ( n12004 & n19918 ) | ( n12004 & n35930 ) | ( n19918 & n35930 ) ;
  assign n50887 = n3493 | n22655 ;
  assign n50888 = ( n4961 & n16981 ) | ( n4961 & n50887 ) | ( n16981 & n50887 ) ;
  assign n50889 = ~n25713 & n50888 ;
  assign n50890 = ( n15178 & n28870 ) | ( n15178 & ~n50889 ) | ( n28870 & ~n50889 ) ;
  assign n50891 = n50890 ^ n42474 ^ n11478 ;
  assign n50892 = ( n16748 & ~n19215 ) | ( n16748 & n43723 ) | ( ~n19215 & n43723 ) ;
  assign n50893 = ( n11194 & ~n11247 ) | ( n11194 & n14682 ) | ( ~n11247 & n14682 ) ;
  assign n50894 = n11999 & ~n50893 ;
  assign n50895 = ~n15848 & n50894 ;
  assign n50896 = n50895 ^ n27913 ^ 1'b0 ;
  assign n50897 = n20303 | n50896 ;
  assign n50898 = n50892 & ~n50897 ;
  assign n50899 = ( n10428 & n16071 ) | ( n10428 & n49977 ) | ( n16071 & n49977 ) ;
  assign n50900 = ( n18256 & n20787 ) | ( n18256 & n50899 ) | ( n20787 & n50899 ) ;
  assign n50901 = n43641 ^ n16506 ^ n11287 ;
  assign n50902 = n31264 ^ n16451 ^ n4908 ;
  assign n50903 = n50902 ^ n24604 ^ n5352 ;
  assign n50904 = n41200 ^ n13703 ^ n9001 ;
  assign n50905 = n50904 ^ n16709 ^ n8553 ;
  assign n50906 = n27730 ^ n10114 ^ n5963 ;
  assign n50907 = ( n46106 & n50905 ) | ( n46106 & n50906 ) | ( n50905 & n50906 ) ;
  assign n50908 = n2404 & ~n50907 ;
  assign n50909 = n10578 | n26255 ;
  assign n50910 = n7963 & ~n50909 ;
  assign n50911 = n50910 ^ n22788 ^ n13191 ;
  assign n50912 = n48232 | n50911 ;
  assign n50913 = n27394 ^ n16708 ^ n11887 ;
  assign n50914 = ( n30835 & ~n37667 ) | ( n30835 & n50913 ) | ( ~n37667 & n50913 ) ;
  assign n50915 = n13741 | n50914 ;
  assign n50916 = x249 & n3735 ;
  assign n50917 = n50916 ^ n36144 ^ n809 ;
  assign n50918 = n15115 & n50917 ;
  assign n50919 = ( n13694 & ~n41849 ) | ( n13694 & n50918 ) | ( ~n41849 & n50918 ) ;
  assign n50920 = ( n15122 & n17518 ) | ( n15122 & ~n49993 ) | ( n17518 & ~n49993 ) ;
  assign n50921 = n32241 ^ n6492 ^ n1351 ;
  assign n50922 = n50921 ^ n14597 ^ n3235 ;
  assign n50924 = n2213 & ~n12815 ;
  assign n50923 = n47322 ^ n44566 ^ n28980 ;
  assign n50925 = n50924 ^ n50923 ^ n31452 ;
  assign n50926 = n47368 ^ n5400 ^ 1'b0 ;
  assign n50927 = ( ~n13296 & n35353 ) | ( ~n13296 & n50068 ) | ( n35353 & n50068 ) ;
  assign n50928 = ( n33409 & n50926 ) | ( n33409 & n50927 ) | ( n50926 & n50927 ) ;
  assign n50929 = n31143 ^ n23084 ^ n20807 ;
  assign n50931 = n6670 & ~n10712 ;
  assign n50930 = n8584 & ~n32543 ;
  assign n50932 = n50931 ^ n50930 ^ 1'b0 ;
  assign n50934 = n43062 ^ n15909 ^ n310 ;
  assign n50935 = n50934 ^ n17384 ^ 1'b0 ;
  assign n50933 = ~n2559 & n23857 ;
  assign n50936 = n50935 ^ n50933 ^ 1'b0 ;
  assign n50937 = n12555 & ~n24634 ;
  assign n50938 = ( ~n9062 & n16072 ) | ( ~n9062 & n25970 ) | ( n16072 & n25970 ) ;
  assign n50939 = ( n4430 & ~n6214 ) | ( n4430 & n50938 ) | ( ~n6214 & n50938 ) ;
  assign n50940 = ( n793 & ~n6143 ) | ( n793 & n50939 ) | ( ~n6143 & n50939 ) ;
  assign n50941 = ~n2331 & n9040 ;
  assign n50942 = n50941 ^ n31568 ^ 1'b0 ;
  assign n50943 = n50942 ^ n30845 ^ n16500 ;
  assign n50944 = n49810 ^ n34951 ^ n3308 ;
  assign n50945 = n34369 & ~n35058 ;
  assign n50946 = n33261 ^ n30095 ^ n12171 ;
  assign n50947 = n50946 ^ n41766 ^ n24798 ;
  assign n50948 = n27329 ^ n20474 ^ 1'b0 ;
  assign n50949 = n622 & n50948 ;
  assign n50950 = ( ~n19274 & n23351 ) | ( ~n19274 & n50949 ) | ( n23351 & n50949 ) ;
  assign n50951 = ( n24411 & n28189 ) | ( n24411 & n34802 ) | ( n28189 & n34802 ) ;
  assign n50952 = n10253 & n46733 ;
  assign n50953 = ~n45447 & n50952 ;
  assign n50954 = n21780 ^ n14344 ^ n12689 ;
  assign n50955 = ( n4068 & n8013 ) | ( n4068 & n42035 ) | ( n8013 & n42035 ) ;
  assign n50956 = n50955 ^ n11739 ^ n6117 ;
  assign n50957 = n16532 ^ n7685 ^ n792 ;
  assign n50958 = ( n26623 & n28536 ) | ( n26623 & ~n50957 ) | ( n28536 & ~n50957 ) ;
  assign n50959 = n50958 ^ n35868 ^ n34419 ;
  assign n50960 = ( ~n50954 & n50956 ) | ( ~n50954 & n50959 ) | ( n50956 & n50959 ) ;
  assign n50961 = ( n2520 & n7820 ) | ( n2520 & n15898 ) | ( n7820 & n15898 ) ;
  assign n50962 = n10645 ^ n869 ^ 1'b0 ;
  assign n50963 = n26025 ^ n12332 ^ n3916 ;
  assign n50964 = ( ~n23290 & n48816 ) | ( ~n23290 & n50963 ) | ( n48816 & n50963 ) ;
  assign n50965 = n49768 ^ n15463 ^ n14383 ;
  assign n50966 = n12467 ^ n1068 ^ 1'b0 ;
  assign n50967 = n3603 | n50966 ;
  assign n50968 = ( n4749 & n12328 ) | ( n4749 & n50967 ) | ( n12328 & n50967 ) ;
  assign n50969 = n50968 ^ n46874 ^ 1'b0 ;
  assign n50970 = ( ~n2222 & n18599 ) | ( ~n2222 & n50969 ) | ( n18599 & n50969 ) ;
  assign n50971 = n50970 ^ n10607 ^ n5117 ;
  assign n50972 = n50266 ^ n17992 ^ 1'b0 ;
  assign n50973 = n35299 ^ n27492 ^ n9360 ;
  assign n50974 = ~n8345 & n23951 ;
  assign n50975 = ~n50973 & n50974 ;
  assign n50976 = ( ~n27349 & n32468 ) | ( ~n27349 & n50975 ) | ( n32468 & n50975 ) ;
  assign n50977 = n16017 | n26713 ;
  assign n50978 = n20096 | n50977 ;
  assign n50979 = n42264 ^ n342 ^ 1'b0 ;
  assign n50980 = n35253 & ~n50979 ;
  assign n50981 = n25138 ^ n6492 ^ 1'b0 ;
  assign n50982 = n41856 ^ n4338 ^ 1'b0 ;
  assign n50983 = ( n1177 & ~n12652 ) | ( n1177 & n41859 ) | ( ~n12652 & n41859 ) ;
  assign n50984 = ( n1744 & n20715 ) | ( n1744 & n43769 ) | ( n20715 & n43769 ) ;
  assign n50985 = ( n6352 & ~n19426 ) | ( n6352 & n27243 ) | ( ~n19426 & n27243 ) ;
  assign n50986 = n45806 ^ n27739 ^ n2210 ;
  assign n50987 = ( n38183 & n50985 ) | ( n38183 & n50986 ) | ( n50985 & n50986 ) ;
  assign n50990 = n40430 ^ n10638 ^ 1'b0 ;
  assign n50988 = ~n1896 & n26843 ;
  assign n50989 = ~n11377 & n50988 ;
  assign n50991 = n50990 ^ n50989 ^ n34014 ;
  assign n50992 = n8548 & ~n45523 ;
  assign n50993 = n50992 ^ n21235 ^ 1'b0 ;
  assign n50994 = n28294 ^ n15670 ^ 1'b0 ;
  assign n50995 = ~n22143 & n50994 ;
  assign n50996 = n13939 & n45543 ;
  assign n50997 = n3671 | n13474 ;
  assign n50998 = n24687 & ~n50997 ;
  assign n50999 = n50998 ^ n46071 ^ n1990 ;
  assign n51000 = n13925 ^ n11181 ^ n8528 ;
  assign n51001 = n51000 ^ n18069 ^ n8935 ;
  assign n51002 = n51001 ^ n40406 ^ n30478 ;
  assign n51003 = ( ~n37402 & n41386 ) | ( ~n37402 & n51002 ) | ( n41386 & n51002 ) ;
  assign n51004 = n50018 ^ n7588 ^ n3659 ;
  assign n51005 = n8383 | n14466 ;
  assign n51006 = n51005 ^ n3993 ^ 1'b0 ;
  assign n51007 = ( n30405 & n51004 ) | ( n30405 & n51006 ) | ( n51004 & n51006 ) ;
  assign n51008 = n28113 ^ n18498 ^ n12921 ;
  assign n51009 = ( ~n5328 & n24491 ) | ( ~n5328 & n39613 ) | ( n24491 & n39613 ) ;
  assign n51010 = ( n31344 & ~n45734 ) | ( n31344 & n51009 ) | ( ~n45734 & n51009 ) ;
  assign n51012 = ~n14673 & n41464 ;
  assign n51013 = n51012 ^ n11779 ^ 1'b0 ;
  assign n51011 = n46795 ^ n1185 ^ 1'b0 ;
  assign n51014 = n51013 ^ n51011 ^ n6970 ;
  assign n51018 = n27300 & ~n36013 ;
  assign n51015 = n14543 & ~n14674 ;
  assign n51016 = n51015 ^ n5441 ^ 1'b0 ;
  assign n51017 = n46211 & ~n51016 ;
  assign n51019 = n51018 ^ n51017 ^ 1'b0 ;
  assign n51020 = n43064 ^ n10765 ^ 1'b0 ;
  assign n51021 = ~n23891 & n51020 ;
  assign n51022 = n12384 | n14354 ;
  assign n51023 = n51022 ^ n18735 ^ 1'b0 ;
  assign n51024 = ( n8112 & n21092 ) | ( n8112 & n51023 ) | ( n21092 & n51023 ) ;
  assign n51025 = n51024 ^ n43287 ^ n3530 ;
  assign n51026 = ( ~n26070 & n26882 ) | ( ~n26070 & n51025 ) | ( n26882 & n51025 ) ;
  assign n51027 = ( n14852 & ~n16257 ) | ( n14852 & n51026 ) | ( ~n16257 & n51026 ) ;
  assign n51028 = n48357 ^ n22335 ^ 1'b0 ;
  assign n51029 = ( n18551 & ~n36363 ) | ( n18551 & n51028 ) | ( ~n36363 & n51028 ) ;
  assign n51030 = n38267 ^ n27987 ^ n2583 ;
  assign n51031 = n26319 ^ n23361 ^ n21261 ;
  assign n51032 = n34550 ^ n22749 ^ n6881 ;
  assign n51033 = ( n37079 & n37174 ) | ( n37079 & n48760 ) | ( n37174 & n48760 ) ;
  assign n51034 = n23123 & ~n51033 ;
  assign n51035 = ( n6632 & ~n35866 ) | ( n6632 & n51034 ) | ( ~n35866 & n51034 ) ;
  assign n51038 = n40885 ^ n36541 ^ n21479 ;
  assign n51036 = ~n10656 & n32388 ;
  assign n51037 = n51036 ^ n7007 ^ 1'b0 ;
  assign n51039 = n51038 ^ n51037 ^ n1656 ;
  assign n51040 = ~n7651 & n17217 ;
  assign n51041 = n15768 | n48726 ;
  assign n51042 = n51041 ^ n14316 ^ 1'b0 ;
  assign n51043 = n51042 ^ n13776 ^ n9055 ;
  assign n51044 = n42654 ^ n38071 ^ n14376 ;
  assign n51045 = n51044 ^ n14563 ^ 1'b0 ;
  assign n51046 = n51043 & ~n51045 ;
  assign n51047 = n17727 ^ n17221 ^ 1'b0 ;
  assign n51048 = n27312 ^ n23299 ^ 1'b0 ;
  assign n51049 = n51047 | n51048 ;
  assign n51050 = n33603 ^ n26273 ^ 1'b0 ;
  assign n51051 = n50211 ^ n2384 ^ 1'b0 ;
  assign n51052 = ( ~n3929 & n11662 ) | ( ~n3929 & n13481 ) | ( n11662 & n13481 ) ;
  assign n51053 = ( n26803 & n37438 ) | ( n26803 & ~n51052 ) | ( n37438 & ~n51052 ) ;
  assign n51054 = n24888 ^ n2629 ^ 1'b0 ;
  assign n51055 = n15723 ^ n2966 ^ n1326 ;
  assign n51056 = n46711 ^ n22671 ^ 1'b0 ;
  assign n51057 = n26599 & n40221 ;
  assign n51058 = ~n9347 & n26643 ;
  assign n51059 = n51058 ^ n5580 ^ 1'b0 ;
  assign n51060 = n6226 & n42258 ;
  assign n51061 = n51060 ^ n1936 ^ 1'b0 ;
  assign n51062 = ( n22346 & n22761 ) | ( n22346 & n27641 ) | ( n22761 & n27641 ) ;
  assign n51063 = n51062 ^ n24207 ^ n16602 ;
  assign n51064 = ~n12376 & n36568 ;
  assign n51065 = n21684 ^ n18378 ^ 1'b0 ;
  assign n51066 = n9246 ^ n6470 ^ 1'b0 ;
  assign n51067 = n25940 | n51066 ;
  assign n51068 = n51067 ^ n47433 ^ n3181 ;
  assign n51069 = n5161 ^ x28 ^ 1'b0 ;
  assign n51070 = n51068 & ~n51069 ;
  assign n51071 = ( ~n19296 & n51065 ) | ( ~n19296 & n51070 ) | ( n51065 & n51070 ) ;
  assign n51072 = ( n1371 & ~n15941 ) | ( n1371 & n50686 ) | ( ~n15941 & n50686 ) ;
  assign n51074 = ( n2046 & n30394 ) | ( n2046 & n46435 ) | ( n30394 & n46435 ) ;
  assign n51073 = ~n2027 & n15869 ;
  assign n51075 = n51074 ^ n51073 ^ 1'b0 ;
  assign n51076 = n31006 ^ n22553 ^ n13381 ;
  assign n51077 = ( n35651 & n51075 ) | ( n35651 & ~n51076 ) | ( n51075 & ~n51076 ) ;
  assign n51078 = ~n2081 & n20576 ;
  assign n51079 = n51078 ^ n34589 ^ n7896 ;
  assign n51080 = ~n20473 & n22034 ;
  assign n51081 = n51080 ^ n31907 ^ 1'b0 ;
  assign n51082 = n18452 | n39632 ;
  assign n51083 = n9640 | n51082 ;
  assign n51084 = n39028 ^ n20484 ^ n14613 ;
  assign n51085 = ( n2566 & n42162 ) | ( n2566 & ~n43159 ) | ( n42162 & ~n43159 ) ;
  assign n51086 = n51085 ^ n42405 ^ 1'b0 ;
  assign n51087 = ~n38932 & n47531 ;
  assign n51088 = n4132 & ~n20449 ;
  assign n51089 = n26689 ^ n9857 ^ n9326 ;
  assign n51090 = n24712 ^ n15238 ^ 1'b0 ;
  assign n51091 = n26824 | n51090 ;
  assign n51092 = ( n27494 & ~n51089 ) | ( n27494 & n51091 ) | ( ~n51089 & n51091 ) ;
  assign n51093 = n16076 ^ n8386 ^ n1881 ;
  assign n51094 = n14457 ^ n7531 ^ 1'b0 ;
  assign n51095 = ( n39250 & n39636 ) | ( n39250 & n51094 ) | ( n39636 & n51094 ) ;
  assign n51097 = n25288 & n44015 ;
  assign n51098 = n51097 ^ n10022 ^ 1'b0 ;
  assign n51099 = n51098 ^ n20199 ^ n8611 ;
  assign n51096 = n44873 & ~n50679 ;
  assign n51100 = n51099 ^ n51096 ^ 1'b0 ;
  assign n51101 = n40131 ^ n8045 ^ 1'b0 ;
  assign n51102 = ~n8667 & n51101 ;
  assign n51103 = n8903 & ~n23623 ;
  assign n51104 = n51103 ^ n36734 ^ 1'b0 ;
  assign n51105 = n3412 | n37439 ;
  assign n51106 = n51105 ^ n31029 ^ 1'b0 ;
  assign n51107 = n51106 ^ n50382 ^ n28764 ;
  assign n51108 = n47001 ^ n17805 ^ n905 ;
  assign n51109 = n2394 & ~n3453 ;
  assign n51110 = n51109 ^ n5916 ^ 1'b0 ;
  assign n51111 = n38563 & n51110 ;
  assign n51112 = ( n5134 & n51108 ) | ( n5134 & n51111 ) | ( n51108 & n51111 ) ;
  assign n51113 = ( n6971 & n41335 ) | ( n6971 & ~n43759 ) | ( n41335 & ~n43759 ) ;
  assign n51114 = n51113 ^ n39527 ^ n29093 ;
  assign n51115 = n23821 ^ n2102 ^ 1'b0 ;
  assign n51116 = n11245 & ~n15675 ;
  assign n51117 = n51116 ^ n4802 ^ 1'b0 ;
  assign n51118 = n51117 ^ n19927 ^ n12648 ;
  assign n51119 = n26371 & n51118 ;
  assign n51120 = ~n29905 & n51119 ;
  assign n51121 = n51120 ^ n49982 ^ n13982 ;
  assign n51122 = n35126 ^ n18066 ^ n4357 ;
  assign n51123 = ( ~n10111 & n31881 ) | ( ~n10111 & n51122 ) | ( n31881 & n51122 ) ;
  assign n51124 = n47371 ^ n1482 ^ 1'b0 ;
  assign n51125 = ~n38237 & n51124 ;
  assign n51127 = n32832 ^ n5257 ^ 1'b0 ;
  assign n51128 = n11890 & ~n51127 ;
  assign n51129 = ~n27489 & n51128 ;
  assign n51130 = n51129 ^ n21980 ^ 1'b0 ;
  assign n51126 = n3329 | n48492 ;
  assign n51131 = n51130 ^ n51126 ^ 1'b0 ;
  assign n51132 = ~n6353 & n43803 ;
  assign n51133 = n51132 ^ n25093 ^ 1'b0 ;
  assign n51134 = ( ~n16836 & n50604 ) | ( ~n16836 & n51133 ) | ( n50604 & n51133 ) ;
  assign n51135 = ( ~n15230 & n38427 ) | ( ~n15230 & n47858 ) | ( n38427 & n47858 ) ;
  assign n51136 = ( n11680 & ~n15024 ) | ( n11680 & n33343 ) | ( ~n15024 & n33343 ) ;
  assign n51137 = ( n983 & ~n4062 ) | ( n983 & n50883 ) | ( ~n4062 & n50883 ) ;
  assign n51138 = n20668 ^ n12468 ^ n10430 ;
  assign n51139 = ( ~n874 & n28103 ) | ( ~n874 & n51138 ) | ( n28103 & n51138 ) ;
  assign n51140 = n51139 ^ n9263 ^ 1'b0 ;
  assign n51141 = ~n50806 & n51140 ;
  assign n51142 = n51141 ^ n33908 ^ n700 ;
  assign n51143 = n25429 ^ n22847 ^ n14092 ;
  assign n51144 = ( n8310 & ~n11991 ) | ( n8310 & n26029 ) | ( ~n11991 & n26029 ) ;
  assign n51145 = ( ~n31089 & n51143 ) | ( ~n31089 & n51144 ) | ( n51143 & n51144 ) ;
  assign n51146 = n51145 ^ n625 ^ 1'b0 ;
  assign n51147 = n34444 ^ n28014 ^ n25250 ;
  assign n51148 = n51147 ^ n29946 ^ n8442 ;
  assign n51149 = n21650 | n47961 ;
  assign n51150 = ( n6034 & n8183 ) | ( n6034 & n17849 ) | ( n8183 & n17849 ) ;
  assign n51151 = n51150 ^ n1825 ^ 1'b0 ;
  assign n51152 = n11709 & ~n51151 ;
  assign n51153 = n15864 & n17629 ;
  assign n51154 = n23234 ^ n14902 ^ n2558 ;
  assign n51155 = ( n1872 & n20814 ) | ( n1872 & n51154 ) | ( n20814 & n51154 ) ;
  assign n51156 = n18183 & ~n22943 ;
  assign n51157 = ~n51155 & n51156 ;
  assign n51158 = ( n6044 & ~n7259 ) | ( n6044 & n26724 ) | ( ~n7259 & n26724 ) ;
  assign n51159 = n51158 ^ n47053 ^ n19373 ;
  assign n51160 = n6215 | n51159 ;
  assign n51161 = ( n16348 & ~n51157 ) | ( n16348 & n51160 ) | ( ~n51157 & n51160 ) ;
  assign n51162 = ( n35666 & n51153 ) | ( n35666 & n51161 ) | ( n51153 & n51161 ) ;
  assign n51163 = n26402 ^ n10118 ^ n5024 ;
  assign n51164 = ( n15775 & ~n36103 ) | ( n15775 & n51163 ) | ( ~n36103 & n51163 ) ;
  assign n51165 = n44202 ^ n31524 ^ 1'b0 ;
  assign n51166 = n48819 ^ n18195 ^ n5900 ;
  assign n51167 = n21418 ^ n16096 ^ n15618 ;
  assign n51168 = n51167 ^ n25128 ^ n17337 ;
  assign n51169 = n44925 ^ n41930 ^ n4500 ;
  assign n51170 = ( n7059 & n14550 ) | ( n7059 & ~n51169 ) | ( n14550 & ~n51169 ) ;
  assign n51171 = ~n11044 & n31521 ;
  assign n51172 = n26477 & n51171 ;
  assign n51174 = ( ~n8719 & n34667 ) | ( ~n8719 & n47663 ) | ( n34667 & n47663 ) ;
  assign n51175 = n51174 ^ n36009 ^ n9850 ;
  assign n51173 = ( n689 & ~n10650 ) | ( n689 & n11101 ) | ( ~n10650 & n11101 ) ;
  assign n51176 = n51175 ^ n51173 ^ n41387 ;
  assign n51177 = n28229 ^ n14196 ^ n12786 ;
  assign n51178 = n23517 | n51177 ;
  assign n51179 = ( n1126 & ~n14847 ) | ( n1126 & n15256 ) | ( ~n14847 & n15256 ) ;
  assign n51180 = n51179 ^ n25840 ^ n5088 ;
  assign n51181 = n46013 ^ n29677 ^ n1365 ;
  assign n51182 = n6486 & n23870 ;
  assign n51183 = ( ~n47084 & n51181 ) | ( ~n47084 & n51182 ) | ( n51181 & n51182 ) ;
  assign n51184 = n34917 ^ n15564 ^ n10646 ;
  assign n51185 = ( n14357 & n50532 ) | ( n14357 & ~n51184 ) | ( n50532 & ~n51184 ) ;
  assign n51186 = ~n4190 & n14153 ;
  assign n51187 = n15430 & n51186 ;
  assign n51188 = n51187 ^ n46032 ^ n10949 ;
  assign n51189 = ( ~n14295 & n19945 ) | ( ~n14295 & n37967 ) | ( n19945 & n37967 ) ;
  assign n51190 = n36270 | n51189 ;
  assign n51191 = n6374 | n51190 ;
  assign n51192 = n43108 ^ n19876 ^ n17313 ;
  assign n51193 = n41621 ^ n16372 ^ 1'b0 ;
  assign n51194 = ~n31981 & n51193 ;
  assign n51195 = n51194 ^ n37308 ^ 1'b0 ;
  assign n51196 = n16902 ^ n13200 ^ n6737 ;
  assign n51197 = n46638 ^ n10366 ^ 1'b0 ;
  assign n51198 = n21603 ^ n16928 ^ n8364 ;
  assign n51199 = n14317 ^ n8724 ^ 1'b0 ;
  assign n51200 = n14490 & ~n51199 ;
  assign n51201 = n990 & n32930 ;
  assign n51202 = n11181 & n51201 ;
  assign n51203 = n51202 ^ n15953 ^ n6105 ;
  assign n51204 = n51203 ^ n45113 ^ n35151 ;
  assign n51205 = ( n4570 & n51200 ) | ( n4570 & n51204 ) | ( n51200 & n51204 ) ;
  assign n51206 = n44592 ^ n19008 ^ 1'b0 ;
  assign n51207 = n36908 & n51206 ;
  assign n51208 = x92 & ~n16275 ;
  assign n51209 = n51208 ^ n24643 ^ 1'b0 ;
  assign n51210 = n1837 | n8918 ;
  assign n51211 = n46033 | n51210 ;
  assign n51212 = n37017 ^ n14817 ^ n9339 ;
  assign n51213 = n33011 ^ n32812 ^ 1'b0 ;
  assign n51220 = ( n10330 & n36056 ) | ( n10330 & ~n50465 ) | ( n36056 & ~n50465 ) ;
  assign n51214 = n4982 & ~n11348 ;
  assign n51215 = ~n10840 & n51214 ;
  assign n51216 = ( n5529 & n22793 ) | ( n5529 & ~n51215 ) | ( n22793 & ~n51215 ) ;
  assign n51217 = ( n10435 & ~n23807 ) | ( n10435 & n51216 ) | ( ~n23807 & n51216 ) ;
  assign n51218 = n3443 & ~n51217 ;
  assign n51219 = n51218 ^ n974 ^ 1'b0 ;
  assign n51221 = n51220 ^ n51219 ^ 1'b0 ;
  assign n51222 = n35502 & n51221 ;
  assign n51223 = n23278 | n36669 ;
  assign n51224 = ( ~n8342 & n25273 ) | ( ~n8342 & n38766 ) | ( n25273 & n38766 ) ;
  assign n51227 = n7025 | n25153 ;
  assign n51228 = n51227 ^ n7415 ^ 1'b0 ;
  assign n51225 = n31964 ^ n5117 ^ 1'b0 ;
  assign n51226 = n51225 ^ n19330 ^ n9328 ;
  assign n51229 = n51228 ^ n51226 ^ n11607 ;
  assign n51230 = ~n905 & n35214 ;
  assign n51231 = n13175 ^ n3517 ^ 1'b0 ;
  assign n51232 = n18671 | n36226 ;
  assign n51233 = n48464 & ~n51232 ;
  assign n51236 = n33719 ^ n28039 ^ n2801 ;
  assign n51234 = ( x9 & ~n1391 ) | ( x9 & n9370 ) | ( ~n1391 & n9370 ) ;
  assign n51235 = ~n47448 & n51234 ;
  assign n51237 = n51236 ^ n51235 ^ 1'b0 ;
  assign n51238 = n33037 ^ n25730 ^ n21974 ;
  assign n51239 = ~n21110 & n26720 ;
  assign n51240 = n51238 & n51239 ;
  assign n51241 = ( n33134 & n34694 ) | ( n33134 & n51240 ) | ( n34694 & n51240 ) ;
  assign n51242 = n31732 ^ n25891 ^ 1'b0 ;
  assign n51243 = ( n29258 & n31150 ) | ( n29258 & ~n51242 ) | ( n31150 & ~n51242 ) ;
  assign n51244 = ( n18394 & n46608 ) | ( n18394 & n51243 ) | ( n46608 & n51243 ) ;
  assign n51245 = ( n620 & n2578 ) | ( n620 & ~n4218 ) | ( n2578 & ~n4218 ) ;
  assign n51246 = ( n12032 & ~n21446 ) | ( n12032 & n51245 ) | ( ~n21446 & n51245 ) ;
  assign n51247 = n51246 ^ n49415 ^ n48000 ;
  assign n51248 = n40051 ^ n36557 ^ n17158 ;
  assign n51249 = n51248 ^ n48169 ^ 1'b0 ;
  assign n51250 = n46610 ^ n31196 ^ n5564 ;
  assign n51251 = n4094 & n11098 ;
  assign n51252 = ~n14379 & n51251 ;
  assign n51253 = ( n583 & n4732 ) | ( n583 & ~n51252 ) | ( n4732 & ~n51252 ) ;
  assign n51254 = ( ~n5302 & n19355 ) | ( ~n5302 & n40134 ) | ( n19355 & n40134 ) ;
  assign n51255 = n18457 | n51254 ;
  assign n51256 = n51255 ^ n34018 ^ 1'b0 ;
  assign n51257 = ( n3574 & n34059 ) | ( n3574 & n51256 ) | ( n34059 & n51256 ) ;
  assign n51258 = ( ~n43711 & n51253 ) | ( ~n43711 & n51257 ) | ( n51253 & n51257 ) ;
  assign n51259 = n32363 ^ n14806 ^ n11181 ;
  assign n51260 = n24214 & n39173 ;
  assign n51261 = n47594 & n51260 ;
  assign n51262 = x136 & ~n20856 ;
  assign n51265 = n5839 & n10381 ;
  assign n51266 = n51265 ^ n10710 ^ 1'b0 ;
  assign n51264 = n10226 & n25189 ;
  assign n51263 = n25120 ^ n14493 ^ n6460 ;
  assign n51267 = n51266 ^ n51264 ^ n51263 ;
  assign n51268 = n51267 ^ n19753 ^ 1'b0 ;
  assign n51269 = ( n2168 & n5035 ) | ( n2168 & ~n9625 ) | ( n5035 & ~n9625 ) ;
  assign n51270 = ( n16813 & n27888 ) | ( n16813 & n35982 ) | ( n27888 & n35982 ) ;
  assign n51271 = ( n1996 & ~n48475 ) | ( n1996 & n51270 ) | ( ~n48475 & n51270 ) ;
  assign n51272 = ( n39550 & ~n51269 ) | ( n39550 & n51271 ) | ( ~n51269 & n51271 ) ;
  assign n51273 = ~n1410 & n13293 ;
  assign n51274 = ( n10804 & n12871 ) | ( n10804 & n51273 ) | ( n12871 & n51273 ) ;
  assign n51275 = n3532 & ~n14332 ;
  assign n51276 = ~n51274 & n51275 ;
  assign n51277 = ( n6179 & ~n50197 ) | ( n6179 & n51276 ) | ( ~n50197 & n51276 ) ;
  assign n51278 = ~n5324 & n36951 ;
  assign n51279 = n15278 & n51278 ;
  assign n51280 = n51279 ^ n13120 ^ n12581 ;
  assign n51281 = ( n19434 & n20089 ) | ( n19434 & n29146 ) | ( n20089 & n29146 ) ;
  assign n51282 = n51281 ^ n40246 ^ n5271 ;
  assign n51283 = n9527 ^ n1544 ^ 1'b0 ;
  assign n51284 = ~n14506 & n51283 ;
  assign n51285 = ( n29696 & ~n37847 ) | ( n29696 & n51284 ) | ( ~n37847 & n51284 ) ;
  assign n51286 = n3327 & n34863 ;
  assign n51287 = n51286 ^ n38386 ^ 1'b0 ;
  assign n51288 = n22309 & n51287 ;
  assign n51289 = ~n19648 & n31081 ;
  assign n51290 = n34771 & n51289 ;
  assign n51291 = n51290 ^ n15645 ^ 1'b0 ;
  assign n51292 = n38130 ^ n14088 ^ n9250 ;
  assign n51293 = ( n12975 & n26409 ) | ( n12975 & n51292 ) | ( n26409 & n51292 ) ;
  assign n51294 = n51293 ^ n37808 ^ n20893 ;
  assign n51295 = ( n12059 & ~n18134 ) | ( n12059 & n22363 ) | ( ~n18134 & n22363 ) ;
  assign n51296 = n51295 ^ n14141 ^ x104 ;
  assign n51297 = n51296 ^ n44343 ^ n12422 ;
  assign n51298 = n9337 ^ x208 ^ 1'b0 ;
  assign n51299 = ( ~n16261 & n29277 ) | ( ~n16261 & n51298 ) | ( n29277 & n51298 ) ;
  assign n51300 = n51299 ^ n35105 ^ n25940 ;
  assign n51301 = n24912 & ~n26881 ;
  assign n51302 = ( n4277 & n51300 ) | ( n4277 & ~n51301 ) | ( n51300 & ~n51301 ) ;
  assign n51303 = n30463 ^ n14534 ^ n2701 ;
  assign n51304 = n51303 ^ n27027 ^ n4576 ;
  assign n51305 = ( n9318 & ~n31112 ) | ( n9318 & n51304 ) | ( ~n31112 & n51304 ) ;
  assign n51306 = n19428 ^ n3512 ^ 1'b0 ;
  assign n51307 = n35232 | n51306 ;
  assign n51308 = ( n34260 & n41267 ) | ( n34260 & n51307 ) | ( n41267 & n51307 ) ;
  assign n51309 = n22218 ^ n22066 ^ 1'b0 ;
  assign n51310 = ( ~n2068 & n10710 ) | ( ~n2068 & n29105 ) | ( n10710 & n29105 ) ;
  assign n51311 = n51310 ^ n37102 ^ n6842 ;
  assign n51312 = ( ~n296 & n9414 ) | ( ~n296 & n19336 ) | ( n9414 & n19336 ) ;
  assign n51313 = n46407 ^ n31901 ^ n27059 ;
  assign n51314 = ( n25310 & n51312 ) | ( n25310 & ~n51313 ) | ( n51312 & ~n51313 ) ;
  assign n51315 = n51314 ^ n18832 ^ n10209 ;
  assign n51316 = n51315 ^ n30086 ^ 1'b0 ;
  assign n51317 = ( n23992 & ~n27985 ) | ( n23992 & n41684 ) | ( ~n27985 & n41684 ) ;
  assign n51318 = n16231 | n51317 ;
  assign n51319 = n8868 | n51318 ;
  assign n51320 = ~n34070 & n46767 ;
  assign n51321 = n51320 ^ n47110 ^ 1'b0 ;
  assign n51322 = n7664 ^ n7624 ^ n4063 ;
  assign n51323 = n51322 ^ n16735 ^ n3874 ;
  assign n51324 = ( ~n1652 & n27991 ) | ( ~n1652 & n41993 ) | ( n27991 & n41993 ) ;
  assign n51325 = n51324 ^ n27941 ^ n7180 ;
  assign n51326 = ( n12514 & n51323 ) | ( n12514 & n51325 ) | ( n51323 & n51325 ) ;
  assign n51327 = n21834 ^ n14888 ^ n12977 ;
  assign n51328 = n27854 ^ n17985 ^ n4513 ;
  assign n51329 = ( ~n6897 & n18539 ) | ( ~n6897 & n51328 ) | ( n18539 & n51328 ) ;
  assign n51330 = ( ~n6964 & n11977 ) | ( ~n6964 & n36613 ) | ( n11977 & n36613 ) ;
  assign n51331 = n51330 ^ n30975 ^ n22687 ;
  assign n51332 = n24675 ^ n1138 ^ 1'b0 ;
  assign n51333 = n39377 & ~n51332 ;
  assign n51334 = ( n7075 & n10145 ) | ( n7075 & n11767 ) | ( n10145 & n11767 ) ;
  assign n51335 = ( n33973 & n51333 ) | ( n33973 & n51334 ) | ( n51333 & n51334 ) ;
  assign n51336 = ( ~n20361 & n40976 ) | ( ~n20361 & n51335 ) | ( n40976 & n51335 ) ;
  assign n51337 = ( n10286 & ~n27223 ) | ( n10286 & n51336 ) | ( ~n27223 & n51336 ) ;
  assign n51338 = ( n25105 & n30299 ) | ( n25105 & ~n31056 ) | ( n30299 & ~n31056 ) ;
  assign n51339 = ( ~n19602 & n21217 ) | ( ~n19602 & n34493 ) | ( n21217 & n34493 ) ;
  assign n51340 = ( n385 & n11517 ) | ( n385 & ~n19975 ) | ( n11517 & ~n19975 ) ;
  assign n51341 = n51340 ^ n36569 ^ n10144 ;
  assign n51342 = n16031 ^ n9659 ^ n5715 ;
  assign n51343 = n51342 ^ n9363 ^ n5166 ;
  assign n51344 = n31136 & n51343 ;
  assign n51345 = ( ~n2903 & n23891 ) | ( ~n2903 & n51344 ) | ( n23891 & n51344 ) ;
  assign n51346 = ( ~n7287 & n10429 ) | ( ~n7287 & n12272 ) | ( n10429 & n12272 ) ;
  assign n51347 = n51345 | n51346 ;
  assign n51348 = n51347 ^ n31034 ^ 1'b0 ;
  assign n51349 = ( n27386 & ~n51341 ) | ( n27386 & n51348 ) | ( ~n51341 & n51348 ) ;
  assign n51350 = ( n15271 & n30115 ) | ( n15271 & n34577 ) | ( n30115 & n34577 ) ;
  assign n51351 = ( ~n3063 & n5757 ) | ( ~n3063 & n19552 ) | ( n5757 & n19552 ) ;
  assign n51352 = n30579 & n51351 ;
  assign n51353 = ~n51350 & n51352 ;
  assign n51354 = ( n5207 & n7605 ) | ( n5207 & n43058 ) | ( n7605 & n43058 ) ;
  assign n51355 = n46622 & n51354 ;
  assign n51356 = ( n1393 & n26920 ) | ( n1393 & n38152 ) | ( n26920 & n38152 ) ;
  assign n51357 = n42525 ^ n1205 ^ 1'b0 ;
  assign n51358 = n34397 | n51357 ;
  assign n51359 = ( n5291 & ~n51356 ) | ( n5291 & n51358 ) | ( ~n51356 & n51358 ) ;
  assign n51360 = n12266 & n22981 ;
  assign n51361 = ( ~n5864 & n6338 ) | ( ~n5864 & n33970 ) | ( n6338 & n33970 ) ;
  assign n51362 = n6380 ^ n2659 ^ x66 ;
  assign n51363 = ( n3060 & n12688 ) | ( n3060 & n51362 ) | ( n12688 & n51362 ) ;
  assign n51364 = ( ~n8867 & n51361 ) | ( ~n8867 & n51363 ) | ( n51361 & n51363 ) ;
  assign n51365 = n34275 ^ n33780 ^ n5679 ;
  assign n51366 = ~n25617 & n51365 ;
  assign n51368 = n10897 ^ n4570 ^ 1'b0 ;
  assign n51367 = n48677 ^ n39504 ^ 1'b0 ;
  assign n51369 = n51368 ^ n51367 ^ 1'b0 ;
  assign n51372 = n10401 ^ n3691 ^ n604 ;
  assign n51373 = n51372 ^ n12713 ^ n7493 ;
  assign n51374 = n51373 ^ n10716 ^ n5094 ;
  assign n51370 = ~n18913 & n36063 ;
  assign n51371 = ~n13363 & n51370 ;
  assign n51375 = n51374 ^ n51371 ^ n8215 ;
  assign n51376 = ~n1664 & n5897 ;
  assign n51377 = n51376 ^ n2879 ^ 1'b0 ;
  assign n51378 = n9209 ^ n8538 ^ n4748 ;
  assign n51379 = ~n6573 & n51378 ;
  assign n51380 = n2182 & n51379 ;
  assign n51381 = n9848 ^ n7797 ^ 1'b0 ;
  assign n51382 = n42901 ^ n39054 ^ n37798 ;
  assign n51383 = n3027 | n8970 ;
  assign n51384 = n33749 & ~n51383 ;
  assign n51385 = n23317 & ~n51384 ;
  assign n51386 = n47715 ^ n37362 ^ n24229 ;
  assign n51387 = n31000 ^ n22456 ^ n17040 ;
  assign n51388 = n9166 ^ n2774 ^ 1'b0 ;
  assign n51389 = n14749 | n51388 ;
  assign n51390 = ( ~n1543 & n8823 ) | ( ~n1543 & n51389 ) | ( n8823 & n51389 ) ;
  assign n51391 = ( n6435 & ~n29333 ) | ( n6435 & n39356 ) | ( ~n29333 & n39356 ) ;
  assign n51392 = ( n16522 & n51390 ) | ( n16522 & n51391 ) | ( n51390 & n51391 ) ;
  assign n51393 = n16566 ^ n15821 ^ 1'b0 ;
  assign n51394 = n4951 | n51393 ;
  assign n51395 = n51394 ^ n37515 ^ n10092 ;
  assign n51396 = n36635 ^ n25624 ^ n14392 ;
  assign n51397 = ( ~n14407 & n51395 ) | ( ~n14407 & n51396 ) | ( n51395 & n51396 ) ;
  assign n51398 = ( n17553 & n21425 ) | ( n17553 & n51397 ) | ( n21425 & n51397 ) ;
  assign n51399 = n35182 ^ n25999 ^ n6062 ;
  assign n51400 = ( ~n9575 & n26942 ) | ( ~n9575 & n51399 ) | ( n26942 & n51399 ) ;
  assign n51401 = ( n20275 & n51398 ) | ( n20275 & n51400 ) | ( n51398 & n51400 ) ;
  assign n51402 = ( n10879 & n21681 ) | ( n10879 & ~n51401 ) | ( n21681 & ~n51401 ) ;
  assign n51404 = ( ~n383 & n4009 ) | ( ~n383 & n19221 ) | ( n4009 & n19221 ) ;
  assign n51405 = n51404 ^ n27376 ^ n473 ;
  assign n51406 = ( n20290 & n38994 ) | ( n20290 & ~n51405 ) | ( n38994 & ~n51405 ) ;
  assign n51403 = n11524 ^ n4082 ^ n3014 ;
  assign n51407 = n51406 ^ n51403 ^ n13998 ;
  assign n51408 = n20684 ^ n4433 ^ 1'b0 ;
  assign n51409 = n5171 & n6119 ;
  assign n51410 = n1450 & n51409 ;
  assign n51411 = n28294 ^ n7062 ^ 1'b0 ;
  assign n51412 = ~n6351 & n51411 ;
  assign n51413 = n29282 ^ n25450 ^ n3305 ;
  assign n51414 = ( n20976 & ~n25320 ) | ( n20976 & n51413 ) | ( ~n25320 & n51413 ) ;
  assign n51415 = ( n4710 & n13231 ) | ( n4710 & ~n40753 ) | ( n13231 & ~n40753 ) ;
  assign n51416 = n24224 ^ n12169 ^ n861 ;
  assign n51417 = ( n13244 & ~n38243 ) | ( n13244 & n51416 ) | ( ~n38243 & n51416 ) ;
  assign n51418 = ( ~n7413 & n31070 ) | ( ~n7413 & n31941 ) | ( n31070 & n31941 ) ;
  assign n51419 = n51418 ^ n12921 ^ 1'b0 ;
  assign n51420 = ( n3936 & n4325 ) | ( n3936 & ~n51419 ) | ( n4325 & ~n51419 ) ;
  assign n51421 = ( n17237 & n27980 ) | ( n17237 & n49188 ) | ( n27980 & n49188 ) ;
  assign n51422 = n51421 ^ n32993 ^ n3783 ;
  assign n51423 = n11645 ^ n8148 ^ 1'b0 ;
  assign n51424 = n2408 & n51423 ;
  assign n51425 = ( n16593 & ~n51422 ) | ( n16593 & n51424 ) | ( ~n51422 & n51424 ) ;
  assign n51426 = n12296 ^ n9204 ^ 1'b0 ;
  assign n51427 = n28460 ^ n5506 ^ 1'b0 ;
  assign n51428 = ~n51426 & n51427 ;
  assign n51429 = n51428 ^ n37931 ^ n17916 ;
  assign n51430 = n46314 ^ n38481 ^ n11061 ;
  assign n51431 = ( n29702 & ~n43719 ) | ( n29702 & n51430 ) | ( ~n43719 & n51430 ) ;
  assign n51432 = ( n4739 & n7806 ) | ( n4739 & n41250 ) | ( n7806 & n41250 ) ;
  assign n51433 = n12133 ^ n9856 ^ 1'b0 ;
  assign n51434 = n33979 | n51433 ;
  assign n51435 = n28973 | n51434 ;
  assign n51436 = n7470 | n51435 ;
  assign n51437 = n11438 & ~n51436 ;
  assign n51438 = n1078 ^ n331 ^ 1'b0 ;
  assign n51439 = ( n8537 & n38527 ) | ( n8537 & ~n39560 ) | ( n38527 & ~n39560 ) ;
  assign n51440 = n11007 ^ n5596 ^ n4062 ;
  assign n51441 = ( n14437 & ~n23595 ) | ( n14437 & n51440 ) | ( ~n23595 & n51440 ) ;
  assign n51442 = n51441 ^ n28278 ^ n15387 ;
  assign n51443 = ( n26137 & n51439 ) | ( n26137 & n51442 ) | ( n51439 & n51442 ) ;
  assign n51444 = n1512 | n19039 ;
  assign n51445 = ( ~n2002 & n23129 ) | ( ~n2002 & n25639 ) | ( n23129 & n25639 ) ;
  assign n51446 = n5961 & ~n36823 ;
  assign n51447 = n51446 ^ n25327 ^ 1'b0 ;
  assign n51448 = ( n14159 & n51445 ) | ( n14159 & ~n51447 ) | ( n51445 & ~n51447 ) ;
  assign n51452 = ~n9647 & n32300 ;
  assign n51449 = n19577 & n23036 ;
  assign n51450 = n51449 ^ n38461 ^ 1'b0 ;
  assign n51451 = ( n4960 & n23367 ) | ( n4960 & n51450 ) | ( n23367 & n51450 ) ;
  assign n51453 = n51452 ^ n51451 ^ n31866 ;
  assign n51454 = n3837 | n19154 ;
  assign n51455 = n51454 ^ n6930 ^ 1'b0 ;
  assign n51456 = ( n12842 & n21257 ) | ( n12842 & ~n51455 ) | ( n21257 & ~n51455 ) ;
  assign n51457 = n51456 ^ n43121 ^ n22287 ;
  assign n51458 = n50828 ^ n10532 ^ n3286 ;
  assign n51459 = n51458 ^ n6345 ^ 1'b0 ;
  assign n51462 = n30696 ^ n7314 ^ n5236 ;
  assign n51460 = n8913 & n20849 ;
  assign n51461 = ~n13903 & n51460 ;
  assign n51463 = n51462 ^ n51461 ^ n18688 ;
  assign n51464 = n31724 ^ n13714 ^ n12880 ;
  assign n51465 = n597 & ~n10024 ;
  assign n51466 = ~n51464 & n51465 ;
  assign n51467 = ( n1629 & n26710 ) | ( n1629 & n27612 ) | ( n26710 & n27612 ) ;
  assign n51468 = n51467 ^ n28586 ^ n27229 ;
  assign n51469 = ( n26296 & n51466 ) | ( n26296 & n51468 ) | ( n51466 & n51468 ) ;
  assign n51470 = n36046 ^ n11591 ^ n7424 ;
  assign n51471 = ( ~n13090 & n24274 ) | ( ~n13090 & n51470 ) | ( n24274 & n51470 ) ;
  assign n51472 = n51471 ^ n12534 ^ n7198 ;
  assign n51473 = n41584 ^ n34822 ^ n5524 ;
  assign n51474 = ( n8945 & ~n13985 ) | ( n8945 & n49315 ) | ( ~n13985 & n49315 ) ;
  assign n51475 = ( n5536 & ~n38673 ) | ( n5536 & n51474 ) | ( ~n38673 & n51474 ) ;
  assign n51476 = n14041 & ~n24956 ;
  assign n51477 = ~n17623 & n22889 ;
  assign n51478 = n51477 ^ n2174 ^ 1'b0 ;
  assign n51479 = ( n21380 & n51476 ) | ( n21380 & ~n51478 ) | ( n51476 & ~n51478 ) ;
  assign n51480 = n21180 & ~n37813 ;
  assign n51481 = n6810 & n24664 ;
  assign n51482 = n51481 ^ n11219 ^ 1'b0 ;
  assign n51483 = n22300 ^ n10309 ^ n2364 ;
  assign n51484 = n51483 ^ n33627 ^ 1'b0 ;
  assign n51485 = n31238 ^ n30980 ^ n5795 ;
  assign n51486 = ( n7314 & n24817 ) | ( n7314 & ~n32545 ) | ( n24817 & ~n32545 ) ;
  assign n51487 = n2157 & ~n22811 ;
  assign n51488 = n37095 ^ n20984 ^ n12604 ;
  assign n51489 = n17947 & ~n26587 ;
  assign n51490 = n20784 & n51489 ;
  assign n51491 = n51490 ^ n5145 ^ 1'b0 ;
  assign n51492 = n24215 | n51491 ;
  assign n51493 = n19988 | n24103 ;
  assign n51494 = n51493 ^ n25880 ^ 1'b0 ;
  assign n51495 = n32570 | n51494 ;
  assign n51496 = ( ~n26945 & n51492 ) | ( ~n26945 & n51495 ) | ( n51492 & n51495 ) ;
  assign n51498 = n23310 ^ n16128 ^ n9533 ;
  assign n51499 = n51498 ^ n31413 ^ x67 ;
  assign n51497 = ( ~n17761 & n28320 ) | ( ~n17761 & n50748 ) | ( n28320 & n50748 ) ;
  assign n51500 = n51499 ^ n51497 ^ n23703 ;
  assign n51504 = ~n13634 & n20872 ;
  assign n51502 = n26236 ^ n2341 ^ 1'b0 ;
  assign n51503 = n905 & ~n51502 ;
  assign n51501 = ( ~n25556 & n38110 ) | ( ~n25556 & n40102 ) | ( n38110 & n40102 ) ;
  assign n51505 = n51504 ^ n51503 ^ n51501 ;
  assign n51506 = ~n2832 & n17862 ;
  assign n51507 = n33163 ^ n6344 ^ 1'b0 ;
  assign n51508 = n13676 | n15381 ;
  assign n51509 = n24200 | n51508 ;
  assign n51510 = n16354 & ~n51509 ;
  assign n51511 = n39943 ^ n11700 ^ n1104 ;
  assign n51512 = ~n3451 & n6258 ;
  assign n51513 = n13935 & n27157 ;
  assign n51514 = n51513 ^ n1370 ^ 1'b0 ;
  assign n51515 = ( n40902 & n51512 ) | ( n40902 & ~n51514 ) | ( n51512 & ~n51514 ) ;
  assign n51516 = n28930 ^ n26713 ^ n4040 ;
  assign n51517 = n29268 ^ n5536 ^ 1'b0 ;
  assign n51518 = n648 & ~n51517 ;
  assign n51519 = ( n11707 & ~n17729 ) | ( n11707 & n51518 ) | ( ~n17729 & n51518 ) ;
  assign n51521 = n27723 ^ n6333 ^ n699 ;
  assign n51522 = n51521 ^ n23841 ^ n20383 ;
  assign n51520 = n34331 | n35165 ;
  assign n51523 = n51522 ^ n51520 ^ n37369 ;
  assign n51524 = n21780 ^ n10539 ^ n8543 ;
  assign n51525 = ( x143 & ~n8431 ) | ( x143 & n40828 ) | ( ~n8431 & n40828 ) ;
  assign n51526 = ( ~n4573 & n14235 ) | ( ~n4573 & n27322 ) | ( n14235 & n27322 ) ;
  assign n51527 = ( n4394 & n10179 ) | ( n4394 & ~n44250 ) | ( n10179 & ~n44250 ) ;
  assign n51528 = ( ~n4547 & n51526 ) | ( ~n4547 & n51527 ) | ( n51526 & n51527 ) ;
  assign n51530 = ( n2440 & n9763 ) | ( n2440 & n38122 ) | ( n9763 & n38122 ) ;
  assign n51529 = n12050 & n23667 ;
  assign n51531 = n51530 ^ n51529 ^ 1'b0 ;
  assign n51532 = n21373 | n27504 ;
  assign n51533 = n6934 & ~n32668 ;
  assign n51534 = n51533 ^ n37060 ^ 1'b0 ;
  assign n51535 = n41115 & n51534 ;
  assign n51536 = ( ~n39851 & n49480 ) | ( ~n39851 & n51535 ) | ( n49480 & n51535 ) ;
  assign n51537 = n26212 ^ n11890 ^ 1'b0 ;
  assign n51538 = n5570 ^ n2076 ^ 1'b0 ;
  assign n51539 = ~n3512 & n22180 ;
  assign n51540 = ( n9750 & n36062 ) | ( n9750 & ~n41711 ) | ( n36062 & ~n41711 ) ;
  assign n51541 = ( n8740 & n11876 ) | ( n8740 & ~n20119 ) | ( n11876 & ~n20119 ) ;
  assign n51542 = ~n8671 & n49771 ;
  assign n51543 = n17516 & n51542 ;
  assign n51544 = n32749 ^ n23626 ^ 1'b0 ;
  assign n51545 = n10158 & ~n51544 ;
  assign n51549 = ( n1161 & ~n1665 ) | ( n1161 & n17028 ) | ( ~n1665 & n17028 ) ;
  assign n51546 = ~n7877 & n27150 ;
  assign n51547 = ~n26121 & n51546 ;
  assign n51548 = n10161 | n51547 ;
  assign n51550 = n51549 ^ n51548 ^ 1'b0 ;
  assign n51551 = ( n4556 & n25297 ) | ( n4556 & ~n29102 ) | ( n25297 & ~n29102 ) ;
  assign n51552 = n34247 & n51551 ;
  assign n51553 = n41404 ^ n7348 ^ 1'b0 ;
  assign n51554 = ( n1181 & ~n45226 ) | ( n1181 & n51553 ) | ( ~n45226 & n51553 ) ;
  assign n51555 = n51554 ^ n39608 ^ n38198 ;
  assign n51556 = n47122 ^ n23860 ^ n3060 ;
  assign n51557 = ( ~n8743 & n16416 ) | ( ~n8743 & n16892 ) | ( n16416 & n16892 ) ;
  assign n51558 = ( n604 & ~n5921 ) | ( n604 & n24723 ) | ( ~n5921 & n24723 ) ;
  assign n51559 = ( n12896 & ~n51557 ) | ( n12896 & n51558 ) | ( ~n51557 & n51558 ) ;
  assign n51560 = ( n3341 & n38794 ) | ( n3341 & n43072 ) | ( n38794 & n43072 ) ;
  assign n51561 = n15554 ^ n14555 ^ n607 ;
  assign n51562 = n5727 | n29273 ;
  assign n51563 = n14450 & ~n51562 ;
  assign n51564 = n51563 ^ n43192 ^ x162 ;
  assign n51565 = n43923 & n51564 ;
  assign n51568 = n44390 ^ n32943 ^ n20295 ;
  assign n51566 = n44968 ^ n34119 ^ n30947 ;
  assign n51567 = ~n30011 & n51566 ;
  assign n51569 = n51568 ^ n51567 ^ 1'b0 ;
  assign n51570 = n41100 ^ n8515 ^ 1'b0 ;
  assign n51571 = n30337 & ~n51570 ;
  assign n51572 = n9543 | n10395 ;
  assign n51573 = n51572 ^ n25341 ^ 1'b0 ;
  assign n51576 = n10492 ^ n10262 ^ n5942 ;
  assign n51577 = ( n13894 & ~n33907 ) | ( n13894 & n51576 ) | ( ~n33907 & n51576 ) ;
  assign n51574 = n7691 & ~n46726 ;
  assign n51575 = ~n1196 & n51574 ;
  assign n51578 = n51577 ^ n51575 ^ n17283 ;
  assign n51579 = ( n9931 & n16138 ) | ( n9931 & n42239 ) | ( n16138 & n42239 ) ;
  assign n51580 = n41412 ^ n35733 ^ n19594 ;
  assign n51581 = n37401 ^ n35300 ^ n30260 ;
  assign n51582 = n26284 ^ n15219 ^ 1'b0 ;
  assign n51583 = n51582 ^ n33194 ^ 1'b0 ;
  assign n51584 = n34467 | n36281 ;
  assign n51585 = n36620 ^ n2972 ^ 1'b0 ;
  assign n51586 = n4403 | n51585 ;
  assign n51587 = n51586 ^ n16429 ^ 1'b0 ;
  assign n51588 = n51587 ^ n47791 ^ n47716 ;
  assign n51589 = n13632 & n31334 ;
  assign n51590 = n51589 ^ n22277 ^ 1'b0 ;
  assign n51591 = n28260 & ~n40916 ;
  assign n51592 = n13412 ^ n11612 ^ n1090 ;
  assign n51593 = n37420 ^ n13651 ^ 1'b0 ;
  assign n51594 = n51593 ^ n20585 ^ n14325 ;
  assign n51595 = n1179 & n36169 ;
  assign n51596 = ~n14392 & n51595 ;
  assign n51597 = ( n16593 & ~n22671 ) | ( n16593 & n51596 ) | ( ~n22671 & n51596 ) ;
  assign n51598 = n40424 ^ n25702 ^ n14509 ;
  assign n51599 = ( n21614 & n51597 ) | ( n21614 & ~n51598 ) | ( n51597 & ~n51598 ) ;
  assign n51601 = n6756 | n7252 ;
  assign n51602 = n22171 & ~n51601 ;
  assign n51600 = n39707 ^ n22841 ^ 1'b0 ;
  assign n51603 = n51602 ^ n51600 ^ n17442 ;
  assign n51604 = ( n8586 & n16448 ) | ( n8586 & n36981 ) | ( n16448 & n36981 ) ;
  assign n51605 = n50879 ^ n33801 ^ n2476 ;
  assign n51606 = n51604 & ~n51605 ;
  assign n51607 = n6771 & ~n9390 ;
  assign n51608 = ( x73 & n1489 ) | ( x73 & ~n51607 ) | ( n1489 & ~n51607 ) ;
  assign n51609 = n51608 ^ n48107 ^ n42645 ;
  assign n51610 = ~n13985 & n17456 ;
  assign n51611 = n51610 ^ n28436 ^ 1'b0 ;
  assign n51612 = ( n22113 & n40036 ) | ( n22113 & n51611 ) | ( n40036 & n51611 ) ;
  assign n51613 = n48632 ^ n24109 ^ n18716 ;
  assign n51614 = n36614 ^ n3136 ^ 1'b0 ;
  assign n51615 = n5996 & n21916 ;
  assign n51616 = n51615 ^ n21192 ^ 1'b0 ;
  assign n51617 = n38339 & n51616 ;
  assign n51618 = n51617 ^ n4328 ^ 1'b0 ;
  assign n51619 = n17155 ^ n5326 ^ n4763 ;
  assign n51620 = ( ~n16131 & n40873 ) | ( ~n16131 & n51619 ) | ( n40873 & n51619 ) ;
  assign n51621 = ( n5044 & ~n27387 ) | ( n5044 & n34987 ) | ( ~n27387 & n34987 ) ;
  assign n51622 = ( n22658 & n29349 ) | ( n22658 & ~n48982 ) | ( n29349 & ~n48982 ) ;
  assign n51623 = n51622 ^ n38767 ^ n17824 ;
  assign n51624 = n22126 ^ n16751 ^ n12533 ;
  assign n51625 = n51624 ^ n13730 ^ n9075 ;
  assign n51626 = n36193 & n51625 ;
  assign n51627 = ~n23765 & n51626 ;
  assign n51628 = n20922 ^ n17165 ^ n5654 ;
  assign n51629 = n41403 ^ n9093 ^ n6534 ;
  assign n51630 = ( n19771 & n51628 ) | ( n19771 & n51629 ) | ( n51628 & n51629 ) ;
  assign n51631 = n21261 ^ n20380 ^ n16202 ;
  assign n51632 = n29400 ^ n4834 ^ 1'b0 ;
  assign n51633 = n26044 & ~n51632 ;
  assign n51634 = ( ~n1484 & n25625 ) | ( ~n1484 & n51633 ) | ( n25625 & n51633 ) ;
  assign n51635 = ( ~n16142 & n36228 ) | ( ~n16142 & n47295 ) | ( n36228 & n47295 ) ;
  assign n51636 = ( n6390 & n8439 ) | ( n6390 & n51635 ) | ( n8439 & n51635 ) ;
  assign n51637 = n12635 & n19852 ;
  assign n51638 = n51637 ^ n45474 ^ 1'b0 ;
  assign n51640 = ~n5959 & n16926 ;
  assign n51641 = ~n22267 & n51640 ;
  assign n51642 = ( ~n25814 & n37851 ) | ( ~n25814 & n51641 ) | ( n37851 & n51641 ) ;
  assign n51639 = n18125 | n33740 ;
  assign n51643 = n51642 ^ n51639 ^ 1'b0 ;
  assign n51644 = ( n14087 & n22892 ) | ( n14087 & ~n29937 ) | ( n22892 & ~n29937 ) ;
  assign n51645 = n18902 ^ n1108 ^ 1'b0 ;
  assign n51646 = n51644 & n51645 ;
  assign n51647 = ( n13072 & ~n15476 ) | ( n13072 & n23158 ) | ( ~n15476 & n23158 ) ;
  assign n51648 = n22395 ^ n1669 ^ 1'b0 ;
  assign n51649 = n5929 & ~n51648 ;
  assign n51650 = n51649 ^ n44638 ^ n12929 ;
  assign n51651 = n17364 ^ n12500 ^ n4379 ;
  assign n51652 = ( n1595 & n15847 ) | ( n1595 & ~n51651 ) | ( n15847 & ~n51651 ) ;
  assign n51653 = ( n6241 & ~n7179 ) | ( n6241 & n51652 ) | ( ~n7179 & n51652 ) ;
  assign n51655 = n26243 ^ n22121 ^ 1'b0 ;
  assign n51656 = n4541 | n51655 ;
  assign n51654 = ( ~n5657 & n17249 ) | ( ~n5657 & n24419 ) | ( n17249 & n24419 ) ;
  assign n51657 = n51656 ^ n51654 ^ n20318 ;
  assign n51658 = ( n3925 & n10428 ) | ( n3925 & n21180 ) | ( n10428 & n21180 ) ;
  assign n51659 = n51658 ^ n38898 ^ 1'b0 ;
  assign n51660 = ( n28096 & n37659 ) | ( n28096 & n51659 ) | ( n37659 & n51659 ) ;
  assign n51661 = ~n51657 & n51660 ;
  assign n51662 = n51661 ^ n31379 ^ 1'b0 ;
  assign n51663 = n51662 ^ n36190 ^ n5448 ;
  assign n51664 = n8516 & n18073 ;
  assign n51665 = n51664 ^ n13473 ^ 1'b0 ;
  assign n51666 = n801 & ~n41547 ;
  assign n51667 = n43819 ^ n1041 ^ 1'b0 ;
  assign n51668 = ( n32957 & n51666 ) | ( n32957 & n51667 ) | ( n51666 & n51667 ) ;
  assign n51669 = ( n27305 & n45374 ) | ( n27305 & n51668 ) | ( n45374 & n51668 ) ;
  assign n51670 = ( n38737 & n38874 ) | ( n38737 & n51669 ) | ( n38874 & n51669 ) ;
  assign n51671 = ( n4287 & n5767 ) | ( n4287 & n19757 ) | ( n5767 & n19757 ) ;
  assign n51672 = ~n47846 & n51671 ;
  assign n51673 = n12975 ^ n10770 ^ n6264 ;
  assign n51674 = ( ~n23982 & n36838 ) | ( ~n23982 & n51673 ) | ( n36838 & n51673 ) ;
  assign n51676 = n19476 ^ n15874 ^ n3141 ;
  assign n51675 = ~n29281 & n42361 ;
  assign n51677 = n51676 ^ n51675 ^ 1'b0 ;
  assign n51678 = ( n7100 & ~n48310 ) | ( n7100 & n49965 ) | ( ~n48310 & n49965 ) ;
  assign n51679 = ( n20684 & n28418 ) | ( n20684 & ~n32606 ) | ( n28418 & ~n32606 ) ;
  assign n51680 = ( n6139 & ~n26250 ) | ( n6139 & n41078 ) | ( ~n26250 & n41078 ) ;
  assign n51681 = n19330 & n36686 ;
  assign n51682 = n51681 ^ n6374 ^ 1'b0 ;
  assign n51683 = n48763 ^ n32425 ^ 1'b0 ;
  assign n51684 = n51683 ^ n19035 ^ n10341 ;
  assign n51685 = n48916 ^ n8941 ^ n6905 ;
  assign n51686 = ( n22376 & n35158 ) | ( n22376 & ~n44268 ) | ( n35158 & ~n44268 ) ;
  assign n51687 = ( ~n4820 & n8104 ) | ( ~n4820 & n28262 ) | ( n8104 & n28262 ) ;
  assign n51688 = ( ~n5411 & n5961 ) | ( ~n5411 & n43343 ) | ( n5961 & n43343 ) ;
  assign n51689 = ~n532 & n51688 ;
  assign n51690 = n41196 & n51689 ;
  assign n51691 = n8687 & n35379 ;
  assign n51692 = n4832 & ~n51691 ;
  assign n51693 = ~n1475 & n11494 ;
  assign n51694 = n51693 ^ n5472 ^ 1'b0 ;
  assign n51695 = ~n40983 & n48418 ;
  assign n51696 = ( ~n3746 & n23945 ) | ( ~n3746 & n51695 ) | ( n23945 & n51695 ) ;
  assign n51697 = n51696 ^ n5486 ^ 1'b0 ;
  assign n51698 = n14838 & ~n51158 ;
  assign n51699 = ~n6529 & n35244 ;
  assign n51700 = ( n7268 & n9218 ) | ( n7268 & ~n24030 ) | ( n9218 & ~n24030 ) ;
  assign n51701 = n51700 ^ n3874 ^ 1'b0 ;
  assign n51702 = n8848 | n51701 ;
  assign n51703 = ( n38195 & ~n45033 ) | ( n38195 & n51702 ) | ( ~n45033 & n51702 ) ;
  assign n51704 = n20144 | n50213 ;
  assign n51709 = ( n4287 & ~n15804 ) | ( n4287 & n22874 ) | ( ~n15804 & n22874 ) ;
  assign n51707 = ( n1659 & n5785 ) | ( n1659 & n11835 ) | ( n5785 & n11835 ) ;
  assign n51708 = n51707 ^ n19854 ^ n11035 ;
  assign n51705 = ( n2250 & n14775 ) | ( n2250 & ~n39153 ) | ( n14775 & ~n39153 ) ;
  assign n51706 = ( n12239 & ~n17407 ) | ( n12239 & n51705 ) | ( ~n17407 & n51705 ) ;
  assign n51710 = n51709 ^ n51708 ^ n51706 ;
  assign n51711 = n6704 & n32468 ;
  assign n51712 = n51711 ^ n21311 ^ 1'b0 ;
  assign n51713 = n51712 ^ n46223 ^ n29745 ;
  assign n51714 = n51713 ^ n1188 ^ 1'b0 ;
  assign n51715 = x158 & n36735 ;
  assign n51716 = n51715 ^ n20710 ^ 1'b0 ;
  assign n51717 = n45826 ^ n22175 ^ n4610 ;
  assign n51718 = n51717 ^ n3385 ^ 1'b0 ;
  assign n51719 = n49117 | n51718 ;
  assign n51720 = n17179 | n51719 ;
  assign n51721 = n51720 ^ n7676 ^ 1'b0 ;
  assign n51723 = n24057 ^ n23443 ^ n5387 ;
  assign n51722 = ( n5198 & ~n29769 ) | ( n5198 & n41151 ) | ( ~n29769 & n41151 ) ;
  assign n51724 = n51723 ^ n51722 ^ 1'b0 ;
  assign n51725 = n3616 & n51724 ;
  assign n51726 = n42262 ^ n30492 ^ 1'b0 ;
  assign n51727 = n11070 & ~n51726 ;
  assign n51728 = ( n1326 & n26186 ) | ( n1326 & ~n51727 ) | ( n26186 & ~n51727 ) ;
  assign n51729 = ( n7479 & n9294 ) | ( n7479 & n51728 ) | ( n9294 & n51728 ) ;
  assign n51730 = n45960 ^ n22795 ^ n803 ;
  assign n51731 = ( n39913 & n46498 ) | ( n39913 & ~n51730 ) | ( n46498 & ~n51730 ) ;
  assign n51732 = n17224 | n47172 ;
  assign n51733 = ( n7358 & n10107 ) | ( n7358 & ~n17954 ) | ( n10107 & ~n17954 ) ;
  assign n51734 = ( n8527 & n14345 ) | ( n8527 & ~n51733 ) | ( n14345 & ~n51733 ) ;
  assign n51735 = n8459 | n24610 ;
  assign n51736 = n51735 ^ n20865 ^ n2988 ;
  assign n51737 = n36192 ^ n14266 ^ n8065 ;
  assign n51738 = n35424 ^ n14368 ^ n3090 ;
  assign n51739 = n34643 & ~n51738 ;
  assign n51740 = n51739 ^ n6964 ^ 1'b0 ;
  assign n51741 = ~n7949 & n25474 ;
  assign n51742 = n24137 & n51741 ;
  assign n51743 = ( x79 & ~n2699 ) | ( x79 & n5577 ) | ( ~n2699 & n5577 ) ;
  assign n51744 = n51743 ^ n3767 ^ 1'b0 ;
  assign n51745 = ~n21921 & n22362 ;
  assign n51746 = n50342 ^ n21806 ^ n7062 ;
  assign n51747 = n47758 ^ n20429 ^ n8425 ;
  assign n51749 = ( ~n26485 & n27983 ) | ( ~n26485 & n42258 ) | ( n27983 & n42258 ) ;
  assign n51748 = ( n4188 & n30630 ) | ( n4188 & ~n31413 ) | ( n30630 & ~n31413 ) ;
  assign n51750 = n51749 ^ n51748 ^ n13955 ;
  assign n51751 = n3446 & n8369 ;
  assign n51752 = ( n21967 & n39426 ) | ( n21967 & n51751 ) | ( n39426 & n51751 ) ;
  assign n51753 = ( ~n2959 & n12409 ) | ( ~n2959 & n36104 ) | ( n12409 & n36104 ) ;
  assign n51754 = n44181 | n51753 ;
  assign n51755 = n10768 | n27013 ;
  assign n51756 = n34742 ^ n13717 ^ 1'b0 ;
  assign n51757 = n15366 & ~n51756 ;
  assign n51758 = ( n7633 & ~n12433 ) | ( n7633 & n15341 ) | ( ~n12433 & n15341 ) ;
  assign n51759 = ~n1626 & n51758 ;
  assign n51760 = n51759 ^ n5689 ^ 1'b0 ;
  assign n51761 = ~n44983 & n51760 ;
  assign n51762 = n51761 ^ n39604 ^ 1'b0 ;
  assign n51763 = n33772 ^ n24649 ^ n4557 ;
  assign n51764 = n5669 ^ n406 ^ 1'b0 ;
  assign n51765 = n7466 & ~n27330 ;
  assign n51766 = n51765 ^ n7617 ^ 1'b0 ;
  assign n51767 = n51766 ^ n34103 ^ x130 ;
  assign n51768 = n51767 ^ n32598 ^ n683 ;
  assign n51769 = n51666 ^ n19657 ^ n7074 ;
  assign n51770 = n34917 ^ n28228 ^ n18455 ;
  assign n51771 = n40313 ^ n36043 ^ 1'b0 ;
  assign n51772 = ( n13950 & n22324 ) | ( n13950 & ~n32417 ) | ( n22324 & ~n32417 ) ;
  assign n51773 = n42472 ^ n18749 ^ n580 ;
  assign n51774 = ( n25354 & ~n46586 ) | ( n25354 & n51773 ) | ( ~n46586 & n51773 ) ;
  assign n51775 = ( n30038 & ~n44428 ) | ( n30038 & n49407 ) | ( ~n44428 & n49407 ) ;
  assign n51776 = ( n34902 & n51774 ) | ( n34902 & ~n51775 ) | ( n51774 & ~n51775 ) ;
  assign n51777 = ~n779 & n21763 ;
  assign n51778 = ~n46983 & n51777 ;
  assign n51779 = n11367 & ~n15439 ;
  assign n51780 = n51779 ^ n43829 ^ 1'b0 ;
  assign n51781 = n46066 ^ n37197 ^ n5686 ;
  assign n51782 = n19227 | n33188 ;
  assign n51783 = n51781 & n51782 ;
  assign n51784 = ( ~n5783 & n8170 ) | ( ~n5783 & n17018 ) | ( n8170 & n17018 ) ;
  assign n51785 = n13858 ^ n9426 ^ 1'b0 ;
  assign n51786 = ~n26275 & n51785 ;
  assign n51787 = n51786 ^ n21890 ^ n5152 ;
  assign n51788 = n51787 ^ n13509 ^ 1'b0 ;
  assign n51789 = n51784 & n51788 ;
  assign n51790 = n51117 ^ n47359 ^ n43834 ;
  assign n51791 = ( n18230 & n51789 ) | ( n18230 & n51790 ) | ( n51789 & n51790 ) ;
  assign n51792 = n43575 ^ n32969 ^ n10901 ;
  assign n51793 = n22972 & ~n51792 ;
  assign n51794 = n51793 ^ n29661 ^ n12025 ;
  assign n51795 = n26930 ^ n8242 ^ n7430 ;
  assign n51796 = ( n2581 & n18141 ) | ( n2581 & ~n51795 ) | ( n18141 & ~n51795 ) ;
  assign n51797 = n41986 ^ n11588 ^ 1'b0 ;
  assign n51798 = n1876 | n51797 ;
  assign n51799 = n51798 ^ n28320 ^ n7829 ;
  assign n51800 = n28174 ^ n4729 ^ 1'b0 ;
  assign n51801 = n15222 & n51800 ;
  assign n51802 = ( n8426 & n10785 ) | ( n8426 & n16098 ) | ( n10785 & n16098 ) ;
  assign n51803 = n51248 ^ n21816 ^ n16280 ;
  assign n51804 = n7191 & n40947 ;
  assign n51805 = n51803 & n51804 ;
  assign n51806 = n35533 ^ n25772 ^ n15431 ;
  assign n51807 = ( n18498 & n32192 ) | ( n18498 & n41056 ) | ( n32192 & n41056 ) ;
  assign n51808 = ( n956 & ~n4481 ) | ( n956 & n8873 ) | ( ~n4481 & n8873 ) ;
  assign n51809 = ( n4530 & n39052 ) | ( n4530 & n40245 ) | ( n39052 & n40245 ) ;
  assign n51810 = n27657 ^ n26368 ^ n22327 ;
  assign n51811 = n51810 ^ n25578 ^ n16019 ;
  assign n51812 = ( n32980 & n51312 ) | ( n32980 & ~n51811 ) | ( n51312 & ~n51811 ) ;
  assign n51813 = n12253 ^ n1695 ^ 1'b0 ;
  assign n51814 = n9034 | n51813 ;
  assign n51815 = n51814 ^ n8316 ^ 1'b0 ;
  assign n51816 = ( ~n7522 & n46803 ) | ( ~n7522 & n51815 ) | ( n46803 & n51815 ) ;
  assign n51820 = n50587 ^ n27386 ^ n6354 ;
  assign n51817 = n17985 ^ n4728 ^ 1'b0 ;
  assign n51818 = n5527 & n51817 ;
  assign n51819 = ( n3114 & ~n50605 ) | ( n3114 & n51818 ) | ( ~n50605 & n51818 ) ;
  assign n51821 = n51820 ^ n51819 ^ n49313 ;
  assign n51822 = ( n332 & n2156 ) | ( n332 & ~n10720 ) | ( n2156 & ~n10720 ) ;
  assign n51823 = n51822 ^ n11573 ^ n5978 ;
  assign n51824 = ~n18903 & n24962 ;
  assign n51825 = n51824 ^ n22670 ^ 1'b0 ;
  assign n51826 = n5639 ^ n4586 ^ 1'b0 ;
  assign n51827 = n6432 & n51826 ;
  assign n51828 = ~n14704 & n19625 ;
  assign n51829 = ~n51827 & n51828 ;
  assign n51831 = n14589 | n33269 ;
  assign n51832 = n20718 | n51831 ;
  assign n51830 = n303 | n901 ;
  assign n51833 = n51832 ^ n51830 ^ n20120 ;
  assign n51834 = n48186 ^ n7612 ^ n3927 ;
  assign n51835 = n3060 | n21583 ;
  assign n51836 = n37536 ^ n35397 ^ 1'b0 ;
  assign n51837 = n51836 ^ n36677 ^ n8048 ;
  assign n51838 = ( ~n39582 & n51835 ) | ( ~n39582 & n51837 ) | ( n51835 & n51837 ) ;
  assign n51839 = n18496 ^ n3353 ^ 1'b0 ;
  assign n51840 = ~n17382 & n51839 ;
  assign n51841 = ( n16477 & ~n26715 ) | ( n16477 & n35332 ) | ( ~n26715 & n35332 ) ;
  assign n51842 = ( ~x224 & n11347 ) | ( ~x224 & n48797 ) | ( n11347 & n48797 ) ;
  assign n51843 = n371 & ~n25757 ;
  assign n51844 = n51843 ^ n25778 ^ 1'b0 ;
  assign n51845 = n9498 ^ n7135 ^ 1'b0 ;
  assign n51846 = n49293 & n51845 ;
  assign n51847 = n7750 & ~n33082 ;
  assign n51848 = n37185 & n51847 ;
  assign n51851 = n10705 & ~n13833 ;
  assign n51849 = n20396 ^ n8332 ^ n5906 ;
  assign n51850 = n24430 & n51849 ;
  assign n51852 = n51851 ^ n51850 ^ n18609 ;
  assign n51853 = n43802 ^ n19209 ^ n8732 ;
  assign n51854 = ( n18296 & n19008 ) | ( n18296 & n38502 ) | ( n19008 & n38502 ) ;
  assign n51855 = n7844 & ~n51854 ;
  assign n51856 = ~n46394 & n51855 ;
  assign n51857 = ( n1670 & ~n24929 ) | ( n1670 & n51856 ) | ( ~n24929 & n51856 ) ;
  assign n51858 = ( n1987 & n3096 ) | ( n1987 & n14775 ) | ( n3096 & n14775 ) ;
  assign n51859 = n51858 ^ n31301 ^ n2693 ;
  assign n51860 = n50686 ^ n48753 ^ 1'b0 ;
  assign n51861 = ( n18878 & ~n37851 ) | ( n18878 & n44325 ) | ( ~n37851 & n44325 ) ;
  assign n51862 = ( ~n27414 & n36528 ) | ( ~n27414 & n51861 ) | ( n36528 & n51861 ) ;
  assign n51863 = ( ~n8138 & n20360 ) | ( ~n8138 & n33464 ) | ( n20360 & n33464 ) ;
  assign n51864 = n51863 ^ n4321 ^ 1'b0 ;
  assign n51865 = n14749 ^ n8972 ^ n8055 ;
  assign n51866 = ( n14151 & n22691 ) | ( n14151 & n29455 ) | ( n22691 & n29455 ) ;
  assign n51867 = n27201 ^ n24710 ^ n18865 ;
  assign n51868 = n31168 ^ n7384 ^ 1'b0 ;
  assign n51869 = n16033 ^ n11989 ^ n6129 ;
  assign n51870 = ( n6132 & n33009 ) | ( n6132 & n51869 ) | ( n33009 & n51869 ) ;
  assign n51871 = ( x182 & n51868 ) | ( x182 & n51870 ) | ( n51868 & n51870 ) ;
  assign n51872 = ~n3500 & n8059 ;
  assign n51873 = n36280 ^ n32164 ^ n26842 ;
  assign n51874 = ( n14595 & n17881 ) | ( n14595 & n24167 ) | ( n17881 & n24167 ) ;
  assign n51875 = n51874 ^ n41975 ^ n22294 ;
  assign n51876 = n15564 ^ n14183 ^ n1863 ;
  assign n51877 = n51876 ^ n43569 ^ n22983 ;
  assign n51878 = ( n28382 & n40571 ) | ( n28382 & n51877 ) | ( n40571 & n51877 ) ;
  assign n51879 = n22951 ^ n15141 ^ 1'b0 ;
  assign n51880 = ~n16396 & n51879 ;
  assign n51881 = ~n966 & n28262 ;
  assign n51882 = n3811 & ~n51881 ;
  assign n51883 = ~n47129 & n51882 ;
  assign n51884 = n51883 ^ n41348 ^ 1'b0 ;
  assign n51885 = ~n6533 & n42822 ;
  assign n51886 = n51885 ^ n2959 ^ 1'b0 ;
  assign n51891 = n37523 ^ n5815 ^ n4877 ;
  assign n51889 = ( n3366 & ~n8386 ) | ( n3366 & n32253 ) | ( ~n8386 & n32253 ) ;
  assign n51887 = ( n10884 & n15697 ) | ( n10884 & ~n31888 ) | ( n15697 & ~n31888 ) ;
  assign n51888 = n51887 ^ n22969 ^ n13049 ;
  assign n51890 = n51889 ^ n51888 ^ n42418 ;
  assign n51892 = n51891 ^ n51890 ^ n3296 ;
  assign n51893 = n48617 ^ n46687 ^ n37134 ;
  assign n51894 = ( n4168 & n23637 ) | ( n4168 & ~n25615 ) | ( n23637 & ~n25615 ) ;
  assign n51895 = ( n8227 & n31473 ) | ( n8227 & ~n51894 ) | ( n31473 & ~n51894 ) ;
  assign n51896 = ( n5985 & n36043 ) | ( n5985 & n49944 ) | ( n36043 & n49944 ) ;
  assign n51897 = n40634 ^ n35120 ^ n9166 ;
  assign n51898 = ( ~n8038 & n28117 ) | ( ~n8038 & n45210 ) | ( n28117 & n45210 ) ;
  assign n51899 = n51898 ^ n44612 ^ n12661 ;
  assign n51900 = n10215 & ~n11243 ;
  assign n51901 = n51900 ^ n7262 ^ n1294 ;
  assign n51902 = n20689 ^ n859 ^ 1'b0 ;
  assign n51903 = n51902 ^ n27717 ^ n16440 ;
  assign n51904 = ( n14857 & n27638 ) | ( n14857 & ~n51903 ) | ( n27638 & ~n51903 ) ;
  assign n51905 = n51904 ^ n41483 ^ n36247 ;
  assign n51906 = ~n11511 & n12081 ;
  assign n51907 = n51906 ^ n13599 ^ 1'b0 ;
  assign n51908 = ~n13194 & n26340 ;
  assign n51909 = n41085 & n51908 ;
  assign n51910 = n22429 ^ n11787 ^ n1564 ;
  assign n51911 = n51910 ^ n34217 ^ n8851 ;
  assign n51912 = n47331 ^ n1629 ^ 1'b0 ;
  assign n51913 = ( n5135 & n51911 ) | ( n5135 & n51912 ) | ( n51911 & n51912 ) ;
  assign n51914 = ( n2919 & n21405 ) | ( n2919 & ~n40888 ) | ( n21405 & ~n40888 ) ;
  assign n51915 = n10551 ^ n1585 ^ 1'b0 ;
  assign n51916 = n51915 ^ n26278 ^ n7467 ;
  assign n51917 = ( n25358 & ~n51914 ) | ( n25358 & n51916 ) | ( ~n51914 & n51916 ) ;
  assign n51918 = n27800 & ~n28285 ;
  assign n51919 = n51918 ^ n3053 ^ 1'b0 ;
  assign n51920 = ( n9910 & n32112 ) | ( n9910 & n51919 ) | ( n32112 & n51919 ) ;
  assign n51921 = n27862 ^ n16208 ^ n3326 ;
  assign n51922 = ( ~n35721 & n38513 ) | ( ~n35721 & n51921 ) | ( n38513 & n51921 ) ;
  assign n51923 = ( ~n1713 & n7991 ) | ( ~n1713 & n43014 ) | ( n7991 & n43014 ) ;
  assign n51924 = n4403 & ~n51923 ;
  assign n51925 = n51924 ^ n33271 ^ 1'b0 ;
  assign n51926 = n51925 ^ n30499 ^ 1'b0 ;
  assign n51927 = n23166 | n41657 ;
  assign n51928 = n34129 | n51927 ;
  assign n51929 = n11737 | n51928 ;
  assign n51930 = n51929 ^ n44558 ^ n11619 ;
  assign n51931 = ( n923 & ~n30338 ) | ( n923 & n48993 ) | ( ~n30338 & n48993 ) ;
  assign n51932 = n31043 ^ n10671 ^ n9610 ;
  assign n51933 = n19256 & n51932 ;
  assign n51934 = ( n5398 & n26570 ) | ( n5398 & n27327 ) | ( n26570 & n27327 ) ;
  assign n51935 = n18803 ^ n9879 ^ n9448 ;
  assign n51936 = ( ~n18644 & n29493 ) | ( ~n18644 & n40477 ) | ( n29493 & n40477 ) ;
  assign n51937 = ( n5379 & n8823 ) | ( n5379 & n18223 ) | ( n8823 & n18223 ) ;
  assign n51938 = ( n8982 & n51936 ) | ( n8982 & n51937 ) | ( n51936 & n51937 ) ;
  assign n51939 = ( ~n11053 & n51935 ) | ( ~n11053 & n51938 ) | ( n51935 & n51938 ) ;
  assign n51940 = ~n44829 & n51939 ;
  assign n51941 = n51940 ^ n22623 ^ 1'b0 ;
  assign n51944 = n1143 & ~n17665 ;
  assign n51945 = n51944 ^ n19882 ^ 1'b0 ;
  assign n51942 = n9555 ^ n625 ^ 1'b0 ;
  assign n51943 = n48956 | n51942 ;
  assign n51946 = n51945 ^ n51943 ^ n746 ;
  assign n51947 = n51946 ^ n37292 ^ 1'b0 ;
  assign n51948 = ( n1405 & ~n16525 ) | ( n1405 & n42134 ) | ( ~n16525 & n42134 ) ;
  assign n51949 = n46112 ^ n6781 ^ 1'b0 ;
  assign n51950 = ( n10335 & n17218 ) | ( n10335 & ~n25379 ) | ( n17218 & ~n25379 ) ;
  assign n51951 = ( n26077 & n35968 ) | ( n26077 & n45223 ) | ( n35968 & n45223 ) ;
  assign n51952 = ( n32582 & n37810 ) | ( n32582 & ~n48431 ) | ( n37810 & ~n48431 ) ;
  assign n51953 = n30665 ^ n16859 ^ n16180 ;
  assign n51954 = ( n1038 & n2876 ) | ( n1038 & n11867 ) | ( n2876 & n11867 ) ;
  assign n51955 = ( n7658 & ~n38219 ) | ( n7658 & n51954 ) | ( ~n38219 & n51954 ) ;
  assign n51956 = n42134 ^ n37778 ^ n3687 ;
  assign n51957 = n34862 ^ n19666 ^ 1'b0 ;
  assign n51958 = n51957 ^ n24615 ^ n20793 ;
  assign n51959 = ( n10661 & n51956 ) | ( n10661 & n51958 ) | ( n51956 & n51958 ) ;
  assign n51960 = ( n51953 & n51955 ) | ( n51953 & ~n51959 ) | ( n51955 & ~n51959 ) ;
  assign n51961 = n9413 | n14555 ;
  assign n51962 = n51961 ^ n27354 ^ 1'b0 ;
  assign n51963 = ( n15613 & ~n20728 ) | ( n15613 & n47606 ) | ( ~n20728 & n47606 ) ;
  assign n51964 = n51963 ^ n43628 ^ n35597 ;
  assign n51965 = ( n4005 & n6461 ) | ( n4005 & ~n17007 ) | ( n6461 & ~n17007 ) ;
  assign n51966 = ( x133 & n35126 ) | ( x133 & ~n51965 ) | ( n35126 & ~n51965 ) ;
  assign n51967 = ( n37894 & n41054 ) | ( n37894 & n43176 ) | ( n41054 & n43176 ) ;
  assign n51968 = n29264 ^ n8240 ^ 1'b0 ;
  assign n51969 = n51968 ^ n37912 ^ n1134 ;
  assign n51970 = n51969 ^ n37007 ^ 1'b0 ;
  assign n51971 = n39918 | n51970 ;
  assign n51972 = n44541 | n51971 ;
  assign n51973 = n32349 & ~n35088 ;
  assign n51974 = n20226 & n51973 ;
  assign n51975 = n51974 ^ n9597 ^ n1976 ;
  assign n51976 = ( n11353 & ~n22063 ) | ( n11353 & n23335 ) | ( ~n22063 & n23335 ) ;
  assign n51977 = n7929 | n8067 ;
  assign n51978 = n51977 ^ n42113 ^ n4708 ;
  assign n51979 = ( n14974 & n24726 ) | ( n14974 & n31695 ) | ( n24726 & n31695 ) ;
  assign n51980 = ( n7483 & n28497 ) | ( n7483 & n51979 ) | ( n28497 & n51979 ) ;
  assign n51981 = ( ~n13325 & n36371 ) | ( ~n13325 & n51980 ) | ( n36371 & n51980 ) ;
  assign n51982 = n31957 ^ n15643 ^ 1'b0 ;
  assign n51983 = n48635 | n51982 ;
  assign n51984 = n32767 ^ n19657 ^ 1'b0 ;
  assign n51985 = n51984 ^ n14922 ^ 1'b0 ;
  assign n51986 = ~n51504 & n51985 ;
  assign n51987 = n51986 ^ n39793 ^ n27695 ;
  assign n51988 = n24843 ^ n8947 ^ n5539 ;
  assign n51989 = n51988 ^ n28403 ^ n20569 ;
  assign n51990 = ( n4550 & n14470 ) | ( n4550 & ~n51989 ) | ( n14470 & ~n51989 ) ;
  assign n51991 = n51990 ^ n41987 ^ n26442 ;
  assign n51992 = n32928 ^ n10690 ^ 1'b0 ;
  assign n51993 = ( ~n829 & n17182 ) | ( ~n829 & n37999 ) | ( n17182 & n37999 ) ;
  assign n51994 = n43970 & ~n51993 ;
  assign n51995 = ( ~n9358 & n27989 ) | ( ~n9358 & n28265 ) | ( n27989 & n28265 ) ;
  assign n51996 = n51995 ^ n24886 ^ n10401 ;
  assign n51998 = n23229 ^ n6915 ^ n5095 ;
  assign n51999 = n8856 ^ n3388 ^ 1'b0 ;
  assign n52000 = n51998 & ~n51999 ;
  assign n51997 = ( n3894 & n31884 ) | ( n3894 & ~n36133 ) | ( n31884 & ~n36133 ) ;
  assign n52001 = n52000 ^ n51997 ^ n21244 ;
  assign n52002 = n52001 ^ n44252 ^ n33071 ;
  assign n52003 = n34055 ^ n33743 ^ n21205 ;
  assign n52004 = n52003 ^ n32628 ^ n17308 ;
  assign n52005 = ( n4574 & ~n5842 ) | ( n4574 & n52004 ) | ( ~n5842 & n52004 ) ;
  assign n52006 = n52005 ^ n51877 ^ n23014 ;
  assign n52007 = ( n1972 & n9627 ) | ( n1972 & ~n27384 ) | ( n9627 & ~n27384 ) ;
  assign n52008 = n39384 ^ n4202 ^ 1'b0 ;
  assign n52009 = ~n13888 & n27425 ;
  assign n52010 = n35498 & n52009 ;
  assign n52015 = n16831 ^ n14664 ^ n4096 ;
  assign n52012 = ( x139 & n8330 ) | ( x139 & n8709 ) | ( n8330 & n8709 ) ;
  assign n52013 = n1613 | n24375 ;
  assign n52014 = n52012 | n52013 ;
  assign n52011 = ( n7030 & n34393 ) | ( n7030 & n37890 ) | ( n34393 & n37890 ) ;
  assign n52016 = n52015 ^ n52014 ^ n52011 ;
  assign n52017 = ( n16193 & n34302 ) | ( n16193 & n40325 ) | ( n34302 & n40325 ) ;
  assign n52018 = ( n2545 & n37672 ) | ( n2545 & ~n47973 ) | ( n37672 & ~n47973 ) ;
  assign n52019 = n3750 ^ n3686 ^ n2824 ;
  assign n52020 = n52019 ^ n11088 ^ 1'b0 ;
  assign n52021 = n42291 & n52020 ;
  assign n52022 = ( n5940 & n43160 ) | ( n5940 & n52021 ) | ( n43160 & n52021 ) ;
  assign n52023 = ( n6494 & n40596 ) | ( n6494 & ~n51365 ) | ( n40596 & ~n51365 ) ;
  assign n52024 = ( n6836 & ~n34243 ) | ( n6836 & n42168 ) | ( ~n34243 & n42168 ) ;
  assign n52025 = n52024 ^ n10363 ^ 1'b0 ;
  assign n52026 = n16805 ^ n14808 ^ 1'b0 ;
  assign n52027 = ~n19539 & n52026 ;
  assign n52028 = n13347 | n34259 ;
  assign n52029 = n52028 ^ n1561 ^ 1'b0 ;
  assign n52030 = ( n2171 & ~n49458 ) | ( n2171 & n52029 ) | ( ~n49458 & n52029 ) ;
  assign n52031 = ~n51840 & n52030 ;
  assign n52032 = n52031 ^ n44919 ^ 1'b0 ;
  assign n52033 = ( n9447 & n24016 ) | ( n9447 & n28384 ) | ( n24016 & n28384 ) ;
  assign n52034 = ( ~n6172 & n16574 ) | ( ~n6172 & n52033 ) | ( n16574 & n52033 ) ;
  assign n52035 = ( n14445 & n24621 ) | ( n14445 & ~n30421 ) | ( n24621 & ~n30421 ) ;
  assign n52036 = n30608 ^ n28517 ^ 1'b0 ;
  assign n52037 = n25569 ^ n11040 ^ n6061 ;
  assign n52038 = n23446 & n25614 ;
  assign n52039 = n10271 & n22485 ;
  assign n52040 = ~n52038 & n52039 ;
  assign n52041 = n52040 ^ n39168 ^ n3922 ;
  assign n52042 = ~n39144 & n43711 ;
  assign n52043 = n24125 ^ n8895 ^ 1'b0 ;
  assign n52044 = n15853 & n52043 ;
  assign n52045 = n13210 ^ n1324 ^ 1'b0 ;
  assign n52046 = n38544 | n52045 ;
  assign n52047 = n48492 ^ n28952 ^ 1'b0 ;
  assign n52048 = n11457 ^ n1564 ^ 1'b0 ;
  assign n52049 = n52048 ^ n48076 ^ n18780 ;
  assign n52050 = n38113 ^ n31107 ^ n4460 ;
  assign n52051 = ( n4957 & n27381 ) | ( n4957 & n52050 ) | ( n27381 & n52050 ) ;
  assign n52052 = n33372 ^ n27335 ^ n23859 ;
  assign n52053 = n47949 ^ n13173 ^ n4769 ;
  assign n52054 = n52053 ^ n46817 ^ n3231 ;
  assign n52055 = n43777 ^ n2938 ^ 1'b0 ;
  assign n52056 = ( n28873 & ~n42615 ) | ( n28873 & n50924 ) | ( ~n42615 & n50924 ) ;
  assign n52057 = n50025 ^ n15887 ^ n2260 ;
  assign n52058 = n10711 ^ n6576 ^ n1522 ;
  assign n52059 = n52058 ^ n44693 ^ n27215 ;
  assign n52060 = n52057 | n52059 ;
  assign n52061 = n52060 ^ n20386 ^ 1'b0 ;
  assign n52062 = ( ~n19131 & n26368 ) | ( ~n19131 & n41711 ) | ( n26368 & n41711 ) ;
  assign n52063 = n52062 ^ n40806 ^ n26844 ;
  assign n52064 = n52063 ^ n13579 ^ 1'b0 ;
  assign n52065 = ~n32075 & n52064 ;
  assign n52066 = ( ~n12927 & n32147 ) | ( ~n12927 & n35188 ) | ( n32147 & n35188 ) ;
  assign n52067 = n9034 ^ x67 ^ 1'b0 ;
  assign n52068 = ( n399 & n3788 ) | ( n399 & n14788 ) | ( n3788 & n14788 ) ;
  assign n52069 = ( n41547 & n43073 ) | ( n41547 & ~n52068 ) | ( n43073 & ~n52068 ) ;
  assign n52070 = n52069 ^ n38088 ^ n33652 ;
  assign n52071 = ~n3254 & n29383 ;
  assign n52072 = n12256 & n52071 ;
  assign n52073 = n21663 | n22730 ;
  assign n52074 = n52073 ^ n36204 ^ 1'b0 ;
  assign n52075 = n52074 ^ n44958 ^ n12951 ;
  assign n52076 = ( n1246 & ~n52072 ) | ( n1246 & n52075 ) | ( ~n52072 & n52075 ) ;
  assign n52077 = ( n5602 & n7880 ) | ( n5602 & n25445 ) | ( n7880 & n25445 ) ;
  assign n52078 = n45485 ^ n18230 ^ n11217 ;
  assign n52079 = ( n14113 & n23640 ) | ( n14113 & n52078 ) | ( n23640 & n52078 ) ;
  assign n52080 = n52079 ^ n41046 ^ n31167 ;
  assign n52081 = n5158 & n47154 ;
  assign n52082 = ( n33032 & n34270 ) | ( n33032 & ~n52081 ) | ( n34270 & ~n52081 ) ;
  assign n52083 = n40722 ^ n32325 ^ n19240 ;
  assign n52084 = n52083 ^ n21637 ^ 1'b0 ;
  assign n52085 = n49668 ^ n30720 ^ 1'b0 ;
  assign n52086 = n1211 | n52085 ;
  assign n52087 = n6745 | n10262 ;
  assign n52088 = ~n8887 & n18069 ;
  assign n52089 = n52087 & n52088 ;
  assign n52090 = n38195 ^ n24728 ^ n17790 ;
  assign n52091 = ( n2421 & ~n17792 ) | ( n2421 & n40787 ) | ( ~n17792 & n40787 ) ;
  assign n52092 = ( n42251 & n43020 ) | ( n42251 & n45084 ) | ( n43020 & n45084 ) ;
  assign n52093 = n30326 ^ n18299 ^ 1'b0 ;
  assign n52094 = n7238 & ~n49241 ;
  assign n52095 = n30050 & n52094 ;
  assign n52096 = n41023 ^ n24552 ^ n17159 ;
  assign n52097 = n52096 ^ n36142 ^ n5777 ;
  assign n52098 = n30002 ^ n27802 ^ n25711 ;
  assign n52099 = n52098 ^ n37709 ^ n7333 ;
  assign n52101 = n46827 ^ n37218 ^ n4951 ;
  assign n52100 = n44379 ^ n38520 ^ n3908 ;
  assign n52102 = n52101 ^ n52100 ^ n42235 ;
  assign n52103 = ( ~n4000 & n23210 ) | ( ~n4000 & n39692 ) | ( n23210 & n39692 ) ;
  assign n52104 = n17344 & ~n52103 ;
  assign n52105 = ( n12068 & n44971 ) | ( n12068 & ~n47144 ) | ( n44971 & ~n47144 ) ;
  assign n52106 = n35600 ^ n1364 ^ 1'b0 ;
  assign n52107 = ~n52105 & n52106 ;
  assign n52108 = n7397 & ~n42277 ;
  assign n52109 = n52108 ^ n23876 ^ 1'b0 ;
  assign n52110 = n16785 & n51723 ;
  assign n52111 = ( n25709 & n34566 ) | ( n25709 & n40732 ) | ( n34566 & n40732 ) ;
  assign n52112 = n3627 | n52111 ;
  assign n52113 = n39102 & ~n52112 ;
  assign n52114 = n52113 ^ n9937 ^ n821 ;
  assign n52115 = n35503 ^ n34848 ^ n8794 ;
  assign n52116 = ( n1846 & n20378 ) | ( n1846 & n25694 ) | ( n20378 & n25694 ) ;
  assign n52117 = n23267 & n52116 ;
  assign n52119 = n43231 ^ n5393 ^ 1'b0 ;
  assign n52120 = ( n6783 & n16354 ) | ( n6783 & ~n52119 ) | ( n16354 & ~n52119 ) ;
  assign n52118 = ( n7945 & n24704 ) | ( n7945 & ~n39164 ) | ( n24704 & ~n39164 ) ;
  assign n52121 = n52120 ^ n52118 ^ n5168 ;
  assign n52122 = ( n2632 & n22542 ) | ( n2632 & ~n29958 ) | ( n22542 & ~n29958 ) ;
  assign n52123 = n50244 & n52122 ;
  assign n52124 = ( n4650 & n12648 ) | ( n4650 & ~n25443 ) | ( n12648 & ~n25443 ) ;
  assign n52125 = ( ~n15803 & n34962 ) | ( ~n15803 & n43711 ) | ( n34962 & n43711 ) ;
  assign n52126 = n28571 ^ n8802 ^ 1'b0 ;
  assign n52127 = ~n7975 & n52126 ;
  assign n52128 = n6349 & ~n18940 ;
  assign n52129 = n47103 & n52128 ;
  assign n52130 = n47417 ^ n20610 ^ 1'b0 ;
  assign n52131 = ~n10858 & n52130 ;
  assign n52132 = n52131 ^ n50631 ^ n2922 ;
  assign n52134 = ( ~n1024 & n17295 ) | ( ~n1024 & n20688 ) | ( n17295 & n20688 ) ;
  assign n52133 = n48272 ^ n34630 ^ 1'b0 ;
  assign n52135 = n52134 ^ n52133 ^ n34425 ;
  assign n52136 = n39624 ^ n25637 ^ n6257 ;
  assign n52137 = ( n4310 & n10416 ) | ( n4310 & ~n16113 ) | ( n10416 & ~n16113 ) ;
  assign n52138 = n48391 ^ n19053 ^ n18012 ;
  assign n52139 = ( ~n51990 & n52137 ) | ( ~n51990 & n52138 ) | ( n52137 & n52138 ) ;
  assign n52140 = n52139 ^ n45059 ^ n9055 ;
  assign n52141 = ( n28981 & n33092 ) | ( n28981 & n52140 ) | ( n33092 & n52140 ) ;
  assign n52142 = ( ~n18041 & n28943 ) | ( ~n18041 & n40629 ) | ( n28943 & n40629 ) ;
  assign n52143 = ( n1944 & n21520 ) | ( n1944 & ~n29435 ) | ( n21520 & ~n29435 ) ;
  assign n52144 = ( ~n24329 & n50875 ) | ( ~n24329 & n52143 ) | ( n50875 & n52143 ) ;
  assign n52145 = n36632 ^ n22331 ^ n14644 ;
  assign n52146 = n4073 ^ n542 ^ 1'b0 ;
  assign n52147 = ( n1212 & ~n25462 ) | ( n1212 & n52146 ) | ( ~n25462 & n52146 ) ;
  assign n52148 = n20801 ^ n7817 ^ n3860 ;
  assign n52149 = ( n2856 & n13825 ) | ( n2856 & ~n52148 ) | ( n13825 & ~n52148 ) ;
  assign n52150 = n12857 & ~n30058 ;
  assign n52151 = ~n19863 & n52150 ;
  assign n52152 = ( n6023 & ~n14345 ) | ( n6023 & n52151 ) | ( ~n14345 & n52151 ) ;
  assign n52153 = ( n52147 & ~n52149 ) | ( n52147 & n52152 ) | ( ~n52149 & n52152 ) ;
  assign n52154 = n36410 ^ n7106 ^ 1'b0 ;
  assign n52155 = n41938 | n52154 ;
  assign n52157 = n1179 & n1652 ;
  assign n52158 = ( n10313 & ~n39530 ) | ( n10313 & n52157 ) | ( ~n39530 & n52157 ) ;
  assign n52156 = n25863 ^ n13317 ^ n644 ;
  assign n52159 = n52158 ^ n52156 ^ n15256 ;
  assign n52161 = ( x12 & n9462 ) | ( x12 & n16503 ) | ( n9462 & n16503 ) ;
  assign n52162 = n1696 & ~n5377 ;
  assign n52163 = ~n52161 & n52162 ;
  assign n52160 = n31705 ^ n9447 ^ 1'b0 ;
  assign n52164 = n52163 ^ n52160 ^ n44389 ;
  assign n52165 = n49004 ^ n25533 ^ n23717 ;
  assign n52166 = ( n1935 & ~n12508 ) | ( n1935 & n34892 ) | ( ~n12508 & n34892 ) ;
  assign n52167 = n52166 ^ n42665 ^ n37578 ;
  assign n52169 = n48096 ^ n39930 ^ n2829 ;
  assign n52168 = ( n4011 & n10683 ) | ( n4011 & ~n14470 ) | ( n10683 & ~n14470 ) ;
  assign n52170 = n52169 ^ n52168 ^ n50506 ;
  assign n52172 = n21014 & n25848 ;
  assign n52171 = ~n6882 & n18720 ;
  assign n52173 = n52172 ^ n52171 ^ 1'b0 ;
  assign n52174 = n52173 ^ n48731 ^ n31241 ;
  assign n52175 = n50661 ^ n45181 ^ n35549 ;
  assign n52176 = ~n13126 & n20227 ;
  assign n52180 = n48098 ^ n27591 ^ 1'b0 ;
  assign n52181 = n41954 ^ n27691 ^ 1'b0 ;
  assign n52182 = n2008 & n52181 ;
  assign n52183 = ( n26773 & n52180 ) | ( n26773 & ~n52182 ) | ( n52180 & ~n52182 ) ;
  assign n52177 = ( n1742 & ~n7696 ) | ( n1742 & n14651 ) | ( ~n7696 & n14651 ) ;
  assign n52178 = n41359 ^ n30873 ^ n25210 ;
  assign n52179 = ( ~n6222 & n52177 ) | ( ~n6222 & n52178 ) | ( n52177 & n52178 ) ;
  assign n52184 = n52183 ^ n52179 ^ n594 ;
  assign n52185 = ~n22935 & n28262 ;
  assign n52186 = n33088 & ~n52185 ;
  assign n52187 = n52186 ^ n7828 ^ 1'b0 ;
  assign n52188 = ( n16460 & n27345 ) | ( n16460 & ~n52187 ) | ( n27345 & ~n52187 ) ;
  assign n52189 = n44718 ^ n36593 ^ 1'b0 ;
  assign n52190 = n51052 ^ n39843 ^ n2262 ;
  assign n52191 = ( ~n17359 & n21719 ) | ( ~n17359 & n36958 ) | ( n21719 & n36958 ) ;
  assign n52193 = n15797 ^ n8505 ^ n892 ;
  assign n52194 = n52193 ^ n27015 ^ n10999 ;
  assign n52195 = n20610 | n34504 ;
  assign n52196 = n52194 | n52195 ;
  assign n52192 = n27350 ^ n22137 ^ n1622 ;
  assign n52197 = n52196 ^ n52192 ^ n10447 ;
  assign n52199 = n40808 ^ n14956 ^ n1963 ;
  assign n52198 = ( n9984 & n22459 ) | ( n9984 & n46289 ) | ( n22459 & n46289 ) ;
  assign n52200 = n52199 ^ n52198 ^ n3451 ;
  assign n52201 = n39193 ^ n3693 ^ 1'b0 ;
  assign n52202 = n5918 | n18280 ;
  assign n52203 = n52202 ^ n3521 ^ 1'b0 ;
  assign n52204 = n31584 & ~n52203 ;
  assign n52205 = n14577 ^ n12566 ^ 1'b0 ;
  assign n52206 = n41274 & ~n52205 ;
  assign n52207 = n37561 ^ n26226 ^ n6021 ;
  assign n52208 = n21909 & ~n52207 ;
  assign n52209 = ( n3377 & n17777 ) | ( n3377 & ~n44614 ) | ( n17777 & ~n44614 ) ;
  assign n52210 = ( n3547 & n29575 ) | ( n3547 & n52209 ) | ( n29575 & n52209 ) ;
  assign n52211 = n50496 ^ n18095 ^ 1'b0 ;
  assign n52212 = n46653 ^ n24439 ^ 1'b0 ;
  assign n52213 = n42403 ^ n24524 ^ n11069 ;
  assign n52214 = n19201 ^ n17841 ^ n6854 ;
  assign n52215 = ( n1429 & n52213 ) | ( n1429 & n52214 ) | ( n52213 & n52214 ) ;
  assign n52216 = ( n1002 & n23580 ) | ( n1002 & ~n24524 ) | ( n23580 & ~n24524 ) ;
  assign n52217 = ( n2176 & n52215 ) | ( n2176 & ~n52216 ) | ( n52215 & ~n52216 ) ;
  assign n52218 = n21798 ^ n10245 ^ n390 ;
  assign n52219 = ~n21081 & n27743 ;
  assign n52220 = n52219 ^ n41368 ^ n32218 ;
  assign n52221 = n52220 ^ n13694 ^ n6777 ;
  assign n52222 = n45672 & ~n51461 ;
  assign n52223 = n45829 & n52222 ;
  assign n52224 = ( n5175 & n6306 ) | ( n5175 & ~n12452 ) | ( n6306 & ~n12452 ) ;
  assign n52225 = n12743 ^ n6590 ^ n6261 ;
  assign n52226 = ( ~n22417 & n23643 ) | ( ~n22417 & n43845 ) | ( n23643 & n43845 ) ;
  assign n52227 = x246 & n52226 ;
  assign n52228 = ~n52225 & n52227 ;
  assign n52229 = ( n34207 & n43758 ) | ( n34207 & n52228 ) | ( n43758 & n52228 ) ;
  assign n52230 = n42868 ^ n5440 ^ 1'b0 ;
  assign n52231 = ~n30262 & n52230 ;
  assign n52232 = n52231 ^ n28591 ^ 1'b0 ;
  assign n52233 = n32190 ^ n26168 ^ n22126 ;
  assign n52234 = ~n25414 & n36242 ;
  assign n52235 = n29878 ^ n12352 ^ n8083 ;
  assign n52236 = ( n5466 & n5751 ) | ( n5466 & ~n8938 ) | ( n5751 & ~n8938 ) ;
  assign n52237 = n19396 & ~n33743 ;
  assign n52238 = n3640 | n12748 ;
  assign n52239 = n52238 ^ n5253 ^ 1'b0 ;
  assign n52240 = n9249 ^ n3960 ^ 1'b0 ;
  assign n52241 = ~n20547 & n52240 ;
  assign n52242 = n6044 | n22375 ;
  assign n52243 = n52242 ^ n29823 ^ 1'b0 ;
  assign n52244 = ( n11969 & n23655 ) | ( n11969 & n24110 ) | ( n23655 & n24110 ) ;
  assign n52245 = ( n4055 & ~n25559 ) | ( n4055 & n33069 ) | ( ~n25559 & n33069 ) ;
  assign n52246 = n15178 ^ n14062 ^ n9875 ;
  assign n52247 = ( ~n32674 & n43439 ) | ( ~n32674 & n52246 ) | ( n43439 & n52246 ) ;
  assign n52248 = ( x6 & n823 ) | ( x6 & ~n16149 ) | ( n823 & ~n16149 ) ;
  assign n52249 = n47742 ^ n27512 ^ n18046 ;
  assign n52250 = n52249 ^ n11689 ^ n7515 ;
  assign n52251 = ( ~n16912 & n17878 ) | ( ~n16912 & n52250 ) | ( n17878 & n52250 ) ;
  assign n52252 = n6257 | n21759 ;
  assign n52253 = ( n3536 & n15692 ) | ( n3536 & ~n33849 ) | ( n15692 & ~n33849 ) ;
  assign n52254 = n581 | n52253 ;
  assign n52255 = n36823 ^ n24952 ^ n12090 ;
  assign n52256 = n16889 & ~n20392 ;
  assign n52257 = ~n33075 & n52256 ;
  assign n52258 = n38781 ^ n5332 ^ 1'b0 ;
  assign n52259 = n829 & ~n52258 ;
  assign n52260 = n20558 | n37134 ;
  assign n52261 = ( n1669 & ~n2108 ) | ( n1669 & n2446 ) | ( ~n2108 & n2446 ) ;
  assign n52262 = ( ~n10664 & n32904 ) | ( ~n10664 & n34907 ) | ( n32904 & n34907 ) ;
  assign n52263 = n3521 | n41295 ;
  assign n52264 = n21318 & n32165 ;
  assign n52265 = n52263 & ~n52264 ;
  assign n52266 = n9684 ^ n9668 ^ 1'b0 ;
  assign n52267 = n40789 ^ n9012 ^ n1008 ;
  assign n52272 = n22655 ^ n17362 ^ n10545 ;
  assign n52269 = ( ~n7864 & n12281 ) | ( ~n7864 & n37659 ) | ( n12281 & n37659 ) ;
  assign n52270 = ( ~n24000 & n29307 ) | ( ~n24000 & n52269 ) | ( n29307 & n52269 ) ;
  assign n52271 = ( n16340 & ~n20767 ) | ( n16340 & n52270 ) | ( ~n20767 & n52270 ) ;
  assign n52268 = n27905 ^ n13896 ^ n10363 ;
  assign n52273 = n52272 ^ n52271 ^ n52268 ;
  assign n52274 = n23806 ^ n9036 ^ n1390 ;
  assign n52275 = n36909 ^ n19446 ^ n2602 ;
  assign n52276 = ( ~n4343 & n14162 ) | ( ~n4343 & n21573 ) | ( n14162 & n21573 ) ;
  assign n52277 = n52276 ^ n42053 ^ n25521 ;
  assign n52278 = n2646 & ~n20315 ;
  assign n52279 = ~n4016 & n52278 ;
  assign n52280 = n52279 ^ n49360 ^ n35145 ;
  assign n52282 = n15153 ^ n11236 ^ n5935 ;
  assign n52283 = n52282 ^ n20419 ^ 1'b0 ;
  assign n52281 = ( n17082 & n34017 ) | ( n17082 & ~n39198 ) | ( n34017 & ~n39198 ) ;
  assign n52284 = n52283 ^ n52281 ^ n939 ;
  assign n52288 = n3111 & ~n6421 ;
  assign n52287 = n21244 ^ n12792 ^ n6445 ;
  assign n52285 = n3580 | n28497 ;
  assign n52286 = n52285 ^ n50131 ^ 1'b0 ;
  assign n52289 = n52288 ^ n52287 ^ n52286 ;
  assign n52290 = ( n11362 & n34896 ) | ( n11362 & n52289 ) | ( n34896 & n52289 ) ;
  assign n52291 = n49687 ^ n30339 ^ n13428 ;
  assign n52292 = n34398 ^ n25961 ^ n4840 ;
  assign n52293 = n42690 ^ n24432 ^ 1'b0 ;
  assign n52294 = ~n37843 & n52293 ;
  assign n52295 = n8914 & ~n17899 ;
  assign n52296 = ~n9083 & n52295 ;
  assign n52297 = n2312 & n7851 ;
  assign n52298 = n52297 ^ n35342 ^ 1'b0 ;
  assign n52299 = ( n11767 & n22431 ) | ( n11767 & n35596 ) | ( n22431 & n35596 ) ;
  assign n52300 = n52299 ^ n44919 ^ n33598 ;
  assign n52301 = n15723 & ~n26300 ;
  assign n52302 = n30449 ^ n26527 ^ n12241 ;
  assign n52303 = ( n7260 & ~n25879 ) | ( n7260 & n44986 ) | ( ~n25879 & n44986 ) ;
  assign n52304 = n28358 ^ n17378 ^ 1'b0 ;
  assign n52305 = n23236 & ~n52304 ;
  assign n52306 = n52305 ^ n13775 ^ n4648 ;
  assign n52308 = n12701 ^ n11355 ^ n5341 ;
  assign n52309 = n52308 ^ n37489 ^ n8104 ;
  assign n52307 = n12146 & ~n28179 ;
  assign n52310 = n52309 ^ n52307 ^ 1'b0 ;
  assign n52311 = n52310 ^ n5425 ^ n448 ;
  assign n52312 = n44588 ^ n12673 ^ n5875 ;
  assign n52313 = n52312 ^ n18412 ^ n12833 ;
  assign n52314 = ( ~n7361 & n28762 ) | ( ~n7361 & n52313 ) | ( n28762 & n52313 ) ;
  assign n52315 = n3367 & n28870 ;
  assign n52316 = ~n24684 & n52315 ;
  assign n52317 = n9515 | n52316 ;
  assign n52318 = n37330 | n44135 ;
  assign n52319 = n52318 ^ n50244 ^ 1'b0 ;
  assign n52320 = n9367 | n33794 ;
  assign n52321 = n12560 & ~n52320 ;
  assign n52324 = ( x54 & n12680 ) | ( x54 & n46076 ) | ( n12680 & n46076 ) ;
  assign n52322 = n2834 | n23965 ;
  assign n52323 = n52322 ^ n21533 ^ 1'b0 ;
  assign n52325 = n52324 ^ n52323 ^ n22593 ;
  assign n52327 = ~n3947 & n3967 ;
  assign n52326 = n40240 ^ n23842 ^ n18245 ;
  assign n52328 = n52327 ^ n52326 ^ n49664 ;
  assign n52332 = n42967 ^ n15600 ^ n2454 ;
  assign n52330 = n43757 ^ n27789 ^ n13961 ;
  assign n52329 = n32398 ^ n16079 ^ n11391 ;
  assign n52331 = n52330 ^ n52329 ^ n43946 ;
  assign n52333 = n52332 ^ n52331 ^ n16238 ;
  assign n52334 = n18610 ^ n11155 ^ n6270 ;
  assign n52335 = ( n13293 & ~n27542 ) | ( n13293 & n52334 ) | ( ~n27542 & n52334 ) ;
  assign n52336 = ( n43814 & n50868 ) | ( n43814 & ~n52335 ) | ( n50868 & ~n52335 ) ;
  assign n52338 = n2574 ^ n1481 ^ n1478 ;
  assign n52337 = ( n11017 & n26065 ) | ( n11017 & n32878 ) | ( n26065 & n32878 ) ;
  assign n52339 = n52338 ^ n52337 ^ n43674 ;
  assign n52340 = n16670 ^ n9471 ^ n5278 ;
  assign n52341 = n52340 ^ n1067 ^ x150 ;
  assign n52342 = n52341 ^ n29204 ^ n342 ;
  assign n52343 = ( n26306 & n36908 ) | ( n26306 & ~n52342 ) | ( n36908 & ~n52342 ) ;
  assign n52344 = n5411 & n22298 ;
  assign n52345 = n4574 | n51699 ;
  assign n52346 = n52345 ^ n34476 ^ 1'b0 ;
  assign n52347 = n34182 & n34922 ;
  assign n52348 = n48854 & n52347 ;
  assign n52349 = n26073 ^ n22392 ^ 1'b0 ;
  assign n52350 = n4196 & ~n52349 ;
  assign n52351 = ( ~n7392 & n20650 ) | ( ~n7392 & n52350 ) | ( n20650 & n52350 ) ;
  assign n52352 = n37770 ^ n32809 ^ n31502 ;
  assign n52353 = n52352 ^ n13657 ^ n12408 ;
  assign n52354 = n41576 ^ n21898 ^ n6937 ;
  assign n52355 = n50959 ^ n25205 ^ 1'b0 ;
  assign n52358 = ( n9391 & ~n15913 ) | ( n9391 & n26112 ) | ( ~n15913 & n26112 ) ;
  assign n52356 = ~n7871 & n17998 ;
  assign n52357 = n25073 & n52356 ;
  assign n52359 = n52358 ^ n52357 ^ n30640 ;
  assign n52360 = ~n39438 & n41685 ;
  assign n52361 = ( n9521 & n10598 ) | ( n9521 & n14457 ) | ( n10598 & n14457 ) ;
  assign n52362 = ~n525 & n41063 ;
  assign n52363 = n8322 & n52362 ;
  assign n52364 = n6290 & n42731 ;
  assign n52365 = n19382 & n52364 ;
  assign n52366 = ( n2059 & ~n19278 ) | ( n2059 & n22384 ) | ( ~n19278 & n22384 ) ;
  assign n52367 = n37271 & n52366 ;
  assign n52368 = n14523 & n52367 ;
  assign n52369 = n7633 ^ n4836 ^ n2717 ;
  assign n52370 = ( ~n26099 & n49937 ) | ( ~n26099 & n52369 ) | ( n49937 & n52369 ) ;
  assign n52371 = n1212 & n2211 ;
  assign n52372 = n52371 ^ n26128 ^ 1'b0 ;
  assign n52373 = n52372 ^ n27207 ^ n16622 ;
  assign n52374 = ( n32948 & n33849 ) | ( n32948 & ~n52373 ) | ( n33849 & ~n52373 ) ;
  assign n52375 = n5916 ^ n2136 ^ n275 ;
  assign n52376 = ( n20526 & n26050 ) | ( n20526 & ~n52375 ) | ( n26050 & ~n52375 ) ;
  assign n52377 = n49482 ^ n18730 ^ 1'b0 ;
  assign n52378 = ( n27929 & n34686 ) | ( n27929 & n37717 ) | ( n34686 & n37717 ) ;
  assign n52379 = n37535 | n52378 ;
  assign n52380 = n17426 ^ n15296 ^ n12641 ;
  assign n52381 = n52380 ^ n12116 ^ 1'b0 ;
  assign n52382 = ~n33585 & n52381 ;
  assign n52383 = ( ~n6959 & n7635 ) | ( ~n6959 & n52382 ) | ( n7635 & n52382 ) ;
  assign n52384 = ( ~n636 & n12550 ) | ( ~n636 & n41711 ) | ( n12550 & n41711 ) ;
  assign n52386 = n39138 ^ n37137 ^ n17530 ;
  assign n52385 = ( n7583 & n17199 ) | ( n7583 & ~n38971 ) | ( n17199 & ~n38971 ) ;
  assign n52387 = n52386 ^ n52385 ^ n42737 ;
  assign n52388 = n17532 ^ n9437 ^ 1'b0 ;
  assign n52389 = ~n46410 & n52388 ;
  assign n52390 = n18060 ^ n17657 ^ n12089 ;
  assign n52391 = n52390 ^ n47940 ^ 1'b0 ;
  assign n52392 = n32948 & ~n52391 ;
  assign n52393 = ( ~n14338 & n32787 ) | ( ~n14338 & n33484 ) | ( n32787 & n33484 ) ;
  assign n52394 = n33242 ^ n21626 ^ n17040 ;
  assign n52395 = n50213 ^ n29094 ^ n23377 ;
  assign n52396 = n10651 & n16169 ;
  assign n52397 = n34737 & n52396 ;
  assign n52398 = ( n1890 & ~n45748 ) | ( n1890 & n52397 ) | ( ~n45748 & n52397 ) ;
  assign n52399 = n41848 ^ n6491 ^ x141 ;
  assign n52400 = ( n8628 & ~n11579 ) | ( n8628 & n37615 ) | ( ~n11579 & n37615 ) ;
  assign n52401 = ( ~n20576 & n48037 ) | ( ~n20576 & n52400 ) | ( n48037 & n52400 ) ;
  assign n52402 = ( n10643 & n19710 ) | ( n10643 & n52401 ) | ( n19710 & n52401 ) ;
  assign n52403 = n39895 ^ n8656 ^ 1'b0 ;
  assign n52404 = n24115 & ~n52403 ;
  assign n52405 = n3111 & n8019 ;
  assign n52406 = ~n19360 & n52405 ;
  assign n52407 = ( n829 & n48260 ) | ( n829 & n52406 ) | ( n48260 & n52406 ) ;
  assign n52408 = n48210 ^ n32518 ^ n19111 ;
  assign n52409 = n52408 ^ n1805 ^ 1'b0 ;
  assign n52410 = n8829 & ~n28385 ;
  assign n52411 = n42090 ^ n26386 ^ n25907 ;
  assign n52412 = ( n6636 & n19192 ) | ( n6636 & n23187 ) | ( n19192 & n23187 ) ;
  assign n52413 = ( n8303 & n8458 ) | ( n8303 & ~n33066 ) | ( n8458 & ~n33066 ) ;
  assign n52414 = n38439 ^ n21410 ^ n17372 ;
  assign n52415 = ( n10516 & n31411 ) | ( n10516 & ~n52414 ) | ( n31411 & ~n52414 ) ;
  assign n52416 = n24668 ^ n8268 ^ 1'b0 ;
  assign n52417 = n19477 ^ n10400 ^ 1'b0 ;
  assign n52418 = ~n52416 & n52417 ;
  assign n52419 = n33825 ^ n21431 ^ n20750 ;
  assign n52420 = ( n892 & n29693 ) | ( n892 & n52419 ) | ( n29693 & n52419 ) ;
  assign n52421 = n52420 ^ n51344 ^ 1'b0 ;
  assign n52422 = n8123 | n39975 ;
  assign n52423 = n52422 ^ n17684 ^ 1'b0 ;
  assign n52424 = ( n6669 & n24016 ) | ( n6669 & ~n32721 ) | ( n24016 & ~n32721 ) ;
  assign n52425 = n2670 & ~n24472 ;
  assign n52426 = ( n4806 & n47154 ) | ( n4806 & ~n52425 ) | ( n47154 & ~n52425 ) ;
  assign n52427 = n24215 ^ n17142 ^ 1'b0 ;
  assign n52428 = ( n1050 & ~n19906 ) | ( n1050 & n41073 ) | ( ~n19906 & n41073 ) ;
  assign n52429 = n52428 ^ n44515 ^ n1252 ;
  assign n52430 = n29083 ^ n18634 ^ 1'b0 ;
  assign n52431 = ( ~n14536 & n29299 ) | ( ~n14536 & n52094 ) | ( n29299 & n52094 ) ;
  assign n52432 = n36604 ^ n25229 ^ n15024 ;
  assign n52433 = n52432 ^ n43971 ^ n42162 ;
  assign n52434 = n49944 ^ n16122 ^ 1'b0 ;
  assign n52435 = n4630 & ~n36537 ;
  assign n52436 = ~n24396 & n52435 ;
  assign n52437 = ( n22740 & n41830 ) | ( n22740 & n46655 ) | ( n41830 & n46655 ) ;
  assign n52438 = n20849 ^ n8925 ^ 1'b0 ;
  assign n52439 = ~n8447 & n52438 ;
  assign n52440 = ( ~n19470 & n34511 ) | ( ~n19470 & n52439 ) | ( n34511 & n52439 ) ;
  assign n52441 = ( ~n9933 & n26053 ) | ( ~n9933 & n41171 ) | ( n26053 & n41171 ) ;
  assign n52442 = ( n13070 & n34156 ) | ( n13070 & n40621 ) | ( n34156 & n40621 ) ;
  assign n52443 = ( n1673 & n5429 ) | ( n1673 & ~n11654 ) | ( n5429 & ~n11654 ) ;
  assign n52444 = n52443 ^ n41258 ^ n26114 ;
  assign n52445 = n33401 & n41521 ;
  assign n52446 = ( n10040 & ~n15112 ) | ( n10040 & n52445 ) | ( ~n15112 & n52445 ) ;
  assign n52447 = n44632 ^ n30254 ^ n15303 ;
  assign n52448 = n3935 | n52447 ;
  assign n52449 = n52448 ^ n33196 ^ n19567 ;
  assign n52450 = n7110 | n13779 ;
  assign n52451 = n52450 ^ n1200 ^ 1'b0 ;
  assign n52452 = n31042 & ~n52451 ;
  assign n52453 = n52452 ^ n47849 ^ 1'b0 ;
  assign n52454 = n17820 & n52453 ;
  assign n52455 = ( n2604 & n20739 ) | ( n2604 & ~n38511 ) | ( n20739 & ~n38511 ) ;
  assign n52456 = ( n32156 & n41278 ) | ( n32156 & ~n49266 ) | ( n41278 & ~n49266 ) ;
  assign n52460 = ( n8061 & n18084 ) | ( n8061 & ~n22336 ) | ( n18084 & ~n22336 ) ;
  assign n52457 = ( n2586 & ~n4710 ) | ( n2586 & n27638 ) | ( ~n4710 & n27638 ) ;
  assign n52458 = n40576 ^ n7856 ^ 1'b0 ;
  assign n52459 = ~n52457 & n52458 ;
  assign n52461 = n52460 ^ n52459 ^ n4090 ;
  assign n52462 = n17988 & n26428 ;
  assign n52463 = n8919 & n52462 ;
  assign n52464 = n34567 ^ n30214 ^ n13615 ;
  assign n52465 = n31423 ^ n20774 ^ 1'b0 ;
  assign n52466 = ~n39215 & n52465 ;
  assign n52467 = ( ~n12471 & n42843 ) | ( ~n12471 & n52466 ) | ( n42843 & n52466 ) ;
  assign n52468 = n52467 ^ n13634 ^ n8617 ;
  assign n52469 = ( n10608 & n19800 ) | ( n10608 & n34801 ) | ( n19800 & n34801 ) ;
  assign n52471 = ( n469 & n3678 ) | ( n469 & ~n3699 ) | ( n3678 & ~n3699 ) ;
  assign n52472 = n52471 ^ n50018 ^ n12833 ;
  assign n52470 = n5625 & n8207 ;
  assign n52473 = n52472 ^ n52470 ^ 1'b0 ;
  assign n52474 = ~n2238 & n31656 ;
  assign n52475 = n52474 ^ n19034 ^ 1'b0 ;
  assign n52476 = n27131 ^ n5290 ^ 1'b0 ;
  assign n52477 = n19132 & ~n52476 ;
  assign n52478 = ( ~n17104 & n18784 ) | ( ~n17104 & n44955 ) | ( n18784 & n44955 ) ;
  assign n52479 = n29993 ^ n25954 ^ n20699 ;
  assign n52480 = n52479 ^ n9649 ^ n4778 ;
  assign n52486 = n7768 ^ n2637 ^ 1'b0 ;
  assign n52483 = n30424 ^ n11507 ^ 1'b0 ;
  assign n52484 = n52483 ^ n24517 ^ n514 ;
  assign n52482 = n14112 & n36934 ;
  assign n52485 = n52484 ^ n52482 ^ 1'b0 ;
  assign n52487 = n52486 ^ n52485 ^ n19596 ;
  assign n52481 = ( ~n11220 & n27681 ) | ( ~n11220 & n46000 ) | ( n27681 & n46000 ) ;
  assign n52488 = n52487 ^ n52481 ^ n22754 ;
  assign n52489 = n47233 ^ n31057 ^ n13554 ;
  assign n52490 = ( n928 & ~n6809 ) | ( n928 & n7025 ) | ( ~n6809 & n7025 ) ;
  assign n52491 = n38808 ^ n23071 ^ n18736 ;
  assign n52492 = ( n17663 & ~n52490 ) | ( n17663 & n52491 ) | ( ~n52490 & n52491 ) ;
  assign n52493 = ( n10722 & n20857 ) | ( n10722 & ~n52492 ) | ( n20857 & ~n52492 ) ;
  assign n52497 = n9658 ^ n6577 ^ n2727 ;
  assign n52495 = n16237 ^ n4198 ^ n2485 ;
  assign n52496 = n52495 ^ n37920 ^ 1'b0 ;
  assign n52494 = n15986 & ~n47624 ;
  assign n52498 = n52497 ^ n52496 ^ n52494 ;
  assign n52499 = ( n11989 & n43767 ) | ( n11989 & n52498 ) | ( n43767 & n52498 ) ;
  assign n52500 = ~n30859 & n41364 ;
  assign n52501 = n31455 & n36773 ;
  assign n52502 = n833 & n9473 ;
  assign n52503 = ~n3915 & n52502 ;
  assign n52504 = n48834 ^ n46951 ^ n3851 ;
  assign n52505 = n40261 ^ n28533 ^ n1264 ;
  assign n52506 = n44516 & ~n46519 ;
  assign n52507 = ( n13587 & n15351 ) | ( n13587 & n27648 ) | ( n15351 & n27648 ) ;
  assign n52508 = n42748 ^ n40881 ^ n1085 ;
  assign n52509 = n13935 ^ n4343 ^ 1'b0 ;
  assign n52510 = n30893 ^ n21557 ^ n17723 ;
  assign n52511 = n29606 | n49875 ;
  assign n52512 = x174 | n367 ;
  assign n52513 = ( n8982 & n21909 ) | ( n8982 & n51889 ) | ( n21909 & n51889 ) ;
  assign n52514 = ( n51491 & ~n52512 ) | ( n51491 & n52513 ) | ( ~n52512 & n52513 ) ;
  assign n52515 = n46489 ^ n28329 ^ n15029 ;
  assign n52516 = n11088 ^ n1745 ^ 1'b0 ;
  assign n52517 = ( n743 & n3517 ) | ( n743 & ~n52516 ) | ( n3517 & ~n52516 ) ;
  assign n52518 = n17438 & n52517 ;
  assign n52519 = n15521 ^ n3336 ^ 1'b0 ;
  assign n52520 = n50018 ^ n30455 ^ n1204 ;
  assign n52521 = n52520 ^ n32514 ^ 1'b0 ;
  assign n52522 = n35372 & n52521 ;
  assign n52523 = n52519 & n52522 ;
  assign n52524 = n16366 ^ n14359 ^ n7080 ;
  assign n52525 = n52283 ^ n28285 ^ 1'b0 ;
  assign n52526 = n29741 & n52525 ;
  assign n52527 = ( n18659 & ~n31517 ) | ( n18659 & n52526 ) | ( ~n31517 & n52526 ) ;
  assign n52528 = ( n4469 & n27988 ) | ( n4469 & n52527 ) | ( n27988 & n52527 ) ;
  assign n52529 = n44124 ^ n42798 ^ n7385 ;
  assign n52530 = n48916 ^ n10077 ^ n9905 ;
  assign n52531 = n33095 ^ n27145 ^ n22829 ;
  assign n52532 = n52531 ^ n1636 ^ 1'b0 ;
  assign n52533 = n23686 & n52532 ;
  assign n52534 = ~n22399 & n51220 ;
  assign n52535 = ~n13688 & n52534 ;
  assign n52536 = n36008 ^ n32123 ^ n30818 ;
  assign n52537 = n52536 ^ n15356 ^ n8297 ;
  assign n52538 = ~n13959 & n30350 ;
  assign n52539 = ~n3683 & n52538 ;
  assign n52540 = n52539 ^ n39901 ^ n8342 ;
  assign n52541 = n33541 ^ n6066 ^ 1'b0 ;
  assign n52547 = n49298 ^ n28039 ^ n7422 ;
  assign n52544 = ~n23287 & n38099 ;
  assign n52545 = n34018 & n52544 ;
  assign n52546 = n52545 ^ n47819 ^ n16479 ;
  assign n52542 = n6327 & n10720 ;
  assign n52543 = ~n21097 & n52542 ;
  assign n52548 = n52547 ^ n52546 ^ n52543 ;
  assign n52549 = ( n418 & n6910 ) | ( n418 & n27892 ) | ( n6910 & n27892 ) ;
  assign n52550 = ( n15619 & ~n18595 ) | ( n15619 & n37165 ) | ( ~n18595 & n37165 ) ;
  assign n52551 = n23998 ^ n1009 ^ 1'b0 ;
  assign n52552 = ( n45517 & n52550 ) | ( n45517 & ~n52551 ) | ( n52550 & ~n52551 ) ;
  assign n52553 = n9661 ^ n2682 ^ 1'b0 ;
  assign n52554 = n39926 ^ n31998 ^ n31109 ;
  assign n52555 = ( n31006 & n52553 ) | ( n31006 & n52554 ) | ( n52553 & n52554 ) ;
  assign n52556 = n23767 & ~n46348 ;
  assign n52557 = n52556 ^ n16138 ^ 1'b0 ;
  assign n52558 = n20761 ^ n10217 ^ 1'b0 ;
  assign n52559 = n27243 | n52558 ;
  assign n52560 = ( ~n5596 & n12791 ) | ( ~n5596 & n15287 ) | ( n12791 & n15287 ) ;
  assign n52561 = n52560 ^ n31150 ^ n13775 ;
  assign n52562 = n2081 | n52561 ;
  assign n52563 = n52562 ^ n4238 ^ 1'b0 ;
  assign n52564 = n25158 ^ n11020 ^ n1613 ;
  assign n52565 = ( ~n10678 & n11037 ) | ( ~n10678 & n11523 ) | ( n11037 & n11523 ) ;
  assign n52566 = ( n4896 & n6270 ) | ( n4896 & n52565 ) | ( n6270 & n52565 ) ;
  assign n52567 = ( n7084 & n8874 ) | ( n7084 & n47225 ) | ( n8874 & n47225 ) ;
  assign n52568 = n33724 & ~n45353 ;
  assign n52569 = n29724 ^ n18866 ^ n8100 ;
  assign n52570 = ( n16270 & ~n47495 ) | ( n16270 & n52569 ) | ( ~n47495 & n52569 ) ;
  assign n52571 = n52570 ^ n29953 ^ 1'b0 ;
  assign n52572 = ( n5132 & n41835 ) | ( n5132 & ~n52571 ) | ( n41835 & ~n52571 ) ;
  assign n52573 = n51345 ^ n49316 ^ 1'b0 ;
  assign n52574 = ( n6536 & n6656 ) | ( n6536 & ~n31143 ) | ( n6656 & ~n31143 ) ;
  assign n52575 = n52574 ^ n34252 ^ n12350 ;
  assign n52576 = n17672 ^ n2726 ^ n963 ;
  assign n52577 = n52576 ^ n22575 ^ n3930 ;
  assign n52578 = n37158 & n42861 ;
  assign n52579 = n52578 ^ n1039 ^ 1'b0 ;
  assign n52580 = n4679 | n22600 ;
  assign n52581 = n52580 ^ n24476 ^ 1'b0 ;
  assign n52582 = n31179 ^ n26009 ^ n16538 ;
  assign n52583 = n29036 ^ n4929 ^ 1'b0 ;
  assign n52584 = ( ~n40999 & n45841 ) | ( ~n40999 & n52583 ) | ( n45841 & n52583 ) ;
  assign n52585 = ~n29874 & n36593 ;
  assign n52586 = n15384 & n52585 ;
  assign n52587 = n7163 | n20354 ;
  assign n52588 = n52587 ^ n9351 ^ 1'b0 ;
  assign n52589 = n52588 ^ n47688 ^ n32211 ;
  assign n52590 = ( n12669 & n16272 ) | ( n12669 & ~n23403 ) | ( n16272 & ~n23403 ) ;
  assign n52591 = ( n23829 & n37845 ) | ( n23829 & ~n52590 ) | ( n37845 & ~n52590 ) ;
  assign n52592 = n19721 ^ n16222 ^ n7906 ;
  assign n52593 = ~n10036 & n52592 ;
  assign n52594 = n46034 ^ n38680 ^ n26886 ;
  assign n52595 = n51361 ^ n26197 ^ n21628 ;
  assign n52596 = ( ~n11277 & n19961 ) | ( ~n11277 & n35117 ) | ( n19961 & n35117 ) ;
  assign n52597 = n39800 | n52596 ;
  assign n52598 = n37545 | n49168 ;
  assign n52599 = ( n9017 & n25538 ) | ( n9017 & n36034 ) | ( n25538 & n36034 ) ;
  assign n52602 = n7353 ^ n4565 ^ n2342 ;
  assign n52600 = n34529 ^ n15231 ^ 1'b0 ;
  assign n52601 = ~n10391 & n52600 ;
  assign n52603 = n52602 ^ n52601 ^ n23126 ;
  assign n52604 = n45616 ^ n32712 ^ n3236 ;
  assign n52605 = n52604 ^ n38318 ^ x72 ;
  assign n52606 = ~n5467 & n23885 ;
  assign n52607 = n6258 & n52606 ;
  assign n52608 = n52607 ^ n33206 ^ n4612 ;
  assign n52609 = n4293 & ~n16120 ;
  assign n52610 = ~n41892 & n52609 ;
  assign n52611 = ( n12274 & ~n35088 ) | ( n12274 & n52610 ) | ( ~n35088 & n52610 ) ;
  assign n52612 = ( n16405 & ~n17401 ) | ( n16405 & n43394 ) | ( ~n17401 & n43394 ) ;
  assign n52613 = n52612 ^ n14867 ^ n9096 ;
  assign n52614 = ~n1500 & n5725 ;
  assign n52615 = n26925 ^ n21386 ^ n1761 ;
  assign n52616 = n23047 & n52615 ;
  assign n52617 = n9857 & ~n50434 ;
  assign n52618 = n30179 | n47457 ;
  assign n52619 = n52617 | n52618 ;
  assign n52620 = n4432 & ~n22773 ;
  assign n52621 = ( ~n28021 & n31790 ) | ( ~n28021 & n49407 ) | ( n31790 & n49407 ) ;
  assign n52622 = n24390 & ~n52621 ;
  assign n52623 = ~n52620 & n52622 ;
  assign n52624 = ( n3366 & n27608 ) | ( n3366 & ~n43704 ) | ( n27608 & ~n43704 ) ;
  assign n52625 = ( ~n11487 & n22955 ) | ( ~n11487 & n52624 ) | ( n22955 & n52624 ) ;
  assign n52626 = ( n17227 & n40462 ) | ( n17227 & ~n49929 ) | ( n40462 & ~n49929 ) ;
  assign n52627 = ( ~n12014 & n47464 ) | ( ~n12014 & n52626 ) | ( n47464 & n52626 ) ;
  assign n52628 = n17675 ^ n5349 ^ 1'b0 ;
  assign n52629 = n52628 ^ n42759 ^ n15057 ;
  assign n52630 = n52629 ^ n12168 ^ n4513 ;
  assign n52631 = ( n8792 & ~n36178 ) | ( n8792 & n42150 ) | ( ~n36178 & n42150 ) ;
  assign n52632 = n1212 & ~n13996 ;
  assign n52633 = n52632 ^ n13092 ^ 1'b0 ;
  assign n52634 = n52633 ^ n18742 ^ n1928 ;
  assign n52635 = n34890 ^ n9620 ^ n4896 ;
  assign n52636 = n30667 ^ n5021 ^ 1'b0 ;
  assign n52637 = ~n2983 & n52636 ;
  assign n52638 = ( ~n26899 & n52635 ) | ( ~n26899 & n52637 ) | ( n52635 & n52637 ) ;
  assign n52639 = n19608 & ~n33483 ;
  assign n52640 = n52639 ^ n37537 ^ 1'b0 ;
  assign n52641 = n52640 ^ n28703 ^ 1'b0 ;
  assign n52642 = n24839 ^ n20270 ^ 1'b0 ;
  assign n52643 = n22457 & ~n52642 ;
  assign n52644 = n3877 & n52643 ;
  assign n52645 = n52644 ^ n37174 ^ 1'b0 ;
  assign n52646 = n17450 ^ n5814 ^ 1'b0 ;
  assign n52647 = n33231 & ~n52646 ;
  assign n52648 = ~n19914 & n28751 ;
  assign n52649 = ( n4623 & n15468 ) | ( n4623 & ~n30984 ) | ( n15468 & ~n30984 ) ;
  assign n52650 = ( n11438 & n46638 ) | ( n11438 & ~n52649 ) | ( n46638 & ~n52649 ) ;
  assign n52651 = n47101 ^ n30093 ^ 1'b0 ;
  assign n52652 = n52651 ^ n35736 ^ n2914 ;
  assign n52653 = n4978 & n33794 ;
  assign n52654 = n31126 ^ n18718 ^ 1'b0 ;
  assign n52655 = n48299 ^ n21972 ^ 1'b0 ;
  assign n52656 = n30599 ^ n9199 ^ 1'b0 ;
  assign n52657 = n52655 & ~n52656 ;
  assign n52659 = n36425 ^ n20296 ^ n5071 ;
  assign n52658 = ( n28669 & ~n34877 ) | ( n28669 & n36655 ) | ( ~n34877 & n36655 ) ;
  assign n52660 = n52659 ^ n52658 ^ n35896 ;
  assign n52661 = n35114 ^ n16263 ^ n15902 ;
  assign n52662 = n24055 ^ n5509 ^ 1'b0 ;
  assign n52663 = n36499 & ~n52662 ;
  assign n52667 = n31386 & n51549 ;
  assign n52668 = n52667 ^ n21843 ^ 1'b0 ;
  assign n52664 = n20343 ^ n9214 ^ 1'b0 ;
  assign n52665 = n13974 & ~n52664 ;
  assign n52666 = ( ~n33962 & n50596 ) | ( ~n33962 & n52665 ) | ( n50596 & n52665 ) ;
  assign n52669 = n52668 ^ n52666 ^ n1204 ;
  assign n52670 = ( n9877 & ~n18961 ) | ( n9877 & n22280 ) | ( ~n18961 & n22280 ) ;
  assign n52671 = ( ~n37031 & n37578 ) | ( ~n37031 & n39975 ) | ( n37578 & n39975 ) ;
  assign n52672 = ( n38528 & ~n52670 ) | ( n38528 & n52671 ) | ( ~n52670 & n52671 ) ;
  assign n52673 = n50506 ^ n32464 ^ n15080 ;
  assign n52674 = n17931 | n26739 ;
  assign n52675 = n9413 & ~n52674 ;
  assign n52676 = ( n13117 & n41748 ) | ( n13117 & ~n52675 ) | ( n41748 & ~n52675 ) ;
  assign n52677 = ( n7536 & n39504 ) | ( n7536 & n52676 ) | ( n39504 & n52676 ) ;
  assign n52678 = ( n3978 & ~n6930 ) | ( n3978 & n24794 ) | ( ~n6930 & n24794 ) ;
  assign n52679 = n52678 ^ n8637 ^ n5229 ;
  assign n52680 = n35702 ^ n10610 ^ 1'b0 ;
  assign n52681 = n10332 & n52680 ;
  assign n52682 = ( n26683 & ~n52679 ) | ( n26683 & n52681 ) | ( ~n52679 & n52681 ) ;
  assign n52683 = ( n2629 & n22586 ) | ( n2629 & n47672 ) | ( n22586 & n47672 ) ;
  assign n52684 = n33723 ^ n26617 ^ n14748 ;
  assign n52685 = n52684 ^ n44181 ^ n8901 ;
  assign n52686 = n5064 ^ n2490 ^ 1'b0 ;
  assign n52687 = n52686 ^ n7781 ^ n5219 ;
  assign n52688 = n1255 & ~n12127 ;
  assign n52689 = n9831 & n52688 ;
  assign n52690 = ~n17473 & n23221 ;
  assign n52691 = n49928 & n52690 ;
  assign n52692 = n48677 ^ n39472 ^ n2485 ;
  assign n52693 = ~n6820 & n52692 ;
  assign n52694 = n31363 ^ n20006 ^ n7058 ;
  assign n52695 = n22766 & ~n29192 ;
  assign n52696 = ~n44867 & n52695 ;
  assign n52697 = n52696 ^ n27309 ^ n3949 ;
  assign n52698 = ( ~n3379 & n10237 ) | ( ~n3379 & n14488 ) | ( n10237 & n14488 ) ;
  assign n52699 = ( n19183 & ~n24537 ) | ( n19183 & n51518 ) | ( ~n24537 & n51518 ) ;
  assign n52700 = ( n38566 & ~n47373 ) | ( n38566 & n48015 ) | ( ~n47373 & n48015 ) ;
  assign n52701 = ( ~n3805 & n9738 ) | ( ~n3805 & n17205 ) | ( n9738 & n17205 ) ;
  assign n52702 = n29278 ^ n19628 ^ 1'b0 ;
  assign n52703 = n26423 & n52702 ;
  assign n52704 = ( n522 & n10042 ) | ( n522 & n52703 ) | ( n10042 & n52703 ) ;
  assign n52706 = n5494 & n15214 ;
  assign n52705 = n20267 | n27309 ;
  assign n52707 = n52706 ^ n52705 ^ 1'b0 ;
  assign n52708 = n36056 ^ n3248 ^ 1'b0 ;
  assign n52709 = n14021 ^ n8450 ^ 1'b0 ;
  assign n52710 = n52709 ^ n33557 ^ 1'b0 ;
  assign n52711 = ( n11435 & ~n24319 ) | ( n11435 & n26217 ) | ( ~n24319 & n26217 ) ;
  assign n52712 = n52711 ^ n12173 ^ n887 ;
  assign n52713 = n52712 ^ n43465 ^ n12793 ;
  assign n52714 = ( n13018 & n36131 ) | ( n13018 & ~n45266 ) | ( n36131 & ~n45266 ) ;
  assign n52715 = n52714 ^ n34877 ^ n18836 ;
  assign n52716 = n49160 ^ n26031 ^ n18910 ;
  assign n52718 = n4920 & n31062 ;
  assign n52717 = ( ~n4596 & n6397 ) | ( ~n4596 & n27035 ) | ( n6397 & n27035 ) ;
  assign n52719 = n52718 ^ n52717 ^ n18236 ;
  assign n52720 = n26591 & n40135 ;
  assign n52721 = n35546 ^ n16699 ^ n10982 ;
  assign n52722 = n52721 ^ n17796 ^ 1'b0 ;
  assign n52724 = n31610 ^ n10260 ^ n1898 ;
  assign n52723 = ( n13398 & n16154 ) | ( n13398 & ~n22892 ) | ( n16154 & ~n22892 ) ;
  assign n52725 = n52724 ^ n52723 ^ n29970 ;
  assign n52726 = n7079 & ~n23367 ;
  assign n52727 = n52726 ^ n36209 ^ 1'b0 ;
  assign n52728 = n30005 ^ n6959 ^ n1366 ;
  assign n52729 = n1274 | n12089 ;
  assign n52730 = ( ~n24577 & n52728 ) | ( ~n24577 & n52729 ) | ( n52728 & n52729 ) ;
  assign n52731 = n43010 & n52730 ;
  assign n52732 = n52731 ^ n26392 ^ 1'b0 ;
  assign n52733 = n1977 & n34729 ;
  assign n52734 = ~n18596 & n52733 ;
  assign n52735 = n9165 ^ n6796 ^ 1'b0 ;
  assign n52736 = ~n11881 & n52735 ;
  assign n52737 = n26789 ^ n25279 ^ n15116 ;
  assign n52738 = ( n26544 & n52736 ) | ( n26544 & n52737 ) | ( n52736 & n52737 ) ;
  assign n52739 = n10412 ^ n8230 ^ n5458 ;
  assign n52740 = ( n6828 & ~n16228 ) | ( n6828 & n23603 ) | ( ~n16228 & n23603 ) ;
  assign n52741 = ( ~n6395 & n13580 ) | ( ~n6395 & n52740 ) | ( n13580 & n52740 ) ;
  assign n52742 = n39930 ^ n20242 ^ n7262 ;
  assign n52744 = ~n9067 & n42967 ;
  assign n52743 = n51717 ^ n35073 ^ n6330 ;
  assign n52745 = n52744 ^ n52743 ^ n12980 ;
  assign n52746 = n47854 ^ n13004 ^ n10871 ;
  assign n52747 = ( n11918 & ~n30802 ) | ( n11918 & n48099 ) | ( ~n30802 & n48099 ) ;
  assign n52748 = n5692 & ~n47335 ;
  assign n52749 = ~n12641 & n52748 ;
  assign n52750 = ~n7930 & n45666 ;
  assign n52751 = ( n12262 & n24622 ) | ( n12262 & n41388 ) | ( n24622 & n41388 ) ;
  assign n52752 = ( ~n24013 & n36012 ) | ( ~n24013 & n37824 ) | ( n36012 & n37824 ) ;
  assign n52753 = ( ~n4629 & n27311 ) | ( ~n4629 & n34194 ) | ( n27311 & n34194 ) ;
  assign n52754 = ( n14842 & ~n25699 ) | ( n14842 & n52753 ) | ( ~n25699 & n52753 ) ;
  assign n52755 = n12604 | n20309 ;
  assign n52756 = n30311 | n52755 ;
  assign n52757 = ~n13558 & n15704 ;
  assign n52758 = n34278 & n52757 ;
  assign n52759 = ( n41213 & n52756 ) | ( n41213 & ~n52758 ) | ( n52756 & ~n52758 ) ;
  assign n52760 = ( n50243 & ~n52754 ) | ( n50243 & n52759 ) | ( ~n52754 & n52759 ) ;
  assign n52761 = n5040 ^ n4006 ^ 1'b0 ;
  assign n52762 = n16290 & n52761 ;
  assign n52763 = n5014 & ~n10442 ;
  assign n52764 = ( ~n47645 & n52762 ) | ( ~n47645 & n52763 ) | ( n52762 & n52763 ) ;
  assign n52765 = ( n4748 & ~n27982 ) | ( n4748 & n52764 ) | ( ~n27982 & n52764 ) ;
  assign n52766 = ( n4080 & n26698 ) | ( n4080 & n40134 ) | ( n26698 & n40134 ) ;
  assign n52767 = ~n12025 & n51984 ;
  assign n52768 = n23268 ^ n10702 ^ n7109 ;
  assign n52769 = n52768 ^ n3154 ^ 1'b0 ;
  assign n52770 = n52769 ^ n17518 ^ n283 ;
  assign n52771 = n37915 ^ n15642 ^ n7842 ;
  assign n52772 = n22979 & ~n49925 ;
  assign n52773 = ~n2227 & n52772 ;
  assign n52775 = n2619 & n33870 ;
  assign n52776 = n22033 & n52775 ;
  assign n52774 = ~n1955 & n9210 ;
  assign n52777 = n52776 ^ n52774 ^ 1'b0 ;
  assign n52778 = n25517 | n52777 ;
  assign n52779 = n18911 ^ n13151 ^ n10430 ;
  assign n52780 = ( n8130 & n31062 ) | ( n8130 & ~n52779 ) | ( n31062 & ~n52779 ) ;
  assign n52781 = n52780 ^ n4288 ^ 1'b0 ;
  assign n52782 = n2582 | n52781 ;
  assign n52783 = n10543 ^ n10438 ^ 1'b0 ;
  assign n52784 = n35036 ^ n2265 ^ x141 ;
  assign n52785 = ( n6926 & ~n39273 ) | ( n6926 & n52784 ) | ( ~n39273 & n52784 ) ;
  assign n52786 = ( ~n48247 & n50470 ) | ( ~n48247 & n52785 ) | ( n50470 & n52785 ) ;
  assign n52787 = n51238 ^ n21450 ^ n8807 ;
  assign n52789 = n45719 ^ n28435 ^ n549 ;
  assign n52788 = n12005 ^ n8945 ^ 1'b0 ;
  assign n52790 = n52789 ^ n52788 ^ n23567 ;
  assign n52791 = n52790 ^ n52068 ^ 1'b0 ;
  assign n52797 = ( n8378 & ~n15765 ) | ( n8378 & n16670 ) | ( ~n15765 & n16670 ) ;
  assign n52795 = n17815 & ~n48373 ;
  assign n52796 = n51242 & n52795 ;
  assign n52792 = ( ~n10606 & n22705 ) | ( ~n10606 & n33538 ) | ( n22705 & n33538 ) ;
  assign n52793 = n52792 ^ n13245 ^ 1'b0 ;
  assign n52794 = n40787 | n52793 ;
  assign n52798 = n52797 ^ n52796 ^ n52794 ;
  assign n52799 = ~n12526 & n32678 ;
  assign n52800 = n26465 ^ n21632 ^ n1102 ;
  assign n52801 = ( ~n18230 & n47240 ) | ( ~n18230 & n52800 ) | ( n47240 & n52800 ) ;
  assign n52802 = n12987 ^ n9837 ^ 1'b0 ;
  assign n52803 = ~n27540 & n52802 ;
  assign n52804 = n28379 ^ n24150 ^ 1'b0 ;
  assign n52805 = ( n1159 & n3685 ) | ( n1159 & ~n15282 ) | ( n3685 & ~n15282 ) ;
  assign n52806 = n52805 ^ n10711 ^ 1'b0 ;
  assign n52807 = n52804 & n52806 ;
  assign n52808 = n40971 ^ n39209 ^ n1823 ;
  assign n52809 = ( ~n9821 & n47778 ) | ( ~n9821 & n52808 ) | ( n47778 & n52808 ) ;
  assign n52810 = ~n2681 & n21932 ;
  assign n52811 = n42008 & n52810 ;
  assign n52812 = n52716 & ~n52811 ;
  assign n52813 = ~n52809 & n52812 ;
  assign n52814 = ( n17975 & n38023 ) | ( n17975 & n38994 ) | ( n38023 & n38994 ) ;
  assign n52815 = n52814 ^ n30984 ^ n24433 ;
  assign n52816 = n13305 ^ n12827 ^ n7749 ;
  assign n52817 = n52816 ^ n23318 ^ n21606 ;
  assign n52819 = ( n5244 & n14610 ) | ( n5244 & ~n21113 ) | ( n14610 & ~n21113 ) ;
  assign n52818 = ( n1556 & n9819 ) | ( n1556 & ~n41948 ) | ( n9819 & ~n41948 ) ;
  assign n52820 = n52819 ^ n52818 ^ n44922 ;
  assign n52821 = n52820 ^ n20402 ^ 1'b0 ;
  assign n52822 = n14361 ^ n558 ^ 1'b0 ;
  assign n52823 = n50699 ^ n35764 ^ n8087 ;
  assign n52824 = n52823 ^ n32014 ^ n4575 ;
  assign n52825 = ( ~n12272 & n52822 ) | ( ~n12272 & n52824 ) | ( n52822 & n52824 ) ;
  assign n52826 = n32192 ^ n30914 ^ n25360 ;
  assign n52827 = ( n3640 & n7157 ) | ( n3640 & ~n8281 ) | ( n7157 & ~n8281 ) ;
  assign n52828 = n28788 & ~n51323 ;
  assign n52829 = ( n37007 & n52827 ) | ( n37007 & ~n52828 ) | ( n52827 & ~n52828 ) ;
  assign n52830 = ( n2004 & n17745 ) | ( n2004 & n24808 ) | ( n17745 & n24808 ) ;
  assign n52831 = n29995 ^ n3132 ^ 1'b0 ;
  assign n52832 = n52830 & n52831 ;
  assign n52833 = ( ~n8442 & n17476 ) | ( ~n8442 & n52832 ) | ( n17476 & n52832 ) ;
  assign n52834 = ( n30279 & n41275 ) | ( n30279 & n45955 ) | ( n41275 & n45955 ) ;
  assign n52835 = n52834 ^ n28796 ^ 1'b0 ;
  assign n52836 = n28670 ^ n22628 ^ x16 ;
  assign n52837 = n24329 ^ n10285 ^ 1'b0 ;
  assign n52838 = n52836 | n52837 ;
  assign n52839 = ( n7863 & n28848 ) | ( n7863 & ~n31301 ) | ( n28848 & ~n31301 ) ;
  assign n52840 = n24786 ^ n8691 ^ 1'b0 ;
  assign n52841 = n21773 ^ n12408 ^ n12152 ;
  assign n52842 = n52841 ^ n17974 ^ n6566 ;
  assign n52843 = n45694 ^ n30187 ^ 1'b0 ;
  assign n52849 = n20961 ^ n18997 ^ n3114 ;
  assign n52850 = n52849 ^ n32380 ^ n31602 ;
  assign n52846 = n32682 ^ n13637 ^ n2048 ;
  assign n52847 = ( n3174 & n32003 ) | ( n3174 & n52846 ) | ( n32003 & n52846 ) ;
  assign n52844 = n16670 & n43388 ;
  assign n52845 = n52844 ^ n12662 ^ 1'b0 ;
  assign n52848 = n52847 ^ n52845 ^ n26856 ;
  assign n52851 = n52850 ^ n52848 ^ n28781 ;
  assign n52852 = ( n26836 & ~n46543 ) | ( n26836 & n52851 ) | ( ~n46543 & n52851 ) ;
  assign n52853 = n31180 ^ n11170 ^ 1'b0 ;
  assign n52854 = n49815 ^ n27369 ^ 1'b0 ;
  assign n52855 = n27817 | n36395 ;
  assign n52856 = ( n13940 & n17518 ) | ( n13940 & ~n52855 ) | ( n17518 & ~n52855 ) ;
  assign n52857 = n52157 & n52856 ;
  assign n52858 = ( n796 & ~n2567 ) | ( n796 & n19450 ) | ( ~n2567 & n19450 ) ;
  assign n52859 = n5551 & ~n52858 ;
  assign n52860 = ( n5792 & n9307 ) | ( n5792 & n41356 ) | ( n9307 & n41356 ) ;
  assign n52861 = n23013 ^ n12824 ^ n11602 ;
  assign n52862 = n37734 ^ n14852 ^ n4017 ;
  assign n52863 = ( n4049 & ~n4166 ) | ( n4049 & n52862 ) | ( ~n4166 & n52862 ) ;
  assign n52864 = ( n14992 & ~n33375 ) | ( n14992 & n38166 ) | ( ~n33375 & n38166 ) ;
  assign n52865 = ( ~n18725 & n35621 ) | ( ~n18725 & n39984 ) | ( n35621 & n39984 ) ;
  assign n52866 = ( n8168 & ~n52864 ) | ( n8168 & n52865 ) | ( ~n52864 & n52865 ) ;
  assign n52867 = ( n3123 & n4557 ) | ( n3123 & ~n5914 ) | ( n4557 & ~n5914 ) ;
  assign n52868 = ( n6553 & n6684 ) | ( n6553 & n50963 ) | ( n6684 & n50963 ) ;
  assign n52869 = ( n7303 & ~n40429 ) | ( n7303 & n52868 ) | ( ~n40429 & n52868 ) ;
  assign n52870 = n4399 ^ n4072 ^ n482 ;
  assign n52871 = ~n1826 & n10828 ;
  assign n52872 = n11869 | n24215 ;
  assign n52873 = n52871 & ~n52872 ;
  assign n52874 = n52873 ^ n46629 ^ 1'b0 ;
  assign n52875 = ~n2541 & n21466 ;
  assign n52876 = n52875 ^ n16584 ^ 1'b0 ;
  assign n52877 = ( n4431 & ~n8293 ) | ( n4431 & n52876 ) | ( ~n8293 & n52876 ) ;
  assign n52878 = n16741 & ~n52877 ;
  assign n52879 = ~n10111 & n52878 ;
  assign n52880 = n933 | n45482 ;
  assign n52881 = n20857 & ~n52880 ;
  assign n52882 = n3384 | n46334 ;
  assign n52883 = n42981 & ~n52882 ;
  assign n52884 = n25441 ^ n5493 ^ n5100 ;
  assign n52885 = ( n34327 & n34965 ) | ( n34327 & ~n52884 ) | ( n34965 & ~n52884 ) ;
  assign n52886 = n6587 | n24343 ;
  assign n52887 = n26811 ^ n14428 ^ n11957 ;
  assign n52888 = n52887 ^ n26587 ^ n12332 ;
  assign n52889 = n9586 & ~n52888 ;
  assign n52890 = ( ~n28399 & n37907 ) | ( ~n28399 & n52889 ) | ( n37907 & n52889 ) ;
  assign n52891 = ~n10785 & n42348 ;
  assign n52892 = ~n3218 & n52891 ;
  assign n52893 = ( n5982 & n15074 ) | ( n5982 & ~n18349 ) | ( n15074 & ~n18349 ) ;
  assign n52894 = n52893 ^ n48343 ^ n15715 ;
  assign n52895 = n35501 ^ n15724 ^ 1'b0 ;
  assign n52896 = n19476 & ~n28540 ;
  assign n52897 = ( n4187 & n17594 ) | ( n4187 & ~n52896 ) | ( n17594 & ~n52896 ) ;
  assign n52898 = n32417 ^ n13848 ^ n9000 ;
  assign n52899 = n52898 ^ n5357 ^ n2951 ;
  assign n52900 = n1075 | n51016 ;
  assign n52901 = n22257 | n52900 ;
  assign n52902 = ( n6907 & n36173 ) | ( n6907 & ~n50571 ) | ( n36173 & ~n50571 ) ;
  assign n52903 = ( n9302 & n22805 ) | ( n9302 & ~n24699 ) | ( n22805 & ~n24699 ) ;
  assign n52904 = n52903 ^ n45519 ^ n20983 ;
  assign n52905 = n29438 ^ n17388 ^ n7335 ;
  assign n52906 = n52905 ^ n39837 ^ n33467 ;
  assign n52908 = ( n2415 & n18476 ) | ( n2415 & ~n49125 ) | ( n18476 & ~n49125 ) ;
  assign n52907 = n17307 | n26428 ;
  assign n52909 = n52908 ^ n52907 ^ n34393 ;
  assign n52910 = n31772 ^ n17916 ^ n8765 ;
  assign n52911 = ( n12129 & ~n15811 ) | ( n12129 & n52910 ) | ( ~n15811 & n52910 ) ;
  assign n52912 = n52911 ^ n32546 ^ n21528 ;
  assign n52913 = n52912 ^ n22570 ^ n20883 ;
  assign n52914 = n52913 ^ n38744 ^ 1'b0 ;
  assign n52915 = n45616 ^ n40854 ^ n31588 ;
  assign n52916 = n43080 ^ n18908 ^ n8567 ;
  assign n52918 = n38879 ^ n25030 ^ n24472 ;
  assign n52917 = ~n16026 & n29249 ;
  assign n52919 = n52918 ^ n52917 ^ 1'b0 ;
  assign n52920 = n52919 ^ n51067 ^ n49938 ;
  assign n52921 = ( ~n8959 & n52916 ) | ( ~n8959 & n52920 ) | ( n52916 & n52920 ) ;
  assign n52922 = ( n21966 & n52915 ) | ( n21966 & ~n52921 ) | ( n52915 & ~n52921 ) ;
  assign n52923 = n42363 ^ n21813 ^ n18907 ;
  assign n52924 = n26235 & ~n30111 ;
  assign n52925 = n47948 ^ n30914 ^ 1'b0 ;
  assign n52926 = n1600 & n52925 ;
  assign n52927 = ( n4538 & n19939 ) | ( n4538 & ~n52926 ) | ( n19939 & ~n52926 ) ;
  assign n52928 = n5338 & ~n23732 ;
  assign n52929 = ~n52927 & n52928 ;
  assign n52930 = n3095 & ~n4865 ;
  assign n52931 = n50931 & n52930 ;
  assign n52932 = ( n3390 & n16879 ) | ( n3390 & n23676 ) | ( n16879 & n23676 ) ;
  assign n52933 = ( x179 & n32025 ) | ( x179 & ~n52932 ) | ( n32025 & ~n52932 ) ;
  assign n52934 = n51782 ^ n24109 ^ n3668 ;
  assign n52935 = n31799 ^ n12668 ^ 1'b0 ;
  assign n52936 = n16968 ^ n2562 ^ 1'b0 ;
  assign n52937 = ~n4600 & n52936 ;
  assign n52938 = n52935 & ~n52937 ;
  assign n52939 = n27406 ^ n24496 ^ n7063 ;
  assign n52940 = n48742 ^ n45758 ^ n34766 ;
  assign n52941 = n19012 & ~n27503 ;
  assign n52942 = n52941 ^ n34498 ^ 1'b0 ;
  assign n52943 = ( n21023 & n23964 ) | ( n21023 & n32005 ) | ( n23964 & n32005 ) ;
  assign n52944 = ( n29255 & n52942 ) | ( n29255 & n52943 ) | ( n52942 & n52943 ) ;
  assign n52945 = n24770 ^ n12056 ^ 1'b0 ;
  assign n52946 = ( n15360 & n30321 ) | ( n15360 & ~n34183 ) | ( n30321 & ~n34183 ) ;
  assign n52947 = n16250 ^ n15488 ^ n11557 ;
  assign n52948 = n52947 ^ n14134 ^ 1'b0 ;
  assign n52949 = n52946 & ~n52948 ;
  assign n52950 = n15303 & n52949 ;
  assign n52951 = ~n346 & n52950 ;
  assign n52952 = n944 | n21286 ;
  assign n52953 = n52952 ^ n869 ^ 1'b0 ;
  assign n52954 = n52953 ^ n37660 ^ n19267 ;
  assign n52955 = n14226 & n42626 ;
  assign n52956 = n52955 ^ n39598 ^ n10378 ;
  assign n52957 = n17079 ^ n16125 ^ n2835 ;
  assign n52958 = ( n8153 & ~n15260 ) | ( n8153 & n52957 ) | ( ~n15260 & n52957 ) ;
  assign n52959 = ( n11124 & ~n15192 ) | ( n11124 & n44273 ) | ( ~n15192 & n44273 ) ;
  assign n52960 = ( ~n427 & n51869 ) | ( ~n427 & n52959 ) | ( n51869 & n52959 ) ;
  assign n52961 = ( n34601 & n51712 ) | ( n34601 & n52960 ) | ( n51712 & n52960 ) ;
  assign n52962 = ( n20619 & ~n52958 ) | ( n20619 & n52961 ) | ( ~n52958 & n52961 ) ;
  assign n52963 = n30687 ^ n27218 ^ n16273 ;
  assign n52964 = n52963 ^ n35394 ^ n7433 ;
  assign n52965 = ( n5622 & n7457 ) | ( n5622 & ~n10516 ) | ( n7457 & ~n10516 ) ;
  assign n52966 = n26467 ^ n21735 ^ n8896 ;
  assign n52967 = ( n30354 & n52965 ) | ( n30354 & n52966 ) | ( n52965 & n52966 ) ;
  assign n52969 = n10441 ^ n9718 ^ 1'b0 ;
  assign n52970 = n35513 & ~n52969 ;
  assign n52968 = ( n16855 & n19155 ) | ( n16855 & n43649 ) | ( n19155 & n43649 ) ;
  assign n52971 = n52970 ^ n52968 ^ n22219 ;
  assign n52972 = n19819 ^ n14048 ^ n7599 ;
  assign n52973 = ( n23196 & n52740 ) | ( n23196 & ~n52972 ) | ( n52740 & ~n52972 ) ;
  assign n52974 = n5001 & ~n27294 ;
  assign n52975 = n52974 ^ n26377 ^ 1'b0 ;
  assign n52976 = n52975 ^ n15840 ^ n9213 ;
  assign n52982 = n6751 ^ n648 ^ 1'b0 ;
  assign n52983 = n1656 | n52982 ;
  assign n52981 = n43029 ^ n29264 ^ n16004 ;
  assign n52977 = n27447 & ~n40512 ;
  assign n52978 = n52977 ^ n6480 ^ 1'b0 ;
  assign n52979 = n52978 ^ n11145 ^ 1'b0 ;
  assign n52980 = n45045 & n52979 ;
  assign n52984 = n52983 ^ n52981 ^ n52980 ;
  assign n52988 = ~n15706 & n32892 ;
  assign n52989 = n52988 ^ n31689 ^ 1'b0 ;
  assign n52985 = n28979 & n46019 ;
  assign n52986 = ~n10944 & n52985 ;
  assign n52987 = n52986 ^ n8569 ^ 1'b0 ;
  assign n52990 = n52989 ^ n52987 ^ n13098 ;
  assign n52991 = n47443 ^ n18685 ^ 1'b0 ;
  assign n52992 = n52991 ^ n43803 ^ n10619 ;
  assign n52993 = ( n810 & n9403 ) | ( n810 & ~n37820 ) | ( n9403 & ~n37820 ) ;
  assign n52994 = n1616 & n9415 ;
  assign n52995 = ( n1430 & n50500 ) | ( n1430 & ~n52994 ) | ( n50500 & ~n52994 ) ;
  assign n52996 = n52995 ^ n37523 ^ n33429 ;
  assign n52997 = ( ~n17313 & n28714 ) | ( ~n17313 & n36657 ) | ( n28714 & n36657 ) ;
  assign n52998 = n52997 ^ n20321 ^ n7349 ;
  assign n52999 = n29630 ^ n4460 ^ n4014 ;
  assign n53001 = ( ~n5806 & n29209 ) | ( ~n5806 & n31575 ) | ( n29209 & n31575 ) ;
  assign n53002 = n53001 ^ n28299 ^ n2032 ;
  assign n53000 = n15073 & n29172 ;
  assign n53003 = n53002 ^ n53000 ^ 1'b0 ;
  assign n53004 = n31291 ^ n25988 ^ n8596 ;
  assign n53005 = ~n11038 & n53004 ;
  assign n53006 = n53005 ^ n8414 ^ 1'b0 ;
  assign n53007 = ~n8050 & n28357 ;
  assign n53008 = ~n47659 & n53007 ;
  assign n53009 = ( n6730 & n18071 ) | ( n6730 & n27940 ) | ( n18071 & n27940 ) ;
  assign n53010 = n3108 | n10984 ;
  assign n53011 = n53009 & ~n53010 ;
  assign n53012 = n53011 ^ n13559 ^ n5832 ;
  assign n53014 = n30170 ^ n27893 ^ n10395 ;
  assign n53013 = n11726 ^ n4833 ^ n1420 ;
  assign n53015 = n53014 ^ n53013 ^ 1'b0 ;
  assign n53016 = n53015 ^ n14212 ^ 1'b0 ;
  assign n53017 = n50716 ^ n24543 ^ n14308 ;
  assign n53018 = ( n19686 & n23284 ) | ( n19686 & n29773 ) | ( n23284 & n29773 ) ;
  assign n53019 = n22866 & n31057 ;
  assign n53020 = n47433 ^ n22889 ^ n15995 ;
  assign n53021 = ( x37 & n16765 ) | ( x37 & n20437 ) | ( n16765 & n20437 ) ;
  assign n53022 = ( n13687 & n19948 ) | ( n13687 & n53021 ) | ( n19948 & n53021 ) ;
  assign n53023 = n7485 & ~n37402 ;
  assign n53024 = ~n23017 & n53023 ;
  assign n53025 = n53024 ^ n24342 ^ n11494 ;
  assign n53026 = n12226 | n15488 ;
  assign n53027 = n15718 | n53026 ;
  assign n53028 = n18091 ^ n5544 ^ 1'b0 ;
  assign n53029 = ~n21660 & n53028 ;
  assign n53030 = ( ~n35890 & n44330 ) | ( ~n35890 & n53029 ) | ( n44330 & n53029 ) ;
  assign n53031 = n30141 ^ n8364 ^ 1'b0 ;
  assign n53032 = n39644 ^ n17742 ^ n16015 ;
  assign n53033 = ( n30739 & n46378 ) | ( n30739 & n53032 ) | ( n46378 & n53032 ) ;
  assign n53034 = n53033 ^ n36497 ^ n9666 ;
  assign n53035 = ( n397 & ~n17055 ) | ( n397 & n35918 ) | ( ~n17055 & n35918 ) ;
  assign n53036 = ( n11269 & n12754 ) | ( n11269 & ~n53035 ) | ( n12754 & ~n53035 ) ;
  assign n53037 = n4630 & ~n34127 ;
  assign n53038 = ( n2240 & ~n8457 ) | ( n2240 & n53037 ) | ( ~n8457 & n53037 ) ;
  assign n53039 = ( n14664 & n31724 ) | ( n14664 & ~n53038 ) | ( n31724 & ~n53038 ) ;
  assign n53040 = n34782 ^ n28494 ^ n5415 ;
  assign n53041 = ( n368 & n1591 ) | ( n368 & ~n9651 ) | ( n1591 & ~n9651 ) ;
  assign n53042 = n53041 ^ n32728 ^ 1'b0 ;
  assign n53043 = ~n24705 & n53042 ;
  assign n53044 = n53043 ^ n51622 ^ n36897 ;
  assign n53045 = n2307 & n25355 ;
  assign n53046 = ( n1142 & n6380 ) | ( n1142 & n53045 ) | ( n6380 & n53045 ) ;
  assign n53047 = n23676 | n27237 ;
  assign n53048 = n53047 ^ n6904 ^ 1'b0 ;
  assign n53049 = n53048 ^ n44873 ^ 1'b0 ;
  assign n53050 = n10604 & ~n53049 ;
  assign n53051 = n8378 | n13433 ;
  assign n53052 = n53051 ^ n50103 ^ 1'b0 ;
  assign n53053 = n4209 | n53052 ;
  assign n53054 = n53053 ^ n8402 ^ 1'b0 ;
  assign n53055 = n8566 & ~n24577 ;
  assign n53056 = n18730 & n53055 ;
  assign n53057 = n42513 ^ n7540 ^ 1'b0 ;
  assign n53058 = n23084 & ~n53057 ;
  assign n53059 = ( n13519 & ~n52958 ) | ( n13519 & n53058 ) | ( ~n52958 & n53058 ) ;
  assign n53060 = ( n1902 & n2100 ) | ( n1902 & ~n13361 ) | ( n2100 & ~n13361 ) ;
  assign n53061 = n15523 ^ x8 ^ 1'b0 ;
  assign n53062 = ( n9710 & n10651 ) | ( n9710 & ~n53061 ) | ( n10651 & ~n53061 ) ;
  assign n53063 = ( n33071 & n53060 ) | ( n33071 & n53062 ) | ( n53060 & n53062 ) ;
  assign n53064 = n51645 ^ n19915 ^ n904 ;
  assign n53065 = ( n7263 & ~n20723 ) | ( n7263 & n24950 ) | ( ~n20723 & n24950 ) ;
  assign n53066 = n53065 ^ n13032 ^ n12950 ;
  assign n53067 = ( n18381 & n53064 ) | ( n18381 & n53066 ) | ( n53064 & n53066 ) ;
  assign n53068 = ( n28019 & n30358 ) | ( n28019 & n53067 ) | ( n30358 & n53067 ) ;
  assign n53071 = ( ~n5724 & n8016 ) | ( ~n5724 & n19612 ) | ( n8016 & n19612 ) ;
  assign n53070 = ( n3109 & n4293 ) | ( n3109 & ~n8510 ) | ( n4293 & ~n8510 ) ;
  assign n53069 = n44157 ^ n27928 ^ n9993 ;
  assign n53072 = n53071 ^ n53070 ^ n53069 ;
  assign n53073 = n28345 ^ n27326 ^ n24164 ;
  assign n53074 = ( n17606 & n31418 ) | ( n17606 & ~n42205 ) | ( n31418 & ~n42205 ) ;
  assign n53075 = n53074 ^ n38962 ^ n4045 ;
  assign n53076 = n11399 | n39688 ;
  assign n53077 = n53076 ^ n6594 ^ 1'b0 ;
  assign n53078 = ( n7306 & n45352 ) | ( n7306 & ~n45967 ) | ( n45352 & ~n45967 ) ;
  assign n53079 = n53078 ^ n26006 ^ 1'b0 ;
  assign n53080 = n4257 & n53079 ;
  assign n53081 = n37573 ^ n9543 ^ n9305 ;
  assign n53082 = ( ~n6875 & n16429 ) | ( ~n6875 & n43008 ) | ( n16429 & n43008 ) ;
  assign n53083 = ~n53081 & n53082 ;
  assign n53084 = n53083 ^ n16006 ^ 1'b0 ;
  assign n53085 = ( n923 & ~n27264 ) | ( n923 & n49063 ) | ( ~n27264 & n49063 ) ;
  assign n53086 = n19682 ^ n12409 ^ n6804 ;
  assign n53087 = n18720 & n22382 ;
  assign n53088 = n53086 & n53087 ;
  assign n53089 = ( ~n19110 & n46619 ) | ( ~n19110 & n53088 ) | ( n46619 & n53088 ) ;
  assign n53090 = n42614 ^ n14798 ^ n11893 ;
  assign n53091 = n10515 & n25047 ;
  assign n53092 = ~n53090 & n53091 ;
  assign n53093 = ( n25601 & n34635 ) | ( n25601 & n43808 ) | ( n34635 & n43808 ) ;
  assign n53094 = ( n29402 & n53092 ) | ( n29402 & n53093 ) | ( n53092 & n53093 ) ;
  assign n53095 = n26625 ^ n21851 ^ n20487 ;
  assign n53096 = n53095 ^ n36365 ^ n3747 ;
  assign n53097 = ( n5707 & n6986 ) | ( n5707 & n43704 ) | ( n6986 & n43704 ) ;
  assign n53098 = n53097 ^ n10118 ^ n4825 ;
  assign n53099 = ( n23013 & n53096 ) | ( n23013 & ~n53098 ) | ( n53096 & ~n53098 ) ;
  assign n53100 = ( ~n7514 & n30938 ) | ( ~n7514 & n37153 ) | ( n30938 & n37153 ) ;
  assign n53101 = n30691 ^ n3753 ^ 1'b0 ;
  assign n53102 = ~n4726 & n6930 ;
  assign n53103 = ( n34157 & n52910 ) | ( n34157 & ~n53102 ) | ( n52910 & ~n53102 ) ;
  assign n53104 = n11330 ^ n4648 ^ 1'b0 ;
  assign n53105 = n44088 & ~n53104 ;
  assign n53106 = n1293 & ~n43626 ;
  assign n53107 = n53106 ^ n15701 ^ 1'b0 ;
  assign n53108 = n11676 & n37068 ;
  assign n53109 = n53108 ^ n48341 ^ 1'b0 ;
  assign n53111 = ( n8517 & n25611 ) | ( n8517 & ~n33921 ) | ( n25611 & ~n33921 ) ;
  assign n53110 = n24417 | n45815 ;
  assign n53112 = n53111 ^ n53110 ^ 1'b0 ;
  assign n53113 = n47799 & n53112 ;
  assign n53116 = n1028 & n25769 ;
  assign n53117 = n53116 ^ n2687 ^ 1'b0 ;
  assign n53118 = ( n806 & ~n14349 ) | ( n806 & n53117 ) | ( ~n14349 & n53117 ) ;
  assign n53114 = n22376 ^ n10848 ^ n3054 ;
  assign n53115 = n53114 ^ n46303 ^ n5621 ;
  assign n53119 = n53118 ^ n53115 ^ 1'b0 ;
  assign n53120 = n24510 ^ n17849 ^ n15553 ;
  assign n53121 = ( n12200 & ~n44716 ) | ( n12200 & n53120 ) | ( ~n44716 & n53120 ) ;
  assign n53122 = n53121 ^ n16204 ^ 1'b0 ;
  assign n53123 = ~n50543 & n53122 ;
  assign n53124 = ( n8806 & n18683 ) | ( n8806 & n53123 ) | ( n18683 & n53123 ) ;
  assign n53125 = ( n10692 & ~n40383 ) | ( n10692 & n52805 ) | ( ~n40383 & n52805 ) ;
  assign n53126 = n47696 ^ n12995 ^ n5615 ;
  assign n53127 = n52768 ^ n18654 ^ x198 ;
  assign n53128 = ( ~n3052 & n22630 ) | ( ~n3052 & n38560 ) | ( n22630 & n38560 ) ;
  assign n53129 = ( n5910 & n18327 ) | ( n5910 & ~n36853 ) | ( n18327 & ~n36853 ) ;
  assign n53130 = n35613 ^ n10570 ^ n9278 ;
  assign n53131 = ( n25228 & ~n27062 ) | ( n25228 & n53130 ) | ( ~n27062 & n53130 ) ;
  assign n53132 = n12830 & ~n21606 ;
  assign n53133 = n53131 & n53132 ;
  assign n53134 = n40494 ^ n33536 ^ n27213 ;
  assign n53135 = n14482 | n53134 ;
  assign n53136 = n53135 ^ n11746 ^ 1'b0 ;
  assign n53137 = n23120 ^ n4327 ^ n2862 ;
  assign n53138 = ( ~n692 & n17762 ) | ( ~n692 & n41166 ) | ( n17762 & n41166 ) ;
  assign n53139 = ~n28048 & n53138 ;
  assign n53140 = ( n21047 & n28669 ) | ( n21047 & n50508 ) | ( n28669 & n50508 ) ;
  assign n53141 = n18269 ^ n17088 ^ n8028 ;
  assign n53142 = n48430 ^ n20133 ^ n10153 ;
  assign n53143 = n53142 ^ n23496 ^ 1'b0 ;
  assign n53144 = ( n5271 & n53141 ) | ( n5271 & n53143 ) | ( n53141 & n53143 ) ;
  assign n53145 = ( n3033 & n22432 ) | ( n3033 & ~n22845 ) | ( n22432 & ~n22845 ) ;
  assign n53146 = ( n8168 & n16948 ) | ( n8168 & ~n53145 ) | ( n16948 & ~n53145 ) ;
  assign n53147 = n35911 ^ n25725 ^ n5188 ;
  assign n53148 = ( ~n9510 & n33827 ) | ( ~n9510 & n51328 ) | ( n33827 & n51328 ) ;
  assign n53149 = ( n1561 & n8980 ) | ( n1561 & n53148 ) | ( n8980 & n53148 ) ;
  assign n53152 = ( n10702 & n22907 ) | ( n10702 & ~n25970 ) | ( n22907 & ~n25970 ) ;
  assign n53150 = n26264 ^ n14924 ^ n11340 ;
  assign n53151 = ( n19822 & ~n25447 ) | ( n19822 & n53150 ) | ( ~n25447 & n53150 ) ;
  assign n53153 = n53152 ^ n53151 ^ n13022 ;
  assign n53154 = ( n18559 & n43065 ) | ( n18559 & ~n53153 ) | ( n43065 & ~n53153 ) ;
  assign n53155 = ( ~n3640 & n18022 ) | ( ~n3640 & n43376 ) | ( n18022 & n43376 ) ;
  assign n53156 = ~n46639 & n53155 ;
  assign n53157 = n53156 ^ n13521 ^ 1'b0 ;
  assign n53158 = ( n19782 & n24241 ) | ( n19782 & n44820 ) | ( n24241 & n44820 ) ;
  assign n53159 = n20229 ^ n9435 ^ n6054 ;
  assign n53160 = n3639 | n7605 ;
  assign n53161 = n53160 ^ n32855 ^ 1'b0 ;
  assign n53163 = ~n7988 & n43558 ;
  assign n53162 = n34321 ^ n12532 ^ n7887 ;
  assign n53164 = n53163 ^ n53162 ^ n17000 ;
  assign n53165 = ( n15152 & n27005 ) | ( n15152 & n29257 ) | ( n27005 & n29257 ) ;
  assign n53166 = n53165 ^ n31263 ^ n15862 ;
  assign n53167 = n44752 ^ n33442 ^ n8322 ;
  assign n53169 = n4779 | n8450 ;
  assign n53170 = n53169 ^ n16894 ^ 1'b0 ;
  assign n53171 = ~n24833 & n53170 ;
  assign n53172 = n13702 & n53171 ;
  assign n53168 = n34254 ^ n31673 ^ n12215 ;
  assign n53173 = n53172 ^ n53168 ^ n1980 ;
  assign n53174 = ( n8566 & n38049 ) | ( n8566 & ~n52910 ) | ( n38049 & ~n52910 ) ;
  assign n53175 = n11143 & n11689 ;
  assign n53176 = n53175 ^ n695 ^ 1'b0 ;
  assign n53177 = n53176 ^ n16435 ^ 1'b0 ;
  assign n53178 = n2231 & n53177 ;
  assign n53179 = n53174 & n53178 ;
  assign n53181 = n24192 ^ n7995 ^ x13 ;
  assign n53180 = n5267 & ~n5316 ;
  assign n53182 = n53181 ^ n53180 ^ 1'b0 ;
  assign n53184 = ~n6073 & n10508 ;
  assign n53183 = n21932 & ~n47895 ;
  assign n53185 = n53184 ^ n53183 ^ n15492 ;
  assign n53186 = ~n3071 & n15426 ;
  assign n53187 = n53186 ^ n20484 ^ 1'b0 ;
  assign n53188 = n35603 ^ n26051 ^ n13785 ;
  assign n53189 = ( n11490 & n17608 ) | ( n11490 & n19308 ) | ( n17608 & n19308 ) ;
  assign n53190 = ( ~n33474 & n36876 ) | ( ~n33474 & n53189 ) | ( n36876 & n53189 ) ;
  assign n53191 = n26950 ^ n17929 ^ 1'b0 ;
  assign n53192 = n26437 ^ n11416 ^ 1'b0 ;
  assign n53193 = n51406 ^ n4085 ^ 1'b0 ;
  assign n53194 = n17180 ^ n14466 ^ 1'b0 ;
  assign n53195 = ~n8811 & n53194 ;
  assign n53196 = n9363 & n53195 ;
  assign n53197 = n30521 ^ n9573 ^ n5277 ;
  assign n53198 = ( n4946 & n53196 ) | ( n4946 & n53197 ) | ( n53196 & n53197 ) ;
  assign n53199 = n53198 ^ n51611 ^ 1'b0 ;
  assign n53200 = ( n8893 & ~n11826 ) | ( n8893 & n21492 ) | ( ~n11826 & n21492 ) ;
  assign n53201 = ~n5249 & n34662 ;
  assign n53202 = n38036 & n53201 ;
  assign n53203 = n35793 ^ n28616 ^ n1042 ;
  assign n53204 = n32703 ^ n24661 ^ n4163 ;
  assign n53205 = n53204 ^ n34275 ^ n12223 ;
  assign n53206 = ( ~n8657 & n11140 ) | ( ~n8657 & n46624 ) | ( n11140 & n46624 ) ;
  assign n53207 = n53206 ^ n46915 ^ n4034 ;
  assign n53208 = ( n3788 & ~n8007 ) | ( n3788 & n18093 ) | ( ~n8007 & n18093 ) ;
  assign n53209 = ( n3153 & n17204 ) | ( n3153 & ~n53208 ) | ( n17204 & ~n53208 ) ;
  assign n53210 = n20349 & ~n45805 ;
  assign n53211 = ( x107 & ~n50942 ) | ( x107 & n53210 ) | ( ~n50942 & n53210 ) ;
  assign n53213 = ( ~n265 & n11582 ) | ( ~n265 & n22063 ) | ( n11582 & n22063 ) ;
  assign n53212 = n7655 ^ n5584 ^ n2525 ;
  assign n53214 = n53213 ^ n53212 ^ n43003 ;
  assign n53218 = n37940 ^ n1873 ^ 1'b0 ;
  assign n53219 = n1387 & ~n53218 ;
  assign n53220 = ( n34022 & n42095 ) | ( n34022 & ~n53219 ) | ( n42095 & ~n53219 ) ;
  assign n53215 = n46591 ^ n9109 ^ 1'b0 ;
  assign n53216 = n1968 & ~n53215 ;
  assign n53217 = n40151 & n53216 ;
  assign n53221 = n53220 ^ n53217 ^ n40829 ;
  assign n53222 = ( n8101 & n23012 ) | ( n8101 & n50439 ) | ( n23012 & n50439 ) ;
  assign n53223 = n3543 ^ n708 ^ x78 ;
  assign n53224 = ( n10167 & n31439 ) | ( n10167 & n48388 ) | ( n31439 & n48388 ) ;
  assign n53225 = n53224 ^ n25489 ^ 1'b0 ;
  assign n53226 = n53223 & n53225 ;
  assign n53227 = ( n1112 & n39346 ) | ( n1112 & ~n44093 ) | ( n39346 & ~n44093 ) ;
  assign n53228 = n1859 & n39701 ;
  assign n53229 = ~n53227 & n53228 ;
  assign n53230 = ( n18490 & ~n34503 ) | ( n18490 & n36705 ) | ( ~n34503 & n36705 ) ;
  assign n53231 = n30649 ^ n12980 ^ 1'b0 ;
  assign n53232 = ( n15758 & n38815 ) | ( n15758 & ~n53231 ) | ( n38815 & ~n53231 ) ;
  assign n53233 = ( ~n23737 & n46568 ) | ( ~n23737 & n53232 ) | ( n46568 & n53232 ) ;
  assign n53235 = n14854 & n22340 ;
  assign n53234 = ( n8414 & n38787 ) | ( n8414 & n45667 ) | ( n38787 & n45667 ) ;
  assign n53236 = n53235 ^ n53234 ^ n2730 ;
  assign n53237 = n53236 ^ n17156 ^ n6933 ;
  assign n53238 = n28648 ^ n19813 ^ n2100 ;
  assign n53239 = ( ~n6815 & n8283 ) | ( ~n6815 & n53238 ) | ( n8283 & n53238 ) ;
  assign n53240 = n40090 ^ n39429 ^ n38316 ;
  assign n53241 = ~n20822 & n21973 ;
  assign n53242 = ( n24349 & n53240 ) | ( n24349 & n53241 ) | ( n53240 & n53241 ) ;
  assign n53249 = n16845 ^ n14426 ^ n14349 ;
  assign n53246 = n28961 | n36335 ;
  assign n53247 = n2064 & ~n53246 ;
  assign n53248 = n53247 ^ n20199 ^ n9623 ;
  assign n53243 = n17424 ^ n11424 ^ n2599 ;
  assign n53244 = n22468 ^ n16041 ^ 1'b0 ;
  assign n53245 = ~n53243 & n53244 ;
  assign n53250 = n53249 ^ n53248 ^ n53245 ;
  assign n53251 = ( n11008 & n18650 ) | ( n11008 & ~n22865 ) | ( n18650 & ~n22865 ) ;
  assign n53254 = n18656 ^ n8239 ^ 1'b0 ;
  assign n53255 = ~n2914 & n53254 ;
  assign n53256 = ( x254 & n25845 ) | ( x254 & n53255 ) | ( n25845 & n53255 ) ;
  assign n53253 = n19087 ^ n7538 ^ n5664 ;
  assign n53257 = n53256 ^ n53253 ^ n43819 ;
  assign n53258 = n53257 ^ n7920 ^ 1'b0 ;
  assign n53259 = ~n42454 & n53258 ;
  assign n53252 = n15216 & n23749 ;
  assign n53260 = n53259 ^ n53252 ^ 1'b0 ;
  assign n53261 = n19190 ^ n4662 ^ 1'b0 ;
  assign n53262 = n53261 ^ n47778 ^ n16102 ;
  assign n53263 = n53262 ^ n49533 ^ n29670 ;
  assign n53264 = n37174 ^ n16058 ^ n5872 ;
  assign n53265 = n53264 ^ n36046 ^ n5441 ;
  assign n53266 = ( n3843 & ~n20359 ) | ( n3843 & n36384 ) | ( ~n20359 & n36384 ) ;
  assign n53269 = n13394 ^ n7177 ^ n4861 ;
  assign n53267 = n10831 & ~n13259 ;
  assign n53268 = n22589 | n53267 ;
  assign n53270 = n53269 ^ n53268 ^ n18025 ;
  assign n53271 = n53269 ^ n41539 ^ n19062 ;
  assign n53272 = n53271 ^ n41986 ^ n8487 ;
  assign n53273 = n7442 & ~n53272 ;
  assign n53274 = n26405 ^ n15454 ^ n3870 ;
  assign n53275 = n14339 & ~n20514 ;
  assign n53276 = ~n35394 & n53275 ;
  assign n53277 = ~n39487 & n53276 ;
  assign n53278 = n5373 | n7248 ;
  assign n53279 = n53278 ^ n23682 ^ 1'b0 ;
  assign n53280 = n53279 ^ n45329 ^ n19271 ;
  assign n53281 = ( n9020 & n26833 ) | ( n9020 & ~n53280 ) | ( n26833 & ~n53280 ) ;
  assign n53286 = n34386 ^ n22876 ^ n10522 ;
  assign n53287 = n53286 ^ n29997 ^ 1'b0 ;
  assign n53283 = ( n272 & n9976 ) | ( n272 & ~n33882 ) | ( n9976 & ~n33882 ) ;
  assign n53284 = ( n23705 & ~n52686 ) | ( n23705 & n53283 ) | ( ~n52686 & n53283 ) ;
  assign n53282 = n16283 ^ n13973 ^ n2187 ;
  assign n53285 = n53284 ^ n53282 ^ n23013 ;
  assign n53288 = n53287 ^ n53285 ^ n24063 ;
  assign n53289 = n2559 | n6034 ;
  assign n53290 = n26877 | n53289 ;
  assign n53291 = n23992 ^ n8124 ^ n7548 ;
  assign n53292 = ( n30039 & n53290 ) | ( n30039 & n53291 ) | ( n53290 & n53291 ) ;
  assign n53293 = n14858 & ~n51787 ;
  assign n53294 = ~n32027 & n53293 ;
  assign n53295 = n53294 ^ n36178 ^ 1'b0 ;
  assign n53296 = n19143 ^ n13335 ^ n445 ;
  assign n53297 = ( n31339 & n31637 ) | ( n31339 & ~n45571 ) | ( n31637 & ~n45571 ) ;
  assign n53298 = ( n28951 & n34413 ) | ( n28951 & n51445 ) | ( n34413 & n51445 ) ;
  assign n53299 = n10018 | n53298 ;
  assign n53300 = n33422 ^ n13022 ^ n1412 ;
  assign n53301 = ( n2766 & n26533 ) | ( n2766 & n53300 ) | ( n26533 & n53300 ) ;
  assign n53302 = n34869 & ~n44716 ;
  assign n53303 = ~n53301 & n53302 ;
  assign n53304 = n28130 ^ n4716 ^ 1'b0 ;
  assign n53305 = ( ~n8825 & n34940 ) | ( ~n8825 & n53304 ) | ( n34940 & n53304 ) ;
  assign n53306 = n23364 ^ n4712 ^ x66 ;
  assign n53307 = n34654 | n53306 ;
  assign n53308 = n19883 ^ n7299 ^ n543 ;
  assign n53309 = n36150 ^ n13136 ^ 1'b0 ;
  assign n53310 = n5969 & n21446 ;
  assign n53314 = n32150 ^ n5287 ^ n1463 ;
  assign n53311 = ~n1271 & n51830 ;
  assign n53312 = n53311 ^ n17045 ^ 1'b0 ;
  assign n53313 = ( n10881 & ~n48244 ) | ( n10881 & n53312 ) | ( ~n48244 & n53312 ) ;
  assign n53315 = n53314 ^ n53313 ^ n542 ;
  assign n53316 = n23371 ^ n21319 ^ n5394 ;
  assign n53317 = n49214 ^ n7334 ^ 1'b0 ;
  assign n53318 = n32545 | n53317 ;
  assign n53319 = n9444 | n11463 ;
  assign n53320 = n3461 | n53319 ;
  assign n53321 = n47217 ^ n11872 ^ 1'b0 ;
  assign n53322 = n24391 & n53321 ;
  assign n53323 = n32366 ^ n5730 ^ 1'b0 ;
  assign n53324 = ( n28220 & n28631 ) | ( n28220 & ~n53323 ) | ( n28631 & ~n53323 ) ;
  assign n53325 = n22391 ^ n14150 ^ n9739 ;
  assign n53326 = ( n3528 & n45781 ) | ( n3528 & ~n53325 ) | ( n45781 & ~n53325 ) ;
  assign n53327 = ( n10043 & ~n28871 ) | ( n10043 & n49098 ) | ( ~n28871 & n49098 ) ;
  assign n53328 = ( n19855 & n30392 ) | ( n19855 & n32946 ) | ( n30392 & n32946 ) ;
  assign n53329 = ( n10421 & n29675 ) | ( n10421 & ~n33292 ) | ( n29675 & ~n33292 ) ;
  assign n53330 = n4762 & n41505 ;
  assign n53331 = n53330 ^ n41766 ^ n19800 ;
  assign n53332 = n5658 & ~n22156 ;
  assign n53333 = n53332 ^ n25603 ^ 1'b0 ;
  assign n53334 = ( ~n12180 & n19241 ) | ( ~n12180 & n53333 ) | ( n19241 & n53333 ) ;
  assign n53335 = ( n2396 & n36408 ) | ( n2396 & n53334 ) | ( n36408 & n53334 ) ;
  assign n53336 = ( ~n22874 & n28233 ) | ( ~n22874 & n53335 ) | ( n28233 & n53335 ) ;
  assign n53337 = n30525 & ~n46310 ;
  assign n53338 = n18391 ^ n12147 ^ n9606 ;
  assign n53339 = n53338 ^ n20272 ^ n3675 ;
  assign n53340 = n28540 ^ n15724 ^ n3857 ;
  assign n53341 = n53340 ^ n37100 ^ 1'b0 ;
  assign n53342 = ( n21611 & n52406 ) | ( n21611 & n53341 ) | ( n52406 & n53341 ) ;
  assign n53343 = n53342 ^ n21310 ^ 1'b0 ;
  assign n53344 = n53339 & n53343 ;
  assign n53345 = n14590 & n27833 ;
  assign n53346 = n53345 ^ n50092 ^ 1'b0 ;
  assign n53347 = ( n7002 & ~n18039 ) | ( n7002 & n27687 ) | ( ~n18039 & n27687 ) ;
  assign n53348 = n53347 ^ n39555 ^ n2839 ;
  assign n53349 = n53348 ^ n43244 ^ n16330 ;
  assign n53350 = n10113 | n23663 ;
  assign n53351 = n39465 ^ n28885 ^ n12369 ;
  assign n53352 = n53351 ^ n16997 ^ n1459 ;
  assign n53354 = n25493 ^ n5898 ^ 1'b0 ;
  assign n53355 = n7364 & n53354 ;
  assign n53353 = n16519 & ~n16865 ;
  assign n53356 = n53355 ^ n53353 ^ 1'b0 ;
  assign n53357 = n53356 ^ n52947 ^ n48861 ;
  assign n53358 = n19454 ^ n4570 ^ 1'b0 ;
  assign n53359 = n11229 ^ n9825 ^ n287 ;
  assign n53360 = ( n5988 & ~n29510 ) | ( n5988 & n36312 ) | ( ~n29510 & n36312 ) ;
  assign n53361 = n53359 & ~n53360 ;
  assign n53362 = ( n10955 & ~n18621 ) | ( n10955 & n33541 ) | ( ~n18621 & n33541 ) ;
  assign n53363 = n7094 & n20907 ;
  assign n53364 = n53363 ^ n35852 ^ n29838 ;
  assign n53365 = n53364 ^ n12084 ^ 1'b0 ;
  assign n53366 = n32196 ^ n19099 ^ 1'b0 ;
  assign n53367 = n33538 | n53366 ;
  assign n53369 = ~n12858 & n15875 ;
  assign n53370 = ( n28406 & ~n42645 ) | ( n28406 & n53369 ) | ( ~n42645 & n53369 ) ;
  assign n53368 = n31556 & ~n53078 ;
  assign n53371 = n53370 ^ n53368 ^ 1'b0 ;
  assign n53372 = n49759 ^ n16905 ^ 1'b0 ;
  assign n53373 = n28489 & n53372 ;
  assign n53374 = n1984 & n19798 ;
  assign n53375 = n23244 & n53374 ;
  assign n53376 = n41257 | n53375 ;
  assign n53377 = n53376 ^ n38008 ^ 1'b0 ;
  assign n53378 = ( n3670 & n16990 ) | ( n3670 & n53377 ) | ( n16990 & n53377 ) ;
  assign n53379 = n53378 ^ n31441 ^ n17903 ;
  assign n53380 = ( ~n8188 & n16715 ) | ( ~n8188 & n35787 ) | ( n16715 & n35787 ) ;
  assign n53381 = n39167 ^ n18859 ^ n8216 ;
  assign n53382 = n53381 ^ n51557 ^ n16017 ;
  assign n53383 = n53382 ^ n32295 ^ 1'b0 ;
  assign n53384 = n27922 ^ n13165 ^ 1'b0 ;
  assign n53385 = n7596 & n53384 ;
  assign n53386 = ( n24439 & n32186 ) | ( n24439 & ~n53385 ) | ( n32186 & ~n53385 ) ;
  assign n53387 = n52072 ^ n37336 ^ n8031 ;
  assign n53388 = ( n5143 & n15776 ) | ( n5143 & n26173 ) | ( n15776 & n26173 ) ;
  assign n53389 = n53388 ^ n47955 ^ n12439 ;
  assign n53390 = n53389 ^ n33332 ^ n18648 ;
  assign n53393 = n46107 ^ n1325 ^ n1211 ;
  assign n53394 = n53393 ^ n24733 ^ n13531 ;
  assign n53395 = ( n27573 & ~n51312 ) | ( n27573 & n53394 ) | ( ~n51312 & n53394 ) ;
  assign n53391 = n14822 ^ n10068 ^ n6335 ;
  assign n53392 = ( n17063 & ~n28687 ) | ( n17063 & n53391 ) | ( ~n28687 & n53391 ) ;
  assign n53396 = n53395 ^ n53392 ^ n9100 ;
  assign n53397 = ( ~x98 & n26291 ) | ( ~x98 & n31470 ) | ( n26291 & n31470 ) ;
  assign n53398 = ~n916 & n2912 ;
  assign n53399 = n53398 ^ n7410 ^ 1'b0 ;
  assign n53400 = n53399 ^ n19613 ^ n9174 ;
  assign n53401 = ~n4668 & n53400 ;
  assign n53402 = n53397 & n53401 ;
  assign n53403 = ( n2315 & ~n9368 ) | ( n2315 & n40019 ) | ( ~n9368 & n40019 ) ;
  assign n53404 = n32714 | n51242 ;
  assign n53405 = n53404 ^ n34917 ^ 1'b0 ;
  assign n53406 = n53403 & ~n53405 ;
  assign n53407 = n53406 ^ n17387 ^ 1'b0 ;
  assign n53409 = ~n2376 & n5833 ;
  assign n53410 = n14985 & n53409 ;
  assign n53408 = ~n15832 & n27116 ;
  assign n53411 = n53410 ^ n53408 ^ n8489 ;
  assign n53413 = n11862 ^ n10887 ^ 1'b0 ;
  assign n53414 = n22382 & n53413 ;
  assign n53412 = n48083 ^ n17769 ^ x151 ;
  assign n53415 = n53414 ^ n53412 ^ n20178 ;
  assign n53416 = ( n12422 & ~n18777 ) | ( n12422 & n29855 ) | ( ~n18777 & n29855 ) ;
  assign n53417 = n53416 ^ n51346 ^ n16811 ;
  assign n53421 = n19382 ^ n8920 ^ 1'b0 ;
  assign n53418 = n28117 ^ n9517 ^ 1'b0 ;
  assign n53419 = ( ~n26549 & n45155 ) | ( ~n26549 & n53418 ) | ( n45155 & n53418 ) ;
  assign n53420 = n53419 ^ n22986 ^ n20090 ;
  assign n53422 = n53421 ^ n53420 ^ n10835 ;
  assign n53424 = n17963 ^ n11747 ^ n7819 ;
  assign n53423 = n46508 ^ n25685 ^ n3144 ;
  assign n53425 = n53424 ^ n53423 ^ n14787 ;
  assign n53426 = ( ~n9226 & n19407 ) | ( ~n9226 & n34206 ) | ( n19407 & n34206 ) ;
  assign n53427 = n34208 ^ n6824 ^ 1'b0 ;
  assign n53428 = ( n29148 & n53426 ) | ( n29148 & ~n53427 ) | ( n53426 & ~n53427 ) ;
  assign n53429 = n53428 ^ n25069 ^ n12704 ;
  assign n53430 = ( n8237 & n30445 ) | ( n8237 & n53429 ) | ( n30445 & n53429 ) ;
  assign n53431 = n7549 ^ n6044 ^ n317 ;
  assign n53432 = n21728 & ~n36228 ;
  assign n53433 = n39824 & n53432 ;
  assign n53434 = n53433 ^ n13948 ^ n6512 ;
  assign n53435 = ( n12243 & n53431 ) | ( n12243 & n53434 ) | ( n53431 & n53434 ) ;
  assign n53436 = n3860 & n4632 ;
  assign n53437 = n7175 & n53436 ;
  assign n53438 = n53437 ^ n4062 ^ 1'b0 ;
  assign n53439 = ( ~n14212 & n27731 ) | ( ~n14212 & n47916 ) | ( n27731 & n47916 ) ;
  assign n53440 = n1233 & n19590 ;
  assign n53441 = ~n53439 & n53440 ;
  assign n53442 = n43842 ^ n15052 ^ x240 ;
  assign n53443 = ( n3284 & ~n12649 ) | ( n3284 & n36996 ) | ( ~n12649 & n36996 ) ;
  assign n53444 = ( ~n18342 & n37489 ) | ( ~n18342 & n44471 ) | ( n37489 & n44471 ) ;
  assign n53445 = n53444 ^ n33798 ^ n14356 ;
  assign n53446 = n53445 ^ n41137 ^ n4503 ;
  assign n53447 = n27912 ^ n13072 ^ n6184 ;
  assign n53448 = ( ~n18955 & n39915 ) | ( ~n18955 & n53447 ) | ( n39915 & n53447 ) ;
  assign n53449 = ( n21226 & n32297 ) | ( n21226 & n37444 ) | ( n32297 & n37444 ) ;
  assign n53450 = n15498 ^ n8792 ^ n4697 ;
  assign n53451 = n12854 | n21533 ;
  assign n53452 = n29401 ^ n28199 ^ n11731 ;
  assign n53453 = n53452 ^ n23774 ^ n17578 ;
  assign n53454 = ~n8707 & n53453 ;
  assign n53455 = ~n4565 & n53454 ;
  assign n53456 = n5384 & ~n23658 ;
  assign n53457 = ~n25750 & n53456 ;
  assign n53458 = ( ~n18661 & n35644 ) | ( ~n18661 & n47461 ) | ( n35644 & n47461 ) ;
  assign n53460 = n33723 ^ n1204 ^ 1'b0 ;
  assign n53459 = ( ~n4122 & n6658 ) | ( ~n4122 & n44455 ) | ( n6658 & n44455 ) ;
  assign n53461 = n53460 ^ n53459 ^ n4165 ;
  assign n53462 = ( n7209 & n9938 ) | ( n7209 & ~n13809 ) | ( n9938 & ~n13809 ) ;
  assign n53463 = n16502 ^ n8337 ^ 1'b0 ;
  assign n53464 = ( n17891 & n25073 ) | ( n17891 & ~n53463 ) | ( n25073 & ~n53463 ) ;
  assign n53465 = ( n20205 & n53462 ) | ( n20205 & n53464 ) | ( n53462 & n53464 ) ;
  assign n53466 = n4894 & n51700 ;
  assign n53467 = n53466 ^ n34371 ^ n28498 ;
  assign n53468 = ~n15898 & n35132 ;
  assign n53469 = ( ~n20244 & n38974 ) | ( ~n20244 & n53468 ) | ( n38974 & n53468 ) ;
  assign n53470 = n18631 ^ n16380 ^ n1282 ;
  assign n53471 = n53470 ^ n53290 ^ n18510 ;
  assign n53472 = n53471 ^ n27655 ^ n11111 ;
  assign n53473 = n38918 ^ n37808 ^ n31699 ;
  assign n53474 = ( n8237 & n9297 ) | ( n8237 & n12595 ) | ( n9297 & n12595 ) ;
  assign n53475 = n53474 ^ n38097 ^ 1'b0 ;
  assign n53476 = n53475 ^ n47813 ^ 1'b0 ;
  assign n53477 = n53227 ^ n42817 ^ 1'b0 ;
  assign n53478 = n45541 | n53477 ;
  assign n53479 = ( n4509 & n5142 ) | ( n4509 & n16220 ) | ( n5142 & n16220 ) ;
  assign n53480 = n53479 ^ n49010 ^ n14473 ;
  assign n53481 = n42967 ^ n40113 ^ n8016 ;
  assign n53482 = ( n33073 & n36939 ) | ( n33073 & n37298 ) | ( n36939 & n37298 ) ;
  assign n53483 = ( ~n4508 & n9510 ) | ( ~n4508 & n53482 ) | ( n9510 & n53482 ) ;
  assign n53484 = n38917 ^ n29884 ^ n26782 ;
  assign n53485 = n25861 ^ n25472 ^ n19828 ;
  assign n53486 = n43991 & ~n53485 ;
  assign n53487 = ~n6980 & n9214 ;
  assign n53488 = n7887 & n53487 ;
  assign n53489 = n1094 & ~n53488 ;
  assign n53490 = ( ~n30574 & n33284 ) | ( ~n30574 & n45477 ) | ( n33284 & n45477 ) ;
  assign n53491 = ( ~n11743 & n28445 ) | ( ~n11743 & n53490 ) | ( n28445 & n53490 ) ;
  assign n53492 = ( n432 & ~n53489 ) | ( n432 & n53491 ) | ( ~n53489 & n53491 ) ;
  assign n53493 = n21612 & ~n27077 ;
  assign n53494 = n53493 ^ n39494 ^ 1'b0 ;
  assign n53495 = n53494 ^ n32093 ^ n18292 ;
  assign n53496 = n9711 ^ n5625 ^ n4384 ;
  assign n53497 = ~n27867 & n30244 ;
  assign n53498 = n16998 ^ n7269 ^ 1'b0 ;
  assign n53499 = ( ~n928 & n13647 ) | ( ~n928 & n36405 ) | ( n13647 & n36405 ) ;
  assign n53500 = ( ~n8541 & n14785 ) | ( ~n8541 & n15465 ) | ( n14785 & n15465 ) ;
  assign n53501 = n53500 ^ n17193 ^ n5855 ;
  assign n53502 = n53501 ^ n3576 ^ n1961 ;
  assign n53503 = n8150 | n45773 ;
  assign n53504 = ( n15269 & ~n22369 ) | ( n15269 & n53503 ) | ( ~n22369 & n53503 ) ;
  assign n53505 = n7816 | n43518 ;
  assign n53506 = n36402 ^ n27310 ^ n13280 ;
  assign n53507 = n22770 ^ n7794 ^ n5912 ;
  assign n53508 = ~n25849 & n34922 ;
  assign n53509 = n53508 ^ n35207 ^ 1'b0 ;
  assign n53510 = ~n2226 & n29859 ;
  assign n53511 = n53510 ^ n1556 ^ 1'b0 ;
  assign n53512 = n1462 & ~n15752 ;
  assign n53513 = n53512 ^ n26613 ^ 1'b0 ;
  assign n53514 = ( n20348 & ~n29204 ) | ( n20348 & n33200 ) | ( ~n29204 & n33200 ) ;
  assign n53515 = n14714 ^ n12551 ^ n1609 ;
  assign n53516 = ( n4364 & ~n32755 ) | ( n4364 & n53515 ) | ( ~n32755 & n53515 ) ;
  assign n53517 = ( ~n15178 & n43334 ) | ( ~n15178 & n53516 ) | ( n43334 & n53516 ) ;
  assign n53518 = n11508 & ~n17329 ;
  assign n53519 = ( ~n10510 & n26512 ) | ( ~n10510 & n53518 ) | ( n26512 & n53518 ) ;
  assign n53520 = ( n4699 & n34885 ) | ( n4699 & n53519 ) | ( n34885 & n53519 ) ;
  assign n53521 = ( n19338 & n33889 ) | ( n19338 & n53520 ) | ( n33889 & n53520 ) ;
  assign n53522 = ( n7693 & n14433 ) | ( n7693 & ~n48300 ) | ( n14433 & ~n48300 ) ;
  assign n53523 = n47029 ^ n24959 ^ n4074 ;
  assign n53524 = n46090 ^ n16338 ^ n9000 ;
  assign n53525 = n53524 ^ n29066 ^ n23762 ;
  assign n53526 = ( n15953 & n16651 ) | ( n15953 & n50904 ) | ( n16651 & n50904 ) ;
  assign n53527 = n53526 ^ n44731 ^ n18420 ;
  assign n53528 = n19691 ^ n10925 ^ n9836 ;
  assign n53529 = ( n36738 & n47953 ) | ( n36738 & ~n53528 ) | ( n47953 & ~n53528 ) ;
  assign n53530 = n6022 ^ n4281 ^ 1'b0 ;
  assign n53531 = n53530 ^ n18884 ^ 1'b0 ;
  assign n53532 = n28622 ^ n26544 ^ n8157 ;
  assign n53533 = n40065 & n53532 ;
  assign n53534 = n40328 ^ n12881 ^ n1249 ;
  assign n53535 = ( n47774 & n49442 ) | ( n47774 & ~n51405 ) | ( n49442 & ~n51405 ) ;
  assign n53536 = ( n7934 & n25041 ) | ( n7934 & ~n37326 ) | ( n25041 & ~n37326 ) ;
  assign n53537 = n40036 ^ n29758 ^ n13670 ;
  assign n53538 = n53537 ^ n4209 ^ 1'b0 ;
  assign n53539 = n53538 ^ n52015 ^ n37986 ;
  assign n53540 = ( n26149 & n53536 ) | ( n26149 & n53539 ) | ( n53536 & n53539 ) ;
  assign n53541 = n48901 ^ n26873 ^ n18231 ;
  assign n53542 = n6539 & ~n41706 ;
  assign n53543 = n24214 & ~n30561 ;
  assign n53546 = n1649 | n17122 ;
  assign n53547 = n53546 ^ n13664 ^ n8977 ;
  assign n53544 = n49938 ^ n14520 ^ n11421 ;
  assign n53545 = ( n2979 & ~n36870 ) | ( n2979 & n53544 ) | ( ~n36870 & n53544 ) ;
  assign n53548 = n53547 ^ n53545 ^ n53138 ;
  assign n53549 = ~n13099 & n20432 ;
  assign n53550 = n53549 ^ n45036 ^ 1'b0 ;
  assign n53551 = ( n10879 & n18302 ) | ( n10879 & ~n42269 ) | ( n18302 & ~n42269 ) ;
  assign n53552 = n50183 ^ n47953 ^ n707 ;
  assign n53553 = n4965 ^ x165 ^ 1'b0 ;
  assign n53554 = n46816 ^ n3376 ^ n517 ;
  assign n53555 = n7268 & ~n53554 ;
  assign n53558 = n23660 ^ n5927 ^ 1'b0 ;
  assign n53556 = n31141 ^ n19347 ^ 1'b0 ;
  assign n53557 = ~n16451 & n53556 ;
  assign n53559 = n53558 ^ n53557 ^ n35452 ;
  assign n53560 = ( n9743 & n12356 ) | ( n9743 & n28368 ) | ( n12356 & n28368 ) ;
  assign n53563 = n33078 ^ n12337 ^ n1509 ;
  assign n53561 = n41016 ^ n38341 ^ n7373 ;
  assign n53562 = n53561 ^ n12988 ^ n2743 ;
  assign n53564 = n53563 ^ n53562 ^ n28478 ;
  assign n53565 = n33478 ^ n28113 ^ 1'b0 ;
  assign n53566 = ( n6138 & n10977 ) | ( n6138 & ~n34260 ) | ( n10977 & ~n34260 ) ;
  assign n53567 = ( n2710 & ~n53565 ) | ( n2710 & n53566 ) | ( ~n53565 & n53566 ) ;
  assign n53568 = n33978 ^ n23555 ^ n2916 ;
  assign n53569 = n1303 & n45253 ;
  assign n53570 = ~n53568 & n53569 ;
  assign n53571 = n35377 ^ n34948 ^ 1'b0 ;
  assign n53572 = n34678 & n53571 ;
  assign n53573 = ( ~n38744 & n43239 ) | ( ~n38744 & n53395 ) | ( n43239 & n53395 ) ;
  assign n53574 = ( n1626 & n12476 ) | ( n1626 & n28410 ) | ( n12476 & n28410 ) ;
  assign n53580 = n3163 & n7191 ;
  assign n53581 = ~n6493 & n53580 ;
  assign n53577 = ( ~n2159 & n3223 ) | ( ~n2159 & n7567 ) | ( n3223 & n7567 ) ;
  assign n53576 = ( n3004 & ~n13413 ) | ( n3004 & n21334 ) | ( ~n13413 & n21334 ) ;
  assign n53575 = n45675 ^ n30705 ^ n4319 ;
  assign n53578 = n53577 ^ n53576 ^ n53575 ;
  assign n53579 = n53578 ^ n5381 ^ 1'b0 ;
  assign n53582 = n53581 ^ n53579 ^ n3185 ;
  assign n53583 = n53582 ^ n26318 ^ n17270 ;
  assign n53584 = n53583 ^ n36702 ^ n17692 ;
  assign n53585 = ( n7165 & n25472 ) | ( n7165 & n32958 ) | ( n25472 & n32958 ) ;
  assign n53586 = n36909 ^ n16642 ^ n2100 ;
  assign n53587 = n5577 | n13930 ;
  assign n53588 = n38707 & n53587 ;
  assign n53589 = n30000 ^ n27681 ^ 1'b0 ;
  assign n53590 = ~n15256 & n23519 ;
  assign n53591 = ( n15274 & ~n28009 ) | ( n15274 & n53590 ) | ( ~n28009 & n53590 ) ;
  assign n53592 = n53591 ^ n3264 ^ 1'b0 ;
  assign n53593 = n35257 | n53592 ;
  assign n53594 = n32751 | n33459 ;
  assign n53595 = n53594 ^ n31173 ^ 1'b0 ;
  assign n53596 = ( n20688 & n36257 ) | ( n20688 & ~n37885 ) | ( n36257 & ~n37885 ) ;
  assign n53597 = n51299 ^ n18095 ^ 1'b0 ;
  assign n53598 = n6425 | n53597 ;
  assign n53599 = ( ~x238 & n31021 ) | ( ~x238 & n53598 ) | ( n31021 & n53598 ) ;
  assign n53600 = ( n19449 & n21139 ) | ( n19449 & n22307 ) | ( n21139 & n22307 ) ;
  assign n53601 = ( n9235 & n9691 ) | ( n9235 & n42296 ) | ( n9691 & n42296 ) ;
  assign n53602 = n50220 ^ n30221 ^ n662 ;
  assign n53603 = n44526 ^ n9432 ^ 1'b0 ;
  assign n53604 = n47791 ^ n19887 ^ n14254 ;
  assign n53605 = n4832 | n27983 ;
  assign n53606 = n53605 ^ n6622 ^ 1'b0 ;
  assign n53607 = ~n10278 & n53606 ;
  assign n53608 = n50448 & n53607 ;
  assign n53609 = ( n9273 & n53604 ) | ( n9273 & ~n53608 ) | ( n53604 & ~n53608 ) ;
  assign n53611 = n31619 ^ n20664 ^ n6699 ;
  assign n53612 = n53611 ^ n16785 ^ n10325 ;
  assign n53610 = ( ~n7244 & n27233 ) | ( ~n7244 & n32033 ) | ( n27233 & n32033 ) ;
  assign n53613 = n53612 ^ n53610 ^ n9825 ;
  assign n53614 = n32399 ^ x180 ^ 1'b0 ;
  assign n53615 = n47716 & n53614 ;
  assign n53622 = ~n11172 & n14590 ;
  assign n53616 = ~n7676 & n25577 ;
  assign n53617 = ~n13489 & n53616 ;
  assign n53618 = ( n5483 & n15390 ) | ( n5483 & ~n19652 ) | ( n15390 & ~n19652 ) ;
  assign n53619 = ( n45876 & n53617 ) | ( n45876 & n53618 ) | ( n53617 & n53618 ) ;
  assign n53620 = n51902 | n53619 ;
  assign n53621 = n53620 ^ n30658 ^ 1'b0 ;
  assign n53623 = n53622 ^ n53621 ^ n12501 ;
  assign n53624 = n53623 ^ n13258 ^ 1'b0 ;
  assign n53625 = n42773 ^ n15742 ^ n4653 ;
  assign n53626 = n981 & ~n37129 ;
  assign n53627 = n39789 | n48673 ;
  assign n53628 = n1248 & ~n53627 ;
  assign n53629 = n22234 | n53628 ;
  assign n53630 = n4496 & ~n53629 ;
  assign n53631 = ( ~n5691 & n30380 ) | ( ~n5691 & n39012 ) | ( n30380 & n39012 ) ;
  assign n53632 = n53631 ^ n42960 ^ 1'b0 ;
  assign n53633 = ~n53630 & n53632 ;
  assign n53634 = ~n23492 & n53633 ;
  assign n53635 = n3973 | n10471 ;
  assign n53636 = n53635 ^ n8787 ^ 1'b0 ;
  assign n53637 = ( n21439 & ~n31919 ) | ( n21439 & n53636 ) | ( ~n31919 & n53636 ) ;
  assign n53638 = ( n14586 & n26183 ) | ( n14586 & n40471 ) | ( n26183 & n40471 ) ;
  assign n53639 = ( n22202 & n45061 ) | ( n22202 & n53638 ) | ( n45061 & n53638 ) ;
  assign n53640 = n53227 ^ n26451 ^ n13905 ;
  assign n53641 = ( n50696 & ~n53639 ) | ( n50696 & n53640 ) | ( ~n53639 & n53640 ) ;
  assign n53644 = ( n2190 & n4161 ) | ( n2190 & ~n11766 ) | ( n4161 & ~n11766 ) ;
  assign n53642 = ( x235 & n2080 ) | ( x235 & n13384 ) | ( n2080 & n13384 ) ;
  assign n53643 = n53642 ^ n51955 ^ n659 ;
  assign n53645 = n53644 ^ n53643 ^ n34566 ;
  assign n53646 = n41181 ^ n40897 ^ n25287 ;
  assign n53647 = ( ~n11772 & n47200 ) | ( ~n11772 & n53646 ) | ( n47200 & n53646 ) ;
  assign n53648 = n16684 ^ n13541 ^ 1'b0 ;
  assign n53649 = n16100 | n32323 ;
  assign n53650 = n53649 ^ n35439 ^ 1'b0 ;
  assign n53651 = n21071 & ~n23905 ;
  assign n53652 = n30869 ^ n27989 ^ n7215 ;
  assign n53653 = n30071 ^ n7481 ^ 1'b0 ;
  assign n53654 = ( n29751 & ~n49057 ) | ( n29751 & n53653 ) | ( ~n49057 & n53653 ) ;
  assign n53655 = n6640 & ~n13532 ;
  assign n53656 = ~n3095 & n53655 ;
  assign n53657 = ( n2604 & n28388 ) | ( n2604 & n53656 ) | ( n28388 & n53656 ) ;
  assign n53658 = ( n18766 & n36145 ) | ( n18766 & n38906 ) | ( n36145 & n38906 ) ;
  assign n53659 = n10445 ^ n4544 ^ n2258 ;
  assign n53660 = ( n18685 & ~n35585 ) | ( n18685 & n53659 ) | ( ~n35585 & n53659 ) ;
  assign n53661 = n53660 ^ n24575 ^ n10902 ;
  assign n53662 = n53661 ^ n20269 ^ n10941 ;
  assign n53663 = n53662 ^ n48424 ^ n6129 ;
  assign n53664 = ( n6946 & ~n14908 ) | ( n6946 & n28932 ) | ( ~n14908 & n28932 ) ;
  assign n53665 = n16155 ^ n5399 ^ 1'b0 ;
  assign n53666 = n53475 ^ n18206 ^ 1'b0 ;
  assign n53667 = n26620 & ~n53666 ;
  assign n53668 = n6444 & ~n32556 ;
  assign n53669 = ( ~n286 & n11053 ) | ( ~n286 & n31261 ) | ( n11053 & n31261 ) ;
  assign n53670 = n32703 ^ n3097 ^ n1042 ;
  assign n53671 = n53670 ^ n25371 ^ n12438 ;
  assign n53672 = n52057 ^ n20810 ^ 1'b0 ;
  assign n53673 = ( n8852 & ~n8869 ) | ( n8852 & n20238 ) | ( ~n8869 & n20238 ) ;
  assign n53674 = ( n33682 & n37040 ) | ( n33682 & n53673 ) | ( n37040 & n53673 ) ;
  assign n53675 = n16153 ^ n9349 ^ n4671 ;
  assign n53676 = n53675 ^ n48600 ^ n40551 ;
  assign n53677 = n28031 ^ n17988 ^ n8401 ;
  assign n53678 = n6698 & n37521 ;
  assign n53679 = n53678 ^ n32134 ^ 1'b0 ;
  assign n53680 = ~n36001 & n53679 ;
  assign n53681 = ( n14111 & ~n39430 ) | ( n14111 & n53680 ) | ( ~n39430 & n53680 ) ;
  assign n53683 = n26784 ^ n20630 ^ n17614 ;
  assign n53684 = ( n44448 & n51868 ) | ( n44448 & ~n53683 ) | ( n51868 & ~n53683 ) ;
  assign n53682 = n7609 | n19082 ;
  assign n53685 = n53684 ^ n53682 ^ 1'b0 ;
  assign n53687 = n15844 ^ n11716 ^ 1'b0 ;
  assign n53688 = ( n11607 & n48995 ) | ( n11607 & ~n53687 ) | ( n48995 & ~n53687 ) ;
  assign n53686 = n4719 & n16066 ;
  assign n53689 = n53688 ^ n53686 ^ 1'b0 ;
  assign n53690 = ~n636 & n4286 ;
  assign n53691 = n27131 ^ n25232 ^ 1'b0 ;
  assign n53692 = ~n53690 & n53691 ;
  assign n53693 = n53692 ^ n4179 ^ 1'b0 ;
  assign n53694 = n2632 & ~n53693 ;
  assign n53695 = ( n15804 & ~n17463 ) | ( n15804 & n22884 ) | ( ~n17463 & n22884 ) ;
  assign n53696 = ( n31922 & ~n40683 ) | ( n31922 & n53695 ) | ( ~n40683 & n53695 ) ;
  assign n53697 = n35142 ^ n19671 ^ n10917 ;
  assign n53698 = n9979 & n13653 ;
  assign n53699 = ( n5966 & n23885 ) | ( n5966 & ~n41291 ) | ( n23885 & ~n41291 ) ;
  assign n53700 = ( n53697 & n53698 ) | ( n53697 & n53699 ) | ( n53698 & n53699 ) ;
  assign n53701 = ( n2801 & n53696 ) | ( n2801 & ~n53700 ) | ( n53696 & ~n53700 ) ;
  assign n53702 = n51371 ^ n22602 ^ 1'b0 ;
  assign n53703 = ~n19519 & n24711 ;
  assign n53704 = ( ~n31829 & n53702 ) | ( ~n31829 & n53703 ) | ( n53702 & n53703 ) ;
  assign n53705 = n33986 ^ n26557 ^ n15818 ;
  assign n53706 = n53705 ^ n39028 ^ n37824 ;
  assign n53707 = n10532 & ~n53706 ;
  assign n53708 = n49262 ^ n48538 ^ n14496 ;
  assign n53709 = ( n11302 & n49919 ) | ( n11302 & n53708 ) | ( n49919 & n53708 ) ;
  assign n53710 = ( n13812 & n26050 ) | ( n13812 & ~n31943 ) | ( n26050 & ~n31943 ) ;
  assign n53711 = n53710 ^ n37165 ^ n6940 ;
  assign n53712 = ( n28065 & n37737 ) | ( n28065 & ~n53711 ) | ( n37737 & ~n53711 ) ;
  assign n53713 = ~n16008 & n17087 ;
  assign n53714 = n53713 ^ n27359 ^ n8454 ;
  assign n53715 = ( n10059 & n12655 ) | ( n10059 & ~n14594 ) | ( n12655 & ~n14594 ) ;
  assign n53716 = n23095 ^ n2392 ^ n1174 ;
  assign n53717 = n53716 ^ n30650 ^ n16358 ;
  assign n53718 = ( n5272 & n53715 ) | ( n5272 & n53717 ) | ( n53715 & n53717 ) ;
  assign n53719 = n30277 ^ n7141 ^ n1302 ;
  assign n53720 = n10566 & n53719 ;
  assign n53721 = n53720 ^ n48213 ^ n19376 ;
  assign n53722 = n31279 & n45555 ;
  assign n53723 = ( ~n16429 & n18913 ) | ( ~n16429 & n53341 ) | ( n18913 & n53341 ) ;
  assign n53724 = n25297 ^ n12230 ^ n11872 ;
  assign n53725 = n39926 ^ n35866 ^ n23306 ;
  assign n53726 = ( n958 & n10189 ) | ( n958 & n14504 ) | ( n10189 & n14504 ) ;
  assign n53727 = ( n19484 & n44576 ) | ( n19484 & n53726 ) | ( n44576 & n53726 ) ;
  assign n53728 = ~n6835 & n31921 ;
  assign n53729 = n53728 ^ n52744 ^ n37662 ;
  assign n53730 = ( n6776 & n6993 ) | ( n6776 & n38535 ) | ( n6993 & n38535 ) ;
  assign n53731 = ~n8389 & n15354 ;
  assign n53732 = n53731 ^ n6569 ^ 1'b0 ;
  assign n53733 = n53732 ^ n46011 ^ n17406 ;
  assign n53734 = n10138 & n13629 ;
  assign n53735 = ( n2558 & ~n23758 ) | ( n2558 & n30005 ) | ( ~n23758 & n30005 ) ;
  assign n53736 = n53735 ^ n36880 ^ 1'b0 ;
  assign n53737 = n24496 & ~n53736 ;
  assign n53738 = n5297 & n22709 ;
  assign n53739 = n25650 & n53738 ;
  assign n53740 = ( n20033 & n29365 ) | ( n20033 & ~n39145 ) | ( n29365 & ~n39145 ) ;
  assign n53741 = n49622 ^ n7361 ^ n3494 ;
  assign n53742 = n28985 ^ n11155 ^ 1'b0 ;
  assign n53743 = ( n44382 & n53741 ) | ( n44382 & n53742 ) | ( n53741 & n53742 ) ;
  assign n53744 = ( n5255 & n25707 ) | ( n5255 & ~n30384 ) | ( n25707 & ~n30384 ) ;
  assign n53745 = n47318 ^ n44339 ^ n13337 ;
  assign n53746 = ( ~n346 & n11836 ) | ( ~n346 & n28054 ) | ( n11836 & n28054 ) ;
  assign n53747 = ( n13521 & ~n20940 ) | ( n13521 & n32158 ) | ( ~n20940 & n32158 ) ;
  assign n53748 = n53747 ^ n47931 ^ n6323 ;
  assign n53749 = n49098 ^ n15897 ^ n1122 ;
  assign n53750 = n2750 ^ n2072 ^ 1'b0 ;
  assign n53751 = ~n8367 & n33410 ;
  assign n53752 = ( ~n260 & n4563 ) | ( ~n260 & n13536 ) | ( n4563 & n13536 ) ;
  assign n53753 = ~n35027 & n53752 ;
  assign n53754 = ~n14924 & n53753 ;
  assign n53755 = n1110 & n12741 ;
  assign n53756 = n695 & n14379 ;
  assign n53757 = ~n53755 & n53756 ;
  assign n53758 = ( n8989 & ~n25514 ) | ( n8989 & n37720 ) | ( ~n25514 & n37720 ) ;
  assign n53759 = ( ~n3584 & n7241 ) | ( ~n3584 & n12097 ) | ( n7241 & n12097 ) ;
  assign n53760 = ( n7532 & n50154 ) | ( n7532 & ~n52675 ) | ( n50154 & ~n52675 ) ;
  assign n53761 = n53760 ^ n19829 ^ n12992 ;
  assign n53762 = ( ~n17159 & n21279 ) | ( ~n17159 & n49708 ) | ( n21279 & n49708 ) ;
  assign n53763 = ~n25133 & n52005 ;
  assign n53764 = ~n44962 & n53763 ;
  assign n53765 = n53764 ^ n48430 ^ n21176 ;
  assign n53766 = n53765 ^ n15106 ^ n10055 ;
  assign n53767 = ( n38544 & n38824 ) | ( n38544 & n43171 ) | ( n38824 & n43171 ) ;
  assign n53769 = n23530 | n27022 ;
  assign n53768 = n47459 ^ n45051 ^ n18439 ;
  assign n53770 = n53769 ^ n53768 ^ n26069 ;
  assign n53771 = n10722 ^ n873 ^ 1'b0 ;
  assign n53772 = n12592 & ~n53771 ;
  assign n53773 = ( ~n7074 & n22998 ) | ( ~n7074 & n53772 ) | ( n22998 & n53772 ) ;
  assign n53774 = n15952 | n53773 ;
  assign n53775 = n28126 | n53774 ;
  assign n53776 = n53617 ^ n44610 ^ n15398 ;
  assign n53777 = n29463 ^ n15506 ^ n13524 ;
  assign n53778 = n53777 ^ n19269 ^ n5407 ;
  assign n53779 = n53778 ^ n53070 ^ n30378 ;
  assign n53780 = ( n3803 & n34487 ) | ( n3803 & n46989 ) | ( n34487 & n46989 ) ;
  assign n53781 = n53780 ^ n51342 ^ 1'b0 ;
  assign n53782 = ( n21174 & n31245 ) | ( n21174 & n53781 ) | ( n31245 & n53781 ) ;
  assign n53783 = n44463 ^ n34810 ^ n28760 ;
  assign n53784 = ( ~n491 & n15857 ) | ( ~n491 & n48256 ) | ( n15857 & n48256 ) ;
  assign n53785 = ( n7071 & ~n44211 ) | ( n7071 & n53784 ) | ( ~n44211 & n53784 ) ;
  assign n53786 = n10382 & ~n18580 ;
  assign n53787 = n53786 ^ n40780 ^ n27879 ;
  assign n53788 = n53787 ^ n1694 ^ 1'b0 ;
  assign n53789 = n31044 ^ n19746 ^ n1839 ;
  assign n53790 = n53789 ^ n40135 ^ 1'b0 ;
  assign n53791 = ( ~n1711 & n16209 ) | ( ~n1711 & n41695 ) | ( n16209 & n41695 ) ;
  assign n53792 = n11790 | n14750 ;
  assign n53793 = n24391 | n53792 ;
  assign n53794 = n53793 ^ n45389 ^ 1'b0 ;
  assign n53795 = n50316 | n53794 ;
  assign n53796 = n18227 | n19207 ;
  assign n53797 = n47827 & ~n53796 ;
  assign n53799 = n21700 ^ n7338 ^ n6795 ;
  assign n53798 = n32252 ^ n27025 ^ n9229 ;
  assign n53800 = n53799 ^ n53798 ^ n41377 ;
  assign n53801 = n53800 ^ n32033 ^ n12980 ;
  assign n53802 = n43937 ^ n16125 ^ 1'b0 ;
  assign n53803 = n45409 ^ n20199 ^ n3936 ;
  assign n53804 = ( ~n1840 & n21355 ) | ( ~n1840 & n51810 ) | ( n21355 & n51810 ) ;
  assign n53805 = n26464 ^ n20047 ^ n17352 ;
  assign n53806 = n11939 ^ n7986 ^ n5610 ;
  assign n53807 = ( ~n4301 & n11849 ) | ( ~n4301 & n53806 ) | ( n11849 & n53806 ) ;
  assign n53808 = ( n22069 & n38301 ) | ( n22069 & n53807 ) | ( n38301 & n53807 ) ;
  assign n53809 = n22280 & n45317 ;
  assign n53810 = ~n26267 & n53809 ;
  assign n53811 = n23519 ^ n6142 ^ 1'b0 ;
  assign n53812 = ( n14606 & n18376 ) | ( n14606 & ~n28110 ) | ( n18376 & ~n28110 ) ;
  assign n53813 = ( n5967 & ~n49641 ) | ( n5967 & n53812 ) | ( ~n49641 & n53812 ) ;
  assign n53814 = n14195 | n53813 ;
  assign n53815 = n53811 | n53814 ;
  assign n53816 = ( n16405 & n20783 ) | ( n16405 & n28597 ) | ( n20783 & n28597 ) ;
  assign n53817 = n43550 ^ n10908 ^ n6215 ;
  assign n53818 = n40753 ^ n40220 ^ 1'b0 ;
  assign n53819 = n29404 ^ n21898 ^ n18484 ;
  assign n53820 = n27040 ^ n17824 ^ 1'b0 ;
  assign n53821 = ( n3410 & ~n9108 ) | ( n3410 & n53820 ) | ( ~n9108 & n53820 ) ;
  assign n53822 = n48083 ^ n38288 ^ n10504 ;
  assign n53823 = ( n17307 & n30931 ) | ( n17307 & n40144 ) | ( n30931 & n40144 ) ;
  assign n53824 = ( n7102 & n10273 ) | ( n7102 & n23408 ) | ( n10273 & n23408 ) ;
  assign n53825 = n17587 ^ n12286 ^ 1'b0 ;
  assign n53826 = n50868 | n53825 ;
  assign n53827 = n31716 ^ n2082 ^ 1'b0 ;
  assign n53828 = ( ~n12352 & n14551 ) | ( ~n12352 & n42123 ) | ( n14551 & n42123 ) ;
  assign n53829 = n46085 ^ n21054 ^ n15017 ;
  assign n53830 = ( n8829 & n12335 ) | ( n8829 & n37979 ) | ( n12335 & n37979 ) ;
  assign n53831 = ( n13334 & n25011 ) | ( n13334 & n40022 ) | ( n25011 & n40022 ) ;
  assign n53832 = n27953 ^ n16149 ^ n2628 ;
  assign n53833 = n53832 ^ n26685 ^ n20894 ;
  assign n53834 = n11016 | n53833 ;
  assign n53835 = ~n16328 & n36854 ;
  assign n53836 = n32755 & n53835 ;
  assign n53837 = ( ~n10606 & n21201 ) | ( ~n10606 & n38465 ) | ( n21201 & n38465 ) ;
  assign n53838 = ( n643 & n53836 ) | ( n643 & n53837 ) | ( n53836 & n53837 ) ;
  assign n53839 = n39359 ^ n32197 ^ n24214 ;
  assign n53840 = n26956 & ~n47444 ;
  assign n53841 = n2892 & ~n16250 ;
  assign n53842 = n53841 ^ n21652 ^ 1'b0 ;
  assign n53843 = n5952 | n24616 ;
  assign n53844 = n39677 & ~n53843 ;
  assign n53845 = n53844 ^ n43078 ^ n30889 ;
  assign n53846 = ~n40135 & n51289 ;
  assign n53847 = ~n53845 & n53846 ;
  assign n53852 = ( n3369 & n5359 ) | ( n3369 & n31876 ) | ( n5359 & n31876 ) ;
  assign n53853 = n53536 ^ n1767 ^ 1'b0 ;
  assign n53854 = ~n53852 & n53853 ;
  assign n53848 = n11652 | n19195 ;
  assign n53849 = n11475 | n53848 ;
  assign n53850 = n53849 ^ n22139 ^ n14722 ;
  assign n53851 = ( n5088 & n46129 ) | ( n5088 & n53850 ) | ( n46129 & n53850 ) ;
  assign n53855 = n53854 ^ n53851 ^ n25595 ;
  assign n53856 = n49893 ^ n18037 ^ n14002 ;
  assign n53857 = ( n32000 & ~n46644 ) | ( n32000 & n53856 ) | ( ~n46644 & n53856 ) ;
  assign n53858 = n42763 ^ n2159 ^ n868 ;
  assign n53859 = ~n7554 & n41711 ;
  assign n53860 = n37174 & n53859 ;
  assign n53861 = n53860 ^ n32412 ^ n17607 ;
  assign n53862 = ( n8969 & n13546 ) | ( n8969 & ~n22415 ) | ( n13546 & ~n22415 ) ;
  assign n53863 = ( n4422 & n7405 ) | ( n4422 & ~n11379 ) | ( n7405 & ~n11379 ) ;
  assign n53864 = n53695 ^ n4168 ^ 1'b0 ;
  assign n53865 = n48695 ^ n28870 ^ n21460 ;
  assign n53866 = n20089 ^ n7821 ^ 1'b0 ;
  assign n53867 = ~n38413 & n53866 ;
  assign n53868 = n48623 ^ n5156 ^ 1'b0 ;
  assign n53869 = n3093 | n53868 ;
  assign n53870 = n33116 & n39071 ;
  assign n53871 = n53870 ^ n9566 ^ 1'b0 ;
  assign n53872 = n53871 ^ n24205 ^ n3126 ;
  assign n53873 = n13394 ^ n7079 ^ n3143 ;
  assign n53874 = n26218 ^ n16194 ^ n1547 ;
  assign n53875 = n33858 ^ n23578 ^ n2133 ;
  assign n53876 = ( n14851 & ~n52827 ) | ( n14851 & n53875 ) | ( ~n52827 & n53875 ) ;
  assign n53877 = ~n24847 & n53876 ;
  assign n53878 = n53877 ^ n5954 ^ 1'b0 ;
  assign n53879 = n53878 ^ n50673 ^ n31413 ;
  assign n53880 = n39691 ^ n24162 ^ 1'b0 ;
  assign n53881 = n46378 ^ n45013 ^ n24038 ;
  assign n53882 = n47284 ^ n44574 ^ n7006 ;
  assign n53883 = n4787 & ~n14296 ;
  assign n53884 = n9055 & n53883 ;
  assign n53885 = n53884 ^ n2630 ^ 1'b0 ;
  assign n53886 = n48399 ^ n43063 ^ 1'b0 ;
  assign n53887 = n5590 | n53886 ;
  assign n53888 = ( n5329 & ~n18810 ) | ( n5329 & n22939 ) | ( ~n18810 & n22939 ) ;
  assign n53889 = n53888 ^ n32025 ^ n16019 ;
  assign n53890 = ( n3315 & n22410 ) | ( n3315 & ~n53889 ) | ( n22410 & ~n53889 ) ;
  assign n53891 = n1832 | n3450 ;
  assign n53892 = n53561 & ~n53891 ;
  assign n53893 = n40600 ^ n17621 ^ n15745 ;
  assign n53894 = ( ~n23238 & n33969 ) | ( ~n23238 & n49189 ) | ( n33969 & n49189 ) ;
  assign n53895 = n37942 ^ n8427 ^ x171 ;
  assign n53896 = ( n15241 & n23737 ) | ( n15241 & ~n36902 ) | ( n23737 & ~n36902 ) ;
  assign n53897 = n47182 | n48647 ;
  assign n53898 = n53896 | n53897 ;
  assign n53899 = n53898 ^ n41914 ^ n8646 ;
  assign n53900 = n19518 & ~n53899 ;
  assign n53902 = ( n12848 & n18466 ) | ( n12848 & n39129 ) | ( n18466 & n39129 ) ;
  assign n53901 = n46274 ^ n43261 ^ n9605 ;
  assign n53903 = n53902 ^ n53901 ^ n52646 ;
  assign n53904 = n26046 ^ n17173 ^ 1'b0 ;
  assign n53905 = x224 & ~n21171 ;
  assign n53906 = n53904 & n53905 ;
  assign n53907 = n2936 | n7130 ;
  assign n53909 = ~n5302 & n24351 ;
  assign n53910 = ~n24351 & n53909 ;
  assign n53911 = n7660 & ~n53910 ;
  assign n53912 = n53911 ^ n47694 ^ n34160 ;
  assign n53913 = n12768 & ~n53912 ;
  assign n53914 = n22074 & n53913 ;
  assign n53908 = ~n10626 & n35144 ;
  assign n53915 = n53914 ^ n53908 ^ 1'b0 ;
  assign n53918 = ( n31061 & n40285 ) | ( n31061 & ~n47711 ) | ( n40285 & ~n47711 ) ;
  assign n53916 = n9024 | n17503 ;
  assign n53917 = n53916 ^ n21533 ^ n6740 ;
  assign n53919 = n53918 ^ n53917 ^ n1444 ;
  assign n53920 = n45183 ^ n38823 ^ n10219 ;
  assign n53921 = ( n16662 & ~n17513 ) | ( n16662 & n53920 ) | ( ~n17513 & n53920 ) ;
  assign n53922 = ~n7032 & n37804 ;
  assign n53923 = ~n14026 & n31175 ;
  assign n53924 = ~n20900 & n28266 ;
  assign n53926 = ( n13049 & n22887 ) | ( n13049 & ~n29195 ) | ( n22887 & ~n29195 ) ;
  assign n53925 = ( n17536 & ~n23476 ) | ( n17536 & n24377 ) | ( ~n23476 & n24377 ) ;
  assign n53927 = n53926 ^ n53925 ^ n15111 ;
  assign n53928 = ( n11969 & n37390 ) | ( n11969 & n38343 ) | ( n37390 & n38343 ) ;
  assign n53929 = n53928 ^ n9628 ^ n4629 ;
  assign n53933 = n44446 ^ n26074 ^ n5277 ;
  assign n53930 = n43692 ^ n13697 ^ n10170 ;
  assign n53931 = n5439 & n8837 ;
  assign n53932 = ~n53930 & n53931 ;
  assign n53934 = n53933 ^ n53932 ^ n20132 ;
  assign n53935 = ~n36624 & n50473 ;
  assign n53936 = n26478 & n53935 ;
  assign n53937 = n42310 ^ n36431 ^ 1'b0 ;
  assign n53938 = ( n5952 & n7593 ) | ( n5952 & n42705 ) | ( n7593 & n42705 ) ;
  assign n53939 = ( n6766 & n45374 ) | ( n6766 & ~n52814 ) | ( n45374 & ~n52814 ) ;
  assign n53940 = ( ~n6804 & n11812 ) | ( ~n6804 & n28280 ) | ( n11812 & n28280 ) ;
  assign n53941 = n45163 ^ n19463 ^ n7747 ;
  assign n53942 = ( n347 & n9092 ) | ( n347 & ~n15350 ) | ( n9092 & ~n15350 ) ;
  assign n53943 = n51798 ^ n7551 ^ 1'b0 ;
  assign n53944 = n53942 | n53943 ;
  assign n53945 = ( n20170 & n27682 ) | ( n20170 & n53944 ) | ( n27682 & n53944 ) ;
  assign n53946 = ( ~n16275 & n31177 ) | ( ~n16275 & n37588 ) | ( n31177 & n37588 ) ;
  assign n53947 = n53946 ^ n44705 ^ n13330 ;
  assign n53948 = n47185 ^ n32806 ^ n2974 ;
  assign n53949 = ~n2546 & n2887 ;
  assign n53950 = n53949 ^ n31887 ^ 1'b0 ;
  assign n53951 = n50723 ^ n13545 ^ n9336 ;
  assign n53952 = ( n43826 & ~n45140 ) | ( n43826 & n53951 ) | ( ~n45140 & n53951 ) ;
  assign n53953 = ( n29469 & n53950 ) | ( n29469 & n53952 ) | ( n53950 & n53952 ) ;
  assign n53954 = n23113 ^ n20841 ^ 1'b0 ;
  assign n53955 = ( ~n2032 & n7337 ) | ( ~n2032 & n12597 ) | ( n7337 & n12597 ) ;
  assign n53956 = n40618 ^ n26209 ^ n10858 ;
  assign n53957 = n45649 ^ n43356 ^ n20175 ;
  assign n53958 = n48427 ^ n43050 ^ 1'b0 ;
  assign n53959 = n13013 & n53958 ;
  assign n53960 = ( n7268 & n34528 ) | ( n7268 & ~n53959 ) | ( n34528 & ~n53959 ) ;
  assign n53961 = ( n11164 & n11930 ) | ( n11164 & ~n39027 ) | ( n11930 & ~n39027 ) ;
  assign n53962 = n53961 ^ n21358 ^ n16411 ;
  assign n53963 = ( ~n7302 & n9509 ) | ( ~n7302 & n42314 ) | ( n9509 & n42314 ) ;
  assign n53964 = ~n13444 & n29427 ;
  assign n53966 = n22984 ^ n17408 ^ 1'b0 ;
  assign n53965 = ( ~n7176 & n28827 ) | ( ~n7176 & n29849 ) | ( n28827 & n29849 ) ;
  assign n53967 = n53966 ^ n53965 ^ n4275 ;
  assign n53968 = n14066 | n21439 ;
  assign n53969 = ( n19188 & ~n53967 ) | ( n19188 & n53968 ) | ( ~n53967 & n53968 ) ;
  assign n53970 = ~n6549 & n25366 ;
  assign n53971 = ~n35909 & n53970 ;
  assign n53972 = n19955 ^ n19157 ^ 1'b0 ;
  assign n53973 = n19719 & n53972 ;
  assign n53974 = n53973 ^ n11360 ^ 1'b0 ;
  assign n53975 = n39136 | n53974 ;
  assign n53976 = n53975 ^ n48894 ^ 1'b0 ;
  assign n53977 = ~n53971 & n53976 ;
  assign n53978 = n45977 ^ n35063 ^ n28223 ;
  assign n53979 = ( n7783 & n15213 ) | ( n7783 & ~n53978 ) | ( n15213 & ~n53978 ) ;
  assign n53980 = n39628 ^ n32626 ^ n9441 ;
  assign n53981 = n17631 ^ n15433 ^ n5167 ;
  assign n53982 = n16782 & n53981 ;
  assign n53984 = ~n3526 & n30043 ;
  assign n53985 = ~n25871 & n53984 ;
  assign n53983 = n41871 & n48492 ;
  assign n53986 = n53985 ^ n53983 ^ n20523 ;
  assign n53987 = n53986 ^ n25025 ^ n8281 ;
  assign n53988 = n42251 ^ n30171 ^ n8180 ;
  assign n53989 = ( n8992 & n10886 ) | ( n8992 & n27075 ) | ( n10886 & n27075 ) ;
  assign n53990 = ( n5184 & n30006 ) | ( n5184 & ~n53989 ) | ( n30006 & ~n53989 ) ;
  assign n53991 = ( ~n4348 & n15669 ) | ( ~n4348 & n51461 ) | ( n15669 & n51461 ) ;
  assign n53992 = n24925 ^ n18396 ^ n9761 ;
  assign n53993 = n2056 & n21694 ;
  assign n53994 = n22319 & n53993 ;
  assign n53995 = n8597 & ~n36320 ;
  assign n53996 = n24669 ^ n11656 ^ n10896 ;
  assign n53997 = ( n793 & n25913 ) | ( n793 & n27035 ) | ( n25913 & n27035 ) ;
  assign n53998 = ( n27506 & ~n53996 ) | ( n27506 & n53997 ) | ( ~n53996 & n53997 ) ;
  assign n53999 = n53998 ^ n39289 ^ n15058 ;
  assign n54000 = n42403 ^ x227 ^ 1'b0 ;
  assign n54001 = n54000 ^ n34949 ^ n30339 ;
  assign n54002 = n3379 & n11828 ;
  assign n54003 = n49994 ^ n21541 ^ n9100 ;
  assign n54006 = ( n14824 & n20898 ) | ( n14824 & n29286 ) | ( n20898 & n29286 ) ;
  assign n54004 = ( n11395 & n22540 ) | ( n11395 & n36782 ) | ( n22540 & n36782 ) ;
  assign n54005 = ( n11621 & ~n24127 ) | ( n11621 & n54004 ) | ( ~n24127 & n54004 ) ;
  assign n54007 = n54006 ^ n54005 ^ n17113 ;
  assign n54008 = n26466 ^ n23164 ^ 1'b0 ;
  assign n54009 = n24074 & ~n54008 ;
  assign n54010 = ( n17478 & ~n38642 ) | ( n17478 & n54009 ) | ( ~n38642 & n54009 ) ;
  assign n54011 = n47671 ^ n35229 ^ n33062 ;
  assign n54012 = n40153 ^ n25765 ^ n7463 ;
  assign n54013 = ( n1770 & n36963 ) | ( n1770 & ~n54012 ) | ( n36963 & ~n54012 ) ;
  assign n54014 = n21585 | n25138 ;
  assign n54015 = n28996 | n54014 ;
  assign n54016 = n47699 ^ n2891 ^ 1'b0 ;
  assign n54017 = ~n13329 & n54016 ;
  assign n54018 = ( n2901 & ~n9422 ) | ( n2901 & n39837 ) | ( ~n9422 & n39837 ) ;
  assign n54019 = n2167 | n31789 ;
  assign n54020 = n54019 ^ n4503 ^ 1'b0 ;
  assign n54021 = n54020 ^ n12701 ^ n6454 ;
  assign n54022 = ( n2142 & ~n8463 ) | ( n2142 & n11471 ) | ( ~n8463 & n11471 ) ;
  assign n54023 = n54022 ^ n36425 ^ n13507 ;
  assign n54024 = ( n9257 & n9739 ) | ( n9257 & n25001 ) | ( n9739 & n25001 ) ;
  assign n54025 = ( n13494 & ~n15649 ) | ( n13494 & n54024 ) | ( ~n15649 & n54024 ) ;
  assign n54026 = ~n47014 & n54025 ;
  assign n54027 = n7044 & n13879 ;
  assign n54028 = n54027 ^ n13954 ^ 1'b0 ;
  assign n54029 = ( n8042 & ~n29964 ) | ( n8042 & n36415 ) | ( ~n29964 & n36415 ) ;
  assign n54030 = n54029 ^ n14584 ^ n13116 ;
  assign n54031 = ( ~n35956 & n40626 ) | ( ~n35956 & n54030 ) | ( n40626 & n54030 ) ;
  assign n54032 = ( ~n18674 & n54028 ) | ( ~n18674 & n54031 ) | ( n54028 & n54031 ) ;
  assign n54034 = ~n9836 & n24373 ;
  assign n54035 = n54034 ^ n46397 ^ 1'b0 ;
  assign n54033 = n39012 ^ n31381 ^ n18753 ;
  assign n54036 = n54035 ^ n54033 ^ n12157 ;
  assign n54037 = n49562 ^ n9066 ^ n445 ;
  assign n54038 = n12807 | n21171 ;
  assign n54039 = n54038 ^ n22249 ^ 1'b0 ;
  assign n54040 = n54039 ^ n34369 ^ 1'b0 ;
  assign n54041 = n7711 & n35894 ;
  assign n54042 = n54041 ^ n2832 ^ 1'b0 ;
  assign n54043 = n35118 & ~n51410 ;
  assign n54044 = n32900 & n54043 ;
  assign n54045 = n12416 ^ n10494 ^ 1'b0 ;
  assign n54046 = ~n21027 & n54045 ;
  assign n54047 = ( ~n4529 & n22527 ) | ( ~n4529 & n37384 ) | ( n22527 & n37384 ) ;
  assign n54048 = ( n17583 & n47058 ) | ( n17583 & ~n54047 ) | ( n47058 & ~n54047 ) ;
  assign n54049 = n39896 ^ n15399 ^ n14372 ;
  assign n54050 = n41533 ^ n22938 ^ n12278 ;
  assign n54051 = ( ~n50899 & n54049 ) | ( ~n50899 & n54050 ) | ( n54049 & n54050 ) ;
  assign n54052 = ( n14644 & n18972 ) | ( n14644 & n51881 ) | ( n18972 & n51881 ) ;
  assign n54054 = n9844 ^ n7195 ^ n3742 ;
  assign n54053 = n49500 ^ n24708 ^ n20350 ;
  assign n54055 = n54054 ^ n54053 ^ n21484 ;
  assign n54056 = n33861 ^ n25183 ^ n14359 ;
  assign n54057 = n54056 ^ n33772 ^ n28932 ;
  assign n54061 = n35483 & ~n41194 ;
  assign n54058 = n18441 & ~n33210 ;
  assign n54059 = n54058 ^ n37940 ^ 1'b0 ;
  assign n54060 = ( n26801 & ~n39758 ) | ( n26801 & n54059 ) | ( ~n39758 & n54059 ) ;
  assign n54062 = n54061 ^ n54060 ^ n7796 ;
  assign n54063 = n44372 ^ n42603 ^ n19404 ;
  assign n54064 = ( n16890 & n23479 ) | ( n16890 & ~n32226 ) | ( n23479 & ~n32226 ) ;
  assign n54065 = n11737 & ~n17393 ;
  assign n54066 = n25466 & n37401 ;
  assign n54067 = n25832 | n54066 ;
  assign n54068 = n4060 & ~n54067 ;
  assign n54069 = n32093 & ~n35074 ;
  assign n54070 = n23089 & n54069 ;
  assign n54071 = n16486 ^ n8249 ^ n7919 ;
  assign n54072 = ( n1270 & n19211 ) | ( n1270 & n54071 ) | ( n19211 & n54071 ) ;
  assign n54073 = ~n342 & n30454 ;
  assign n54074 = n54073 ^ n14918 ^ 1'b0 ;
  assign n54075 = n54074 ^ n49131 ^ n35403 ;
  assign n54076 = ( ~n38998 & n51619 ) | ( ~n38998 & n54075 ) | ( n51619 & n54075 ) ;
  assign n54079 = n22134 | n37605 ;
  assign n54080 = n54079 ^ n3794 ^ 1'b0 ;
  assign n54077 = n5145 | n44095 ;
  assign n54078 = n25317 & ~n54077 ;
  assign n54081 = n54080 ^ n54078 ^ n41637 ;
  assign n54082 = n38994 | n39265 ;
  assign n54085 = ( n1366 & n48279 ) | ( n1366 & ~n50697 ) | ( n48279 & ~n50697 ) ;
  assign n54083 = n34772 ^ n33400 ^ 1'b0 ;
  assign n54084 = ( n4311 & n15734 ) | ( n4311 & n54083 ) | ( n15734 & n54083 ) ;
  assign n54086 = n54085 ^ n54084 ^ n42246 ;
  assign n54087 = n34383 | n46396 ;
  assign n54088 = ( n15807 & n32010 ) | ( n15807 & ~n54087 ) | ( n32010 & ~n54087 ) ;
  assign n54089 = ( n35495 & ~n39829 ) | ( n35495 & n45825 ) | ( ~n39829 & n45825 ) ;
  assign n54090 = n47131 ^ n22057 ^ n8569 ;
  assign n54091 = n641 | n54090 ;
  assign n54092 = n53710 | n54091 ;
  assign n54093 = n30752 ^ n9227 ^ n7862 ;
  assign n54094 = n32323 | n39232 ;
  assign n54095 = n54093 | n54094 ;
  assign n54096 = ~n8681 & n52849 ;
  assign n54097 = n54096 ^ n12168 ^ 1'b0 ;
  assign n54098 = n22952 ^ n7152 ^ 1'b0 ;
  assign n54099 = ( ~n14023 & n19276 ) | ( ~n14023 & n54098 ) | ( n19276 & n54098 ) ;
  assign n54100 = ~n2495 & n3707 ;
  assign n54101 = ( n12662 & n17021 ) | ( n12662 & n54100 ) | ( n17021 & n54100 ) ;
  assign n54102 = n53013 ^ n36782 ^ n490 ;
  assign n54103 = ( n25452 & ~n41898 ) | ( n25452 & n53719 ) | ( ~n41898 & n53719 ) ;
  assign n54104 = n13139 ^ n9319 ^ n2036 ;
  assign n54105 = n20718 ^ n17362 ^ n16493 ;
  assign n54106 = ( ~n10737 & n39348 ) | ( ~n10737 & n54105 ) | ( n39348 & n54105 ) ;
  assign n54107 = ( n16998 & n40442 ) | ( n16998 & ~n54106 ) | ( n40442 & ~n54106 ) ;
  assign n54108 = n49533 ^ n27939 ^ n6131 ;
  assign n54109 = ( x26 & ~n10452 ) | ( x26 & n14935 ) | ( ~n10452 & n14935 ) ;
  assign n54110 = n33838 & ~n54109 ;
  assign n54111 = n54108 & n54110 ;
  assign n54112 = ~n16073 & n21381 ;
  assign n54113 = n54112 ^ n41485 ^ 1'b0 ;
  assign n54114 = ( n1707 & n26190 ) | ( n1707 & ~n33607 ) | ( n26190 & ~n33607 ) ;
  assign n54115 = n8719 & n54114 ;
  assign n54116 = n54115 ^ n1467 ^ 1'b0 ;
  assign n54117 = n54113 | n54116 ;
  assign n54118 = ~n1295 & n26002 ;
  assign n54119 = ( n2201 & ~n17018 ) | ( n2201 & n33541 ) | ( ~n17018 & n33541 ) ;
  assign n54120 = ( ~n23192 & n30187 ) | ( ~n23192 & n54119 ) | ( n30187 & n54119 ) ;
  assign n54121 = ( n31708 & n54118 ) | ( n31708 & n54120 ) | ( n54118 & n54120 ) ;
  assign n54122 = n38887 ^ n38270 ^ n461 ;
  assign n54123 = n12433 | n34602 ;
  assign n54124 = n53876 ^ n28280 ^ n8342 ;
  assign n54128 = n33024 ^ n10362 ^ n1012 ;
  assign n54125 = n53410 ^ n697 ^ n338 ;
  assign n54126 = n31778 ^ n3333 ^ 1'b0 ;
  assign n54127 = n54125 & n54126 ;
  assign n54129 = n54128 ^ n54127 ^ 1'b0 ;
  assign n54130 = ( n8959 & n30732 ) | ( n8959 & n37796 ) | ( n30732 & n37796 ) ;
  assign n54131 = ( ~n27269 & n30905 ) | ( ~n27269 & n54130 ) | ( n30905 & n54130 ) ;
  assign n54132 = ( n3576 & n15396 ) | ( n3576 & ~n54131 ) | ( n15396 & ~n54131 ) ;
  assign n54134 = ( ~n14419 & n21726 ) | ( ~n14419 & n36108 ) | ( n21726 & n36108 ) ;
  assign n54133 = n29357 ^ n17922 ^ n17795 ;
  assign n54135 = n54134 ^ n54133 ^ n40043 ;
  assign n54136 = ~n3679 & n33986 ;
  assign n54137 = ~n33484 & n54136 ;
  assign n54138 = ( n21346 & ~n39059 ) | ( n21346 & n54137 ) | ( ~n39059 & n54137 ) ;
  assign n54139 = n44957 ^ n19774 ^ 1'b0 ;
  assign n54140 = n15344 & ~n54139 ;
  assign n54142 = n37619 ^ n19121 ^ 1'b0 ;
  assign n54141 = n849 | n34434 ;
  assign n54143 = n54142 ^ n54141 ^ 1'b0 ;
  assign n54144 = n5095 & n43018 ;
  assign n54145 = n6569 & ~n54144 ;
  assign n54146 = n54145 ^ n11664 ^ 1'b0 ;
  assign n54147 = n3063 & ~n20487 ;
  assign n54148 = ( n14449 & n14551 ) | ( n14449 & ~n33401 ) | ( n14551 & ~n33401 ) ;
  assign n54149 = n54148 ^ n745 ^ 1'b0 ;
  assign n54150 = n54147 | n54149 ;
  assign n54151 = n39196 | n54150 ;
  assign n54152 = n33343 ^ n23564 ^ n15370 ;
  assign n54153 = n19346 ^ n2042 ^ 1'b0 ;
  assign n54154 = n54153 ^ n33390 ^ n22872 ;
  assign n54155 = ( x152 & ~n19640 ) | ( x152 & n54154 ) | ( ~n19640 & n54154 ) ;
  assign n54156 = ( n35930 & n40018 ) | ( n35930 & ~n54155 ) | ( n40018 & ~n54155 ) ;
  assign n54157 = n17808 & ~n48251 ;
  assign n54158 = n54156 & n54157 ;
  assign n54159 = ( ~n34235 & n54152 ) | ( ~n34235 & n54158 ) | ( n54152 & n54158 ) ;
  assign n54160 = n21609 ^ n7045 ^ n3231 ;
  assign n54161 = n54160 ^ n14715 ^ n7008 ;
  assign n54163 = n6897 & n27255 ;
  assign n54162 = n37340 ^ n28433 ^ n2485 ;
  assign n54164 = n54163 ^ n54162 ^ n2054 ;
  assign n54165 = ( ~n13745 & n54161 ) | ( ~n13745 & n54164 ) | ( n54161 & n54164 ) ;
  assign n54166 = n38875 ^ n23166 ^ n19200 ;
  assign n54167 = n4334 | n29160 ;
  assign n54168 = n9353 & ~n11020 ;
  assign n54169 = ( ~n3082 & n25555 ) | ( ~n3082 & n54168 ) | ( n25555 & n54168 ) ;
  assign n54170 = ( n36976 & n51988 ) | ( n36976 & n54169 ) | ( n51988 & n54169 ) ;
  assign n54171 = ( ~n16350 & n54167 ) | ( ~n16350 & n54170 ) | ( n54167 & n54170 ) ;
  assign n54172 = ( n20354 & n22309 ) | ( n20354 & n41043 ) | ( n22309 & n41043 ) ;
  assign n54173 = n41404 ^ n11157 ^ n3324 ;
  assign n54174 = ~n2524 & n15535 ;
  assign n54175 = n54174 ^ n12813 ^ 1'b0 ;
  assign n54176 = n37757 ^ n34240 ^ 1'b0 ;
  assign n54177 = ~n47582 & n54176 ;
  assign n54178 = n54177 ^ n16765 ^ 1'b0 ;
  assign n54179 = n37813 & n54178 ;
  assign n54180 = n54179 ^ n18241 ^ 1'b0 ;
  assign n54181 = n17750 ^ n5557 ^ 1'b0 ;
  assign n54182 = ~n45094 & n54181 ;
  assign n54183 = n48801 ^ n35026 ^ n28523 ;
  assign n54184 = n26152 ^ n25592 ^ n15510 ;
  assign n54185 = ~n16627 & n18382 ;
  assign n54186 = n54184 & n54185 ;
  assign n54187 = ( n19156 & n39028 ) | ( n19156 & ~n41945 ) | ( n39028 & ~n41945 ) ;
  assign n54188 = ( n29668 & n54186 ) | ( n29668 & n54187 ) | ( n54186 & n54187 ) ;
  assign n54189 = n42085 ^ n28601 ^ n2806 ;
  assign n54190 = ( n6092 & n22506 ) | ( n6092 & n25801 ) | ( n22506 & n25801 ) ;
  assign n54191 = n34074 ^ n13282 ^ n1655 ;
  assign n54192 = ( n6582 & ~n16120 ) | ( n6582 & n33736 ) | ( ~n16120 & n33736 ) ;
  assign n54193 = n11409 ^ n10084 ^ n5376 ;
  assign n54195 = n40934 ^ n26521 ^ n4130 ;
  assign n54196 = ( ~n17613 & n27617 ) | ( ~n17613 & n54195 ) | ( n27617 & n54195 ) ;
  assign n54194 = ~n4824 & n8454 ;
  assign n54197 = n54196 ^ n54194 ^ 1'b0 ;
  assign n54198 = n28307 & ~n49013 ;
  assign n54199 = n21425 ^ n15934 ^ 1'b0 ;
  assign n54200 = ( n8379 & ~n20035 ) | ( n8379 & n54199 ) | ( ~n20035 & n54199 ) ;
  assign n54201 = n47872 ^ n21063 ^ n11813 ;
  assign n54202 = n23101 ^ n10479 ^ 1'b0 ;
  assign n54203 = n47018 ^ n36624 ^ n27392 ;
  assign n54204 = n19013 ^ n12565 ^ n11547 ;
  assign n54205 = ( ~n22308 & n24075 ) | ( ~n22308 & n54204 ) | ( n24075 & n54204 ) ;
  assign n54206 = ( n11058 & n25761 ) | ( n11058 & ~n54205 ) | ( n25761 & ~n54205 ) ;
  assign n54207 = ( n10928 & ~n14794 ) | ( n10928 & n25603 ) | ( ~n14794 & n25603 ) ;
  assign n54208 = ( n1717 & n2492 ) | ( n1717 & n54207 ) | ( n2492 & n54207 ) ;
  assign n54209 = ( n18410 & ~n39266 ) | ( n18410 & n51854 ) | ( ~n39266 & n51854 ) ;
  assign n54214 = ( n3399 & n8686 ) | ( n3399 & ~n9902 ) | ( n8686 & ~n9902 ) ;
  assign n54210 = n11039 ^ n5457 ^ n1015 ;
  assign n54211 = n54210 ^ n579 ^ 1'b0 ;
  assign n54212 = n5880 & n54211 ;
  assign n54213 = n18263 & n54212 ;
  assign n54215 = n54214 ^ n54213 ^ x225 ;
  assign n54216 = ( n30337 & ~n46494 ) | ( n30337 & n54215 ) | ( ~n46494 & n54215 ) ;
  assign n54217 = ~n6467 & n44071 ;
  assign n54218 = n54217 ^ n18145 ^ 1'b0 ;
  assign n54219 = n35031 ^ n25337 ^ 1'b0 ;
  assign n54220 = ~n22114 & n54219 ;
  assign n54221 = n15674 ^ n2565 ^ 1'b0 ;
  assign n54222 = ( n28857 & n34148 ) | ( n28857 & n51815 ) | ( n34148 & n51815 ) ;
  assign n54223 = ( ~n8942 & n45001 ) | ( ~n8942 & n54222 ) | ( n45001 & n54222 ) ;
  assign n54224 = n8178 ^ n1822 ^ 1'b0 ;
  assign n54225 = n545 | n23389 ;
  assign n54226 = ( n17515 & n49045 ) | ( n17515 & ~n54225 ) | ( n49045 & ~n54225 ) ;
  assign n54229 = ( n757 & ~n6098 ) | ( n757 & n17376 ) | ( ~n6098 & n17376 ) ;
  assign n54227 = n30526 & n36882 ;
  assign n54228 = ~n8007 & n54227 ;
  assign n54230 = n54229 ^ n54228 ^ n27602 ;
  assign n54231 = n49446 ^ n23618 ^ 1'b0 ;
  assign n54232 = n27326 ^ n639 ^ 1'b0 ;
  assign n54233 = ( n3282 & ~n5372 ) | ( n3282 & n35502 ) | ( ~n5372 & n35502 ) ;
  assign n54234 = n20918 | n48524 ;
  assign n54235 = n54234 ^ n29618 ^ 1'b0 ;
  assign n54236 = n9672 & n22431 ;
  assign n54237 = n27075 & n54236 ;
  assign n54238 = n54237 ^ n468 ^ 1'b0 ;
  assign n54239 = n33880 & n54238 ;
  assign n54240 = ~n1926 & n14800 ;
  assign n54241 = ( n2096 & ~n33682 ) | ( n2096 & n54240 ) | ( ~n33682 & n54240 ) ;
  assign n54242 = n29643 ^ n21217 ^ 1'b0 ;
  assign n54243 = ~n6336 & n24118 ;
  assign n54244 = ( n7640 & n19978 ) | ( n7640 & ~n37267 ) | ( n19978 & ~n37267 ) ;
  assign n54245 = n54244 ^ n17019 ^ n12093 ;
  assign n54246 = ( ~n13844 & n29558 ) | ( ~n13844 & n38415 ) | ( n29558 & n38415 ) ;
  assign n54247 = n2444 & n15919 ;
  assign n54248 = ( ~n16565 & n47334 ) | ( ~n16565 & n54247 ) | ( n47334 & n54247 ) ;
  assign n54249 = ( ~n7187 & n8965 ) | ( ~n7187 & n20144 ) | ( n8965 & n20144 ) ;
  assign n54250 = n54249 ^ n46489 ^ n9572 ;
  assign n54251 = n27443 ^ n5903 ^ n1217 ;
  assign n54252 = n42524 & n54251 ;
  assign n54253 = n54252 ^ n21599 ^ 1'b0 ;
  assign n54254 = n20073 ^ n4583 ^ 1'b0 ;
  assign n54255 = ( n569 & ~n18390 ) | ( n569 & n37110 ) | ( ~n18390 & n37110 ) ;
  assign n54256 = n18973 ^ n14340 ^ n2804 ;
  assign n54257 = n53178 ^ n12278 ^ 1'b0 ;
  assign n54258 = n6709 & ~n9361 ;
  assign n54259 = n9307 & ~n34058 ;
  assign n54260 = ~n9882 & n26667 ;
  assign n54261 = n35949 ^ n22015 ^ 1'b0 ;
  assign n54262 = ~n28344 & n54261 ;
  assign n54263 = ( n11917 & n54260 ) | ( n11917 & ~n54262 ) | ( n54260 & ~n54262 ) ;
  assign n54264 = ~n9819 & n24706 ;
  assign n54265 = ~n3427 & n54264 ;
  assign n54266 = n270 & ~n27075 ;
  assign n54267 = n54266 ^ n33226 ^ 1'b0 ;
  assign n54268 = ( n3359 & ~n23746 ) | ( n3359 & n25259 ) | ( ~n23746 & n25259 ) ;
  assign n54269 = ~n23793 & n29419 ;
  assign n54270 = ( ~n633 & n17070 ) | ( ~n633 & n44897 ) | ( n17070 & n44897 ) ;
  assign n54271 = ( ~n18122 & n54269 ) | ( ~n18122 & n54270 ) | ( n54269 & n54270 ) ;
  assign n54272 = ( ~n16707 & n18072 ) | ( ~n16707 & n54271 ) | ( n18072 & n54271 ) ;
  assign n54273 = n34184 & ~n49682 ;
  assign n54274 = ( ~n18318 & n23636 ) | ( ~n18318 & n28073 ) | ( n23636 & n28073 ) ;
  assign n54275 = n20350 & ~n54274 ;
  assign n54276 = n54275 ^ n33623 ^ n9029 ;
  assign n54283 = n42223 ^ n23305 ^ n21967 ;
  assign n54277 = n32665 ^ n12834 ^ 1'b0 ;
  assign n54278 = n7342 & n39898 ;
  assign n54279 = ~n6429 & n54278 ;
  assign n54280 = ( n10543 & n22777 ) | ( n10543 & ~n54279 ) | ( n22777 & ~n54279 ) ;
  assign n54281 = ( n10242 & n49643 ) | ( n10242 & n54280 ) | ( n49643 & n54280 ) ;
  assign n54282 = ( n22255 & ~n54277 ) | ( n22255 & n54281 ) | ( ~n54277 & n54281 ) ;
  assign n54284 = n54283 ^ n54282 ^ n2525 ;
  assign n54285 = ( ~n8009 & n37861 ) | ( ~n8009 & n40028 ) | ( n37861 & n40028 ) ;
  assign n54286 = n38341 ^ n5910 ^ x213 ;
  assign n54287 = n54286 ^ n39423 ^ n9003 ;
  assign n54288 = ~n51389 & n54287 ;
  assign n54289 = n17505 ^ n11007 ^ 1'b0 ;
  assign n54290 = n25378 & n54289 ;
  assign n54291 = n54290 ^ n33146 ^ n23016 ;
  assign n54292 = n17080 | n31147 ;
  assign n54293 = n54292 ^ n13317 ^ n5841 ;
  assign n54294 = ( n16565 & ~n16765 ) | ( n16565 & n54293 ) | ( ~n16765 & n54293 ) ;
  assign n54295 = ( n54288 & n54291 ) | ( n54288 & ~n54294 ) | ( n54291 & ~n54294 ) ;
  assign n54296 = ( ~n388 & n13824 ) | ( ~n388 & n53515 ) | ( n13824 & n53515 ) ;
  assign n54297 = ( n17275 & n39083 ) | ( n17275 & n54296 ) | ( n39083 & n54296 ) ;
  assign n54298 = ( n2258 & n29975 ) | ( n2258 & ~n54297 ) | ( n29975 & ~n54297 ) ;
  assign n54299 = n4657 & ~n18657 ;
  assign n54300 = n52198 & n54299 ;
  assign n54301 = n22172 & ~n47861 ;
  assign n54302 = n54301 ^ n34141 ^ n33911 ;
  assign n54303 = n23370 & ~n54302 ;
  assign n54304 = n21652 ^ n14114 ^ 1'b0 ;
  assign n54305 = n41067 | n54304 ;
  assign n54306 = n54305 ^ n53851 ^ n27468 ;
  assign n54307 = n32310 ^ n20857 ^ n1972 ;
  assign n54308 = n54307 ^ n54211 ^ n13753 ;
  assign n54309 = ( n16757 & n34739 ) | ( n16757 & ~n41782 ) | ( n34739 & ~n41782 ) ;
  assign n54310 = ( ~n3433 & n5527 ) | ( ~n3433 & n54309 ) | ( n5527 & n54309 ) ;
  assign n54311 = n35051 ^ n30670 ^ 1'b0 ;
  assign n54312 = ( ~n16950 & n19846 ) | ( ~n16950 & n44668 ) | ( n19846 & n44668 ) ;
  assign n54313 = n25020 ^ n498 ^ 1'b0 ;
  assign n54314 = ( ~n7177 & n31057 ) | ( ~n7177 & n54313 ) | ( n31057 & n54313 ) ;
  assign n54315 = n35768 ^ n22785 ^ n20449 ;
  assign n54316 = n1316 & n11955 ;
  assign n54317 = n54316 ^ n46011 ^ 1'b0 ;
  assign n54318 = ( n11536 & ~n54315 ) | ( n11536 & n54317 ) | ( ~n54315 & n54317 ) ;
  assign n54319 = n30180 ^ n17657 ^ 1'b0 ;
  assign n54320 = n42078 ^ n12542 ^ n10053 ;
  assign n54321 = ( n32886 & n54319 ) | ( n32886 & n54320 ) | ( n54319 & n54320 ) ;
  assign n54322 = n53134 ^ n365 ^ 1'b0 ;
  assign n54323 = n19801 & n54322 ;
  assign n54324 = n5920 & n14910 ;
  assign n54325 = n54324 ^ n7249 ^ 1'b0 ;
  assign n54326 = ~n22298 & n42508 ;
  assign n54327 = ~n54325 & n54326 ;
  assign n54328 = n54327 ^ n50665 ^ 1'b0 ;
  assign n54329 = ( n5689 & n7394 ) | ( n5689 & n54328 ) | ( n7394 & n54328 ) ;
  assign n54330 = ( n1217 & n39727 ) | ( n1217 & n45377 ) | ( n39727 & n45377 ) ;
  assign n54331 = n54330 ^ n45510 ^ n16751 ;
  assign n54332 = ( n8367 & n9624 ) | ( n8367 & n10445 ) | ( n9624 & n10445 ) ;
  assign n54333 = n54332 ^ n37390 ^ n29419 ;
  assign n54334 = ( n8258 & n19124 ) | ( n8258 & ~n24393 ) | ( n19124 & ~n24393 ) ;
  assign n54335 = n14377 ^ n14308 ^ n10161 ;
  assign n54336 = ( n23369 & ~n23443 ) | ( n23369 & n37562 ) | ( ~n23443 & n37562 ) ;
  assign n54337 = n21152 ^ n15933 ^ n5899 ;
  assign n54338 = ( n51666 & n52131 ) | ( n51666 & ~n54337 ) | ( n52131 & ~n54337 ) ;
  assign n54339 = n44375 ^ n25747 ^ n5918 ;
  assign n54340 = n54339 ^ n46239 ^ n7093 ;
  assign n54341 = ( n25888 & n33134 ) | ( n25888 & n54340 ) | ( n33134 & n54340 ) ;
  assign n54342 = n7927 & n52728 ;
  assign n54343 = n54342 ^ n9760 ^ 1'b0 ;
  assign n54347 = n11398 ^ n9104 ^ n8394 ;
  assign n54348 = n54347 ^ n35025 ^ 1'b0 ;
  assign n54344 = n18010 ^ n16432 ^ n2319 ;
  assign n54345 = n54344 ^ n27947 ^ n4823 ;
  assign n54346 = n5347 | n54345 ;
  assign n54349 = n54348 ^ n54346 ^ 1'b0 ;
  assign n54350 = ( n5900 & n15550 ) | ( n5900 & ~n27706 ) | ( n15550 & ~n27706 ) ;
  assign n54352 = n14296 ^ n4763 ^ n460 ;
  assign n54351 = n31589 ^ n15749 ^ n4984 ;
  assign n54353 = n54352 ^ n54351 ^ n37389 ;
  assign n54354 = n54353 ^ n35811 ^ n13925 ;
  assign n54355 = n31227 ^ n17519 ^ n3399 ;
  assign n54356 = ( ~n2738 & n5498 ) | ( ~n2738 & n5739 ) | ( n5498 & n5739 ) ;
  assign n54357 = n54356 ^ n34807 ^ n12260 ;
  assign n54358 = ( n1166 & n6578 ) | ( n1166 & n6751 ) | ( n6578 & n6751 ) ;
  assign n54359 = ( ~n19446 & n36330 ) | ( ~n19446 & n54358 ) | ( n36330 & n54358 ) ;
  assign n54360 = n54359 ^ n32737 ^ n13423 ;
  assign n54361 = n12899 & n48362 ;
  assign n54362 = ( n33852 & n38285 ) | ( n33852 & ~n54361 ) | ( n38285 & ~n54361 ) ;
  assign n54363 = n7229 ^ n6915 ^ x198 ;
  assign n54364 = ( n463 & ~n5824 ) | ( n463 & n18536 ) | ( ~n5824 & n18536 ) ;
  assign n54365 = n46600 ^ n31221 ^ n25616 ;
  assign n54366 = ( ~n10567 & n17650 ) | ( ~n10567 & n54365 ) | ( n17650 & n54365 ) ;
  assign n54367 = ( n5115 & n54364 ) | ( n5115 & ~n54366 ) | ( n54364 & ~n54366 ) ;
  assign n54368 = n31370 | n37222 ;
  assign n54369 = n54368 ^ n25584 ^ 1'b0 ;
  assign n54370 = n25764 | n54369 ;
  assign n54371 = n9016 ^ n7894 ^ 1'b0 ;
  assign n54372 = n10832 & n54371 ;
  assign n54373 = n54372 ^ n27116 ^ 1'b0 ;
  assign n54374 = n39860 ^ n4630 ^ 1'b0 ;
  assign n54375 = ( n817 & ~n9858 ) | ( n817 & n54374 ) | ( ~n9858 & n54374 ) ;
  assign n54376 = n16859 ^ n12090 ^ 1'b0 ;
  assign n54377 = ( ~n1149 & n5041 ) | ( ~n1149 & n14006 ) | ( n5041 & n14006 ) ;
  assign n54378 = n54377 ^ n28020 ^ n23996 ;
  assign n54379 = ( n14710 & n18031 ) | ( n14710 & ~n54378 ) | ( n18031 & ~n54378 ) ;
  assign n54387 = n5343 | n6807 ;
  assign n54380 = ( ~n8387 & n15100 ) | ( ~n8387 & n21496 ) | ( n15100 & n21496 ) ;
  assign n54381 = ( n3820 & ~n12980 ) | ( n3820 & n16094 ) | ( ~n12980 & n16094 ) ;
  assign n54382 = ( ~n25599 & n33141 ) | ( ~n25599 & n54381 ) | ( n33141 & n54381 ) ;
  assign n54383 = n9186 & n54382 ;
  assign n54384 = ~n9548 & n54383 ;
  assign n54385 = n28350 & ~n54384 ;
  assign n54386 = ( n46536 & n54380 ) | ( n46536 & n54385 ) | ( n54380 & n54385 ) ;
  assign n54388 = n54387 ^ n54386 ^ 1'b0 ;
  assign n54390 = ( n6114 & ~n19077 ) | ( n6114 & n23746 ) | ( ~n19077 & n23746 ) ;
  assign n54389 = n10088 & n19921 ;
  assign n54391 = n54390 ^ n54389 ^ 1'b0 ;
  assign n54392 = ( n18379 & ~n23443 ) | ( n18379 & n54391 ) | ( ~n23443 & n54391 ) ;
  assign n54393 = n54392 ^ n12648 ^ n4460 ;
  assign n54394 = ( n10124 & n16209 ) | ( n10124 & ~n40919 ) | ( n16209 & ~n40919 ) ;
  assign n54398 = n37173 ^ n11724 ^ n3231 ;
  assign n54399 = n9832 & ~n54398 ;
  assign n54396 = n23885 ^ n13261 ^ n9173 ;
  assign n54395 = n42023 ^ n20623 ^ n6796 ;
  assign n54397 = n54396 ^ n54395 ^ n20783 ;
  assign n54400 = n54399 ^ n54397 ^ n16879 ;
  assign n54401 = n31729 ^ n21084 ^ n17781 ;
  assign n54402 = ~n16382 & n54401 ;
  assign n54403 = n54402 ^ n27474 ^ 1'b0 ;
  assign n54404 = ( ~n1801 & n2201 ) | ( ~n1801 & n25030 ) | ( n2201 & n25030 ) ;
  assign n54405 = n11794 ^ n11604 ^ n4869 ;
  assign n54406 = ( n13132 & n15519 ) | ( n13132 & n50562 ) | ( n15519 & n50562 ) ;
  assign n54407 = ( ~x213 & n31135 ) | ( ~x213 & n54406 ) | ( n31135 & n54406 ) ;
  assign n54408 = ( ~n19971 & n54405 ) | ( ~n19971 & n54407 ) | ( n54405 & n54407 ) ;
  assign n54409 = ( n1679 & n16443 ) | ( n1679 & ~n20473 ) | ( n16443 & ~n20473 ) ;
  assign n54410 = n4280 & ~n54409 ;
  assign n54411 = n54410 ^ n29849 ^ 1'b0 ;
  assign n54412 = ( n4564 & ~n5422 ) | ( n4564 & n54411 ) | ( ~n5422 & n54411 ) ;
  assign n54413 = ( n6524 & n22611 ) | ( n6524 & ~n51348 ) | ( n22611 & ~n51348 ) ;
  assign n54414 = n54287 ^ n42191 ^ n306 ;
  assign n54415 = n34031 ^ n31181 ^ n14337 ;
  assign n54416 = n54415 ^ n11095 ^ 1'b0 ;
  assign n54421 = n2002 & ~n16805 ;
  assign n54422 = n39998 & n54421 ;
  assign n54418 = ~n1532 & n32779 ;
  assign n54419 = ( n4744 & ~n52283 ) | ( n4744 & n54418 ) | ( ~n52283 & n54418 ) ;
  assign n54417 = ( n9176 & n11210 ) | ( n9176 & n14190 ) | ( n11210 & n14190 ) ;
  assign n54420 = n54419 ^ n54417 ^ n1473 ;
  assign n54423 = n54422 ^ n54420 ^ n9859 ;
  assign n54424 = n51518 ^ n40897 ^ n8519 ;
  assign n54425 = ( n13032 & n14716 ) | ( n13032 & ~n54424 ) | ( n14716 & ~n54424 ) ;
  assign n54426 = ~n21127 & n41533 ;
  assign n54427 = n54426 ^ n32192 ^ 1'b0 ;
  assign n54428 = ( n24959 & n28456 ) | ( n24959 & n29609 ) | ( n28456 & n29609 ) ;
  assign n54429 = ~n20035 & n35408 ;
  assign n54430 = n54428 & n54429 ;
  assign n54431 = n46883 ^ n40508 ^ n13068 ;
  assign n54432 = n19602 ^ n13625 ^ n10716 ;
  assign n54433 = n54432 ^ n13712 ^ n4452 ;
  assign n54441 = n25336 ^ n24096 ^ 1'b0 ;
  assign n54435 = n2232 ^ x232 ^ 1'b0 ;
  assign n54436 = n2564 | n54435 ;
  assign n54437 = n54436 ^ n25185 ^ n509 ;
  assign n54438 = n54437 ^ n26877 ^ n22675 ;
  assign n54439 = n18583 ^ n11900 ^ n9444 ;
  assign n54440 = ( n10998 & ~n54438 ) | ( n10998 & n54439 ) | ( ~n54438 & n54439 ) ;
  assign n54434 = n39109 ^ n38458 ^ n18859 ;
  assign n54442 = n54441 ^ n54440 ^ n54434 ;
  assign n54443 = ( n2545 & ~n17396 ) | ( n2545 & n31048 ) | ( ~n17396 & n31048 ) ;
  assign n54444 = n16007 & ~n43016 ;
  assign n54445 = ( n24207 & n34538 ) | ( n24207 & ~n34579 ) | ( n34538 & ~n34579 ) ;
  assign n54446 = n40787 ^ n27444 ^ n7987 ;
  assign n54450 = ( n10139 & n15541 ) | ( n10139 & ~n40010 ) | ( n15541 & ~n40010 ) ;
  assign n54447 = n12476 & ~n24653 ;
  assign n54448 = n54447 ^ n19795 ^ 1'b0 ;
  assign n54449 = n54448 ^ n49264 ^ 1'b0 ;
  assign n54451 = n54450 ^ n54449 ^ n30387 ;
  assign n54453 = n29862 ^ n15666 ^ n2927 ;
  assign n54452 = ( n4017 & ~n4375 ) | ( n4017 & n51642 ) | ( ~n4375 & n51642 ) ;
  assign n54454 = n54453 ^ n54452 ^ n5997 ;
  assign n54455 = n33546 | n35934 ;
  assign n54456 = n54454 | n54455 ;
  assign n54457 = n25129 & n47600 ;
  assign n54458 = n11527 & n54457 ;
  assign n54459 = n52942 ^ n2468 ^ 1'b0 ;
  assign n54460 = n38280 | n54459 ;
  assign n54461 = n54460 ^ n35379 ^ n26250 ;
  assign n54462 = ( ~n4304 & n22324 ) | ( ~n4304 & n37661 ) | ( n22324 & n37661 ) ;
  assign n54463 = n54462 ^ n10390 ^ x231 ;
  assign n54464 = n39906 ^ n32688 ^ 1'b0 ;
  assign n54465 = n6625 & n54464 ;
  assign n54466 = ( n23471 & n51660 ) | ( n23471 & ~n54465 ) | ( n51660 & ~n54465 ) ;
  assign n54467 = n29290 ^ n20743 ^ n8611 ;
  assign n54468 = n30777 ^ n1043 ^ 1'b0 ;
  assign n54469 = n53381 ^ n14546 ^ n7563 ;
  assign n54470 = ( n28097 & ~n54468 ) | ( n28097 & n54469 ) | ( ~n54468 & n54469 ) ;
  assign n54471 = ( n9486 & n25221 ) | ( n9486 & ~n26097 ) | ( n25221 & ~n26097 ) ;
  assign n54472 = n45279 ^ n10938 ^ n4286 ;
  assign n54473 = ( ~n4582 & n27685 ) | ( ~n4582 & n54472 ) | ( n27685 & n54472 ) ;
  assign n54474 = ( n6132 & ~n10212 ) | ( n6132 & n18371 ) | ( ~n10212 & n18371 ) ;
  assign n54475 = n10038 ^ n4276 ^ 1'b0 ;
  assign n54476 = n47871 | n54475 ;
  assign n54477 = n21485 | n54476 ;
  assign n54478 = n32112 ^ n3464 ^ 1'b0 ;
  assign n54479 = n31671 & n54478 ;
  assign n54480 = n34119 ^ n16945 ^ n16172 ;
  assign n54481 = n54480 ^ n51787 ^ n41404 ;
  assign n54482 = ( n14423 & ~n20821 ) | ( n14423 & n39793 ) | ( ~n20821 & n39793 ) ;
  assign n54485 = n26590 ^ n20894 ^ 1'b0 ;
  assign n54483 = n11646 ^ n4420 ^ 1'b0 ;
  assign n54484 = ~n40655 & n54483 ;
  assign n54486 = n54485 ^ n54484 ^ n17199 ;
  assign n54487 = n38500 ^ n8342 ^ n263 ;
  assign n54488 = ( n7948 & n9610 ) | ( n7948 & ~n54487 ) | ( n9610 & ~n54487 ) ;
  assign n54489 = n990 & ~n23074 ;
  assign n54490 = n54489 ^ n24800 ^ 1'b0 ;
  assign n54491 = ( n11079 & ~n40364 ) | ( n11079 & n54490 ) | ( ~n40364 & n54490 ) ;
  assign n54492 = n46510 ^ n23993 ^ 1'b0 ;
  assign n54493 = ~n14197 & n15195 ;
  assign n54494 = n9375 & n54493 ;
  assign n54495 = ( n27428 & ~n54492 ) | ( n27428 & n54494 ) | ( ~n54492 & n54494 ) ;
  assign n54496 = ( ~n24101 & n38660 ) | ( ~n24101 & n49681 ) | ( n38660 & n49681 ) ;
  assign n54497 = ( ~n2396 & n9466 ) | ( ~n2396 & n10794 ) | ( n9466 & n10794 ) ;
  assign n54498 = n54497 ^ n38528 ^ n29300 ;
  assign n54499 = n26387 | n35684 ;
  assign n54500 = n54499 ^ n19327 ^ 1'b0 ;
  assign n54501 = ~n774 & n4471 ;
  assign n54502 = ~n8355 & n54501 ;
  assign n54503 = ( n3891 & ~n23064 ) | ( n3891 & n24756 ) | ( ~n23064 & n24756 ) ;
  assign n54504 = ( n20037 & ~n27978 ) | ( n20037 & n54503 ) | ( ~n27978 & n54503 ) ;
  assign n54505 = ( n17054 & ~n44885 ) | ( n17054 & n48522 ) | ( ~n44885 & n48522 ) ;
  assign n54506 = n54505 ^ n6358 ^ 1'b0 ;
  assign n54507 = n54504 & n54506 ;
  assign n54508 = ( ~n4583 & n11511 ) | ( ~n4583 & n12372 ) | ( n11511 & n12372 ) ;
  assign n54509 = ( ~n9075 & n19463 ) | ( ~n9075 & n54508 ) | ( n19463 & n54508 ) ;
  assign n54510 = ( ~n36244 & n39934 ) | ( ~n36244 & n54509 ) | ( n39934 & n54509 ) ;
  assign n54511 = ~n612 & n25227 ;
  assign n54512 = n47889 & n54511 ;
  assign n54513 = ( n1292 & n28355 ) | ( n1292 & ~n54512 ) | ( n28355 & ~n54512 ) ;
  assign n54514 = n47584 ^ n38767 ^ n38718 ;
  assign n54515 = n54514 ^ n51144 ^ n38477 ;
  assign n54516 = n27005 ^ n17939 ^ n7691 ;
  assign n54517 = n54516 ^ n28548 ^ n13186 ;
  assign n54518 = n27208 ^ n10203 ^ 1'b0 ;
  assign n54519 = ( n7043 & n13583 ) | ( n7043 & ~n19677 ) | ( n13583 & ~n19677 ) ;
  assign n54520 = ( n3419 & n15102 ) | ( n3419 & n15610 ) | ( n15102 & n15610 ) ;
  assign n54521 = ( n1601 & n33780 ) | ( n1601 & n44438 ) | ( n33780 & n44438 ) ;
  assign n54522 = n28909 ^ n19457 ^ 1'b0 ;
  assign n54523 = n17948 & n54522 ;
  assign n54524 = n7581 & ~n12411 ;
  assign n54525 = n31531 & n54524 ;
  assign n54526 = n5615 | n8378 ;
  assign n54527 = n54526 ^ n49571 ^ 1'b0 ;
  assign n54528 = ( n33676 & n42599 ) | ( n33676 & n48262 ) | ( n42599 & n48262 ) ;
  assign n54529 = ( n24826 & n34733 ) | ( n24826 & ~n54528 ) | ( n34733 & ~n54528 ) ;
  assign n54530 = n44240 ^ n18794 ^ n15192 ;
  assign n54531 = ( n3645 & n13051 ) | ( n3645 & ~n54530 ) | ( n13051 & ~n54530 ) ;
  assign n54532 = ( n852 & n15774 ) | ( n852 & ~n32171 ) | ( n15774 & ~n32171 ) ;
  assign n54534 = ~n7816 & n39115 ;
  assign n54535 = ( n11974 & ~n30469 ) | ( n11974 & n54534 ) | ( ~n30469 & n54534 ) ;
  assign n54533 = ( n12725 & n14768 ) | ( n12725 & n24650 ) | ( n14768 & n24650 ) ;
  assign n54536 = n54535 ^ n54533 ^ 1'b0 ;
  assign n54538 = n2148 & ~n16454 ;
  assign n54539 = n7972 & n54538 ;
  assign n54537 = n39926 ^ n5127 ^ 1'b0 ;
  assign n54540 = n54539 ^ n54537 ^ n4389 ;
  assign n54541 = ( ~n34369 & n45946 ) | ( ~n34369 & n49168 ) | ( n45946 & n49168 ) ;
  assign n54542 = n51980 ^ n11734 ^ 1'b0 ;
  assign n54543 = n3456 & n16859 ;
  assign n54544 = n22159 ^ n20672 ^ n11304 ;
  assign n54545 = n10544 & n45809 ;
  assign n54546 = ~n54544 & n54545 ;
  assign n54547 = ( n3412 & n5260 ) | ( n3412 & ~n16006 ) | ( n5260 & ~n16006 ) ;
  assign n54548 = ( n16454 & n36497 ) | ( n16454 & n54547 ) | ( n36497 & n54547 ) ;
  assign n54549 = ( ~n2476 & n8060 ) | ( ~n2476 & n46427 ) | ( n8060 & n46427 ) ;
  assign n54550 = n54549 ^ n31201 ^ n9509 ;
  assign n54551 = ( n49799 & ~n54548 ) | ( n49799 & n54550 ) | ( ~n54548 & n54550 ) ;
  assign n54552 = n36614 ^ n30197 ^ n16359 ;
  assign n54553 = n14665 ^ n4891 ^ n4104 ;
  assign n54554 = n54553 ^ n18027 ^ n592 ;
  assign n54555 = ~n16470 & n49641 ;
  assign n54556 = ( ~n5006 & n16527 ) | ( ~n5006 & n31117 ) | ( n16527 & n31117 ) ;
  assign n54557 = n54556 ^ n39592 ^ n4278 ;
  assign n54558 = n36218 ^ n25371 ^ n18039 ;
  assign n54559 = n51462 ^ n13320 ^ n7567 ;
  assign n54560 = ( ~x251 & n4238 ) | ( ~x251 & n19200 ) | ( n4238 & n19200 ) ;
  assign n54561 = ( n4713 & ~n7086 ) | ( n4713 & n54560 ) | ( ~n7086 & n54560 ) ;
  assign n54562 = n9252 ^ n5086 ^ n2446 ;
  assign n54563 = n9144 ^ n8077 ^ 1'b0 ;
  assign n54564 = n54562 | n54563 ;
  assign n54565 = n18603 ^ n417 ^ 1'b0 ;
  assign n54566 = n48008 & ~n54565 ;
  assign n54567 = ( n5739 & ~n17142 ) | ( n5739 & n29785 ) | ( ~n17142 & n29785 ) ;
  assign n54568 = ( n3332 & n7020 ) | ( n3332 & n14790 ) | ( n7020 & n14790 ) ;
  assign n54569 = n54568 ^ n26945 ^ n19777 ;
  assign n54570 = ~n11359 & n26562 ;
  assign n54571 = n21065 & n54570 ;
  assign n54572 = ( n54567 & n54569 ) | ( n54567 & n54571 ) | ( n54569 & n54571 ) ;
  assign n54573 = ( n37846 & n44901 ) | ( n37846 & n54572 ) | ( n44901 & n54572 ) ;
  assign n54574 = n6050 & ~n54573 ;
  assign n54575 = ( n8036 & n8307 ) | ( n8036 & n38273 ) | ( n8307 & n38273 ) ;
  assign n54576 = ( n29777 & n34530 ) | ( n29777 & ~n54575 ) | ( n34530 & ~n54575 ) ;
  assign n54577 = n34306 ^ n30994 ^ n11249 ;
  assign n54578 = ( n7634 & ~n12315 ) | ( n7634 & n54577 ) | ( ~n12315 & n54577 ) ;
  assign n54579 = ( ~n14676 & n54576 ) | ( ~n14676 & n54578 ) | ( n54576 & n54578 ) ;
  assign n54580 = ( n15575 & n16494 ) | ( n15575 & n27826 ) | ( n16494 & n27826 ) ;
  assign n54581 = ( n37151 & n46957 ) | ( n37151 & ~n54580 ) | ( n46957 & ~n54580 ) ;
  assign n54585 = n23867 ^ n4529 ^ 1'b0 ;
  assign n54586 = ~n29994 & n54585 ;
  assign n54582 = ( ~n10518 & n19315 ) | ( ~n10518 & n42093 ) | ( n19315 & n42093 ) ;
  assign n54583 = ( n705 & n29729 ) | ( n705 & ~n54582 ) | ( n29729 & ~n54582 ) ;
  assign n54584 = ( n12142 & ~n12307 ) | ( n12142 & n54583 ) | ( ~n12307 & n54583 ) ;
  assign n54587 = n54586 ^ n54584 ^ n36569 ;
  assign n54588 = ( n3206 & n32660 ) | ( n3206 & ~n34679 ) | ( n32660 & ~n34679 ) ;
  assign n54589 = n540 & n15853 ;
  assign n54590 = n54589 ^ n21861 ^ 1'b0 ;
  assign n54591 = ( n21047 & n54588 ) | ( n21047 & n54590 ) | ( n54588 & n54590 ) ;
  assign n54592 = n32232 | n34378 ;
  assign n54593 = n54592 ^ n27865 ^ n26611 ;
  assign n54594 = n7904 | n31198 ;
  assign n54595 = n34327 ^ n27725 ^ n14594 ;
  assign n54597 = n522 & n18754 ;
  assign n54598 = ~n32375 & n54597 ;
  assign n54596 = n22829 & n34627 ;
  assign n54599 = n54598 ^ n54596 ^ 1'b0 ;
  assign n54600 = ( ~n7641 & n22811 ) | ( ~n7641 & n23819 ) | ( n22811 & n23819 ) ;
  assign n54601 = n54600 ^ n39285 ^ n32874 ;
  assign n54603 = n2383 ^ n1693 ^ n949 ;
  assign n54602 = n46045 ^ n35702 ^ n11833 ;
  assign n54604 = n54603 ^ n54602 ^ n17879 ;
  assign n54605 = n19333 ^ n13083 ^ n2241 ;
  assign n54606 = ( ~n15565 & n16138 ) | ( ~n15565 & n54605 ) | ( n16138 & n54605 ) ;
  assign n54607 = n32243 ^ n17131 ^ n9970 ;
  assign n54608 = ( n23928 & n50733 ) | ( n23928 & n54607 ) | ( n50733 & n54607 ) ;
  assign n54609 = n2145 & n30760 ;
  assign n54610 = n43510 & n54609 ;
  assign n54611 = n54610 ^ n14420 ^ 1'b0 ;
  assign n54612 = ( n9014 & ~n25015 ) | ( n9014 & n38520 ) | ( ~n25015 & n38520 ) ;
  assign n54613 = n43670 ^ n32967 ^ n31041 ;
  assign n54618 = n14785 ^ n6269 ^ 1'b0 ;
  assign n54619 = n54618 ^ n25971 ^ n17266 ;
  assign n54614 = n3054 & n26400 ;
  assign n54615 = n14608 & n54614 ;
  assign n54616 = n6464 & ~n54615 ;
  assign n54617 = ~n7315 & n54616 ;
  assign n54620 = n54619 ^ n54617 ^ n44453 ;
  assign n54621 = n10879 & n49112 ;
  assign n54622 = n45449 & n54621 ;
  assign n54623 = n12116 ^ n9624 ^ n8787 ;
  assign n54624 = n54623 ^ n14898 ^ n2593 ;
  assign n54625 = n54624 ^ n24331 ^ 1'b0 ;
  assign n54626 = n19628 & n54625 ;
  assign n54627 = ~n25380 & n48514 ;
  assign n54628 = ( n6120 & n26200 ) | ( n6120 & ~n36971 ) | ( n26200 & ~n36971 ) ;
  assign n54629 = n51939 ^ n17142 ^ n10777 ;
  assign n54630 = n2108 | n9410 ;
  assign n54631 = n54630 ^ n48602 ^ n12730 ;
  assign n54632 = n47439 ^ n34975 ^ 1'b0 ;
  assign n54633 = n18322 ^ n16892 ^ n2620 ;
  assign n54634 = n52617 ^ n31359 ^ n7694 ;
  assign n54635 = n54634 ^ n33905 ^ n947 ;
  assign n54636 = ( n54632 & n54633 ) | ( n54632 & ~n54635 ) | ( n54633 & ~n54635 ) ;
  assign n54637 = n43134 ^ n39659 ^ n39076 ;
  assign n54638 = n48334 ^ n29274 ^ n27186 ;
  assign n54639 = n54638 ^ n47537 ^ n22002 ;
  assign n54640 = n54639 ^ n22569 ^ 1'b0 ;
  assign n54641 = ~n17424 & n41762 ;
  assign n54642 = n20955 ^ n15218 ^ n5261 ;
  assign n54643 = n54642 ^ n26029 ^ 1'b0 ;
  assign n54644 = ( n3968 & ~n4710 ) | ( n3968 & n54643 ) | ( ~n4710 & n54643 ) ;
  assign n54645 = n3996 & n54644 ;
  assign n54646 = ( ~n3363 & n7088 ) | ( ~n3363 & n48657 ) | ( n7088 & n48657 ) ;
  assign n54647 = n54646 ^ n667 ^ 1'b0 ;
  assign n54648 = n9097 & n54647 ;
  assign n54649 = n41944 ^ n32267 ^ 1'b0 ;
  assign n54650 = n40350 & n54649 ;
  assign n54651 = ( n11105 & n13918 ) | ( n11105 & ~n25639 ) | ( n13918 & ~n25639 ) ;
  assign n54652 = n54651 ^ n23808 ^ n21773 ;
  assign n54653 = n26501 ^ n8124 ^ n7676 ;
  assign n54654 = n54653 ^ n29066 ^ n8764 ;
  assign n54655 = n27485 ^ n23623 ^ n22018 ;
  assign n54656 = ( n11999 & n22805 ) | ( n11999 & n54655 ) | ( n22805 & n54655 ) ;
  assign n54657 = n54656 ^ n40685 ^ 1'b0 ;
  assign n54658 = ( n6063 & n53081 ) | ( n6063 & n54657 ) | ( n53081 & n54657 ) ;
  assign n54659 = ( ~n6712 & n9401 ) | ( ~n6712 & n10395 ) | ( n9401 & n10395 ) ;
  assign n54660 = n11478 & ~n41782 ;
  assign n54661 = n2211 & ~n44212 ;
  assign n54662 = n27468 & n54661 ;
  assign n54663 = n20603 & ~n45828 ;
  assign n54664 = n24683 & n54663 ;
  assign n54665 = n54664 ^ n46418 ^ 1'b0 ;
  assign n54666 = n34924 ^ n23360 ^ n14989 ;
  assign n54667 = n36014 ^ n27722 ^ n11334 ;
  assign n54668 = ~n3519 & n26374 ;
  assign n54669 = n36576 ^ n35038 ^ n983 ;
  assign n54670 = n11647 & ~n32380 ;
  assign n54671 = n15770 | n21298 ;
  assign n54673 = ( n7169 & ~n12190 ) | ( n7169 & n32742 ) | ( ~n12190 & n32742 ) ;
  assign n54672 = n33832 ^ n28294 ^ n3583 ;
  assign n54674 = n54673 ^ n54672 ^ n4704 ;
  assign n54675 = ( n5848 & n16841 ) | ( n5848 & ~n47983 ) | ( n16841 & ~n47983 ) ;
  assign n54677 = n36490 ^ n27263 ^ 1'b0 ;
  assign n54676 = n8712 | n45275 ;
  assign n54678 = n54677 ^ n54676 ^ 1'b0 ;
  assign n54679 = n54678 ^ n1549 ^ 1'b0 ;
  assign n54680 = ~n20055 & n54679 ;
  assign n54681 = n36443 ^ n30771 ^ 1'b0 ;
  assign n54682 = n18915 & n54681 ;
  assign n54683 = ( n9604 & ~n11719 ) | ( n9604 & n12964 ) | ( ~n11719 & n12964 ) ;
  assign n54684 = ( n5767 & n40281 ) | ( n5767 & ~n54683 ) | ( n40281 & ~n54683 ) ;
  assign n54685 = n43633 ^ n14199 ^ n5447 ;
  assign n54686 = n54685 ^ n33905 ^ 1'b0 ;
  assign n54687 = ( n2919 & ~n8477 ) | ( n2919 & n20139 ) | ( ~n8477 & n20139 ) ;
  assign n54688 = n42644 ^ n31562 ^ n16728 ;
  assign n54689 = n26738 ^ n7199 ^ n3847 ;
  assign n54690 = n54689 ^ n47536 ^ 1'b0 ;
  assign n54691 = n12585 ^ n3941 ^ 1'b0 ;
  assign n54692 = n54691 ^ n35366 ^ 1'b0 ;
  assign n54693 = ~n54690 & n54692 ;
  assign n54694 = ( ~n3738 & n54688 ) | ( ~n3738 & n54693 ) | ( n54688 & n54693 ) ;
  assign n54695 = ( n2559 & ~n41941 ) | ( n2559 & n54694 ) | ( ~n41941 & n54694 ) ;
  assign n54697 = ( ~n11970 & n25308 ) | ( ~n11970 & n28827 ) | ( n25308 & n28827 ) ;
  assign n54696 = ( n11924 & ~n21511 ) | ( n11924 & n40949 ) | ( ~n21511 & n40949 ) ;
  assign n54698 = n54697 ^ n54696 ^ n7940 ;
  assign n54699 = ( n8534 & n17078 ) | ( n8534 & ~n41223 ) | ( n17078 & ~n41223 ) ;
  assign n54700 = n54699 ^ n24055 ^ n20807 ;
  assign n54701 = ( ~n16776 & n20968 ) | ( ~n16776 & n47114 ) | ( n20968 & n47114 ) ;
  assign n54702 = n19165 ^ n271 ^ 1'b0 ;
  assign n54703 = n17886 & ~n54702 ;
  assign n54705 = n30826 & ~n49273 ;
  assign n54704 = ~n551 & n32980 ;
  assign n54706 = n54705 ^ n54704 ^ 1'b0 ;
  assign n54707 = ~n9239 & n40759 ;
  assign n54708 = ~n11760 & n54707 ;
  assign n54709 = n26405 & ~n54708 ;
  assign n54710 = n54709 ^ n37956 ^ 1'b0 ;
  assign n54711 = ( n11246 & n12891 ) | ( n11246 & n50352 ) | ( n12891 & n50352 ) ;
  assign n54712 = n54711 ^ n24564 ^ n6536 ;
  assign n54713 = n54712 ^ n37165 ^ 1'b0 ;
  assign n54714 = n844 | n11345 ;
  assign n54715 = n54714 ^ n13505 ^ 1'b0 ;
  assign n54716 = ( n1369 & n41402 ) | ( n1369 & n54715 ) | ( n41402 & n54715 ) ;
  assign n54717 = ( n34231 & n34493 ) | ( n34231 & n46567 ) | ( n34493 & n46567 ) ;
  assign n54718 = ( n3094 & n20118 ) | ( n3094 & ~n36188 ) | ( n20118 & ~n36188 ) ;
  assign n54719 = ~n31076 & n35904 ;
  assign n54720 = n6909 | n54719 ;
  assign n54721 = n54720 ^ n2665 ^ 1'b0 ;
  assign n54722 = n54721 ^ n52898 ^ n38369 ;
  assign n54723 = n14186 ^ n1514 ^ 1'b0 ;
  assign n54724 = ( ~n4832 & n15455 ) | ( ~n4832 & n54723 ) | ( n15455 & n54723 ) ;
  assign n54725 = n27432 ^ n13512 ^ 1'b0 ;
  assign n54726 = n17958 | n31259 ;
  assign n54727 = n54726 ^ n11207 ^ 1'b0 ;
  assign n54728 = ~n2423 & n50872 ;
  assign n54729 = n54728 ^ n48887 ^ 1'b0 ;
  assign n54730 = ( n8227 & n19376 ) | ( n8227 & ~n21154 ) | ( n19376 & ~n21154 ) ;
  assign n54731 = n47799 ^ n33232 ^ n4563 ;
  assign n54732 = n34999 ^ n14572 ^ n10909 ;
  assign n54733 = ( n16101 & ~n47781 ) | ( n16101 & n48004 ) | ( ~n47781 & n48004 ) ;
  assign n54734 = ( n13745 & ~n20616 ) | ( n13745 & n38643 ) | ( ~n20616 & n38643 ) ;
  assign n54735 = ( n4778 & n43470 ) | ( n4778 & n44710 ) | ( n43470 & n44710 ) ;
  assign n54738 = n43255 ^ n27875 ^ n2210 ;
  assign n54736 = n22642 ^ n8188 ^ n5855 ;
  assign n54737 = n54736 ^ n9194 ^ 1'b0 ;
  assign n54739 = n54738 ^ n54737 ^ n8652 ;
  assign n54740 = n51163 ^ n36943 ^ n4317 ;
  assign n54741 = n32689 ^ n5615 ^ 1'b0 ;
  assign n54742 = n52199 | n54741 ;
  assign n54743 = n8599 & ~n54742 ;
  assign n54744 = n54743 ^ n42429 ^ 1'b0 ;
  assign n54745 = n34206 ^ n26531 ^ n8256 ;
  assign n54746 = ~n24789 & n54745 ;
  assign n54747 = n54746 ^ n11101 ^ 1'b0 ;
  assign n54748 = n4320 ^ n1492 ^ 1'b0 ;
  assign n54749 = n15893 & ~n23558 ;
  assign n54750 = ~n13355 & n16708 ;
  assign n54751 = n54750 ^ n8740 ^ 1'b0 ;
  assign n54752 = ( n50684 & n50735 ) | ( n50684 & n54751 ) | ( n50735 & n54751 ) ;
  assign n54753 = ( ~n54748 & n54749 ) | ( ~n54748 & n54752 ) | ( n54749 & n54752 ) ;
  assign n54754 = n48276 ^ n17687 ^ n9421 ;
  assign n54755 = ( n2602 & n3008 ) | ( n2602 & n16623 ) | ( n3008 & n16623 ) ;
  assign n54756 = ~n7989 & n13225 ;
  assign n54757 = ( n41161 & ~n54553 ) | ( n41161 & n54756 ) | ( ~n54553 & n54756 ) ;
  assign n54758 = n41990 ^ n25549 ^ n783 ;
  assign n54759 = n34398 ^ n26168 ^ n2944 ;
  assign n54760 = ~n8973 & n20139 ;
  assign n54761 = n54760 ^ n41083 ^ 1'b0 ;
  assign n54762 = ( n38636 & ~n47027 ) | ( n38636 & n54761 ) | ( ~n47027 & n54761 ) ;
  assign n54763 = ( n17073 & ~n23072 ) | ( n17073 & n31462 ) | ( ~n23072 & n31462 ) ;
  assign n54764 = n23110 & ~n47559 ;
  assign n54765 = n47537 & n54764 ;
  assign n54766 = n8756 & n53538 ;
  assign n54767 = n54765 & n54766 ;
  assign n54768 = n49561 ^ n27378 ^ n23328 ;
  assign n54769 = n10666 ^ n6122 ^ 1'b0 ;
  assign n54770 = n7468 & ~n54769 ;
  assign n54771 = ( n34910 & n41437 ) | ( n34910 & n54770 ) | ( n41437 & n54770 ) ;
  assign n54772 = n54771 ^ n39536 ^ n28870 ;
  assign n54773 = ( ~n6365 & n54768 ) | ( ~n6365 & n54772 ) | ( n54768 & n54772 ) ;
  assign n54774 = ( n6483 & ~n21298 ) | ( n6483 & n50024 ) | ( ~n21298 & n50024 ) ;
  assign n54775 = n29623 ^ n27024 ^ 1'b0 ;
  assign n54776 = n30707 & n54775 ;
  assign n54777 = ( n9051 & n18689 ) | ( n9051 & n54776 ) | ( n18689 & n54776 ) ;
  assign n54778 = n35757 ^ n29982 ^ n8115 ;
  assign n54779 = ( n2376 & ~n11984 ) | ( n2376 & n35687 ) | ( ~n11984 & n35687 ) ;
  assign n54781 = x160 & n36889 ;
  assign n54782 = n54781 ^ n5413 ^ 1'b0 ;
  assign n54780 = n4163 & ~n31187 ;
  assign n54783 = n54782 ^ n54780 ^ n10703 ;
  assign n54784 = ( n5010 & n10646 ) | ( n5010 & ~n24551 ) | ( n10646 & ~n24551 ) ;
  assign n54785 = n54784 ^ n23907 ^ n7947 ;
  assign n54786 = n54785 ^ n32700 ^ n19264 ;
  assign n54787 = n46619 ^ n7710 ^ n7285 ;
  assign n54788 = n15259 ^ n4677 ^ 1'b0 ;
  assign n54789 = n4110 & n54788 ;
  assign n54790 = n337 & n11256 ;
  assign n54791 = ~n54789 & n54790 ;
  assign n54792 = n10175 | n49475 ;
  assign n54793 = n54792 ^ n44195 ^ 1'b0 ;
  assign n54794 = ~n52210 & n54793 ;
  assign n54795 = n54794 ^ n9262 ^ 1'b0 ;
  assign n54796 = ( n7781 & ~n10469 ) | ( n7781 & n42490 ) | ( ~n10469 & n42490 ) ;
  assign n54797 = n54796 ^ n8408 ^ 1'b0 ;
  assign n54798 = n49643 & ~n54797 ;
  assign n54799 = n10697 | n43544 ;
  assign n54800 = n24619 ^ n9085 ^ n6721 ;
  assign n54801 = n32245 ^ n24468 ^ n1310 ;
  assign n54802 = n2276 ^ n954 ^ 1'b0 ;
  assign n54803 = ( n9931 & n31619 ) | ( n9931 & ~n54802 ) | ( n31619 & ~n54802 ) ;
  assign n54804 = n31723 ^ n19689 ^ 1'b0 ;
  assign n54805 = n44398 & ~n54804 ;
  assign n54806 = ( n7816 & ~n43699 ) | ( n7816 & n54805 ) | ( ~n43699 & n54805 ) ;
  assign n54807 = ( n3812 & n47418 ) | ( n3812 & ~n54806 ) | ( n47418 & ~n54806 ) ;
  assign n54808 = n34207 ^ n17190 ^ n6566 ;
  assign n54809 = n3642 & n12246 ;
  assign n54810 = ( n920 & n17459 ) | ( n920 & n17869 ) | ( n17459 & n17869 ) ;
  assign n54811 = ( n15819 & ~n47882 ) | ( n15819 & n54810 ) | ( ~n47882 & n54810 ) ;
  assign n54812 = n48387 ^ n19749 ^ 1'b0 ;
  assign n54820 = ( n5315 & n35701 ) | ( n5315 & ~n40983 ) | ( n35701 & ~n40983 ) ;
  assign n54821 = n54820 ^ n14966 ^ n4557 ;
  assign n54818 = ~n19689 & n38712 ;
  assign n54819 = n54818 ^ n7509 ^ 1'b0 ;
  assign n54813 = n17867 ^ n8595 ^ n6514 ;
  assign n54814 = n7664 | n8603 ;
  assign n54815 = n1078 & ~n54814 ;
  assign n54816 = ( n7694 & n49273 ) | ( n7694 & n54815 ) | ( n49273 & n54815 ) ;
  assign n54817 = ( n14913 & ~n54813 ) | ( n14913 & n54816 ) | ( ~n54813 & n54816 ) ;
  assign n54822 = n54821 ^ n54819 ^ n54817 ;
  assign n54823 = n45215 ^ n32648 ^ n24814 ;
  assign n54824 = n44606 ^ n2727 ^ 1'b0 ;
  assign n54825 = n10647 & ~n54824 ;
  assign n54826 = ( ~n2704 & n12243 ) | ( ~n2704 & n54825 ) | ( n12243 & n54825 ) ;
  assign n54827 = n54826 ^ n35633 ^ n7545 ;
  assign n54828 = ( n7983 & n10947 ) | ( n7983 & ~n35824 ) | ( n10947 & ~n35824 ) ;
  assign n54829 = ( n5201 & n51916 ) | ( n5201 & n54828 ) | ( n51916 & n54828 ) ;
  assign n54830 = n13068 ^ n7445 ^ 1'b0 ;
  assign n54831 = n12702 & n54830 ;
  assign n54832 = n54831 ^ n12956 ^ 1'b0 ;
  assign n54833 = ( n6330 & n47323 ) | ( n6330 & n54056 ) | ( n47323 & n54056 ) ;
  assign n54834 = n27777 ^ n12620 ^ 1'b0 ;
  assign n54835 = n54834 ^ n21042 ^ 1'b0 ;
  assign n54836 = n36447 ^ n17110 ^ n7473 ;
  assign n54837 = ~n5480 & n54836 ;
  assign n54838 = n9104 & n54837 ;
  assign n54840 = n19629 | n40500 ;
  assign n54839 = n5000 | n36219 ;
  assign n54841 = n54840 ^ n54839 ^ 1'b0 ;
  assign n54842 = ~n14106 & n27051 ;
  assign n54843 = n54842 ^ n18652 ^ 1'b0 ;
  assign n54844 = n54843 ^ n23582 ^ n4092 ;
  assign n54845 = n5114 ^ n1609 ^ n1369 ;
  assign n54846 = n29807 ^ x175 ^ 1'b0 ;
  assign n54847 = ( n25961 & ~n54845 ) | ( n25961 & n54846 ) | ( ~n54845 & n54846 ) ;
  assign n54848 = n3420 | n54847 ;
  assign n54849 = n54844 | n54848 ;
  assign n54850 = ( n2371 & ~n6710 ) | ( n2371 & n26647 ) | ( ~n6710 & n26647 ) ;
  assign n54851 = ~n11249 & n21786 ;
  assign n54852 = n47234 ^ n46826 ^ n34836 ;
  assign n54853 = ( ~n11690 & n22413 ) | ( ~n11690 & n33094 ) | ( n22413 & n33094 ) ;
  assign n54854 = n46246 ^ n33330 ^ 1'b0 ;
  assign n54855 = ( n9384 & n54853 ) | ( n9384 & ~n54854 ) | ( n54853 & ~n54854 ) ;
  assign n54856 = ~n7922 & n29952 ;
  assign n54857 = n44143 ^ n26920 ^ n16367 ;
  assign n54858 = ( n9826 & n10131 ) | ( n9826 & n53618 ) | ( n10131 & n53618 ) ;
  assign n54859 = n44239 ^ n31203 ^ 1'b0 ;
  assign n54860 = ( ~n4859 & n54858 ) | ( ~n4859 & n54859 ) | ( n54858 & n54859 ) ;
  assign n54861 = ( ~n4028 & n5183 ) | ( ~n4028 & n10713 ) | ( n5183 & n10713 ) ;
  assign n54862 = ( n16281 & n42463 ) | ( n16281 & ~n54861 ) | ( n42463 & ~n54861 ) ;
  assign n54863 = n15391 & n54862 ;
  assign n54864 = n53361 ^ n21009 ^ 1'b0 ;
  assign n54865 = ~n54863 & n54864 ;
  assign n54866 = n6353 ^ n1046 ^ 1'b0 ;
  assign n54867 = n21050 & ~n54866 ;
  assign n54868 = ( ~n1666 & n20455 ) | ( ~n1666 & n23415 ) | ( n20455 & n23415 ) ;
  assign n54869 = ( n31793 & n39441 ) | ( n31793 & n54868 ) | ( n39441 & n54868 ) ;
  assign n54870 = ( n16349 & n28812 ) | ( n16349 & ~n47417 ) | ( n28812 & ~n47417 ) ;
  assign n54871 = n52288 ^ n35834 ^ n21718 ;
  assign n54872 = n9678 & n54871 ;
  assign n54873 = n41278 ^ n25538 ^ n14712 ;
  assign n54874 = n39504 ^ n23530 ^ n10221 ;
  assign n54875 = ( n37606 & n54873 ) | ( n37606 & ~n54874 ) | ( n54873 & ~n54874 ) ;
  assign n54876 = ( ~n13459 & n25613 ) | ( ~n13459 & n54875 ) | ( n25613 & n54875 ) ;
  assign n54877 = n2187 & ~n47368 ;
  assign n54878 = n54877 ^ n11168 ^ 1'b0 ;
  assign n54879 = n54878 ^ n39421 ^ n423 ;
  assign n54880 = n42087 ^ n38630 ^ n11513 ;
  assign n54881 = ( n11392 & n16627 ) | ( n11392 & ~n24521 ) | ( n16627 & ~n24521 ) ;
  assign n54882 = n54881 ^ n51498 ^ n1756 ;
  assign n54883 = ( n18396 & n20015 ) | ( n18396 & n54882 ) | ( n20015 & n54882 ) ;
  assign n54884 = n30906 ^ n24339 ^ n17975 ;
  assign n54885 = n47384 ^ n13669 ^ n5057 ;
  assign n54886 = ( n25581 & n28735 ) | ( n25581 & ~n54885 ) | ( n28735 & ~n54885 ) ;
  assign n54887 = n23585 ^ n2341 ^ 1'b0 ;
  assign n54888 = n54886 | n54887 ;
  assign n54889 = ~n9644 & n19037 ;
  assign n54890 = n54889 ^ n13190 ^ 1'b0 ;
  assign n54891 = ( ~n1414 & n4436 ) | ( ~n1414 & n48806 ) | ( n4436 & n48806 ) ;
  assign n54892 = n39676 & n54891 ;
  assign n54893 = n54892 ^ n1085 ^ 1'b0 ;
  assign n54894 = n2909 & ~n32584 ;
  assign n54895 = ( n23280 & n41843 ) | ( n23280 & ~n54894 ) | ( n41843 & ~n54894 ) ;
  assign n54896 = n37628 ^ n24786 ^ n13003 ;
  assign n54897 = ( n5361 & n18449 ) | ( n5361 & n51597 ) | ( n18449 & n51597 ) ;
  assign n54898 = ( n6381 & ~n6442 ) | ( n6381 & n11841 ) | ( ~n6442 & n11841 ) ;
  assign n54899 = n2156 & ~n12496 ;
  assign n54900 = ( n11264 & n12313 ) | ( n11264 & n54899 ) | ( n12313 & n54899 ) ;
  assign n54901 = n15852 ^ n1549 ^ 1'b0 ;
  assign n54902 = n54901 ^ n47140 ^ n34639 ;
  assign n54903 = ( n17639 & n24667 ) | ( n17639 & ~n28785 ) | ( n24667 & ~n28785 ) ;
  assign n54904 = n8997 & n14915 ;
  assign n54905 = x27 & ~n54904 ;
  assign n54906 = n9451 & n54905 ;
  assign n54907 = n54514 ^ n49586 ^ n3039 ;
  assign n54908 = n40031 & n42115 ;
  assign n54909 = n25074 ^ n14381 ^ n12951 ;
  assign n54910 = n13441 & n26004 ;
  assign n54911 = n4242 & n54910 ;
  assign n54912 = n54911 ^ n42622 ^ n4272 ;
  assign n54913 = n25556 ^ n17683 ^ n2585 ;
  assign n54914 = ( n16194 & ~n45374 ) | ( n16194 & n54913 ) | ( ~n45374 & n54913 ) ;
  assign n54915 = n49245 ^ n42317 ^ n7170 ;
  assign n54916 = n46812 ^ n19081 ^ 1'b0 ;
  assign n54917 = n1080 | n17803 ;
  assign n54918 = n44171 | n54917 ;
  assign n54919 = ( n9598 & n31297 ) | ( n9598 & ~n32956 ) | ( n31297 & ~n32956 ) ;
  assign n54920 = n41990 ^ n35420 ^ 1'b0 ;
  assign n54921 = n46118 ^ n9273 ^ n8268 ;
  assign n54922 = ( ~n54919 & n54920 ) | ( ~n54919 & n54921 ) | ( n54920 & n54921 ) ;
  assign n54923 = n54922 ^ n31802 ^ n28180 ;
  assign n54924 = ( n1619 & ~n11465 ) | ( n1619 & n43072 ) | ( ~n11465 & n43072 ) ;
  assign n54925 = n54924 ^ n40982 ^ n24729 ;
  assign n54926 = ( n8766 & ~n23074 ) | ( n8766 & n33947 ) | ( ~n23074 & n33947 ) ;
  assign n54927 = ( x243 & n9920 ) | ( x243 & n54926 ) | ( n9920 & n54926 ) ;
  assign n54928 = n54927 ^ n13297 ^ n6329 ;
  assign n54929 = ( n14183 & n24654 ) | ( n14183 & n39085 ) | ( n24654 & n39085 ) ;
  assign n54930 = ( n17778 & n21433 ) | ( n17778 & n29715 ) | ( n21433 & n29715 ) ;
  assign n54931 = ( n6472 & n37107 ) | ( n6472 & ~n54930 ) | ( n37107 & ~n54930 ) ;
  assign n54932 = n54931 ^ n21381 ^ 1'b0 ;
  assign n54937 = n7748 & n13114 ;
  assign n54934 = n24144 ^ n21113 ^ n2275 ;
  assign n54933 = n9588 & ~n47326 ;
  assign n54935 = n54934 ^ n54933 ^ 1'b0 ;
  assign n54936 = n54935 ^ n8348 ^ 1'b0 ;
  assign n54938 = n54937 ^ n54936 ^ n44198 ;
  assign n54939 = n54938 ^ n41851 ^ 1'b0 ;
  assign n54940 = ( n27497 & n44070 ) | ( n27497 & n54939 ) | ( n44070 & n54939 ) ;
  assign n54941 = ( ~n6290 & n12566 ) | ( ~n6290 & n19887 ) | ( n12566 & n19887 ) ;
  assign n54942 = n54941 ^ n34192 ^ x152 ;
  assign n54943 = ( n11365 & ~n22633 ) | ( n11365 & n54942 ) | ( ~n22633 & n54942 ) ;
  assign n54944 = ( n1657 & n11314 ) | ( n1657 & ~n17707 ) | ( n11314 & ~n17707 ) ;
  assign n54945 = n54944 ^ n54009 ^ n23677 ;
  assign n54946 = n42588 ^ n20894 ^ n4938 ;
  assign n54947 = ( n3183 & n6997 ) | ( n3183 & ~n19887 ) | ( n6997 & ~n19887 ) ;
  assign n54948 = n54947 ^ n22356 ^ 1'b0 ;
  assign n54949 = n54946 | n54948 ;
  assign n54950 = n29979 ^ n2631 ^ 1'b0 ;
  assign n54951 = n4946 & ~n54950 ;
  assign n54952 = ( n4525 & n11859 ) | ( n4525 & ~n17844 ) | ( n11859 & ~n17844 ) ;
  assign n54953 = n4554 | n7080 ;
  assign n54954 = n54953 ^ n7747 ^ x94 ;
  assign n54955 = n15364 ^ n10904 ^ 1'b0 ;
  assign n54956 = ~n54954 & n54955 ;
  assign n54957 = ( n24968 & n54952 ) | ( n24968 & ~n54956 ) | ( n54952 & ~n54956 ) ;
  assign n54958 = n25456 ^ n18891 ^ n7584 ;
  assign n54959 = ( n15725 & n50211 ) | ( n15725 & ~n54958 ) | ( n50211 & ~n54958 ) ;
  assign n54960 = ( n6394 & n22377 ) | ( n6394 & ~n54959 ) | ( n22377 & ~n54959 ) ;
  assign n54961 = n54960 ^ n46802 ^ n24066 ;
  assign n54962 = n41567 ^ n21262 ^ n17139 ;
  assign n54963 = n15554 & ~n30528 ;
  assign n54964 = n48869 ^ n39112 ^ n2325 ;
  assign n54965 = ( n45225 & n54963 ) | ( n45225 & ~n54964 ) | ( n54963 & ~n54964 ) ;
  assign n54966 = ( ~n13460 & n16254 ) | ( ~n13460 & n54965 ) | ( n16254 & n54965 ) ;
  assign n54967 = ( n6118 & ~n28726 ) | ( n6118 & n40962 ) | ( ~n28726 & n40962 ) ;
  assign n54968 = ( n6476 & n40947 ) | ( n6476 & n45829 ) | ( n40947 & n45829 ) ;
  assign n54969 = n34990 ^ n23720 ^ n7284 ;
  assign n54970 = n523 & n54969 ;
  assign n54971 = ( n835 & n3969 ) | ( n835 & n14949 ) | ( n3969 & n14949 ) ;
  assign n54972 = ( ~n30562 & n54970 ) | ( ~n30562 & n54971 ) | ( n54970 & n54971 ) ;
  assign n54973 = ( n4840 & ~n25789 ) | ( n4840 & n40090 ) | ( ~n25789 & n40090 ) ;
  assign n54974 = ( n38500 & ~n53538 ) | ( n38500 & n54973 ) | ( ~n53538 & n54973 ) ;
  assign n54975 = ~n11700 & n39820 ;
  assign n54976 = n54975 ^ n40428 ^ 1'b0 ;
  assign n54977 = ( n12755 & n14034 ) | ( n12755 & ~n48321 ) | ( n14034 & ~n48321 ) ;
  assign n54978 = n46371 ^ n39259 ^ n10232 ;
  assign n54979 = ~n17541 & n31715 ;
  assign n54980 = n54979 ^ n13545 ^ 1'b0 ;
  assign n54981 = n54980 ^ n33645 ^ n16762 ;
  assign n54982 = ( n3372 & ~n5828 ) | ( n3372 & n29847 ) | ( ~n5828 & n29847 ) ;
  assign n54983 = ( n4938 & n40906 ) | ( n4938 & ~n54982 ) | ( n40906 & ~n54982 ) ;
  assign n54984 = n33711 ^ n33372 ^ n24879 ;
  assign n54985 = ( ~n9450 & n31444 ) | ( ~n9450 & n35620 ) | ( n31444 & n35620 ) ;
  assign n54986 = n8207 ^ n2716 ^ 1'b0 ;
  assign n54987 = ( n8795 & n9683 ) | ( n8795 & ~n54986 ) | ( n9683 & ~n54986 ) ;
  assign n54988 = ( ~x243 & n18237 ) | ( ~x243 & n49699 ) | ( n18237 & n49699 ) ;
  assign n54989 = ( n4840 & n6710 ) | ( n4840 & ~n29020 ) | ( n6710 & ~n29020 ) ;
  assign n54990 = ( ~n8107 & n54988 ) | ( ~n8107 & n54989 ) | ( n54988 & n54989 ) ;
  assign n54991 = n32224 ^ n13057 ^ 1'b0 ;
  assign n54992 = ~n20545 & n54991 ;
  assign n54993 = n5420 & n38434 ;
  assign n54994 = ~n14458 & n54993 ;
  assign n54995 = ( ~n27201 & n50043 ) | ( ~n27201 & n54994 ) | ( n50043 & n54994 ) ;
  assign n54996 = ( n810 & ~n24411 ) | ( n810 & n27136 ) | ( ~n24411 & n27136 ) ;
  assign n54997 = ( n6037 & ~n45044 ) | ( n6037 & n51361 ) | ( ~n45044 & n51361 ) ;
  assign n54998 = ( x136 & ~n5014 ) | ( x136 & n38772 ) | ( ~n5014 & n38772 ) ;
  assign n54999 = n25655 | n50846 ;
  assign n55000 = n54999 ^ n29254 ^ 1'b0 ;
  assign n55001 = n28347 ^ n20805 ^ n13054 ;
  assign n55002 = n21095 ^ n17144 ^ n9848 ;
  assign n55003 = ( ~n26764 & n34160 ) | ( ~n26764 & n40585 ) | ( n34160 & n40585 ) ;
  assign n55005 = n1050 & n30693 ;
  assign n55006 = n55005 ^ n26411 ^ n557 ;
  assign n55004 = ( n11669 & n39964 ) | ( n11669 & n47728 ) | ( n39964 & n47728 ) ;
  assign n55007 = n55006 ^ n55004 ^ n25105 ;
  assign n55008 = n55007 ^ n25960 ^ 1'b0 ;
  assign n55011 = n22846 ^ n18348 ^ n6905 ;
  assign n55012 = ( n3366 & n31159 ) | ( n3366 & n55011 ) | ( n31159 & n55011 ) ;
  assign n55009 = n30987 ^ n3578 ^ 1'b0 ;
  assign n55010 = ( n5324 & n45293 ) | ( n5324 & n55009 ) | ( n45293 & n55009 ) ;
  assign n55013 = n55012 ^ n55010 ^ n27935 ;
  assign n55014 = n46898 ^ n2204 ^ n1134 ;
  assign n55015 = n55014 ^ n36354 ^ 1'b0 ;
  assign n55016 = n55015 ^ n2557 ^ 1'b0 ;
  assign n55017 = ( ~n50305 & n53711 ) | ( ~n50305 & n54109 ) | ( n53711 & n54109 ) ;
  assign n55018 = n11074 ^ n4614 ^ x3 ;
  assign n55019 = ( n2542 & n23931 ) | ( n2542 & n55018 ) | ( n23931 & n55018 ) ;
  assign n55021 = n39829 ^ n27419 ^ n8068 ;
  assign n55020 = n4324 & n11949 ;
  assign n55022 = n55021 ^ n55020 ^ n38680 ;
  assign n55023 = n40856 ^ n31942 ^ n19307 ;
  assign n55024 = n15008 ^ n10322 ^ 1'b0 ;
  assign n55025 = n55024 ^ n30550 ^ n315 ;
  assign n55026 = ( n986 & n55023 ) | ( n986 & n55025 ) | ( n55023 & n55025 ) ;
  assign n55027 = n2783 & ~n41945 ;
  assign n55028 = ( n3321 & n32064 ) | ( n3321 & ~n55027 ) | ( n32064 & ~n55027 ) ;
  assign n55029 = ( n1008 & n17356 ) | ( n1008 & n20066 ) | ( n17356 & n20066 ) ;
  assign n55030 = ~n25774 & n52560 ;
  assign n55031 = n55029 & n55030 ;
  assign n55032 = n44872 ^ n34864 ^ 1'b0 ;
  assign n55033 = ~n55031 & n55032 ;
  assign n55034 = n44222 ^ n530 ^ 1'b0 ;
  assign n55035 = ( n22089 & n55033 ) | ( n22089 & ~n55034 ) | ( n55033 & ~n55034 ) ;
  assign n55036 = n55035 ^ n26803 ^ 1'b0 ;
  assign n55037 = ~n8610 & n12587 ;
  assign n55038 = n55037 ^ n21268 ^ 1'b0 ;
  assign n55039 = ( n11722 & n16136 ) | ( n11722 & ~n29790 ) | ( n16136 & ~n29790 ) ;
  assign n55040 = ( x235 & ~n12139 ) | ( x235 & n12907 ) | ( ~n12139 & n12907 ) ;
  assign n55041 = ~n8411 & n55040 ;
  assign n55042 = n55041 ^ n18525 ^ 1'b0 ;
  assign n55043 = ( n8399 & n40710 ) | ( n8399 & n55042 ) | ( n40710 & n55042 ) ;
  assign n55044 = ( n15995 & n37553 ) | ( n15995 & ~n55043 ) | ( n37553 & ~n55043 ) ;
  assign n55045 = ( n55038 & ~n55039 ) | ( n55038 & n55044 ) | ( ~n55039 & n55044 ) ;
  assign n55046 = n55045 ^ n11218 ^ 1'b0 ;
  assign n55047 = ~n54638 & n55046 ;
  assign n55049 = ( n20163 & n26521 ) | ( n20163 & ~n49413 ) | ( n26521 & ~n49413 ) ;
  assign n55048 = n8913 & ~n28401 ;
  assign n55050 = n55049 ^ n55048 ^ 1'b0 ;
  assign n55051 = n4798 | n19875 ;
  assign n55052 = ( ~n822 & n15528 ) | ( ~n822 & n48901 ) | ( n15528 & n48901 ) ;
  assign n55053 = ~n24400 & n55052 ;
  assign n55054 = n54133 ^ n49810 ^ 1'b0 ;
  assign n55055 = n2538 & ~n55054 ;
  assign n55056 = n55055 ^ n36665 ^ n33092 ;
  assign n55057 = ( n17052 & n40636 ) | ( n17052 & ~n55056 ) | ( n40636 & ~n55056 ) ;
  assign n55058 = ( x11 & n7215 ) | ( x11 & ~n7440 ) | ( n7215 & ~n7440 ) ;
  assign n55059 = n55058 ^ n34329 ^ n11197 ;
  assign n55060 = ~n9954 & n25257 ;
  assign n55061 = n55059 & n55060 ;
  assign n55062 = n46350 ^ n39091 ^ n25701 ;
  assign n55063 = n55062 ^ n13984 ^ n5708 ;
  assign n55064 = ( n1240 & ~n55061 ) | ( n1240 & n55063 ) | ( ~n55061 & n55063 ) ;
  assign n55065 = ( n13756 & n25459 ) | ( n13756 & n43646 ) | ( n25459 & n43646 ) ;
  assign n55066 = n55065 ^ n44598 ^ n36717 ;
  assign n55067 = n51292 ^ n25529 ^ n18451 ;
  assign n55068 = n6426 & n25815 ;
  assign n55069 = n55068 ^ n9036 ^ 1'b0 ;
  assign n55070 = ( n9750 & ~n28421 ) | ( n9750 & n28729 ) | ( ~n28421 & n28729 ) ;
  assign n55071 = ( n7062 & n55069 ) | ( n7062 & ~n55070 ) | ( n55069 & ~n55070 ) ;
  assign n55072 = n20900 ^ n18716 ^ 1'b0 ;
  assign n55073 = n25617 | n55072 ;
  assign n55074 = ( ~n17344 & n20872 ) | ( ~n17344 & n45576 ) | ( n20872 & n45576 ) ;
  assign n55075 = ( n5698 & ~n55073 ) | ( n5698 & n55074 ) | ( ~n55073 & n55074 ) ;
  assign n55076 = ( n3259 & ~n5927 ) | ( n3259 & n13264 ) | ( ~n5927 & n13264 ) ;
  assign n55077 = ~n34369 & n55076 ;
  assign n55078 = n43418 ^ n40090 ^ n19208 ;
  assign n55079 = ( n8826 & ~n54820 ) | ( n8826 & n55078 ) | ( ~n54820 & n55078 ) ;
  assign n55080 = n29507 | n55079 ;
  assign n55081 = n26186 | n55080 ;
  assign n55082 = n43929 ^ n42377 ^ n20534 ;
  assign n55083 = n46306 ^ n36198 ^ 1'b0 ;
  assign n55084 = n21067 & n55083 ;
  assign n55085 = n55084 ^ n37357 ^ 1'b0 ;
  assign n55086 = ( ~n1756 & n30050 ) | ( ~n1756 & n55085 ) | ( n30050 & n55085 ) ;
  assign n55087 = n7845 | n11659 ;
  assign n55088 = n55087 ^ n37746 ^ 1'b0 ;
  assign n55089 = n17629 & ~n33117 ;
  assign n55090 = x245 & ~n23159 ;
  assign n55091 = n55089 & n55090 ;
  assign n55092 = n55091 ^ n31430 ^ n29274 ;
  assign n55093 = ( n9521 & n9752 ) | ( n9521 & n23062 ) | ( n9752 & n23062 ) ;
  assign n55094 = n33476 ^ n28285 ^ n23524 ;
  assign n55095 = n20558 ^ n15662 ^ 1'b0 ;
  assign n55097 = n32724 ^ n8267 ^ n2432 ;
  assign n55098 = ( ~n21436 & n28133 ) | ( ~n21436 & n55097 ) | ( n28133 & n55097 ) ;
  assign n55096 = n19321 ^ n14310 ^ n10222 ;
  assign n55099 = n55098 ^ n55096 ^ n7563 ;
  assign n55100 = n55099 ^ n41684 ^ n1604 ;
  assign n55102 = n36209 ^ n32653 ^ x14 ;
  assign n55101 = n44457 & n51624 ;
  assign n55103 = n55102 ^ n55101 ^ 1'b0 ;
  assign n55104 = ( n7349 & n10710 ) | ( n7349 & n15287 ) | ( n10710 & n15287 ) ;
  assign n55105 = n41541 | n55104 ;
  assign n55106 = n3570 | n49771 ;
  assign n55107 = n42750 ^ n7634 ^ 1'b0 ;
  assign n55108 = ( n1962 & n18594 ) | ( n1962 & n28608 ) | ( n18594 & n28608 ) ;
  assign n55109 = ( n19507 & n23650 ) | ( n19507 & n41737 ) | ( n23650 & n41737 ) ;
  assign n55110 = ( n3613 & ~n21855 ) | ( n3613 & n49440 ) | ( ~n21855 & n49440 ) ;
  assign n55113 = n41682 ^ n27744 ^ n19593 ;
  assign n55111 = n15582 ^ n13122 ^ n7153 ;
  assign n55112 = ( n30957 & ~n45188 ) | ( n30957 & n55111 ) | ( ~n45188 & n55111 ) ;
  assign n55114 = n55113 ^ n55112 ^ n40901 ;
  assign n55115 = n38224 ^ n32973 ^ n21437 ;
  assign n55116 = n39533 ^ n32083 ^ n1243 ;
  assign n55117 = n46048 ^ n1967 ^ 1'b0 ;
  assign n55118 = ~n6390 & n55117 ;
  assign n55119 = n34243 ^ n956 ^ 1'b0 ;
  assign n55120 = n2974 | n55119 ;
  assign n55121 = n44035 & ~n55120 ;
  assign n55122 = n53386 ^ n2162 ^ 1'b0 ;
  assign n55123 = n55121 & ~n55122 ;
  assign n55124 = n32564 ^ n3413 ^ 1'b0 ;
  assign n55125 = n26884 & n55124 ;
  assign n55126 = n43692 ^ n21578 ^ n13360 ;
  assign n55127 = ( n20049 & ~n22891 ) | ( n20049 & n55126 ) | ( ~n22891 & n55126 ) ;
  assign n55128 = n16206 & ~n37781 ;
  assign n55129 = ( ~n3491 & n55127 ) | ( ~n3491 & n55128 ) | ( n55127 & n55128 ) ;
  assign n55130 = x100 & n12411 ;
  assign n55131 = ( n13639 & n14757 ) | ( n13639 & n27978 ) | ( n14757 & n27978 ) ;
  assign n55132 = ( n23763 & n34474 ) | ( n23763 & ~n50025 ) | ( n34474 & ~n50025 ) ;
  assign n55133 = n32606 ^ n25112 ^ n23506 ;
  assign n55134 = n50634 ^ n37508 ^ n15972 ;
  assign n55135 = n32886 ^ n15182 ^ 1'b0 ;
  assign n55136 = n55134 | n55135 ;
  assign n55137 = n55136 ^ n40293 ^ n689 ;
  assign n55138 = ( n8730 & ~n20649 ) | ( n8730 & n41322 ) | ( ~n20649 & n41322 ) ;
  assign n55139 = n6148 & ~n55138 ;
  assign n55140 = n42983 ^ n39043 ^ n17916 ;
  assign n55141 = n45371 ^ n4570 ^ 1'b0 ;
  assign n55142 = n498 & ~n55141 ;
  assign n55143 = n28100 ^ n14948 ^ 1'b0 ;
  assign n55144 = n38932 & n55143 ;
  assign n55145 = ~n19362 & n32038 ;
  assign n55146 = ( n2216 & n52014 ) | ( n2216 & n55145 ) | ( n52014 & n55145 ) ;
  assign n55147 = ( x10 & ~n11055 ) | ( x10 & n13580 ) | ( ~n11055 & n13580 ) ;
  assign n55148 = n55147 ^ n18749 ^ n1784 ;
  assign n55149 = n42599 ^ n12188 ^ 1'b0 ;
  assign n55150 = n14405 & n22016 ;
  assign n55151 = n25699 & n55150 ;
  assign n55152 = n55151 ^ n24555 ^ n11740 ;
  assign n55153 = n13891 & n22704 ;
  assign n55154 = ~n8031 & n55153 ;
  assign n55155 = ( ~n12794 & n42463 ) | ( ~n12794 & n55154 ) | ( n42463 & n55154 ) ;
  assign n55156 = ( n18122 & n25140 ) | ( n18122 & ~n55155 ) | ( n25140 & ~n55155 ) ;
  assign n55157 = n37212 ^ n20753 ^ n16768 ;
  assign n55158 = n30062 ^ n25837 ^ n1647 ;
  assign n55159 = n53219 ^ n9054 ^ 1'b0 ;
  assign n55160 = ( n8700 & ~n55158 ) | ( n8700 & n55159 ) | ( ~n55158 & n55159 ) ;
  assign n55161 = ( n55156 & n55157 ) | ( n55156 & ~n55160 ) | ( n55157 & ~n55160 ) ;
  assign n55162 = n31547 ^ n11860 ^ 1'b0 ;
  assign n55163 = n25709 ^ n21425 ^ n11579 ;
  assign n55164 = n32534 ^ n28784 ^ 1'b0 ;
  assign n55165 = n7696 & ~n18972 ;
  assign n55166 = n55165 ^ n3746 ^ 1'b0 ;
  assign n55167 = n46011 ^ n23926 ^ n10502 ;
  assign n55168 = n8166 & ~n55167 ;
  assign n55169 = ~n15972 & n55168 ;
  assign n55170 = n30521 ^ n15000 ^ 1'b0 ;
  assign n55171 = n4454 | n55170 ;
  assign n55172 = n2902 & ~n55171 ;
  assign n55173 = n55172 ^ n2402 ^ 1'b0 ;
  assign n55174 = n31821 ^ n9212 ^ n4204 ;
  assign n55175 = ( n22898 & ~n45611 ) | ( n22898 & n55174 ) | ( ~n45611 & n55174 ) ;
  assign n55176 = n4332 | n18145 ;
  assign n55177 = n55176 ^ n19582 ^ 1'b0 ;
  assign n55178 = n42472 ^ n28679 ^ n9586 ;
  assign n55179 = ( ~n3810 & n39829 ) | ( ~n3810 & n55178 ) | ( n39829 & n55178 ) ;
  assign n55180 = ( n6261 & n55177 ) | ( n6261 & ~n55179 ) | ( n55177 & ~n55179 ) ;
  assign n55181 = n23180 ^ n8751 ^ 1'b0 ;
  assign n55182 = ( n21288 & n40089 ) | ( n21288 & ~n55181 ) | ( n40089 & ~n55181 ) ;
  assign n55183 = ( ~n17778 & n23931 ) | ( ~n17778 & n45664 ) | ( n23931 & n45664 ) ;
  assign n55184 = ( n558 & n33134 ) | ( n558 & n55183 ) | ( n33134 & n55183 ) ;
  assign n55185 = n55184 ^ n45990 ^ n23128 ;
  assign n55186 = n27681 ^ n23757 ^ n793 ;
  assign n55187 = n55186 ^ n29855 ^ n4381 ;
  assign n55188 = n31387 ^ n27657 ^ n20526 ;
  assign n55189 = n49625 ^ n41990 ^ n30064 ;
  assign n55190 = n55188 & n55189 ;
  assign n55191 = ~n1254 & n20832 ;
  assign n55192 = n15656 & n55191 ;
  assign n55193 = ( ~n1790 & n23474 ) | ( ~n1790 & n25814 ) | ( n23474 & n25814 ) ;
  assign n55194 = n55193 ^ n22158 ^ n15421 ;
  assign n55195 = ( n1211 & n55192 ) | ( n1211 & ~n55194 ) | ( n55192 & ~n55194 ) ;
  assign n55196 = n19799 ^ n18271 ^ n4406 ;
  assign n55197 = ( n7315 & ~n16882 ) | ( n7315 & n43971 ) | ( ~n16882 & n43971 ) ;
  assign n55198 = n5777 & n9672 ;
  assign n55199 = ~n55197 & n55198 ;
  assign n55200 = n24488 | n28281 ;
  assign n55201 = n54999 | n55200 ;
  assign n55202 = n42984 ^ n10445 ^ n5658 ;
  assign n55203 = n55202 ^ n13303 ^ 1'b0 ;
  assign n55204 = ~n46264 & n55203 ;
  assign n55205 = n19263 & ~n28114 ;
  assign n55206 = ( n26267 & ~n31742 ) | ( n26267 & n55205 ) | ( ~n31742 & n55205 ) ;
  assign n55207 = n31756 ^ n31170 ^ n23895 ;
  assign n55208 = ( n18192 & n31855 ) | ( n18192 & n32462 ) | ( n31855 & n32462 ) ;
  assign n55210 = ( n8553 & ~n23306 ) | ( n8553 & n49329 ) | ( ~n23306 & n49329 ) ;
  assign n55209 = n40473 ^ n23401 ^ n6995 ;
  assign n55211 = n55210 ^ n55209 ^ n55069 ;
  assign n55212 = ( ~n26948 & n31931 ) | ( ~n26948 & n40705 ) | ( n31931 & n40705 ) ;
  assign n55213 = ~n49449 & n55212 ;
  assign n55214 = ( ~n5756 & n36031 ) | ( ~n5756 & n55213 ) | ( n36031 & n55213 ) ;
  assign n55215 = n32005 ^ n15258 ^ n3851 ;
  assign n55216 = ( ~n16180 & n19609 ) | ( ~n16180 & n27595 ) | ( n19609 & n27595 ) ;
  assign n55217 = n55216 ^ n28053 ^ n15552 ;
  assign n55218 = ( n2245 & n40435 ) | ( n2245 & ~n55217 ) | ( n40435 & ~n55217 ) ;
  assign n55219 = ( n13719 & n30870 ) | ( n13719 & ~n55218 ) | ( n30870 & ~n55218 ) ;
  assign n55220 = ( n1411 & n9876 ) | ( n1411 & ~n55219 ) | ( n9876 & ~n55219 ) ;
  assign n55221 = ~n882 & n21785 ;
  assign n55222 = n55221 ^ n12879 ^ 1'b0 ;
  assign n55223 = ( n18616 & n35470 ) | ( n18616 & n55222 ) | ( n35470 & n55222 ) ;
  assign n55224 = n55223 ^ n35651 ^ n26278 ;
  assign n55225 = ( n24908 & n36259 ) | ( n24908 & n55224 ) | ( n36259 & n55224 ) ;
  assign n55226 = n38653 & n52384 ;
  assign n55227 = n55226 ^ n2746 ^ 1'b0 ;
  assign n55228 = n11726 & n40634 ;
  assign n55229 = n55228 ^ n38225 ^ 1'b0 ;
  assign n55231 = n46484 ^ n39593 ^ n17907 ;
  assign n55230 = ( n8941 & n12146 ) | ( n8941 & n31997 ) | ( n12146 & n31997 ) ;
  assign n55232 = n55231 ^ n55230 ^ n45630 ;
  assign n55233 = n18137 & n31979 ;
  assign n55234 = ( n7097 & n12413 ) | ( n7097 & n55233 ) | ( n12413 & n55233 ) ;
  assign n55235 = ( n13947 & n16399 ) | ( n13947 & n40069 ) | ( n16399 & n40069 ) ;
  assign n55236 = ( n24507 & ~n29830 ) | ( n24507 & n44560 ) | ( ~n29830 & n44560 ) ;
  assign n55237 = n43213 ^ n40797 ^ 1'b0 ;
  assign n55238 = n50465 ^ n7768 ^ x15 ;
  assign n55239 = ( n7619 & n53619 ) | ( n7619 & ~n55238 ) | ( n53619 & ~n55238 ) ;
  assign n55241 = n28254 ^ n13904 ^ n5267 ;
  assign n55240 = n33235 ^ n28618 ^ 1'b0 ;
  assign n55242 = n55241 ^ n55240 ^ n5374 ;
  assign n55243 = ~n24921 & n53333 ;
  assign n55244 = ( n8475 & n16222 ) | ( n8475 & ~n55243 ) | ( n16222 & ~n55243 ) ;
  assign n55245 = n6261 ^ n5592 ^ 1'b0 ;
  assign n55246 = ~n13158 & n52539 ;
  assign n55247 = n24708 ^ n439 ^ 1'b0 ;
  assign n55248 = n55247 ^ n35704 ^ n15419 ;
  assign n55249 = n23476 ^ n10475 ^ 1'b0 ;
  assign n55250 = ~n34953 & n55249 ;
  assign n55251 = n35006 ^ n22873 ^ n8650 ;
  assign n55252 = ( n18484 & n51988 ) | ( n18484 & n55251 ) | ( n51988 & n55251 ) ;
  assign n55253 = n55250 & n55252 ;
  assign n55254 = ( ~n2592 & n20354 ) | ( ~n2592 & n23273 ) | ( n20354 & n23273 ) ;
  assign n55255 = n55254 ^ n48572 ^ n36531 ;
  assign n55256 = ( n22065 & n23478 ) | ( n22065 & n53703 ) | ( n23478 & n53703 ) ;
  assign n55257 = ( n8491 & n17873 ) | ( n8491 & n51076 ) | ( n17873 & n51076 ) ;
  assign n55258 = n36609 ^ n28531 ^ n9777 ;
  assign n55259 = n55258 ^ n11539 ^ n8504 ;
  assign n55260 = ( n2080 & ~n4841 ) | ( n2080 & n55259 ) | ( ~n4841 & n55259 ) ;
  assign n55263 = n37254 ^ n29343 ^ 1'b0 ;
  assign n55261 = n51654 ^ n12314 ^ n4209 ;
  assign n55262 = n55261 ^ n16882 ^ n5980 ;
  assign n55264 = n55263 ^ n55262 ^ n1126 ;
  assign n55268 = ( n9382 & n11134 ) | ( n9382 & n17424 ) | ( n11134 & n17424 ) ;
  assign n55266 = n22724 | n24623 ;
  assign n55267 = n55266 ^ n5189 ^ 1'b0 ;
  assign n55265 = n50391 ^ n7523 ^ n3451 ;
  assign n55269 = n55268 ^ n55267 ^ n55265 ;
  assign n55270 = ~n49046 & n55269 ;
  assign n55271 = n16066 & n35087 ;
  assign n55272 = n55271 ^ n8565 ^ 1'b0 ;
  assign n55273 = n27306 ^ n13023 ^ 1'b0 ;
  assign n55274 = n45202 | n55273 ;
  assign n55275 = ~n16638 & n51840 ;
  assign n55276 = n3401 & n55275 ;
  assign n55277 = ( n5226 & n7241 ) | ( n5226 & n11004 ) | ( n7241 & n11004 ) ;
  assign n55278 = ( n559 & ~n13676 ) | ( n559 & n40495 ) | ( ~n13676 & n40495 ) ;
  assign n55279 = ( n32700 & n55277 ) | ( n32700 & ~n55278 ) | ( n55277 & ~n55278 ) ;
  assign n55281 = n33760 ^ n32705 ^ n6010 ;
  assign n55280 = ( n7065 & ~n17527 ) | ( n7065 & n17757 ) | ( ~n17527 & n17757 ) ;
  assign n55282 = n55281 ^ n55280 ^ n1056 ;
  assign n55283 = n55282 ^ n20012 ^ n17722 ;
  assign n55284 = ( n5692 & n9277 ) | ( n5692 & ~n23444 ) | ( n9277 & ~n23444 ) ;
  assign n55285 = n55284 ^ n42550 ^ n29260 ;
  assign n55286 = n9829 | n34596 ;
  assign n55287 = n41657 ^ n16950 ^ n4365 ;
  assign n55288 = n29147 ^ n17405 ^ 1'b0 ;
  assign n55289 = ( ~n7956 & n21062 ) | ( ~n7956 & n52624 ) | ( n21062 & n52624 ) ;
  assign n55290 = ( n20794 & n21213 ) | ( n20794 & ~n54280 ) | ( n21213 & ~n54280 ) ;
  assign n55291 = n12800 & n14377 ;
  assign n55292 = n55291 ^ n35194 ^ 1'b0 ;
  assign n55293 = n40534 ^ n5856 ^ 1'b0 ;
  assign n55294 = n23772 & n55293 ;
  assign n55295 = n54770 ^ n29737 ^ 1'b0 ;
  assign n55296 = ( ~n18124 & n41207 ) | ( ~n18124 & n55295 ) | ( n41207 & n55295 ) ;
  assign n55297 = n34903 ^ n10629 ^ 1'b0 ;
  assign n55298 = n10532 | n29078 ;
  assign n55299 = ( n45400 & ~n55297 ) | ( n45400 & n55298 ) | ( ~n55297 & n55298 ) ;
  assign n55300 = ( n11809 & n41879 ) | ( n11809 & ~n49639 ) | ( n41879 & ~n49639 ) ;
  assign n55302 = n23740 & n23890 ;
  assign n55303 = n55302 ^ n11836 ^ 1'b0 ;
  assign n55304 = n1122 & ~n55303 ;
  assign n55305 = ~n8224 & n55304 ;
  assign n55306 = n55305 ^ n50778 ^ n9633 ;
  assign n55301 = ( n14546 & n19333 ) | ( n14546 & n34665 ) | ( n19333 & n34665 ) ;
  assign n55307 = n55306 ^ n55301 ^ n16667 ;
  assign n55308 = n50545 ^ n29027 ^ n1128 ;
  assign n55313 = ~n30086 & n35227 ;
  assign n55309 = n1790 & n6421 ;
  assign n55310 = ~n39837 & n55309 ;
  assign n55311 = ( n19024 & n20295 ) | ( n19024 & ~n55310 ) | ( n20295 & ~n55310 ) ;
  assign n55312 = n55311 ^ n5800 ^ n1371 ;
  assign n55314 = n55313 ^ n55312 ^ n16072 ;
  assign n55315 = ( n2800 & n8631 ) | ( n2800 & n12725 ) | ( n8631 & n12725 ) ;
  assign n55316 = n55315 ^ n23582 ^ n5286 ;
  assign n55317 = ( n12109 & n21562 ) | ( n12109 & n42801 ) | ( n21562 & n42801 ) ;
  assign n55318 = n55317 ^ n49342 ^ 1'b0 ;
  assign n55319 = ( n16793 & n20265 ) | ( n16793 & n55318 ) | ( n20265 & n55318 ) ;
  assign n55320 = n26886 ^ n8407 ^ 1'b0 ;
  assign n55321 = ~n7145 & n55320 ;
  assign n55322 = ~n11560 & n15303 ;
  assign n55323 = ~n55321 & n55322 ;
  assign n55324 = n41030 ^ n14266 ^ n1723 ;
  assign n55325 = n55324 ^ n28954 ^ 1'b0 ;
  assign n55326 = n3093 | n55325 ;
  assign n55327 = n21789 ^ n4177 ^ 1'b0 ;
  assign n55328 = n22297 & n37888 ;
  assign n55329 = n55328 ^ n9311 ^ 1'b0 ;
  assign n55330 = n55329 ^ n37746 ^ n16076 ;
  assign n55331 = ( n22987 & n47719 ) | ( n22987 & ~n55330 ) | ( n47719 & ~n55330 ) ;
  assign n55332 = n11607 & ~n13437 ;
  assign n55333 = n55332 ^ n9426 ^ 1'b0 ;
  assign n55334 = n47524 ^ n18233 ^ n15088 ;
  assign n55335 = ( n8919 & n55333 ) | ( n8919 & n55334 ) | ( n55333 & n55334 ) ;
  assign n55337 = ~n2777 & n12718 ;
  assign n55338 = n55337 ^ n6218 ^ 1'b0 ;
  assign n55339 = ( ~n5761 & n9454 ) | ( ~n5761 & n35543 ) | ( n9454 & n35543 ) ;
  assign n55340 = ( n31755 & ~n55338 ) | ( n31755 & n55339 ) | ( ~n55338 & n55339 ) ;
  assign n55336 = ( n10406 & n11135 ) | ( n10406 & ~n48572 ) | ( n11135 & ~n48572 ) ;
  assign n55341 = n55340 ^ n55336 ^ n28414 ;
  assign n55342 = ( n6069 & ~n15153 ) | ( n6069 & n49264 ) | ( ~n15153 & n49264 ) ;
  assign n55343 = ( n37079 & ~n43756 ) | ( n37079 & n55342 ) | ( ~n43756 & n55342 ) ;
  assign n55344 = ( n7947 & ~n11443 ) | ( n7947 & n39707 ) | ( ~n11443 & n39707 ) ;
  assign n55345 = ( ~n6524 & n11952 ) | ( ~n6524 & n40013 ) | ( n11952 & n40013 ) ;
  assign n55346 = ~n14506 & n26022 ;
  assign n55347 = ( n2751 & n22278 ) | ( n2751 & n54861 ) | ( n22278 & n54861 ) ;
  assign n55348 = n33327 & ~n55347 ;
  assign n55349 = ~n9438 & n35815 ;
  assign n55350 = n23643 & n55349 ;
  assign n55352 = n43146 ^ n28638 ^ 1'b0 ;
  assign n55353 = n44972 | n55352 ;
  assign n55351 = n842 | n15451 ;
  assign n55354 = n55353 ^ n55351 ^ 1'b0 ;
  assign n55355 = n30793 ^ n19534 ^ 1'b0 ;
  assign n55356 = ~n16992 & n55355 ;
  assign n55361 = n6555 & n13110 ;
  assign n55357 = n40309 ^ n4528 ^ 1'b0 ;
  assign n55358 = ~n34558 & n55357 ;
  assign n55359 = n39851 ^ n8907 ^ 1'b0 ;
  assign n55360 = ( n37722 & n55358 ) | ( n37722 & ~n55359 ) | ( n55358 & ~n55359 ) ;
  assign n55362 = n55361 ^ n55360 ^ n5244 ;
  assign n55363 = ( ~n856 & n35873 ) | ( ~n856 & n51109 ) | ( n35873 & n51109 ) ;
  assign n55364 = n49930 ^ n47403 ^ n43285 ;
  assign n55365 = n51743 ^ n24100 ^ n19147 ;
  assign n55366 = ( ~n11364 & n29734 ) | ( ~n11364 & n55365 ) | ( n29734 & n55365 ) ;
  assign n55367 = ( ~n19190 & n43055 ) | ( ~n19190 & n55366 ) | ( n43055 & n55366 ) ;
  assign n55368 = ( n8840 & ~n25158 ) | ( n8840 & n42478 ) | ( ~n25158 & n42478 ) ;
  assign n55369 = ( n2422 & n6328 ) | ( n2422 & ~n49749 ) | ( n6328 & ~n49749 ) ;
  assign n55370 = n32534 & n52131 ;
  assign n55371 = ( n4685 & ~n17097 ) | ( n4685 & n29807 ) | ( ~n17097 & n29807 ) ;
  assign n55372 = ( n28742 & ~n49045 ) | ( n28742 & n55371 ) | ( ~n49045 & n55371 ) ;
  assign n55373 = ( n11337 & ~n12085 ) | ( n11337 & n12910 ) | ( ~n12085 & n12910 ) ;
  assign n55374 = n50621 ^ n47501 ^ 1'b0 ;
  assign n55375 = n55373 & n55374 ;
  assign n55376 = n23539 & ~n28345 ;
  assign n55377 = n2177 & n55376 ;
  assign n55378 = n6364 & ~n27410 ;
  assign n55379 = ~n1508 & n18614 ;
  assign n55380 = n55378 & n55379 ;
  assign n55381 = n50353 ^ n49315 ^ n2276 ;
  assign n55382 = n23024 ^ n12398 ^ n8663 ;
  assign n55383 = ( n29198 & ~n41293 ) | ( n29198 & n55382 ) | ( ~n41293 & n55382 ) ;
  assign n55384 = ( n6274 & ~n43904 ) | ( n6274 & n46380 ) | ( ~n43904 & n46380 ) ;
  assign n55385 = n32003 ^ n23354 ^ n2081 ;
  assign n55386 = ( n10837 & n48370 ) | ( n10837 & n55385 ) | ( n48370 & n55385 ) ;
  assign n55387 = n45019 ^ n8700 ^ 1'b0 ;
  assign n55388 = n5660 | n31818 ;
  assign n55389 = n55388 ^ n16450 ^ n14022 ;
  assign n55390 = ( ~n4924 & n11373 ) | ( ~n4924 & n24344 ) | ( n11373 & n24344 ) ;
  assign n55391 = n28352 ^ n16348 ^ 1'b0 ;
  assign n55392 = ( n7071 & ~n55390 ) | ( n7071 & n55391 ) | ( ~n55390 & n55391 ) ;
  assign n55393 = ( n13847 & n50709 ) | ( n13847 & ~n55392 ) | ( n50709 & ~n55392 ) ;
  assign n55394 = n1270 | n4956 ;
  assign n55395 = n55394 ^ n31039 ^ 1'b0 ;
  assign n55396 = ( n1792 & n34195 ) | ( n1792 & n42023 ) | ( n34195 & n42023 ) ;
  assign n55397 = n55396 ^ n51274 ^ n17229 ;
  assign n55398 = n55397 ^ n50612 ^ n10268 ;
  assign n55399 = n30565 ^ n21570 ^ n3229 ;
  assign n55400 = n26003 ^ n22929 ^ n18312 ;
  assign n55401 = ~n41986 & n55400 ;
  assign n55402 = n12507 | n16780 ;
  assign n55403 = n55402 ^ n7512 ^ 1'b0 ;
  assign n55404 = n55403 ^ n5028 ^ n745 ;
  assign n55405 = ( n8222 & n16327 ) | ( n8222 & ~n48821 ) | ( n16327 & ~n48821 ) ;
  assign n55406 = n55405 ^ n19895 ^ n14503 ;
  assign n55407 = ( n24642 & n55404 ) | ( n24642 & ~n55406 ) | ( n55404 & ~n55406 ) ;
  assign n55408 = n47499 ^ n26778 ^ n18306 ;
  assign n55409 = n9629 & ~n16667 ;
  assign n55410 = n46579 ^ n2838 ^ 1'b0 ;
  assign n55411 = n55410 ^ n43487 ^ n39716 ;
  assign n55412 = ( n16320 & ~n22795 ) | ( n16320 & n55411 ) | ( ~n22795 & n55411 ) ;
  assign n55413 = ( n34048 & n34949 ) | ( n34048 & ~n47813 ) | ( n34949 & ~n47813 ) ;
  assign n55414 = n24827 ^ n4333 ^ 1'b0 ;
  assign n55415 = ~n31979 & n55414 ;
  assign n55416 = n23157 ^ n4968 ^ n4877 ;
  assign n55417 = ( n2710 & ~n34704 ) | ( n2710 & n55416 ) | ( ~n34704 & n55416 ) ;
  assign n55418 = n51959 ^ n40655 ^ 1'b0 ;
  assign n55420 = ( n6952 & n21842 ) | ( n6952 & ~n26321 ) | ( n21842 & ~n26321 ) ;
  assign n55419 = n12496 & n41497 ;
  assign n55421 = n55420 ^ n55419 ^ n16848 ;
  assign n55422 = ( n15509 & n34131 ) | ( n15509 & ~n55421 ) | ( n34131 & ~n55421 ) ;
  assign n55423 = n55422 ^ n20333 ^ x203 ;
  assign n55425 = n45308 ^ n11111 ^ n3910 ;
  assign n55424 = ( n19641 & n22778 ) | ( n19641 & n30178 ) | ( n22778 & n30178 ) ;
  assign n55426 = n55425 ^ n55424 ^ n17284 ;
  assign n55427 = ~n40797 & n48891 ;
  assign n55428 = ( n21052 & n25829 ) | ( n21052 & n55427 ) | ( n25829 & n55427 ) ;
  assign n55430 = n26183 ^ n2647 ^ 1'b0 ;
  assign n55429 = ~n2729 & n22107 ;
  assign n55431 = n55430 ^ n55429 ^ n32568 ;
  assign n55432 = n1357 & n28595 ;
  assign n55433 = ( n21315 & n22003 ) | ( n21315 & n55432 ) | ( n22003 & n55432 ) ;
  assign n55434 = ( ~n16486 & n28730 ) | ( ~n16486 & n34508 ) | ( n28730 & n34508 ) ;
  assign n55435 = n42898 ^ n12138 ^ n11501 ;
  assign n55436 = ( ~n1508 & n17257 ) | ( ~n1508 & n55435 ) | ( n17257 & n55435 ) ;
  assign n55437 = n55436 ^ n13550 ^ 1'b0 ;
  assign n55438 = n23987 & n55437 ;
  assign n55439 = n7903 ^ n5171 ^ 1'b0 ;
  assign n55440 = n16928 & n55439 ;
  assign n55441 = n26488 ^ n13308 ^ 1'b0 ;
  assign n55442 = ~n7561 & n23662 ;
  assign n55443 = n15630 & n55442 ;
  assign n55444 = n55443 ^ n33658 ^ n33088 ;
  assign n55445 = n1827 ^ n1238 ^ 1'b0 ;
  assign n55446 = n49524 | n55445 ;
  assign n55447 = n39649 ^ n29299 ^ n1877 ;
  assign n55448 = ( n17869 & n50528 ) | ( n17869 & n55447 ) | ( n50528 & n55447 ) ;
  assign n55450 = n23518 ^ n20778 ^ n6279 ;
  assign n55451 = n55450 ^ n14533 ^ n6167 ;
  assign n55449 = ( ~n7430 & n16405 ) | ( ~n7430 & n39389 ) | ( n16405 & n39389 ) ;
  assign n55452 = n55451 ^ n55449 ^ n37788 ;
  assign n55453 = n49977 ^ n18051 ^ n11495 ;
  assign n55454 = ( ~n13824 & n42703 ) | ( ~n13824 & n55453 ) | ( n42703 & n55453 ) ;
  assign n55455 = n55454 ^ n25609 ^ 1'b0 ;
  assign n55456 = ( n37864 & ~n40021 ) | ( n37864 & n45106 ) | ( ~n40021 & n45106 ) ;
  assign n55457 = ( n24177 & n33185 ) | ( n24177 & n55456 ) | ( n33185 & n55456 ) ;
  assign n55458 = n12261 & n14541 ;
  assign n55459 = n55458 ^ n6632 ^ 1'b0 ;
  assign n55460 = ~n10509 & n11322 ;
  assign n55461 = n55460 ^ n15159 ^ 1'b0 ;
  assign n55462 = ( x153 & ~n6670 ) | ( x153 & n8497 ) | ( ~n6670 & n8497 ) ;
  assign n55463 = ( n2892 & n8678 ) | ( n2892 & ~n55462 ) | ( n8678 & ~n55462 ) ;
  assign n55464 = n8462 ^ n3719 ^ 1'b0 ;
  assign n55465 = n55464 ^ n27796 ^ n10086 ;
  assign n55466 = ( ~n2368 & n16589 ) | ( ~n2368 & n55465 ) | ( n16589 & n55465 ) ;
  assign n55467 = ( n16129 & n55463 ) | ( n16129 & ~n55466 ) | ( n55463 & ~n55466 ) ;
  assign n55468 = ( ~n3612 & n51827 ) | ( ~n3612 & n55396 ) | ( n51827 & n55396 ) ;
  assign n55469 = n12780 ^ n3958 ^ n830 ;
  assign n55470 = n12194 | n55469 ;
  assign n55471 = n55470 ^ n42125 ^ 1'b0 ;
  assign n55472 = n55471 ^ n8240 ^ n3866 ;
  assign n55473 = n31737 ^ n4143 ^ 1'b0 ;
  assign n55474 = n55473 ^ n53262 ^ n2026 ;
  assign n55475 = ( ~n13912 & n28480 ) | ( ~n13912 & n44642 ) | ( n28480 & n44642 ) ;
  assign n55477 = ~n22443 & n25563 ;
  assign n55478 = n55477 ^ n25680 ^ 1'b0 ;
  assign n55476 = ( ~n9094 & n21756 ) | ( ~n9094 & n32064 ) | ( n21756 & n32064 ) ;
  assign n55479 = n55478 ^ n55476 ^ n11381 ;
  assign n55480 = n8154 & ~n16135 ;
  assign n55481 = n55480 ^ n12062 ^ 1'b0 ;
  assign n55482 = ( n9904 & n14078 ) | ( n9904 & n55481 ) | ( n14078 & n55481 ) ;
  assign n55486 = n18822 ^ n3614 ^ n3144 ;
  assign n55484 = ~n36596 & n37824 ;
  assign n55485 = n55484 ^ n29064 ^ 1'b0 ;
  assign n55483 = n39620 ^ n16507 ^ n5365 ;
  assign n55487 = n55486 ^ n55485 ^ n55483 ;
  assign n55488 = n12934 & n30214 ;
  assign n55489 = n55488 ^ n4315 ^ 1'b0 ;
  assign n55490 = ~n3512 & n16034 ;
  assign n55491 = n55489 & n55490 ;
  assign n55492 = n6736 | n34924 ;
  assign n55493 = n29286 & ~n55492 ;
  assign n55494 = n15310 | n55493 ;
  assign n55495 = n55494 ^ n27518 ^ 1'b0 ;
  assign n55496 = n28465 ^ n28181 ^ n3646 ;
  assign n55497 = ( ~n2441 & n8077 ) | ( ~n2441 & n31833 ) | ( n8077 & n31833 ) ;
  assign n55498 = ( n4865 & n19910 ) | ( n4865 & ~n35504 ) | ( n19910 & ~n35504 ) ;
  assign n55499 = ( ~n25715 & n32129 ) | ( ~n25715 & n33235 ) | ( n32129 & n33235 ) ;
  assign n55500 = ~n34942 & n44792 ;
  assign n55501 = n36150 ^ n27419 ^ n7559 ;
  assign n55502 = n20085 ^ n10768 ^ 1'b0 ;
  assign n55503 = ( n37880 & n49208 ) | ( n37880 & ~n55502 ) | ( n49208 & ~n55502 ) ;
  assign n55504 = n38757 ^ n27345 ^ n9260 ;
  assign n55505 = n55504 ^ n21065 ^ n6162 ;
  assign n55507 = n26155 & ~n33134 ;
  assign n55508 = ( ~n23670 & n53474 ) | ( ~n23670 & n55507 ) | ( n53474 & n55507 ) ;
  assign n55506 = n15753 & n32267 ;
  assign n55509 = n55508 ^ n55506 ^ n9571 ;
  assign n55510 = n43553 ^ n34383 ^ 1'b0 ;
  assign n55511 = ~n19011 & n55510 ;
  assign n55512 = n36312 ^ n17962 ^ 1'b0 ;
  assign n55513 = n30738 & ~n55512 ;
  assign n55514 = n51234 ^ n3235 ^ 1'b0 ;
  assign n55515 = n13105 & ~n28183 ;
  assign n55516 = n22559 & n55515 ;
  assign n55517 = n36462 | n55516 ;
  assign n55518 = ( ~n3568 & n7698 ) | ( ~n3568 & n34529 ) | ( n7698 & n34529 ) ;
  assign n55519 = n40930 ^ n32533 ^ 1'b0 ;
  assign n55520 = ( ~n9741 & n14511 ) | ( ~n9741 & n37848 ) | ( n14511 & n37848 ) ;
  assign n55521 = ( n55518 & n55519 ) | ( n55518 & ~n55520 ) | ( n55519 & ~n55520 ) ;
  assign n55522 = ( ~n1074 & n55517 ) | ( ~n1074 & n55521 ) | ( n55517 & n55521 ) ;
  assign n55523 = n24941 ^ n18863 ^ n10789 ;
  assign n55524 = ( n9042 & n24879 ) | ( n9042 & n42487 ) | ( n24879 & n42487 ) ;
  assign n55525 = ( n2095 & n42340 ) | ( n2095 & n55524 ) | ( n42340 & n55524 ) ;
  assign n55526 = ( ~n21544 & n55523 ) | ( ~n21544 & n55525 ) | ( n55523 & n55525 ) ;
  assign n55527 = ( ~n3422 & n11307 ) | ( ~n3422 & n27822 ) | ( n11307 & n27822 ) ;
  assign n55528 = n19711 & ~n21812 ;
  assign n55529 = n55528 ^ n32107 ^ 1'b0 ;
  assign n55530 = ( n18336 & n30288 ) | ( n18336 & n41153 ) | ( n30288 & n41153 ) ;
  assign n55531 = n55530 ^ n51856 ^ n48278 ;
  assign n55532 = n55529 & ~n55531 ;
  assign n55533 = n23491 ^ n7478 ^ 1'b0 ;
  assign n55534 = n4806 & n55533 ;
  assign n55535 = ( n5390 & n39478 ) | ( n5390 & ~n55534 ) | ( n39478 & ~n55534 ) ;
  assign n55536 = n3317 | n28157 ;
  assign n55537 = n55536 ^ n8731 ^ n5550 ;
  assign n55538 = n26803 | n30180 ;
  assign n55539 = n37491 ^ n7347 ^ 1'b0 ;
  assign n55540 = n4315 & n55539 ;
  assign n55541 = ( n14278 & ~n29790 ) | ( n14278 & n55540 ) | ( ~n29790 & n55540 ) ;
  assign n55542 = n55541 ^ n17000 ^ n13875 ;
  assign n55543 = n40220 ^ n11209 ^ n2789 ;
  assign n55544 = ~n12095 & n55543 ;
  assign n55545 = ~n55542 & n55544 ;
  assign n55546 = n26798 ^ n16788 ^ n5846 ;
  assign n55547 = n31390 ^ n21427 ^ 1'b0 ;
  assign n55548 = n1394 & ~n55547 ;
  assign n55549 = ( n33884 & ~n40717 ) | ( n33884 & n55548 ) | ( ~n40717 & n55548 ) ;
  assign n55550 = ( n19988 & n23512 ) | ( n19988 & n36976 ) | ( n23512 & n36976 ) ;
  assign n55551 = n21512 ^ n14595 ^ n9499 ;
  assign n55553 = n9025 ^ n6582 ^ n4428 ;
  assign n55552 = n55281 ^ n19390 ^ n10497 ;
  assign n55554 = n55553 ^ n55552 ^ n15986 ;
  assign n55555 = ~n9801 & n49797 ;
  assign n55556 = n32583 ^ n27834 ^ n26751 ;
  assign n55557 = n55556 ^ n10077 ^ n2541 ;
  assign n55558 = n46672 & ~n51628 ;
  assign n55559 = n49013 ^ n7194 ^ 1'b0 ;
  assign n55560 = n16098 | n55559 ;
  assign n55561 = n53791 ^ n6430 ^ 1'b0 ;
  assign n55562 = n45616 & ~n55561 ;
  assign n55565 = ( n2697 & ~n8120 ) | ( n2697 & n26669 ) | ( ~n8120 & n26669 ) ;
  assign n55566 = ( ~n8690 & n12962 ) | ( ~n8690 & n55565 ) | ( n12962 & n55565 ) ;
  assign n55563 = ~n30942 & n34413 ;
  assign n55564 = n40247 & ~n55563 ;
  assign n55567 = n55566 ^ n55564 ^ 1'b0 ;
  assign n55568 = n17963 ^ n9192 ^ n7715 ;
  assign n55569 = n14039 & ~n49612 ;
  assign n55570 = n55569 ^ n25287 ^ n8935 ;
  assign n55571 = n34394 & ~n55570 ;
  assign n55572 = ( n4424 & ~n47977 ) | ( n4424 & n55571 ) | ( ~n47977 & n55571 ) ;
  assign n55573 = n3379 & n16340 ;
  assign n55574 = n44632 ^ n17774 ^ n17100 ;
  assign n55575 = n55574 ^ n31954 ^ n23218 ;
  assign n55576 = ( n7587 & n15481 ) | ( n7587 & n51979 ) | ( n15481 & n51979 ) ;
  assign n55577 = ( n6886 & n54598 ) | ( n6886 & ~n55576 ) | ( n54598 & ~n55576 ) ;
  assign n55578 = ( n26056 & ~n44057 ) | ( n26056 & n50873 ) | ( ~n44057 & n50873 ) ;
  assign n55579 = ( n2929 & n7685 ) | ( n2929 & n25016 ) | ( n7685 & n25016 ) ;
  assign n55580 = ( n25796 & ~n43667 ) | ( n25796 & n55579 ) | ( ~n43667 & n55579 ) ;
  assign n55581 = ( n7513 & n53141 ) | ( n7513 & ~n55580 ) | ( n53141 & ~n55580 ) ;
  assign n55582 = n24466 ^ n14381 ^ n13669 ;
  assign n55584 = n25599 ^ n6197 ^ 1'b0 ;
  assign n55583 = n2105 & n27174 ;
  assign n55585 = n55584 ^ n55583 ^ 1'b0 ;
  assign n55586 = n38094 ^ n11378 ^ 1'b0 ;
  assign n55587 = ( n16686 & n19615 ) | ( n16686 & n37605 ) | ( n19615 & n37605 ) ;
  assign n55588 = n55587 ^ n11793 ^ 1'b0 ;
  assign n55589 = ~n55586 & n55588 ;
  assign n55590 = n24899 | n29918 ;
  assign n55591 = n41509 & ~n55590 ;
  assign n55592 = n48529 ^ n39279 ^ n22951 ;
  assign n55593 = n2347 & ~n38210 ;
  assign n55594 = ( n42295 & ~n46361 ) | ( n42295 & n55593 ) | ( ~n46361 & n55593 ) ;
  assign n55597 = ( n5839 & n19732 ) | ( n5839 & n20238 ) | ( n19732 & n20238 ) ;
  assign n55595 = n795 & ~n18515 ;
  assign n55596 = n55595 ^ n20845 ^ 1'b0 ;
  assign n55598 = n55597 ^ n55596 ^ n37143 ;
  assign n55599 = ( n16140 & n55594 ) | ( n16140 & ~n55598 ) | ( n55594 & ~n55598 ) ;
  assign n55600 = ( ~n11852 & n11991 ) | ( ~n11852 & n14549 ) | ( n11991 & n14549 ) ;
  assign n55601 = n55600 ^ n24341 ^ n23871 ;
  assign n55602 = n55601 ^ n26160 ^ n26103 ;
  assign n55603 = ( n761 & ~n2211 ) | ( n761 & n2423 ) | ( ~n2211 & n2423 ) ;
  assign n55604 = n37908 ^ n17897 ^ n17701 ;
  assign n55605 = ( n15104 & n55603 ) | ( n15104 & n55604 ) | ( n55603 & n55604 ) ;
  assign n55606 = n25320 ^ n18271 ^ n1727 ;
  assign n55607 = n55606 ^ n25970 ^ n15888 ;
  assign n55608 = n34032 ^ n8366 ^ 1'b0 ;
  assign n55609 = ~n16784 & n33603 ;
  assign n55610 = ~n9670 & n55609 ;
  assign n55611 = n15823 & ~n16827 ;
  assign n55612 = ~n10804 & n55611 ;
  assign n55613 = ( n41165 & ~n55610 ) | ( n41165 & n55612 ) | ( ~n55610 & n55612 ) ;
  assign n55614 = n55613 ^ n12456 ^ 1'b0 ;
  assign n55615 = n10651 & ~n20912 ;
  assign n55616 = n3023 & n23267 ;
  assign n55617 = n55616 ^ n34097 ^ 1'b0 ;
  assign n55618 = n32145 ^ n5219 ^ 1'b0 ;
  assign n55619 = n3259 & n55618 ;
  assign n55620 = n30658 ^ n26661 ^ 1'b0 ;
  assign n55621 = n6329 & ~n55620 ;
  assign n55622 = n54090 ^ n50470 ^ 1'b0 ;
  assign n55623 = n55621 & n55622 ;
  assign n55624 = n10327 & n23017 ;
  assign n55625 = ~n37717 & n41506 ;
  assign n55626 = ~n6258 & n50261 ;
  assign n55627 = n55626 ^ n27613 ^ n15419 ;
  assign n55628 = n42119 ^ n14662 ^ 1'b0 ;
  assign n55629 = n38418 ^ n32243 ^ 1'b0 ;
  assign n55630 = n45155 ^ n43652 ^ n21025 ;
  assign n55631 = ( n39676 & ~n49140 ) | ( n39676 & n55630 ) | ( ~n49140 & n55630 ) ;
  assign n55632 = n18708 | n22022 ;
  assign n55633 = n4404 | n51374 ;
  assign n55634 = n55633 ^ n21107 ^ 1'b0 ;
  assign n55635 = n6368 | n15671 ;
  assign n55636 = n55635 ^ n34304 ^ 1'b0 ;
  assign n55637 = ( n28415 & ~n55634 ) | ( n28415 & n55636 ) | ( ~n55634 & n55636 ) ;
  assign n55638 = n35602 ^ n6001 ^ 1'b0 ;
  assign n55639 = n24476 ^ n385 ^ 1'b0 ;
  assign n55640 = n2143 & n55639 ;
  assign n55641 = n5061 & ~n11650 ;
  assign n55642 = ( n45375 & n55640 ) | ( n45375 & n55641 ) | ( n55640 & n55641 ) ;
  assign n55643 = ( ~n2190 & n36116 ) | ( ~n2190 & n53208 ) | ( n36116 & n53208 ) ;
  assign n55647 = n55613 ^ n40246 ^ n22022 ;
  assign n55645 = n20359 ^ n6822 ^ n4675 ;
  assign n55644 = n25004 ^ n17399 ^ n3720 ;
  assign n55646 = n55645 ^ n55644 ^ n10536 ;
  assign n55648 = n55647 ^ n55646 ^ n3771 ;
  assign n55649 = n55508 ^ n46887 ^ n2335 ;
  assign n55650 = n32589 ^ n12473 ^ n10557 ;
  assign n55651 = ~n12503 & n55650 ;
  assign n55652 = n55651 ^ n17006 ^ n396 ;
  assign n55653 = n2336 | n50606 ;
  assign n55654 = ( ~n6278 & n14398 ) | ( ~n6278 & n42986 ) | ( n14398 & n42986 ) ;
  assign n55655 = ( n12389 & n24682 ) | ( n12389 & n44033 ) | ( n24682 & n44033 ) ;
  assign y0 = x22 ;
  assign y1 = x23 ;
  assign y2 = x44 ;
  assign y3 = x63 ;
  assign y4 = x81 ;
  assign y5 = x89 ;
  assign y6 = x113 ;
  assign y7 = x129 ;
  assign y8 = x134 ;
  assign y9 = x137 ;
  assign y10 = x147 ;
  assign y11 = x154 ;
  assign y12 = x158 ;
  assign y13 = x159 ;
  assign y14 = x160 ;
  assign y15 = x161 ;
  assign y16 = x168 ;
  assign y17 = x185 ;
  assign y18 = x186 ;
  assign y19 = x205 ;
  assign y20 = x227 ;
  assign y21 = x245 ;
  assign y22 = x247 ;
  assign y23 = ~n256 ;
  assign y24 = n259 ;
  assign y25 = n264 ;
  assign y26 = n265 ;
  assign y27 = n269 ;
  assign y28 = ~1'b0 ;
  assign y29 = n271 ;
  assign y30 = ~n273 ;
  assign y31 = ~1'b0 ;
  assign y32 = ~n275 ;
  assign y33 = n277 ;
  assign y34 = ~n278 ;
  assign y35 = n279 ;
  assign y36 = ~n282 ;
  assign y37 = n284 ;
  assign y38 = n287 ;
  assign y39 = ~n288 ;
  assign y40 = ~n290 ;
  assign y41 = ~n294 ;
  assign y42 = n297 ;
  assign y43 = ~n299 ;
  assign y44 = n302 ;
  assign y45 = n304 ;
  assign y46 = n307 ;
  assign y47 = n311 ;
  assign y48 = n313 ;
  assign y49 = ~n316 ;
  assign y50 = ~n318 ;
  assign y51 = ~n321 ;
  assign y52 = ~n323 ;
  assign y53 = ~1'b0 ;
  assign y54 = n327 ;
  assign y55 = n328 ;
  assign y56 = n333 ;
  assign y57 = n335 ;
  assign y58 = ~n342 ;
  assign y59 = n354 ;
  assign y60 = n361 ;
  assign y61 = n364 ;
  assign y62 = ~n365 ;
  assign y63 = n371 ;
  assign y64 = n374 ;
  assign y65 = ~1'b0 ;
  assign y66 = ~1'b0 ;
  assign y67 = n375 ;
  assign y68 = ~1'b0 ;
  assign y69 = ~1'b0 ;
  assign y70 = n379 ;
  assign y71 = ~n380 ;
  assign y72 = n384 ;
  assign y73 = n393 ;
  assign y74 = n394 ;
  assign y75 = ~n400 ;
  assign y76 = n402 ;
  assign y77 = n403 ;
  assign y78 = n405 ;
  assign y79 = ~1'b0 ;
  assign y80 = ~1'b0 ;
  assign y81 = ~n408 ;
  assign y82 = n420 ;
  assign y83 = n428 ;
  assign y84 = n439 ;
  assign y85 = n447 ;
  assign y86 = n453 ;
  assign y87 = ~n455 ;
  assign y88 = ~n460 ;
  assign y89 = n462 ;
  assign y90 = n466 ;
  assign y91 = ~n468 ;
  assign y92 = n469 ;
  assign y93 = ~n479 ;
  assign y94 = x77 ;
  assign y95 = ~n488 ;
  assign y96 = ~1'b0 ;
  assign y97 = ~1'b0 ;
  assign y98 = ~n495 ;
  assign y99 = ~1'b0 ;
  assign y100 = n508 ;
  assign y101 = ~1'b0 ;
  assign y102 = n512 ;
  assign y103 = n523 ;
  assign y104 = n526 ;
  assign y105 = ~n532 ;
  assign y106 = n538 ;
  assign y107 = n548 ;
  assign y108 = ~n551 ;
  assign y109 = n557 ;
  assign y110 = ~n566 ;
  assign y111 = ~n572 ;
  assign y112 = n599 ;
  assign y113 = n602 ;
  assign y114 = ~n606 ;
  assign y115 = ~n612 ;
  assign y116 = n613 ;
  assign y117 = n615 ;
  assign y118 = ~n620 ;
  assign y119 = n628 ;
  assign y120 = ~n632 ;
  assign y121 = ~n641 ;
  assign y122 = n645 ;
  assign y123 = n647 ;
  assign y124 = ~n663 ;
  assign y125 = ~n667 ;
  assign y126 = n670 ;
  assign y127 = n676 ;
  assign y128 = ~n678 ;
  assign y129 = ~n688 ;
  assign y130 = ~n692 ;
  assign y131 = n693 ;
  assign y132 = ~1'b0 ;
  assign y133 = n695 ;
  assign y134 = n696 ;
  assign y135 = n702 ;
  assign y136 = ~n703 ;
  assign y137 = ~1'b0 ;
  assign y138 = n709 ;
  assign y139 = n714 ;
  assign y140 = n721 ;
  assign y141 = ~n732 ;
  assign y142 = n734 ;
  assign y143 = n742 ;
  assign y144 = ~n745 ;
  assign y145 = n757 ;
  assign y146 = ~1'b0 ;
  assign y147 = ~n764 ;
  assign y148 = ~n773 ;
  assign y149 = ~n774 ;
  assign y150 = 1'b0 ;
  assign y151 = ~1'b0 ;
  assign y152 = ~n779 ;
  assign y153 = ~n781 ;
  assign y154 = n785 ;
  assign y155 = n789 ;
  assign y156 = n799 ;
  assign y157 = ~1'b0 ;
  assign y158 = ~n814 ;
  assign y159 = n827 ;
  assign y160 = n833 ;
  assign y161 = ~1'b0 ;
  assign y162 = n836 ;
  assign y163 = ~n842 ;
  assign y164 = ~n855 ;
  assign y165 = ~n858 ;
  assign y166 = n862 ;
  assign y167 = n869 ;
  assign y168 = ~n872 ;
  assign y169 = ~1'b0 ;
  assign y170 = ~n888 ;
  assign y171 = ~1'b0 ;
  assign y172 = ~n889 ;
  assign y173 = ~n903 ;
  assign y174 = n908 ;
  assign y175 = ~n910 ;
  assign y176 = n915 ;
  assign y177 = n924 ;
  assign y178 = ~n933 ;
  assign y179 = n934 ;
  assign y180 = ~n944 ;
  assign y181 = n962 ;
  assign y182 = ~n969 ;
  assign y183 = ~n973 ;
  assign y184 = n977 ;
  assign y185 = n990 ;
  assign y186 = ~n993 ;
  assign y187 = ~n994 ;
  assign y188 = n1005 ;
  assign y189 = ~n1013 ;
  assign y190 = n1018 ;
  assign y191 = n1022 ;
  assign y192 = ~n1026 ;
  assign y193 = ~n1045 ;
  assign y194 = n1048 ;
  assign y195 = n1049 ;
  assign y196 = n1050 ;
  assign y197 = n1052 ;
  assign y198 = ~n1062 ;
  assign y199 = ~n1063 ;
  assign y200 = ~n1067 ;
  assign y201 = n1072 ;
  assign y202 = ~n1075 ;
  assign y203 = ~n1078 ;
  assign y204 = ~n1080 ;
  assign y205 = ~n1081 ;
  assign y206 = n1084 ;
  assign y207 = ~1'b0 ;
  assign y208 = ~n1093 ;
  assign y209 = n1099 ;
  assign y210 = ~n1108 ;
  assign y211 = ~n1111 ;
  assign y212 = n1120 ;
  assign y213 = n1133 ;
  assign y214 = n1135 ;
  assign y215 = n1143 ;
  assign y216 = n1148 ;
  assign y217 = n1152 ;
  assign y218 = n1160 ;
  assign y219 = ~n1165 ;
  assign y220 = n1179 ;
  assign y221 = ~n1187 ;
  assign y222 = ~n1188 ;
  assign y223 = ~1'b0 ;
  assign y224 = n1189 ;
  assign y225 = ~n1190 ;
  assign y226 = ~n1198 ;
  assign y227 = ~1'b0 ;
  assign y228 = ~n1200 ;
  assign y229 = n1203 ;
  assign y230 = ~n1208 ;
  assign y231 = n1213 ;
  assign y232 = ~n1216 ;
  assign y233 = n1221 ;
  assign y234 = ~n1226 ;
  assign y235 = ~1'b0 ;
  assign y236 = ~n1248 ;
  assign y237 = ~n1254 ;
  assign y238 = ~1'b0 ;
  assign y239 = n1256 ;
  assign y240 = n1262 ;
  assign y241 = ~n1272 ;
  assign y242 = n1289 ;
  assign y243 = n1293 ;
  assign y244 = n1302 ;
  assign y245 = n1304 ;
  assign y246 = n1307 ;
  assign y247 = n1308 ;
  assign y248 = n1317 ;
  assign y249 = ~n1318 ;
  assign y250 = ~n1335 ;
  assign y251 = ~1'b0 ;
  assign y252 = n1346 ;
  assign y253 = n1349 ;
  assign y254 = ~n1351 ;
  assign y255 = n1362 ;
  assign y256 = ~n1364 ;
  assign y257 = n1394 ;
  assign y258 = n1427 ;
  assign y259 = ~n1467 ;
  assign y260 = n1470 ;
  assign y261 = ~n1475 ;
  assign y262 = n1482 ;
  assign y263 = ~n1492 ;
  assign y264 = ~n1502 ;
  assign y265 = n1503 ;
  assign y266 = n1519 ;
  assign y267 = n1536 ;
  assign y268 = n1539 ;
  assign y269 = n1544 ;
  assign y270 = ~n1549 ;
  assign y271 = ~1'b0 ;
  assign y272 = ~n1551 ;
  assign y273 = n1565 ;
  assign y274 = ~n1566 ;
  assign y275 = n1576 ;
  assign y276 = n1581 ;
  assign y277 = ~n1588 ;
  assign y278 = n1590 ;
  assign y279 = ~n1610 ;
  assign y280 = ~n1620 ;
  assign y281 = n1621 ;
  assign y282 = ~n1627 ;
  assign y283 = ~n1635 ;
  assign y284 = n1636 ;
  assign y285 = n1648 ;
  assign y286 = ~n1654 ;
  assign y287 = ~n1659 ;
  assign y288 = ~n1678 ;
  assign y289 = n1686 ;
  assign y290 = ~1'b0 ;
  assign y291 = ~n1693 ;
  assign y292 = n1696 ;
  assign y293 = ~n1700 ;
  assign y294 = ~n1706 ;
  assign y295 = n1714 ;
  assign y296 = ~n1729 ;
  assign y297 = ~n1734 ;
  assign y298 = ~n1739 ;
  assign y299 = ~n1741 ;
  assign y300 = n1745 ;
  assign y301 = ~n1751 ;
  assign y302 = ~n1759 ;
  assign y303 = n1775 ;
  assign y304 = n1776 ;
  assign y305 = n1779 ;
  assign y306 = ~n1794 ;
  assign y307 = ~n1796 ;
  assign y308 = ~1'b0 ;
  assign y309 = n1802 ;
  assign y310 = ~n1806 ;
  assign y311 = n1811 ;
  assign y312 = ~n1819 ;
  assign y313 = ~n1825 ;
  assign y314 = ~n1831 ;
  assign y315 = ~n1832 ;
  assign y316 = n1835 ;
  assign y317 = ~1'b0 ;
  assign y318 = ~n1838 ;
  assign y319 = n1846 ;
  assign y320 = n1858 ;
  assign y321 = n1859 ;
  assign y322 = ~n1862 ;
  assign y323 = ~n1883 ;
  assign y324 = n1886 ;
  assign y325 = ~n1888 ;
  assign y326 = ~n1896 ;
  assign y327 = n1900 ;
  assign y328 = n1908 ;
  assign y329 = n1916 ;
  assign y330 = ~n1635 ;
  assign y331 = n1926 ;
  assign y332 = ~n1927 ;
  assign y333 = ~n1932 ;
  assign y334 = n1941 ;
  assign y335 = n1944 ;
  assign y336 = ~n1953 ;
  assign y337 = ~n1960 ;
  assign y338 = ~1'b0 ;
  assign y339 = n1975 ;
  assign y340 = n1983 ;
  assign y341 = n1984 ;
  assign y342 = n1988 ;
  assign y343 = ~1'b0 ;
  assign y344 = ~1'b0 ;
  assign y345 = ~1'b0 ;
  assign y346 = n2002 ;
  assign y347 = n2003 ;
  assign y348 = ~n2004 ;
  assign y349 = ~n2006 ;
  assign y350 = ~n2022 ;
  assign y351 = ~n2029 ;
  assign y352 = ~n2035 ;
  assign y353 = n2037 ;
  assign y354 = ~1'b0 ;
  assign y355 = ~n2039 ;
  assign y356 = ~n2050 ;
  assign y357 = ~n2062 ;
  assign y358 = ~x200 ;
  assign y359 = ~n2065 ;
  assign y360 = n2067 ;
  assign y361 = ~n2074 ;
  assign y362 = n2077 ;
  assign y363 = ~n2081 ;
  assign y364 = ~n2083 ;
  assign y365 = ~n2092 ;
  assign y366 = n2094 ;
  assign y367 = n2097 ;
  assign y368 = n2098 ;
  assign y369 = n2106 ;
  assign y370 = ~n2109 ;
  assign y371 = n2113 ;
  assign y372 = ~n2140 ;
  assign y373 = n2148 ;
  assign y374 = n2150 ;
  assign y375 = n2152 ;
  assign y376 = ~n2167 ;
  assign y377 = n2173 ;
  assign y378 = n2178 ;
  assign y379 = ~1'b0 ;
  assign y380 = n2180 ;
  assign y381 = n2187 ;
  assign y382 = n2191 ;
  assign y383 = ~n2193 ;
  assign y384 = n2199 ;
  assign y385 = ~n2208 ;
  assign y386 = ~1'b0 ;
  assign y387 = n2209 ;
  assign y388 = ~n2223 ;
  assign y389 = ~n2226 ;
  assign y390 = ~1'b0 ;
  assign y391 = n2228 ;
  assign y392 = ~n2235 ;
  assign y393 = ~n2240 ;
  assign y394 = n2247 ;
  assign y395 = ~n2248 ;
  assign y396 = n2272 ;
  assign y397 = ~n2287 ;
  assign y398 = n2290 ;
  assign y399 = n2298 ;
  assign y400 = ~n2299 ;
  assign y401 = ~n2304 ;
  assign y402 = n2305 ;
  assign y403 = n2312 ;
  assign y404 = ~n2319 ;
  assign y405 = n2322 ;
  assign y406 = n2325 ;
  assign y407 = n2326 ;
  assign y408 = n2330 ;
  assign y409 = ~n2331 ;
  assign y410 = ~n2332 ;
  assign y411 = ~n2339 ;
  assign y412 = n2341 ;
  assign y413 = n2354 ;
  assign y414 = ~n2366 ;
  assign y415 = n2369 ;
  assign y416 = n2381 ;
  assign y417 = n2385 ;
  assign y418 = ~n2387 ;
  assign y419 = n2392 ;
  assign y420 = n2404 ;
  assign y421 = ~n2407 ;
  assign y422 = ~n2413 ;
  assign y423 = n2416 ;
  assign y424 = ~n2423 ;
  assign y425 = n2428 ;
  assign y426 = ~n2439 ;
  assign y427 = ~n2448 ;
  assign y428 = ~n2451 ;
  assign y429 = ~n2458 ;
  assign y430 = ~1'b0 ;
  assign y431 = ~n2464 ;
  assign y432 = ~n439 ;
  assign y433 = n2466 ;
  assign y434 = n2468 ;
  assign y435 = n2471 ;
  assign y436 = n2477 ;
  assign y437 = ~n2481 ;
  assign y438 = ~n2488 ;
  assign y439 = n2496 ;
  assign y440 = ~n2497 ;
  assign y441 = n2501 ;
  assign y442 = ~n2514 ;
  assign y443 = n2519 ;
  assign y444 = ~n2524 ;
  assign y445 = n2533 ;
  assign y446 = n2536 ;
  assign y447 = n2538 ;
  assign y448 = ~n2561 ;
  assign y449 = ~1'b0 ;
  assign y450 = n2562 ;
  assign y451 = n2572 ;
  assign y452 = ~n2574 ;
  assign y453 = ~n2575 ;
  assign y454 = n2576 ;
  assign y455 = ~n2580 ;
  assign y456 = n2585 ;
  assign y457 = ~n2587 ;
  assign y458 = n2596 ;
  assign y459 = ~n2597 ;
  assign y460 = ~n2612 ;
  assign y461 = n2613 ;
  assign y462 = ~n2620 ;
  assign y463 = n2638 ;
  assign y464 = n2640 ;
  assign y465 = n2656 ;
  assign y466 = n2661 ;
  assign y467 = ~n2666 ;
  assign y468 = ~n2669 ;
  assign y469 = n2677 ;
  assign y470 = ~n2682 ;
  assign y471 = ~n2688 ;
  assign y472 = ~n2694 ;
  assign y473 = ~1'b0 ;
  assign y474 = n2712 ;
  assign y475 = n2713 ;
  assign y476 = ~1'b0 ;
  assign y477 = n2714 ;
  assign y478 = ~1'b0 ;
  assign y479 = ~n2722 ;
  assign y480 = n2731 ;
  assign y481 = ~n2741 ;
  assign y482 = n2744 ;
  assign y483 = ~n2747 ;
  assign y484 = ~n2763 ;
  assign y485 = ~n2774 ;
  assign y486 = ~n2780 ;
  assign y487 = n2784 ;
  assign y488 = ~n2811 ;
  assign y489 = ~n2826 ;
  assign y490 = ~n2832 ;
  assign y491 = ~n2833 ;
  assign y492 = n2889 ;
  assign y493 = ~n2891 ;
  assign y494 = n2892 ;
  assign y495 = ~1'b0 ;
  assign y496 = n2896 ;
  assign y497 = n2898 ;
  assign y498 = n2902 ;
  assign y499 = n2911 ;
  assign y500 = ~n2927 ;
  assign y501 = ~1'b0 ;
  assign y502 = n2932 ;
  assign y503 = n2948 ;
  assign y504 = ~n2972 ;
  assign y505 = n2992 ;
  assign y506 = ~n3003 ;
  assign y507 = n3005 ;
  assign y508 = n3011 ;
  assign y509 = n3035 ;
  assign y510 = n3045 ;
  assign y511 = ~n3049 ;
  assign y512 = ~n3051 ;
  assign y513 = ~n3056 ;
  assign y514 = ~n2381 ;
  assign y515 = ~n3080 ;
  assign y516 = ~n3085 ;
  assign y517 = n3086 ;
  assign y518 = ~n3090 ;
  assign y519 = n522 ;
  assign y520 = n3095 ;
  assign y521 = n3103 ;
  assign y522 = ~n3107 ;
  assign y523 = ~n3108 ;
  assign y524 = ~n3110 ;
  assign y525 = n3111 ;
  assign y526 = ~n3113 ;
  assign y527 = n3119 ;
  assign y528 = ~n3122 ;
  assign y529 = n3128 ;
  assign y530 = ~n3145 ;
  assign y531 = n3148 ;
  assign y532 = ~1'b0 ;
  assign y533 = ~n3162 ;
  assign y534 = ~n3165 ;
  assign y535 = n3167 ;
  assign y536 = ~n3173 ;
  assign y537 = n3192 ;
  assign y538 = n3194 ;
  assign y539 = ~n3195 ;
  assign y540 = ~n3197 ;
  assign y541 = ~n3199 ;
  assign y542 = ~n3208 ;
  assign y543 = ~n3210 ;
  assign y544 = n3222 ;
  assign y545 = ~n3231 ;
  assign y546 = n3239 ;
  assign y547 = ~n3243 ;
  assign y548 = n3244 ;
  assign y549 = n3248 ;
  assign y550 = ~1'b0 ;
  assign y551 = n3263 ;
  assign y552 = n3264 ;
  assign y553 = ~1'b0 ;
  assign y554 = ~n3274 ;
  assign y555 = ~n3279 ;
  assign y556 = ~n3281 ;
  assign y557 = ~n3292 ;
  assign y558 = n3295 ;
  assign y559 = ~n3297 ;
  assign y560 = ~n3304 ;
  assign y561 = ~n3311 ;
  assign y562 = n3322 ;
  assign y563 = ~n3329 ;
  assign y564 = n3332 ;
  assign y565 = ~1'b0 ;
  assign y566 = ~n3333 ;
  assign y567 = n2646 ;
  assign y568 = n3335 ;
  assign y569 = ~n3337 ;
  assign y570 = n3340 ;
  assign y571 = n3343 ;
  assign y572 = n3359 ;
  assign y573 = n3367 ;
  assign y574 = n3373 ;
  assign y575 = ~n3374 ;
  assign y576 = n3378 ;
  assign y577 = n3385 ;
  assign y578 = n3396 ;
  assign y579 = n3402 ;
  assign y580 = n3403 ;
  assign y581 = ~n3407 ;
  assign y582 = ~n3412 ;
  assign y583 = ~n3413 ;
  assign y584 = ~n3420 ;
  assign y585 = n3435 ;
  assign y586 = ~n3439 ;
  assign y587 = n3443 ;
  assign y588 = ~n3444 ;
  assign y589 = n3447 ;
  assign y590 = ~n3462 ;
  assign y591 = n3464 ;
  assign y592 = n3470 ;
  assign y593 = ~n3473 ;
  assign y594 = n3477 ;
  assign y595 = n3483 ;
  assign y596 = ~1'b0 ;
  assign y597 = ~n3487 ;
  assign y598 = x27 ;
  assign y599 = n3495 ;
  assign y600 = n3498 ;
  assign y601 = ~1'b0 ;
  assign y602 = ~n3503 ;
  assign y603 = ~n3507 ;
  assign y604 = n3511 ;
  assign y605 = ~n3512 ;
  assign y606 = ~n3521 ;
  assign y607 = n3525 ;
  assign y608 = ~n3526 ;
  assign y609 = n3533 ;
  assign y610 = n3538 ;
  assign y611 = n3551 ;
  assign y612 = n3553 ;
  assign y613 = ~n3580 ;
  assign y614 = ~n3581 ;
  assign y615 = ~n3591 ;
  assign y616 = ~n3594 ;
  assign y617 = ~n3597 ;
  assign y618 = ~n3599 ;
  assign y619 = ~n3622 ;
  assign y620 = ~n3624 ;
  assign y621 = n3625 ;
  assign y622 = ~n3627 ;
  assign y623 = ~n3630 ;
  assign y624 = n3631 ;
  assign y625 = n3632 ;
  assign y626 = ~1'b0 ;
  assign y627 = n3641 ;
  assign y628 = ~1'b0 ;
  assign y629 = n3650 ;
  assign y630 = ~n3653 ;
  assign y631 = ~n3660 ;
  assign y632 = n3663 ;
  assign y633 = n3664 ;
  assign y634 = ~n3671 ;
  assign y635 = n3674 ;
  assign y636 = n3676 ;
  assign y637 = ~1'b0 ;
  assign y638 = ~n3681 ;
  assign y639 = n3686 ;
  assign y640 = ~n3690 ;
  assign y641 = n3691 ;
  assign y642 = ~1'b0 ;
  assign y643 = ~n3696 ;
  assign y644 = ~n3697 ;
  assign y645 = n3699 ;
  assign y646 = n3700 ;
  assign y647 = ~n3714 ;
  assign y648 = ~n3717 ;
  assign y649 = ~1'b0 ;
  assign y650 = n3721 ;
  assign y651 = n3722 ;
  assign y652 = n3724 ;
  assign y653 = n3729 ;
  assign y654 = ~n3742 ;
  assign y655 = n3745 ;
  assign y656 = n3758 ;
  assign y657 = n3760 ;
  assign y658 = n3761 ;
  assign y659 = ~n3763 ;
  assign y660 = ~n3773 ;
  assign y661 = ~n3776 ;
  assign y662 = n3787 ;
  assign y663 = ~n3791 ;
  assign y664 = ~1'b0 ;
  assign y665 = ~n3796 ;
  assign y666 = ~1'b0 ;
  assign y667 = n3802 ;
  assign y668 = ~n3808 ;
  assign y669 = ~n3818 ;
  assign y670 = ~n3822 ;
  assign y671 = n3826 ;
  assign y672 = ~n3834 ;
  assign y673 = n3845 ;
  assign y674 = n3854 ;
  assign y675 = n3856 ;
  assign y676 = n3869 ;
  assign y677 = ~n3872 ;
  assign y678 = n3877 ;
  assign y679 = n3883 ;
  assign y680 = ~1'b0 ;
  assign y681 = n3885 ;
  assign y682 = ~n3900 ;
  assign y683 = n3902 ;
  assign y684 = n3909 ;
  assign y685 = ~n3919 ;
  assign y686 = ~n3935 ;
  assign y687 = ~n3938 ;
  assign y688 = ~n3952 ;
  assign y689 = n3955 ;
  assign y690 = n3956 ;
  assign y691 = n3958 ;
  assign y692 = ~1'b0 ;
  assign y693 = ~n3960 ;
  assign y694 = n3967 ;
  assign y695 = n3975 ;
  assign y696 = ~n3980 ;
  assign y697 = n3984 ;
  assign y698 = ~n3987 ;
  assign y699 = ~1'b0 ;
  assign y700 = ~n3991 ;
  assign y701 = n3993 ;
  assign y702 = ~n4010 ;
  assign y703 = n4033 ;
  assign y704 = ~n4035 ;
  assign y705 = n4037 ;
  assign y706 = ~n4038 ;
  assign y707 = n4039 ;
  assign y708 = n4044 ;
  assign y709 = n4047 ;
  assign y710 = n4050 ;
  assign y711 = n4056 ;
  assign y712 = ~n4071 ;
  assign y713 = ~n4081 ;
  assign y714 = ~n4092 ;
  assign y715 = ~n4095 ;
  assign y716 = n4098 ;
  assign y717 = ~n4105 ;
  assign y718 = n4111 ;
  assign y719 = n4115 ;
  assign y720 = n4116 ;
  assign y721 = ~n4141 ;
  assign y722 = n4147 ;
  assign y723 = ~n4148 ;
  assign y724 = n4159 ;
  assign y725 = ~n4179 ;
  assign y726 = ~n4190 ;
  assign y727 = ~n4192 ;
  assign y728 = n4196 ;
  assign y729 = ~n4199 ;
  assign y730 = ~n4203 ;
  assign y731 = ~n4209 ;
  assign y732 = n4215 ;
  assign y733 = n4221 ;
  assign y734 = ~n4224 ;
  assign y735 = ~n4235 ;
  assign y736 = n4239 ;
  assign y737 = ~n4246 ;
  assign y738 = ~n4249 ;
  assign y739 = n4250 ;
  assign y740 = n4251 ;
  assign y741 = ~n4255 ;
  assign y742 = n4260 ;
  assign y743 = ~n4262 ;
  assign y744 = n4265 ;
  assign y745 = ~n4269 ;
  assign y746 = ~n4271 ;
  assign y747 = n4276 ;
  assign y748 = n4280 ;
  assign y749 = ~n4282 ;
  assign y750 = n4287 ;
  assign y751 = n4288 ;
  assign y752 = n4290 ;
  assign y753 = ~n4292 ;
  assign y754 = n4293 ;
  assign y755 = ~1'b0 ;
  assign y756 = n4303 ;
  assign y757 = ~1'b0 ;
  assign y758 = n4312 ;
  assign y759 = n4320 ;
  assign y760 = n4329 ;
  assign y761 = n4333 ;
  assign y762 = n4344 ;
  assign y763 = ~n4349 ;
  assign y764 = n4352 ;
  assign y765 = ~n4369 ;
  assign y766 = ~n4370 ;
  assign y767 = n4372 ;
  assign y768 = n4374 ;
  assign y769 = n4382 ;
  assign y770 = n4391 ;
  assign y771 = n4397 ;
  assign y772 = n4398 ;
  assign y773 = ~n4404 ;
  assign y774 = ~1'b0 ;
  assign y775 = n4407 ;
  assign y776 = n4413 ;
  assign y777 = n4418 ;
  assign y778 = n4420 ;
  assign y779 = n4421 ;
  assign y780 = ~n4429 ;
  assign y781 = n4450 ;
  assign y782 = n4464 ;
  assign y783 = n4466 ;
  assign y784 = ~1'b0 ;
  assign y785 = ~n4467 ;
  assign y786 = ~n4468 ;
  assign y787 = n4472 ;
  assign y788 = ~1'b0 ;
  assign y789 = n4479 ;
  assign y790 = ~n4488 ;
  assign y791 = ~n4498 ;
  assign y792 = n4500 ;
  assign y793 = ~n4503 ;
  assign y794 = n4506 ;
  assign y795 = ~n4518 ;
  assign y796 = n4525 ;
  assign y797 = n4528 ;
  assign y798 = n4529 ;
  assign y799 = n4534 ;
  assign y800 = n4540 ;
  assign y801 = ~n4554 ;
  assign y802 = n4561 ;
  assign y803 = n4568 ;
  assign y804 = n4570 ;
  assign y805 = ~1'b0 ;
  assign y806 = n4575 ;
  assign y807 = n4579 ;
  assign y808 = n4583 ;
  assign y809 = n4586 ;
  assign y810 = n4588 ;
  assign y811 = n4607 ;
  assign y812 = n4614 ;
  assign y813 = n4622 ;
  assign y814 = ~n4623 ;
  assign y815 = n4630 ;
  assign y816 = ~n4633 ;
  assign y817 = n4643 ;
  assign y818 = n4646 ;
  assign y819 = n4647 ;
  assign y820 = n4657 ;
  assign y821 = ~n4668 ;
  assign y822 = n4669 ;
  assign y823 = ~n4679 ;
  assign y824 = ~n4681 ;
  assign y825 = n4689 ;
  assign y826 = n4706 ;
  assign y827 = n4719 ;
  assign y828 = n4722 ;
  assign y829 = n4727 ;
  assign y830 = n4730 ;
  assign y831 = n4733 ;
  assign y832 = n1212 ;
  assign y833 = ~n4734 ;
  assign y834 = ~n4738 ;
  assign y835 = n4756 ;
  assign y836 = n4758 ;
  assign y837 = n4764 ;
  assign y838 = n4777 ;
  assign y839 = ~1'b0 ;
  assign y840 = ~1'b0 ;
  assign y841 = n4781 ;
  assign y842 = n4792 ;
  assign y843 = ~n4795 ;
  assign y844 = n4804 ;
  assign y845 = ~n4809 ;
  assign y846 = ~n4818 ;
  assign y847 = ~n4825 ;
  assign y848 = n4834 ;
  assign y849 = n4839 ;
  assign y850 = ~n4842 ;
  assign y851 = n4852 ;
  assign y852 = n4854 ;
  assign y853 = ~n4857 ;
  assign y854 = n4858 ;
  assign y855 = n4864 ;
  assign y856 = n4875 ;
  assign y857 = ~n4898 ;
  assign y858 = n4905 ;
  assign y859 = ~n4908 ;
  assign y860 = n4928 ;
  assign y861 = n4949 ;
  assign y862 = ~n4956 ;
  assign y863 = n4959 ;
  assign y864 = ~1'b0 ;
  assign y865 = ~n4966 ;
  assign y866 = ~n4999 ;
  assign y867 = n5001 ;
  assign y868 = n5025 ;
  assign y869 = n5027 ;
  assign y870 = n5029 ;
  assign y871 = ~1'b0 ;
  assign y872 = n5032 ;
  assign y873 = ~n5033 ;
  assign y874 = n5054 ;
  assign y875 = n5057 ;
  assign y876 = ~n5062 ;
  assign y877 = ~n5069 ;
  assign y878 = ~1'b0 ;
  assign y879 = n5072 ;
  assign y880 = ~n5078 ;
  assign y881 = n5081 ;
  assign y882 = n5085 ;
  assign y883 = ~1'b0 ;
  assign y884 = ~n5093 ;
  assign y885 = ~n5103 ;
  assign y886 = ~n5106 ;
  assign y887 = n5116 ;
  assign y888 = ~n5117 ;
  assign y889 = n5124 ;
  assign y890 = ~n5126 ;
  assign y891 = n5136 ;
  assign y892 = ~n5138 ;
  assign y893 = n5140 ;
  assign y894 = ~n5145 ;
  assign y895 = ~n5156 ;
  assign y896 = n5158 ;
  assign y897 = n5160 ;
  assign y898 = ~n5165 ;
  assign y899 = ~1'b0 ;
  assign y900 = ~n5166 ;
  assign y901 = n5167 ;
  assign y902 = n5172 ;
  assign y903 = n5177 ;
  assign y904 = ~n5182 ;
  assign y905 = n5185 ;
  assign y906 = ~n5186 ;
  assign y907 = n5190 ;
  assign y908 = n5191 ;
  assign y909 = n5192 ;
  assign y910 = ~n5199 ;
  assign y911 = ~n5200 ;
  assign y912 = n5203 ;
  assign y913 = n5211 ;
  assign y914 = ~n5213 ;
  assign y915 = n5221 ;
  assign y916 = ~n5235 ;
  assign y917 = ~n5240 ;
  assign y918 = n5242 ;
  assign y919 = ~n5243 ;
  assign y920 = ~n5245 ;
  assign y921 = ~n5266 ;
  assign y922 = ~n5273 ;
  assign y923 = n5277 ;
  assign y924 = n5282 ;
  assign y925 = ~n5293 ;
  assign y926 = n5297 ;
  assign y927 = ~n5302 ;
  assign y928 = ~n5311 ;
  assign y929 = ~n5316 ;
  assign y930 = ~n5321 ;
  assign y931 = ~n5336 ;
  assign y932 = ~1'b0 ;
  assign y933 = n5338 ;
  assign y934 = ~n5347 ;
  assign y935 = ~n5350 ;
  assign y936 = ~n5359 ;
  assign y937 = ~n5377 ;
  assign y938 = n5381 ;
  assign y939 = n5384 ;
  assign y940 = ~n5385 ;
  assign y941 = n5393 ;
  assign y942 = n5395 ;
  assign y943 = n5399 ;
  assign y944 = n5400 ;
  assign y945 = n5405 ;
  assign y946 = ~n5407 ;
  assign y947 = ~n5414 ;
  assign y948 = n5416 ;
  assign y949 = n5418 ;
  assign y950 = n5420 ;
  assign y951 = n5427 ;
  assign y952 = n5430 ;
  assign y953 = n5433 ;
  assign y954 = n5439 ;
  assign y955 = ~n5440 ;
  assign y956 = n5443 ;
  assign y957 = n5452 ;
  assign y958 = ~n5464 ;
  assign y959 = ~n5467 ;
  assign y960 = ~n5468 ;
  assign y961 = n5469 ;
  assign y962 = ~n5473 ;
  assign y963 = n5474 ;
  assign y964 = ~n5476 ;
  assign y965 = ~1'b0 ;
  assign y966 = ~n5480 ;
  assign y967 = n5489 ;
  assign y968 = ~n5499 ;
  assign y969 = ~n5501 ;
  assign y970 = ~n5509 ;
  assign y971 = n5525 ;
  assign y972 = n5534 ;
  assign y973 = n5540 ;
  assign y974 = n5547 ;
  assign y975 = ~n5557 ;
  assign y976 = ~n5558 ;
  assign y977 = ~n5568 ;
  assign y978 = ~n5572 ;
  assign y979 = ~n5575 ;
  assign y980 = n5578 ;
  assign y981 = ~1'b0 ;
  assign y982 = ~n5581 ;
  assign y983 = n5598 ;
  assign y984 = ~n5608 ;
  assign y985 = ~n5615 ;
  assign y986 = ~n5624 ;
  assign y987 = ~n5632 ;
  assign y988 = n5656 ;
  assign y989 = ~1'b0 ;
  assign y990 = n5658 ;
  assign y991 = n5663 ;
  assign y992 = ~n5666 ;
  assign y993 = n5678 ;
  assign y994 = ~n5682 ;
  assign y995 = ~n5686 ;
  assign y996 = n5690 ;
  assign y997 = ~1'b0 ;
  assign y998 = n5692 ;
  assign y999 = ~n5697 ;
  assign y1000 = n5703 ;
  assign y1001 = ~n5707 ;
  assign y1002 = ~n5720 ;
  assign y1003 = n5732 ;
  assign y1004 = ~1'b0 ;
  assign y1005 = ~1'b0 ;
  assign y1006 = ~n5740 ;
  assign y1007 = ~n5743 ;
  assign y1008 = ~n5744 ;
  assign y1009 = n5748 ;
  assign y1010 = n5759 ;
  assign y1011 = ~1'b0 ;
  assign y1012 = ~n5769 ;
  assign y1013 = ~n5779 ;
  assign y1014 = n5782 ;
  assign y1015 = n5790 ;
  assign y1016 = ~1'b0 ;
  assign y1017 = ~n5791 ;
  assign y1018 = n5793 ;
  assign y1019 = n5794 ;
  assign y1020 = ~n5796 ;
  assign y1021 = ~n5813 ;
  assign y1022 = ~n5826 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = n5833 ;
  assign y1025 = ~1'b0 ;
  assign y1026 = n5840 ;
  assign y1027 = n5854 ;
  assign y1028 = ~n5856 ;
  assign y1029 = n5862 ;
  assign y1030 = ~n5867 ;
  assign y1031 = ~n5874 ;
  assign y1032 = ~1'b0 ;
  assign y1033 = n5877 ;
  assign y1034 = n5880 ;
  assign y1035 = ~n5888 ;
  assign y1036 = n5897 ;
  assign y1037 = ~1'b0 ;
  assign y1038 = ~n5898 ;
  assign y1039 = ~n5916 ;
  assign y1040 = ~n5925 ;
  assign y1041 = n5948 ;
  assign y1042 = ~n5957 ;
  assign y1043 = ~n5962 ;
  assign y1044 = ~n3794 ;
  assign y1045 = ~n5975 ;
  assign y1046 = n5996 ;
  assign y1047 = ~n5999 ;
  assign y1048 = n6001 ;
  assign y1049 = n6013 ;
  assign y1050 = ~n6017 ;
  assign y1051 = ~n6019 ;
  assign y1052 = n6028 ;
  assign y1053 = ~n6029 ;
  assign y1054 = ~n6036 ;
  assign y1055 = n6040 ;
  assign y1056 = n6048 ;
  assign y1057 = ~n6051 ;
  assign y1058 = ~n6058 ;
  assign y1059 = ~n6060 ;
  assign y1060 = n6061 ;
  assign y1061 = n6070 ;
  assign y1062 = ~n6073 ;
  assign y1063 = ~1'b0 ;
  assign y1064 = ~n6079 ;
  assign y1065 = ~n6081 ;
  assign y1066 = n6084 ;
  assign y1067 = ~n6089 ;
  assign y1068 = n6100 ;
  assign y1069 = ~n6101 ;
  assign y1070 = n6109 ;
  assign y1071 = n6116 ;
  assign y1072 = n6119 ;
  assign y1073 = ~n6136 ;
  assign y1074 = ~1'b0 ;
  assign y1075 = ~n6153 ;
  assign y1076 = ~n6156 ;
  assign y1077 = ~1'b0 ;
  assign y1078 = n6167 ;
  assign y1079 = ~n6174 ;
  assign y1080 = ~n6188 ;
  assign y1081 = n6202 ;
  assign y1082 = ~n6203 ;
  assign y1083 = ~n6205 ;
  assign y1084 = ~n6210 ;
  assign y1085 = ~n6216 ;
  assign y1086 = ~n6219 ;
  assign y1087 = ~n6229 ;
  assign y1088 = n6234 ;
  assign y1089 = n6243 ;
  assign y1090 = n6253 ;
  assign y1091 = n6255 ;
  assign y1092 = n6256 ;
  assign y1093 = n6261 ;
  assign y1094 = n6275 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = ~n6280 ;
  assign y1097 = ~1'b0 ;
  assign y1098 = n6293 ;
  assign y1099 = n6298 ;
  assign y1100 = ~n6300 ;
  assign y1101 = n6310 ;
  assign y1102 = n6325 ;
  assign y1103 = ~n6327 ;
  assign y1104 = ~1'b0 ;
  assign y1105 = n6331 ;
  assign y1106 = ~1'b0 ;
  assign y1107 = ~n6340 ;
  assign y1108 = n6349 ;
  assign y1109 = ~n6353 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = n6356 ;
  assign y1112 = n6358 ;
  assign y1113 = n6362 ;
  assign y1114 = n6369 ;
  assign y1115 = n6373 ;
  assign y1116 = ~n6385 ;
  assign y1117 = ~1'b0 ;
  assign y1118 = ~n6388 ;
  assign y1119 = n6389 ;
  assign y1120 = ~n6392 ;
  assign y1121 = n6398 ;
  assign y1122 = ~n6403 ;
  assign y1123 = n6419 ;
  assign y1124 = n6434 ;
  assign y1125 = ~1'b0 ;
  assign y1126 = ~n6437 ;
  assign y1127 = ~n6449 ;
  assign y1128 = n6455 ;
  assign y1129 = ~n6460 ;
  assign y1130 = n6461 ;
  assign y1131 = ~n6467 ;
  assign y1132 = n6496 ;
  assign y1133 = ~n6505 ;
  assign y1134 = ~n6508 ;
  assign y1135 = n6510 ;
  assign y1136 = n6523 ;
  assign y1137 = ~n6528 ;
  assign y1138 = ~n6533 ;
  assign y1139 = ~1'b0 ;
  assign y1140 = ~n6548 ;
  assign y1141 = n6550 ;
  assign y1142 = ~n6558 ;
  assign y1143 = n6566 ;
  assign y1144 = n6569 ;
  assign y1145 = n6570 ;
  assign y1146 = ~n6573 ;
  assign y1147 = n6581 ;
  assign y1148 = ~n6586 ;
  assign y1149 = n6598 ;
  assign y1150 = ~1'b0 ;
  assign y1151 = n6599 ;
  assign y1152 = ~n6648 ;
  assign y1153 = ~n6652 ;
  assign y1154 = ~n6657 ;
  assign y1155 = ~n6659 ;
  assign y1156 = ~n6668 ;
  assign y1157 = n6674 ;
  assign y1158 = ~n6676 ;
  assign y1159 = ~n6677 ;
  assign y1160 = n6695 ;
  assign y1161 = n6697 ;
  assign y1162 = n6700 ;
  assign y1163 = ~n6702 ;
  assign y1164 = n6703 ;
  assign y1165 = n6704 ;
  assign y1166 = ~n6716 ;
  assign y1167 = n6726 ;
  assign y1168 = n6730 ;
  assign y1169 = ~n6732 ;
  assign y1170 = ~n6736 ;
  assign y1171 = n6741 ;
  assign y1172 = ~1'b0 ;
  assign y1173 = ~n6748 ;
  assign y1174 = ~n6753 ;
  assign y1175 = ~n6755 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = ~n6757 ;
  assign y1178 = n6760 ;
  assign y1179 = n6762 ;
  assign y1180 = ~n6774 ;
  assign y1181 = n6778 ;
  assign y1182 = ~n6780 ;
  assign y1183 = n6782 ;
  assign y1184 = n6797 ;
  assign y1185 = ~n6800 ;
  assign y1186 = n6801 ;
  assign y1187 = n6810 ;
  assign y1188 = ~n6814 ;
  assign y1189 = ~n6816 ;
  assign y1190 = n6820 ;
  assign y1191 = ~1'b0 ;
  assign y1192 = ~n6837 ;
  assign y1193 = ~n6846 ;
  assign y1194 = n6850 ;
  assign y1195 = ~n6851 ;
  assign y1196 = n6853 ;
  assign y1197 = n6865 ;
  assign y1198 = ~1'b0 ;
  assign y1199 = n6868 ;
  assign y1200 = ~1'b0 ;
  assign y1201 = ~n6882 ;
  assign y1202 = n6892 ;
  assign y1203 = ~n6895 ;
  assign y1204 = n6911 ;
  assign y1205 = n6912 ;
  assign y1206 = ~n6914 ;
  assign y1207 = n6920 ;
  assign y1208 = ~n6925 ;
  assign y1209 = n6934 ;
  assign y1210 = n6942 ;
  assign y1211 = n6954 ;
  assign y1212 = ~n6957 ;
  assign y1213 = n6961 ;
  assign y1214 = n6974 ;
  assign y1215 = ~n6980 ;
  assign y1216 = ~n6982 ;
  assign y1217 = ~1'b0 ;
  assign y1218 = n7001 ;
  assign y1219 = ~n7005 ;
  assign y1220 = ~n7015 ;
  assign y1221 = ~n7016 ;
  assign y1222 = ~n7024 ;
  assign y1223 = n7027 ;
  assign y1224 = ~n7028 ;
  assign y1225 = n7030 ;
  assign y1226 = n7036 ;
  assign y1227 = n7041 ;
  assign y1228 = n7044 ;
  assign y1229 = ~n7045 ;
  assign y1230 = n7049 ;
  assign y1231 = ~n7051 ;
  assign y1232 = n7073 ;
  assign y1233 = ~1'b0 ;
  assign y1234 = ~1'b0 ;
  assign y1235 = ~n7081 ;
  assign y1236 = ~1'b0 ;
  assign y1237 = ~n7092 ;
  assign y1238 = ~n7096 ;
  assign y1239 = n7103 ;
  assign y1240 = n7106 ;
  assign y1241 = ~n7108 ;
  assign y1242 = ~n7116 ;
  assign y1243 = n7120 ;
  assign y1244 = ~n7121 ;
  assign y1245 = ~n7126 ;
  assign y1246 = n7133 ;
  assign y1247 = n7135 ;
  assign y1248 = n7147 ;
  assign y1249 = ~n7148 ;
  assign y1250 = ~n7163 ;
  assign y1251 = ~n7174 ;
  assign y1252 = ~n7180 ;
  assign y1253 = n7191 ;
  assign y1254 = ~n7200 ;
  assign y1255 = n7218 ;
  assign y1256 = n7233 ;
  assign y1257 = ~n7242 ;
  assign y1258 = ~n7252 ;
  assign y1259 = ~n7257 ;
  assign y1260 = n7263 ;
  assign y1261 = ~n7265 ;
  assign y1262 = n7269 ;
  assign y1263 = ~n7272 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = n7276 ;
  assign y1266 = ~n7312 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~n7321 ;
  assign y1269 = n7326 ;
  assign y1270 = n7332 ;
  assign y1271 = n7339 ;
  assign y1272 = n7345 ;
  assign y1273 = n7347 ;
  assign y1274 = n7357 ;
  assign y1275 = ~n7360 ;
  assign y1276 = ~n7366 ;
  assign y1277 = n7374 ;
  assign y1278 = ~n7381 ;
  assign y1279 = ~1'b0 ;
  assign y1280 = ~n7391 ;
  assign y1281 = n7397 ;
  assign y1282 = n7398 ;
  assign y1283 = n7409 ;
  assign y1284 = n7413 ;
  assign y1285 = n7420 ;
  assign y1286 = ~n7423 ;
  assign y1287 = ~n7429 ;
  assign y1288 = ~n7435 ;
  assign y1289 = ~n7448 ;
  assign y1290 = ~n7449 ;
  assign y1291 = ~n7452 ;
  assign y1292 = ~n7453 ;
  assign y1293 = n7466 ;
  assign y1294 = ~n7470 ;
  assign y1295 = ~n7481 ;
  assign y1296 = n7496 ;
  assign y1297 = n7501 ;
  assign y1298 = ~n7531 ;
  assign y1299 = n7537 ;
  assign y1300 = ~1'b0 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = n7547 ;
  assign y1303 = n7551 ;
  assign y1304 = ~n7561 ;
  assign y1305 = n7565 ;
  assign y1306 = ~n7569 ;
  assign y1307 = n7581 ;
  assign y1308 = n7590 ;
  assign y1309 = ~n7618 ;
  assign y1310 = n7620 ;
  assign y1311 = ~1'b0 ;
  assign y1312 = n7622 ;
  assign y1313 = n7625 ;
  assign y1314 = ~n7631 ;
  assign y1315 = ~n7637 ;
  assign y1316 = n7642 ;
  assign y1317 = n7644 ;
  assign y1318 = n7653 ;
  assign y1319 = n7657 ;
  assign y1320 = n7659 ;
  assign y1321 = ~n7661 ;
  assign y1322 = n7677 ;
  assign y1323 = ~1'b0 ;
  assign y1324 = n7683 ;
  assign y1325 = n7687 ;
  assign y1326 = n7696 ;
  assign y1327 = ~n7697 ;
  assign y1328 = n7701 ;
  assign y1329 = ~n7703 ;
  assign y1330 = n7711 ;
  assign y1331 = ~n7722 ;
  assign y1332 = n7724 ;
  assign y1333 = n7737 ;
  assign y1334 = n7744 ;
  assign y1335 = n7754 ;
  assign y1336 = n7756 ;
  assign y1337 = ~n7758 ;
  assign y1338 = ~n7779 ;
  assign y1339 = n7805 ;
  assign y1340 = n7809 ;
  assign y1341 = ~n7812 ;
  assign y1342 = ~n7821 ;
  assign y1343 = ~n7822 ;
  assign y1344 = n7824 ;
  assign y1345 = ~n7827 ;
  assign y1346 = n7834 ;
  assign y1347 = n7840 ;
  assign y1348 = n7844 ;
  assign y1349 = n7848 ;
  assign y1350 = ~1'b0 ;
  assign y1351 = n7851 ;
  assign y1352 = ~1'b0 ;
  assign y1353 = ~n7869 ;
  assign y1354 = n7873 ;
  assign y1355 = ~n7877 ;
  assign y1356 = n7882 ;
  assign y1357 = n7890 ;
  assign y1358 = n7900 ;
  assign y1359 = n7903 ;
  assign y1360 = n7908 ;
  assign y1361 = n7920 ;
  assign y1362 = ~1'b0 ;
  assign y1363 = n7923 ;
  assign y1364 = n7927 ;
  assign y1365 = ~n7928 ;
  assign y1366 = ~n7930 ;
  assign y1367 = n7931 ;
  assign y1368 = n7932 ;
  assign y1369 = ~n7934 ;
  assign y1370 = ~1'b0 ;
  assign y1371 = ~n7949 ;
  assign y1372 = ~n7951 ;
  assign y1373 = n7954 ;
  assign y1374 = ~n7959 ;
  assign y1375 = n7969 ;
  assign y1376 = n7971 ;
  assign y1377 = ~n7972 ;
  assign y1378 = n7981 ;
  assign y1379 = ~n7988 ;
  assign y1380 = ~n8000 ;
  assign y1381 = n8029 ;
  assign y1382 = n8041 ;
  assign y1383 = ~n8044 ;
  assign y1384 = ~n8047 ;
  assign y1385 = ~n8050 ;
  assign y1386 = ~n8053 ;
  assign y1387 = n8054 ;
  assign y1388 = ~n8058 ;
  assign y1389 = n8061 ;
  assign y1390 = ~n8062 ;
  assign y1391 = ~1'b0 ;
  assign y1392 = ~n8063 ;
  assign y1393 = n8064 ;
  assign y1394 = ~n8069 ;
  assign y1395 = ~n8070 ;
  assign y1396 = n8072 ;
  assign y1397 = n8075 ;
  assign y1398 = ~n8086 ;
  assign y1399 = ~n8106 ;
  assign y1400 = ~n8111 ;
  assign y1401 = ~n8123 ;
  assign y1402 = n8125 ;
  assign y1403 = n8134 ;
  assign y1404 = n8139 ;
  assign y1405 = ~n8143 ;
  assign y1406 = n8158 ;
  assign y1407 = ~n8165 ;
  assign y1408 = n8166 ;
  assign y1409 = n8171 ;
  assign y1410 = ~n8173 ;
  assign y1411 = n8183 ;
  assign y1412 = n8189 ;
  assign y1413 = ~n8190 ;
  assign y1414 = ~n8196 ;
  assign y1415 = n8207 ;
  assign y1416 = ~n8212 ;
  assign y1417 = ~n8223 ;
  assign y1418 = n8224 ;
  assign y1419 = n8236 ;
  assign y1420 = ~1'b0 ;
  assign y1421 = ~n8246 ;
  assign y1422 = ~1'b0 ;
  assign y1423 = n8261 ;
  assign y1424 = n8266 ;
  assign y1425 = ~n8276 ;
  assign y1426 = ~n8284 ;
  assign y1427 = ~n8291 ;
  assign y1428 = ~n8292 ;
  assign y1429 = n8298 ;
  assign y1430 = ~n8304 ;
  assign y1431 = ~n8307 ;
  assign y1432 = ~n8313 ;
  assign y1433 = ~n8314 ;
  assign y1434 = n8323 ;
  assign y1435 = n8329 ;
  assign y1436 = ~n8337 ;
  assign y1437 = ~n8345 ;
  assign y1438 = n8353 ;
  assign y1439 = ~1'b0 ;
  assign y1440 = ~n8354 ;
  assign y1441 = ~n8360 ;
  assign y1442 = n8367 ;
  assign y1443 = n8370 ;
  assign y1444 = ~n8375 ;
  assign y1445 = n8377 ;
  assign y1446 = n8380 ;
  assign y1447 = ~n8390 ;
  assign y1448 = n8398 ;
  assign y1449 = ~n8406 ;
  assign y1450 = ~n8407 ;
  assign y1451 = n8408 ;
  assign y1452 = ~n8409 ;
  assign y1453 = ~n8411 ;
  assign y1454 = ~n8415 ;
  assign y1455 = ~n8418 ;
  assign y1456 = ~n8421 ;
  assign y1457 = n8423 ;
  assign y1458 = ~1'b0 ;
  assign y1459 = n8449 ;
  assign y1460 = ~n8453 ;
  assign y1461 = n8454 ;
  assign y1462 = ~n8460 ;
  assign y1463 = ~n8476 ;
  assign y1464 = n8478 ;
  assign y1465 = ~n8481 ;
  assign y1466 = n8490 ;
  assign y1467 = ~n8496 ;
  assign y1468 = ~n8498 ;
  assign y1469 = ~1'b0 ;
  assign y1470 = n8499 ;
  assign y1471 = n8500 ;
  assign y1472 = n8510 ;
  assign y1473 = ~n8513 ;
  assign y1474 = ~n8515 ;
  assign y1475 = n8522 ;
  assign y1476 = ~n8525 ;
  assign y1477 = ~n8531 ;
  assign y1478 = n8536 ;
  assign y1479 = n8539 ;
  assign y1480 = ~n8547 ;
  assign y1481 = n8548 ;
  assign y1482 = ~n8549 ;
  assign y1483 = ~n8558 ;
  assign y1484 = n8562 ;
  assign y1485 = n8567 ;
  assign y1486 = n8570 ;
  assign y1487 = n8574 ;
  assign y1488 = ~n8578 ;
  assign y1489 = n8579 ;
  assign y1490 = n8584 ;
  assign y1491 = n8589 ;
  assign y1492 = ~n8594 ;
  assign y1493 = n8597 ;
  assign y1494 = n8598 ;
  assign y1495 = n8601 ;
  assign y1496 = n8616 ;
  assign y1497 = n8622 ;
  assign y1498 = ~n8627 ;
  assign y1499 = n8632 ;
  assign y1500 = ~1'b0 ;
  assign y1501 = n8639 ;
  assign y1502 = ~n8644 ;
  assign y1503 = n8650 ;
  assign y1504 = ~1'b0 ;
  assign y1505 = ~n8656 ;
  assign y1506 = n8658 ;
  assign y1507 = n8661 ;
  assign y1508 = n8663 ;
  assign y1509 = ~n8670 ;
  assign y1510 = ~n8671 ;
  assign y1511 = n8672 ;
  assign y1512 = ~n8673 ;
  assign y1513 = ~n8675 ;
  assign y1514 = ~n8681 ;
  assign y1515 = ~n8685 ;
  assign y1516 = n8704 ;
  assign y1517 = ~n8705 ;
  assign y1518 = ~n8707 ;
  assign y1519 = ~n8712 ;
  assign y1520 = n8715 ;
  assign y1521 = n8722 ;
  assign y1522 = ~n8723 ;
  assign y1523 = ~n8730 ;
  assign y1524 = ~n8751 ;
  assign y1525 = n8752 ;
  assign y1526 = n8753 ;
  assign y1527 = ~1'b0 ;
  assign y1528 = n8756 ;
  assign y1529 = ~n8771 ;
  assign y1530 = ~n8776 ;
  assign y1531 = n8779 ;
  assign y1532 = ~n8793 ;
  assign y1533 = ~n8796 ;
  assign y1534 = ~1'b0 ;
  assign y1535 = ~n8801 ;
  assign y1536 = ~1'b0 ;
  assign y1537 = n8805 ;
  assign y1538 = ~n8811 ;
  assign y1539 = n8817 ;
  assign y1540 = n8821 ;
  assign y1541 = n8832 ;
  assign y1542 = n8843 ;
  assign y1543 = ~n8850 ;
  assign y1544 = n8864 ;
  assign y1545 = ~n8875 ;
  assign y1546 = ~n8880 ;
  assign y1547 = n8883 ;
  assign y1548 = ~n8891 ;
  assign y1549 = ~n8895 ;
  assign y1550 = n8898 ;
  assign y1551 = n8913 ;
  assign y1552 = ~n8918 ;
  assign y1553 = n8923 ;
  assign y1554 = n8925 ;
  assign y1555 = n8936 ;
  assign y1556 = ~n8937 ;
  assign y1557 = n8939 ;
  assign y1558 = n8948 ;
  assign y1559 = n8956 ;
  assign y1560 = n8963 ;
  assign y1561 = ~n8970 ;
  assign y1562 = n8979 ;
  assign y1563 = ~n8987 ;
  assign y1564 = ~n9003 ;
  assign y1565 = ~n9015 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = n9019 ;
  assign y1568 = ~n9028 ;
  assign y1569 = ~n9032 ;
  assign y1570 = n9037 ;
  assign y1571 = ~n9049 ;
  assign y1572 = ~1'b0 ;
  assign y1573 = ~n9050 ;
  assign y1574 = n9056 ;
  assign y1575 = ~n9087 ;
  assign y1576 = ~n9088 ;
  assign y1577 = ~1'b0 ;
  assign y1578 = n9095 ;
  assign y1579 = ~n9099 ;
  assign y1580 = n9101 ;
  assign y1581 = ~1'b0 ;
  assign y1582 = n9102 ;
  assign y1583 = ~n9109 ;
  assign y1584 = n9112 ;
  assign y1585 = n9117 ;
  assign y1586 = ~1'b0 ;
  assign y1587 = ~n9118 ;
  assign y1588 = ~n9127 ;
  assign y1589 = n9133 ;
  assign y1590 = ~n9142 ;
  assign y1591 = ~n9146 ;
  assign y1592 = ~n7470 ;
  assign y1593 = ~n9159 ;
  assign y1594 = ~n9161 ;
  assign y1595 = ~n9165 ;
  assign y1596 = ~n9175 ;
  assign y1597 = ~1'b0 ;
  assign y1598 = ~1'b0 ;
  assign y1599 = ~n9179 ;
  assign y1600 = n9184 ;
  assign y1601 = n9186 ;
  assign y1602 = ~n9200 ;
  assign y1603 = ~n9205 ;
  assign y1604 = ~n9211 ;
  assign y1605 = n9212 ;
  assign y1606 = n9215 ;
  assign y1607 = ~n9225 ;
  assign y1608 = ~n9230 ;
  assign y1609 = n9234 ;
  assign y1610 = ~1'b0 ;
  assign y1611 = ~1'b0 ;
  assign y1612 = n9241 ;
  assign y1613 = n9242 ;
  assign y1614 = ~1'b0 ;
  assign y1615 = ~n9251 ;
  assign y1616 = n9255 ;
  assign y1617 = n9260 ;
  assign y1618 = ~n9263 ;
  assign y1619 = n9275 ;
  assign y1620 = ~n9277 ;
  assign y1621 = n9289 ;
  assign y1622 = ~n9291 ;
  assign y1623 = ~n9293 ;
  assign y1624 = n9317 ;
  assign y1625 = ~n9322 ;
  assign y1626 = ~n9335 ;
  assign y1627 = ~n9336 ;
  assign y1628 = n9346 ;
  assign y1629 = ~n9351 ;
  assign y1630 = ~n9355 ;
  assign y1631 = ~n9367 ;
  assign y1632 = ~n9370 ;
  assign y1633 = ~1'b0 ;
  assign y1634 = ~n9371 ;
  assign y1635 = ~n9373 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = ~n9374 ;
  assign y1638 = ~n9383 ;
  assign y1639 = ~n9390 ;
  assign y1640 = ~n9393 ;
  assign y1641 = n9398 ;
  assign y1642 = ~n9405 ;
  assign y1643 = ~n9413 ;
  assign y1644 = ~n9417 ;
  assign y1645 = n9420 ;
  assign y1646 = ~n9423 ;
  assign y1647 = ~1'b0 ;
  assign y1648 = n9433 ;
  assign y1649 = ~n9442 ;
  assign y1650 = ~n9444 ;
  assign y1651 = ~n9453 ;
  assign y1652 = n9459 ;
  assign y1653 = n9463 ;
  assign y1654 = n9471 ;
  assign y1655 = n9474 ;
  assign y1656 = n9483 ;
  assign y1657 = n9487 ;
  assign y1658 = n9503 ;
  assign y1659 = n9508 ;
  assign y1660 = ~n9513 ;
  assign y1661 = n9519 ;
  assign y1662 = n9525 ;
  assign y1663 = n9528 ;
  assign y1664 = ~n9531 ;
  assign y1665 = n9533 ;
  assign y1666 = n9539 ;
  assign y1667 = ~n9543 ;
  assign y1668 = n9546 ;
  assign y1669 = ~n9554 ;
  assign y1670 = n9561 ;
  assign y1671 = ~n9565 ;
  assign y1672 = n9577 ;
  assign y1673 = ~n9617 ;
  assign y1674 = n9621 ;
  assign y1675 = n9634 ;
  assign y1676 = ~n9636 ;
  assign y1677 = ~n9644 ;
  assign y1678 = n9645 ;
  assign y1679 = n9647 ;
  assign y1680 = n9651 ;
  assign y1681 = n9652 ;
  assign y1682 = n9659 ;
  assign y1683 = ~n9663 ;
  assign y1684 = ~n9669 ;
  assign y1685 = ~n9671 ;
  assign y1686 = ~1'b0 ;
  assign y1687 = n9672 ;
  assign y1688 = ~n9674 ;
  assign y1689 = ~n9679 ;
  assign y1690 = n9686 ;
  assign y1691 = ~n9698 ;
  assign y1692 = n9701 ;
  assign y1693 = n9702 ;
  assign y1694 = ~n9705 ;
  assign y1695 = ~n9708 ;
  assign y1696 = n9709 ;
  assign y1697 = ~1'b0 ;
  assign y1698 = ~n9715 ;
  assign y1699 = ~n9719 ;
  assign y1700 = n9730 ;
  assign y1701 = ~n9731 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = ~n9733 ;
  assign y1704 = ~n9746 ;
  assign y1705 = ~n9749 ;
  assign y1706 = n9755 ;
  assign y1707 = n9759 ;
  assign y1708 = n9762 ;
  assign y1709 = n9770 ;
  assign y1710 = ~n9785 ;
  assign y1711 = n9794 ;
  assign y1712 = ~n9795 ;
  assign y1713 = ~n9800 ;
  assign y1714 = n9806 ;
  assign y1715 = ~n9812 ;
  assign y1716 = n9815 ;
  assign y1717 = ~n9830 ;
  assign y1718 = ~n4735 ;
  assign y1719 = n9832 ;
  assign y1720 = ~n9836 ;
  assign y1721 = n9838 ;
  assign y1722 = ~n9846 ;
  assign y1723 = n9847 ;
  assign y1724 = ~n9856 ;
  assign y1725 = ~n9863 ;
  assign y1726 = ~n9867 ;
  assign y1727 = n9881 ;
  assign y1728 = ~n9889 ;
  assign y1729 = n9909 ;
  assign y1730 = n9916 ;
  assign y1731 = ~n9918 ;
  assign y1732 = ~n9919 ;
  assign y1733 = ~n9921 ;
  assign y1734 = ~n9925 ;
  assign y1735 = n9927 ;
  assign y1736 = n9928 ;
  assign y1737 = n9929 ;
  assign y1738 = n9934 ;
  assign y1739 = n9936 ;
  assign y1740 = ~n9943 ;
  assign y1741 = n9947 ;
  assign y1742 = ~n9950 ;
  assign y1743 = n9973 ;
  assign y1744 = ~n9977 ;
  assign y1745 = n9989 ;
  assign y1746 = ~n9992 ;
  assign y1747 = n9994 ;
  assign y1748 = n9998 ;
  assign y1749 = ~n10003 ;
  assign y1750 = ~n10021 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = n10025 ;
  assign y1753 = ~n10026 ;
  assign y1754 = n10030 ;
  assign y1755 = ~n10039 ;
  assign y1756 = n10041 ;
  assign y1757 = n10056 ;
  assign y1758 = ~n10061 ;
  assign y1759 = ~n10065 ;
  assign y1760 = n10069 ;
  assign y1761 = ~n10081 ;
  assign y1762 = n10088 ;
  assign y1763 = ~n10093 ;
  assign y1764 = n10110 ;
  assign y1765 = ~n10118 ;
  assign y1766 = ~1'b0 ;
  assign y1767 = ~n10127 ;
  assign y1768 = n10138 ;
  assign y1769 = ~n10144 ;
  assign y1770 = ~n10149 ;
  assign y1771 = ~n5814 ;
  assign y1772 = ~n10157 ;
  assign y1773 = n10160 ;
  assign y1774 = ~n10163 ;
  assign y1775 = ~n10164 ;
  assign y1776 = n10165 ;
  assign y1777 = n10166 ;
  assign y1778 = n10178 ;
  assign y1779 = n10180 ;
  assign y1780 = n10185 ;
  assign y1781 = ~n10188 ;
  assign y1782 = ~n10195 ;
  assign y1783 = ~n10207 ;
  assign y1784 = ~n10208 ;
  assign y1785 = n10217 ;
  assign y1786 = n10223 ;
  assign y1787 = n10230 ;
  assign y1788 = ~n10238 ;
  assign y1789 = ~n10254 ;
  assign y1790 = ~n10270 ;
  assign y1791 = n10271 ;
  assign y1792 = ~n10275 ;
  assign y1793 = ~n10278 ;
  assign y1794 = n10285 ;
  assign y1795 = n10291 ;
  assign y1796 = n10293 ;
  assign y1797 = n10304 ;
  assign y1798 = n10308 ;
  assign y1799 = ~n10312 ;
  assign y1800 = n10313 ;
  assign y1801 = ~n10315 ;
  assign y1802 = ~n10318 ;
  assign y1803 = n10324 ;
  assign y1804 = n10331 ;
  assign y1805 = n10333 ;
  assign y1806 = n10342 ;
  assign y1807 = n10346 ;
  assign y1808 = ~n10348 ;
  assign y1809 = n10351 ;
  assign y1810 = n10352 ;
  assign y1811 = ~n10357 ;
  assign y1812 = ~1'b0 ;
  assign y1813 = ~n10370 ;
  assign y1814 = ~n10379 ;
  assign y1815 = n10382 ;
  assign y1816 = ~n10399 ;
  assign y1817 = n10400 ;
  assign y1818 = ~n10405 ;
  assign y1819 = ~1'b0 ;
  assign y1820 = n10410 ;
  assign y1821 = n10415 ;
  assign y1822 = n10420 ;
  assign y1823 = n10422 ;
  assign y1824 = ~n10423 ;
  assign y1825 = ~n10430 ;
  assign y1826 = ~n10432 ;
  assign y1827 = n10441 ;
  assign y1828 = ~n10443 ;
  assign y1829 = ~1'b0 ;
  assign y1830 = ~n10450 ;
  assign y1831 = n10462 ;
  assign y1832 = ~n10468 ;
  assign y1833 = ~n10471 ;
  assign y1834 = ~n10472 ;
  assign y1835 = n10473 ;
  assign y1836 = n10474 ;
  assign y1837 = n10486 ;
  assign y1838 = n10489 ;
  assign y1839 = n10492 ;
  assign y1840 = ~1'b0 ;
  assign y1841 = n10501 ;
  assign y1842 = ~n10507 ;
  assign y1843 = ~n10512 ;
  assign y1844 = ~n10520 ;
  assign y1845 = ~n10527 ;
  assign y1846 = ~n10528 ;
  assign y1847 = ~n10533 ;
  assign y1848 = n10534 ;
  assign y1849 = ~1'b0 ;
  assign y1850 = ~n10546 ;
  assign y1851 = n10553 ;
  assign y1852 = ~n10561 ;
  assign y1853 = n10568 ;
  assign y1854 = n10577 ;
  assign y1855 = n10581 ;
  assign y1856 = ~n10588 ;
  assign y1857 = ~n10599 ;
  assign y1858 = n10602 ;
  assign y1859 = n10610 ;
  assign y1860 = n10611 ;
  assign y1861 = n10613 ;
  assign y1862 = ~n10615 ;
  assign y1863 = n10616 ;
  assign y1864 = n10623 ;
  assign y1865 = ~n10625 ;
  assign y1866 = ~n10626 ;
  assign y1867 = n10635 ;
  assign y1868 = n10641 ;
  assign y1869 = ~1'b0 ;
  assign y1870 = ~n10644 ;
  assign y1871 = n10659 ;
  assign y1872 = ~n10662 ;
  assign y1873 = ~n10666 ;
  assign y1874 = ~n10667 ;
  assign y1875 = ~n10670 ;
  assign y1876 = ~n10675 ;
  assign y1877 = n10676 ;
  assign y1878 = ~n10677 ;
  assign y1879 = n10680 ;
  assign y1880 = ~n10681 ;
  assign y1881 = ~n10693 ;
  assign y1882 = ~n10699 ;
  assign y1883 = ~n10707 ;
  assign y1884 = n10715 ;
  assign y1885 = n10720 ;
  assign y1886 = ~n10729 ;
  assign y1887 = ~n10735 ;
  assign y1888 = n10741 ;
  assign y1889 = n10746 ;
  assign y1890 = ~n10751 ;
  assign y1891 = n10753 ;
  assign y1892 = ~n10757 ;
  assign y1893 = n10770 ;
  assign y1894 = ~n10772 ;
  assign y1895 = ~n10776 ;
  assign y1896 = n10781 ;
  assign y1897 = ~n10788 ;
  assign y1898 = ~n10790 ;
  assign y1899 = n10796 ;
  assign y1900 = n10801 ;
  assign y1901 = ~1'b0 ;
  assign y1902 = n10805 ;
  assign y1903 = ~n10325 ;
  assign y1904 = ~n10807 ;
  assign y1905 = ~n10821 ;
  assign y1906 = n10826 ;
  assign y1907 = n10832 ;
  assign y1908 = ~n10846 ;
  assign y1909 = ~n10847 ;
  assign y1910 = ~n10852 ;
  assign y1911 = ~n10853 ;
  assign y1912 = n10861 ;
  assign y1913 = ~n10872 ;
  assign y1914 = ~1'b0 ;
  assign y1915 = n10879 ;
  assign y1916 = ~n10886 ;
  assign y1917 = n10891 ;
  assign y1918 = n10902 ;
  assign y1919 = n10904 ;
  assign y1920 = n10915 ;
  assign y1921 = n10960 ;
  assign y1922 = ~n10963 ;
  assign y1923 = ~n10965 ;
  assign y1924 = ~n10971 ;
  assign y1925 = n10972 ;
  assign y1926 = n11001 ;
  assign y1927 = n11009 ;
  assign y1928 = n11031 ;
  assign y1929 = n11032 ;
  assign y1930 = ~n11038 ;
  assign y1931 = ~n11041 ;
  assign y1932 = n11042 ;
  assign y1933 = ~n11043 ;
  assign y1934 = n11050 ;
  assign y1935 = ~n11066 ;
  assign y1936 = ~n11080 ;
  assign y1937 = ~n11086 ;
  assign y1938 = n11089 ;
  assign y1939 = ~n11093 ;
  assign y1940 = n11104 ;
  assign y1941 = ~1'b0 ;
  assign y1942 = ~n11110 ;
  assign y1943 = n11116 ;
  assign y1944 = n11118 ;
  assign y1945 = ~n11119 ;
  assign y1946 = ~n11120 ;
  assign y1947 = n11130 ;
  assign y1948 = n11138 ;
  assign y1949 = ~n11145 ;
  assign y1950 = ~n11149 ;
  assign y1951 = ~n11155 ;
  assign y1952 = ~n11156 ;
  assign y1953 = n11162 ;
  assign y1954 = n11171 ;
  assign y1955 = ~n11177 ;
  assign y1956 = n11179 ;
  assign y1957 = n11182 ;
  assign y1958 = ~n11184 ;
  assign y1959 = ~n11186 ;
  assign y1960 = ~1'b0 ;
  assign y1961 = ~1'b0 ;
  assign y1962 = n11190 ;
  assign y1963 = ~n11192 ;
  assign y1964 = n11206 ;
  assign y1965 = n11208 ;
  assign y1966 = n11218 ;
  assign y1967 = n11222 ;
  assign y1968 = ~n11223 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = n11230 ;
  assign y1971 = ~n11234 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = n11238 ;
  assign y1974 = n11240 ;
  assign y1975 = n11245 ;
  assign y1976 = n11246 ;
  assign y1977 = ~n11248 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = ~n11254 ;
  assign y1980 = ~n11255 ;
  assign y1981 = n11256 ;
  assign y1982 = ~n11257 ;
  assign y1983 = n11259 ;
  assign y1984 = n11267 ;
  assign y1985 = ~n11271 ;
  assign y1986 = ~n11279 ;
  assign y1987 = ~n11298 ;
  assign y1988 = n11305 ;
  assign y1989 = n11320 ;
  assign y1990 = n11322 ;
  assign y1991 = n11326 ;
  assign y1992 = ~n11329 ;
  assign y1993 = ~n11330 ;
  assign y1994 = ~n11335 ;
  assign y1995 = n11336 ;
  assign y1996 = ~n11360 ;
  assign y1997 = n11364 ;
  assign y1998 = ~n11366 ;
  assign y1999 = ~n11369 ;
  assign y2000 = n11388 ;
  assign y2001 = ~n11399 ;
  assign y2002 = n11402 ;
  assign y2003 = n11422 ;
  assign y2004 = n11426 ;
  assign y2005 = ~n11445 ;
  assign y2006 = ~n11453 ;
  assign y2007 = n11467 ;
  assign y2008 = n11469 ;
  assign y2009 = n11477 ;
  assign y2010 = ~n11483 ;
  assign y2011 = ~n11485 ;
  assign y2012 = ~n11492 ;
  assign y2013 = ~n11495 ;
  assign y2014 = ~n11498 ;
  assign y2015 = ~1'b0 ;
  assign y2016 = ~n11505 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = ~n11510 ;
  assign y2019 = n11512 ;
  assign y2020 = ~1'b0 ;
  assign y2021 = n11520 ;
  assign y2022 = ~n11522 ;
  assign y2023 = ~n11537 ;
  assign y2024 = ~n11538 ;
  assign y2025 = n11542 ;
  assign y2026 = ~n11545 ;
  assign y2027 = ~n11546 ;
  assign y2028 = ~n11556 ;
  assign y2029 = n11558 ;
  assign y2030 = ~n11560 ;
  assign y2031 = ~1'b0 ;
  assign y2032 = n11563 ;
  assign y2033 = n11569 ;
  assign y2034 = n11587 ;
  assign y2035 = ~n11595 ;
  assign y2036 = ~n11622 ;
  assign y2037 = ~n11623 ;
  assign y2038 = ~n11628 ;
  assign y2039 = n11638 ;
  assign y2040 = ~n11639 ;
  assign y2041 = ~n11640 ;
  assign y2042 = n11643 ;
  assign y2043 = ~1'b0 ;
  assign y2044 = ~1'b0 ;
  assign y2045 = n11649 ;
  assign y2046 = ~n11652 ;
  assign y2047 = ~n11662 ;
  assign y2048 = n11666 ;
  assign y2049 = ~n11669 ;
  assign y2050 = n11670 ;
  assign y2051 = n11676 ;
  assign y2052 = ~n11682 ;
  assign y2053 = n11693 ;
  assign y2054 = ~n11700 ;
  assign y2055 = ~1'b0 ;
  assign y2056 = ~n11710 ;
  assign y2057 = n11713 ;
  assign y2058 = ~n11719 ;
  assign y2059 = ~n11721 ;
  assign y2060 = ~n11725 ;
  assign y2061 = n11726 ;
  assign y2062 = n11731 ;
  assign y2063 = ~1'b0 ;
  assign y2064 = ~n11737 ;
  assign y2065 = n11748 ;
  assign y2066 = ~1'b0 ;
  assign y2067 = n11751 ;
  assign y2068 = n11752 ;
  assign y2069 = n11765 ;
  assign y2070 = ~n11768 ;
  assign y2071 = ~n11771 ;
  assign y2072 = n11774 ;
  assign y2073 = n11777 ;
  assign y2074 = n11779 ;
  assign y2075 = n11782 ;
  assign y2076 = ~n11790 ;
  assign y2077 = ~n11793 ;
  assign y2078 = ~n11795 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = ~n11797 ;
  assign y2081 = ~n11803 ;
  assign y2082 = n11805 ;
  assign y2083 = ~n11811 ;
  assign y2084 = ~n11815 ;
  assign y2085 = ~n11817 ;
  assign y2086 = ~n11827 ;
  assign y2087 = n11831 ;
  assign y2088 = n11837 ;
  assign y2089 = n11843 ;
  assign y2090 = n11844 ;
  assign y2091 = ~n11853 ;
  assign y2092 = n11859 ;
  assign y2093 = ~n11869 ;
  assign y2094 = ~n11870 ;
  assign y2095 = ~n11873 ;
  assign y2096 = n11874 ;
  assign y2097 = ~n11894 ;
  assign y2098 = n11904 ;
  assign y2099 = ~n11905 ;
  assign y2100 = n11913 ;
  assign y2101 = n11920 ;
  assign y2102 = ~1'b0 ;
  assign y2103 = ~n11924 ;
  assign y2104 = ~n11932 ;
  assign y2105 = ~n11938 ;
  assign y2106 = n11946 ;
  assign y2107 = n11955 ;
  assign y2108 = n11956 ;
  assign y2109 = n11959 ;
  assign y2110 = ~n11960 ;
  assign y2111 = ~n11967 ;
  assign y2112 = ~n11975 ;
  assign y2113 = n11981 ;
  assign y2114 = ~1'b0 ;
  assign y2115 = n11986 ;
  assign y2116 = ~n11992 ;
  assign y2117 = ~n11994 ;
  assign y2118 = n11996 ;
  assign y2119 = n11999 ;
  assign y2120 = ~n12000 ;
  assign y2121 = ~n12007 ;
  assign y2122 = ~n12009 ;
  assign y2123 = n12011 ;
  assign y2124 = ~n12016 ;
  assign y2125 = ~n12029 ;
  assign y2126 = n12032 ;
  assign y2127 = n12033 ;
  assign y2128 = n12035 ;
  assign y2129 = n12041 ;
  assign y2130 = n12050 ;
  assign y2131 = ~n12051 ;
  assign y2132 = ~1'b0 ;
  assign y2133 = ~n12058 ;
  assign y2134 = n12061 ;
  assign y2135 = n12075 ;
  assign y2136 = n12081 ;
  assign y2137 = ~n12088 ;
  assign y2138 = ~n12095 ;
  assign y2139 = ~1'b0 ;
  assign y2140 = ~n12098 ;
  assign y2141 = ~n12102 ;
  assign y2142 = n12106 ;
  assign y2143 = ~n12113 ;
  assign y2144 = n12116 ;
  assign y2145 = n12119 ;
  assign y2146 = n12122 ;
  assign y2147 = ~n12127 ;
  assign y2148 = ~n12134 ;
  assign y2149 = n12144 ;
  assign y2150 = ~1'b0 ;
  assign y2151 = ~n12147 ;
  assign y2152 = n12155 ;
  assign y2153 = n12160 ;
  assign y2154 = ~n12161 ;
  assign y2155 = n12164 ;
  assign y2156 = ~n12169 ;
  assign y2157 = ~n12172 ;
  assign y2158 = ~n12175 ;
  assign y2159 = ~n12177 ;
  assign y2160 = n12181 ;
  assign y2161 = n12189 ;
  assign y2162 = ~n12194 ;
  assign y2163 = ~n12197 ;
  assign y2164 = n12206 ;
  assign y2165 = n12209 ;
  assign y2166 = ~n12210 ;
  assign y2167 = ~n12217 ;
  assign y2168 = n12220 ;
  assign y2169 = n12225 ;
  assign y2170 = ~n12226 ;
  assign y2171 = ~n12227 ;
  assign y2172 = n12229 ;
  assign y2173 = n12231 ;
  assign y2174 = ~1'b0 ;
  assign y2175 = n12242 ;
  assign y2176 = ~n12264 ;
  assign y2177 = ~n12270 ;
  assign y2178 = n12275 ;
  assign y2179 = ~n12277 ;
  assign y2180 = ~n12279 ;
  assign y2181 = n12285 ;
  assign y2182 = n12289 ;
  assign y2183 = ~n12297 ;
  assign y2184 = n12298 ;
  assign y2185 = ~n12304 ;
  assign y2186 = n12316 ;
  assign y2187 = ~n12318 ;
  assign y2188 = ~n12327 ;
  assign y2189 = n12328 ;
  assign y2190 = n12330 ;
  assign y2191 = ~n12331 ;
  assign y2192 = ~1'b0 ;
  assign y2193 = ~n12342 ;
  assign y2194 = ~n12354 ;
  assign y2195 = n12359 ;
  assign y2196 = ~n12366 ;
  assign y2197 = ~1'b0 ;
  assign y2198 = ~n12378 ;
  assign y2199 = n12379 ;
  assign y2200 = ~n12380 ;
  assign y2201 = ~n12400 ;
  assign y2202 = n12402 ;
  assign y2203 = n12406 ;
  assign y2204 = ~n12410 ;
  assign y2205 = ~1'b0 ;
  assign y2206 = ~n12415 ;
  assign y2207 = ~n12416 ;
  assign y2208 = n12423 ;
  assign y2209 = ~n12430 ;
  assign y2210 = ~n12435 ;
  assign y2211 = n12440 ;
  assign y2212 = n12442 ;
  assign y2213 = n12446 ;
  assign y2214 = ~n12450 ;
  assign y2215 = ~n12457 ;
  assign y2216 = ~1'b0 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = ~n12459 ;
  assign y2219 = ~n12461 ;
  assign y2220 = n12475 ;
  assign y2221 = n12478 ;
  assign y2222 = ~n12484 ;
  assign y2223 = n12494 ;
  assign y2224 = n12497 ;
  assign y2225 = n12498 ;
  assign y2226 = n12505 ;
  assign y2227 = n12510 ;
  assign y2228 = ~1'b0 ;
  assign y2229 = ~n12512 ;
  assign y2230 = ~n12517 ;
  assign y2231 = n12518 ;
  assign y2232 = ~n12522 ;
  assign y2233 = ~n12524 ;
  assign y2234 = ~n12527 ;
  assign y2235 = n12528 ;
  assign y2236 = ~n12540 ;
  assign y2237 = ~n12548 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = n12553 ;
  assign y2240 = ~n12563 ;
  assign y2241 = ~n12566 ;
  assign y2242 = ~n12586 ;
  assign y2243 = n12625 ;
  assign y2244 = ~n12631 ;
  assign y2245 = n12632 ;
  assign y2246 = n12633 ;
  assign y2247 = n12635 ;
  assign y2248 = ~n12637 ;
  assign y2249 = n12640 ;
  assign y2250 = n12644 ;
  assign y2251 = ~n12650 ;
  assign y2252 = n12658 ;
  assign y2253 = ~n12660 ;
  assign y2254 = ~n12665 ;
  assign y2255 = n12677 ;
  assign y2256 = n12684 ;
  assign y2257 = n12689 ;
  assign y2258 = n12691 ;
  assign y2259 = n12697 ;
  assign y2260 = ~n12698 ;
  assign y2261 = ~n12699 ;
  assign y2262 = ~n12700 ;
  assign y2263 = ~n12705 ;
  assign y2264 = ~1'b0 ;
  assign y2265 = ~n12709 ;
  assign y2266 = ~n12710 ;
  assign y2267 = ~n12712 ;
  assign y2268 = ~1'b0 ;
  assign y2269 = n12729 ;
  assign y2270 = n12734 ;
  assign y2271 = n12736 ;
  assign y2272 = ~n12740 ;
  assign y2273 = ~n12747 ;
  assign y2274 = ~n12748 ;
  assign y2275 = n12756 ;
  assign y2276 = n12763 ;
  assign y2277 = n12765 ;
  assign y2278 = n12768 ;
  assign y2279 = ~n12781 ;
  assign y2280 = n12791 ;
  assign y2281 = ~n12794 ;
  assign y2282 = ~n12796 ;
  assign y2283 = ~1'b0 ;
  assign y2284 = ~1'b0 ;
  assign y2285 = n12797 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = n12799 ;
  assign y2288 = n12803 ;
  assign y2289 = ~n12807 ;
  assign y2290 = n12810 ;
  assign y2291 = ~n12814 ;
  assign y2292 = n12818 ;
  assign y2293 = ~n12823 ;
  assign y2294 = n12829 ;
  assign y2295 = n12830 ;
  assign y2296 = n12837 ;
  assign y2297 = ~n12844 ;
  assign y2298 = ~n12846 ;
  assign y2299 = n12850 ;
  assign y2300 = ~n12860 ;
  assign y2301 = n12870 ;
  assign y2302 = n12875 ;
  assign y2303 = ~n12883 ;
  assign y2304 = n12894 ;
  assign y2305 = ~1'b0 ;
  assign y2306 = n12895 ;
  assign y2307 = n12906 ;
  assign y2308 = n12916 ;
  assign y2309 = n12917 ;
  assign y2310 = n12920 ;
  assign y2311 = n12923 ;
  assign y2312 = n12924 ;
  assign y2313 = n12935 ;
  assign y2314 = ~n12939 ;
  assign y2315 = ~n12946 ;
  assign y2316 = n12952 ;
  assign y2317 = n12953 ;
  assign y2318 = ~n12958 ;
  assign y2319 = ~n12962 ;
  assign y2320 = ~n12968 ;
  assign y2321 = n12969 ;
  assign y2322 = ~n12982 ;
  assign y2323 = ~n12983 ;
  assign y2324 = n12987 ;
  assign y2325 = n12993 ;
  assign y2326 = ~n13009 ;
  assign y2327 = n13011 ;
  assign y2328 = n13016 ;
  assign y2329 = n13020 ;
  assign y2330 = n13023 ;
  assign y2331 = n13024 ;
  assign y2332 = ~n13027 ;
  assign y2333 = ~n13028 ;
  assign y2334 = n13044 ;
  assign y2335 = n13047 ;
  assign y2336 = ~n13057 ;
  assign y2337 = ~n13058 ;
  assign y2338 = n13075 ;
  assign y2339 = n13082 ;
  assign y2340 = ~n13084 ;
  assign y2341 = ~n13093 ;
  assign y2342 = n13094 ;
  assign y2343 = ~n13095 ;
  assign y2344 = n13103 ;
  assign y2345 = n13107 ;
  assign y2346 = ~n13111 ;
  assign y2347 = ~n13124 ;
  assign y2348 = ~n13133 ;
  assign y2349 = n13137 ;
  assign y2350 = ~n13145 ;
  assign y2351 = ~n13149 ;
  assign y2352 = ~n13156 ;
  assign y2353 = ~n13157 ;
  assign y2354 = ~n13158 ;
  assign y2355 = ~n13162 ;
  assign y2356 = ~n13171 ;
  assign y2357 = n13181 ;
  assign y2358 = n13182 ;
  assign y2359 = ~n13194 ;
  assign y2360 = n13197 ;
  assign y2361 = ~n13199 ;
  assign y2362 = ~n13205 ;
  assign y2363 = n13208 ;
  assign y2364 = ~n13210 ;
  assign y2365 = n13217 ;
  assign y2366 = n13219 ;
  assign y2367 = ~n13223 ;
  assign y2368 = ~n13224 ;
  assign y2369 = ~n3495 ;
  assign y2370 = n13226 ;
  assign y2371 = ~n13240 ;
  assign y2372 = ~1'b0 ;
  assign y2373 = ~n13242 ;
  assign y2374 = n13245 ;
  assign y2375 = n13255 ;
  assign y2376 = n13257 ;
  assign y2377 = n13262 ;
  assign y2378 = ~1'b0 ;
  assign y2379 = ~n13264 ;
  assign y2380 = n13271 ;
  assign y2381 = ~n13273 ;
  assign y2382 = ~n13276 ;
  assign y2383 = n13283 ;
  assign y2384 = ~n13285 ;
  assign y2385 = n13287 ;
  assign y2386 = ~1'b0 ;
  assign y2387 = ~n13299 ;
  assign y2388 = ~1'b0 ;
  assign y2389 = ~n13303 ;
  assign y2390 = ~n13304 ;
  assign y2391 = ~n13315 ;
  assign y2392 = ~n13323 ;
  assign y2393 = n13326 ;
  assign y2394 = n13338 ;
  assign y2395 = ~n13342 ;
  assign y2396 = n13345 ;
  assign y2397 = ~n13346 ;
  assign y2398 = n13353 ;
  assign y2399 = ~n13355 ;
  assign y2400 = n13359 ;
  assign y2401 = ~n13361 ;
  assign y2402 = n13365 ;
  assign y2403 = n13368 ;
  assign y2404 = ~n13369 ;
  assign y2405 = n13370 ;
  assign y2406 = ~n13373 ;
  assign y2407 = ~1'b0 ;
  assign y2408 = n13377 ;
  assign y2409 = n13384 ;
  assign y2410 = ~n13391 ;
  assign y2411 = ~n13397 ;
  assign y2412 = ~n6835 ;
  assign y2413 = n13401 ;
  assign y2414 = ~n13402 ;
  assign y2415 = n13414 ;
  assign y2416 = ~n13419 ;
  assign y2417 = ~n13422 ;
  assign y2418 = ~n13434 ;
  assign y2419 = n13436 ;
  assign y2420 = ~n13442 ;
  assign y2421 = n13443 ;
  assign y2422 = n13445 ;
  assign y2423 = ~n13447 ;
  assign y2424 = ~n13448 ;
  assign y2425 = ~n13461 ;
  assign y2426 = ~n13474 ;
  assign y2427 = n13477 ;
  assign y2428 = ~n13483 ;
  assign y2429 = n13485 ;
  assign y2430 = n13488 ;
  assign y2431 = ~n13492 ;
  assign y2432 = ~n13502 ;
  assign y2433 = n13503 ;
  assign y2434 = ~n13509 ;
  assign y2435 = ~n13514 ;
  assign y2436 = ~n13521 ;
  assign y2437 = ~n13523 ;
  assign y2438 = ~n13530 ;
  assign y2439 = ~n13534 ;
  assign y2440 = ~1'b0 ;
  assign y2441 = n13537 ;
  assign y2442 = n13547 ;
  assign y2443 = n13549 ;
  assign y2444 = n13550 ;
  assign y2445 = n13551 ;
  assign y2446 = n13565 ;
  assign y2447 = ~n13572 ;
  assign y2448 = ~n13579 ;
  assign y2449 = ~n13588 ;
  assign y2450 = n13597 ;
  assign y2451 = ~n13602 ;
  assign y2452 = ~n13604 ;
  assign y2453 = ~n13608 ;
  assign y2454 = n13626 ;
  assign y2455 = ~n13628 ;
  assign y2456 = n13631 ;
  assign y2457 = ~n13641 ;
  assign y2458 = ~n13643 ;
  assign y2459 = n13646 ;
  assign y2460 = ~n13650 ;
  assign y2461 = n13651 ;
  assign y2462 = ~n13655 ;
  assign y2463 = n13666 ;
  assign y2464 = ~1'b0 ;
  assign y2465 = ~n13677 ;
  assign y2466 = ~n13678 ;
  assign y2467 = ~1'b0 ;
  assign y2468 = ~n13684 ;
  assign y2469 = n13695 ;
  assign y2470 = n13704 ;
  assign y2471 = ~1'b0 ;
  assign y2472 = ~n13710 ;
  assign y2473 = ~n13711 ;
  assign y2474 = n13716 ;
  assign y2475 = n13723 ;
  assign y2476 = ~n13729 ;
  assign y2477 = ~1'b0 ;
  assign y2478 = n13731 ;
  assign y2479 = ~n13737 ;
  assign y2480 = ~n13738 ;
  assign y2481 = ~n13742 ;
  assign y2482 = n13761 ;
  assign y2483 = ~1'b0 ;
  assign y2484 = ~n13762 ;
  assign y2485 = n13768 ;
  assign y2486 = n13769 ;
  assign y2487 = ~n13771 ;
  assign y2488 = n13773 ;
  assign y2489 = n13774 ;
  assign y2490 = n13782 ;
  assign y2491 = ~1'b0 ;
  assign y2492 = n13788 ;
  assign y2493 = ~n13791 ;
  assign y2494 = ~n13797 ;
  assign y2495 = n13807 ;
  assign y2496 = n13808 ;
  assign y2497 = ~n13810 ;
  assign y2498 = n13813 ;
  assign y2499 = ~n13816 ;
  assign y2500 = n13817 ;
  assign y2501 = n13819 ;
  assign y2502 = n13830 ;
  assign y2503 = n13834 ;
  assign y2504 = n13837 ;
  assign y2505 = n13846 ;
  assign y2506 = ~n13849 ;
  assign y2507 = ~n13850 ;
  assign y2508 = ~n13854 ;
  assign y2509 = n13855 ;
  assign y2510 = ~1'b0 ;
  assign y2511 = ~n13862 ;
  assign y2512 = ~n13866 ;
  assign y2513 = ~n13871 ;
  assign y2514 = ~n13874 ;
  assign y2515 = ~n13876 ;
  assign y2516 = n13886 ;
  assign y2517 = n13891 ;
  assign y2518 = n13892 ;
  assign y2519 = ~n13893 ;
  assign y2520 = n13901 ;
  assign y2521 = ~1'b0 ;
  assign y2522 = ~n13907 ;
  assign y2523 = n13910 ;
  assign y2524 = ~n13915 ;
  assign y2525 = n13916 ;
  assign y2526 = n13920 ;
  assign y2527 = n13934 ;
  assign y2528 = n13937 ;
  assign y2529 = ~n13944 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = n13945 ;
  assign y2532 = ~n13956 ;
  assign y2533 = ~n13959 ;
  assign y2534 = n13964 ;
  assign y2535 = n13970 ;
  assign y2536 = n13972 ;
  assign y2537 = ~n13978 ;
  assign y2538 = ~n13979 ;
  assign y2539 = ~n13981 ;
  assign y2540 = n13986 ;
  assign y2541 = n13993 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = n13999 ;
  assign y2544 = n14001 ;
  assign y2545 = ~n14005 ;
  assign y2546 = ~n14009 ;
  assign y2547 = n14010 ;
  assign y2548 = ~n14014 ;
  assign y2549 = ~n8716 ;
  assign y2550 = ~n14015 ;
  assign y2551 = ~n14019 ;
  assign y2552 = ~n14024 ;
  assign y2553 = ~n14028 ;
  assign y2554 = n14031 ;
  assign y2555 = n14037 ;
  assign y2556 = ~n14043 ;
  assign y2557 = ~n14053 ;
  assign y2558 = n14059 ;
  assign y2559 = n14063 ;
  assign y2560 = n14068 ;
  assign y2561 = ~n14072 ;
  assign y2562 = ~1'b0 ;
  assign y2563 = ~n14074 ;
  assign y2564 = ~n14079 ;
  assign y2565 = n14086 ;
  assign y2566 = ~1'b0 ;
  assign y2567 = ~n14089 ;
  assign y2568 = ~1'b0 ;
  assign y2569 = n14090 ;
  assign y2570 = n14091 ;
  assign y2571 = n14093 ;
  assign y2572 = n14095 ;
  assign y2573 = n14102 ;
  assign y2574 = ~n14106 ;
  assign y2575 = n14112 ;
  assign y2576 = n14113 ;
  assign y2577 = n14120 ;
  assign y2578 = n14126 ;
  assign y2579 = ~n14127 ;
  assign y2580 = ~n14131 ;
  assign y2581 = ~n14134 ;
  assign y2582 = n14135 ;
  assign y2583 = n14139 ;
  assign y2584 = ~n14144 ;
  assign y2585 = ~1'b0 ;
  assign y2586 = ~n14149 ;
  assign y2587 = n14157 ;
  assign y2588 = n14158 ;
  assign y2589 = ~n14169 ;
  assign y2590 = n14171 ;
  assign y2591 = ~n14173 ;
  assign y2592 = ~n14178 ;
  assign y2593 = n14188 ;
  assign y2594 = ~1'b0 ;
  assign y2595 = n14189 ;
  assign y2596 = n14191 ;
  assign y2597 = n14192 ;
  assign y2598 = ~n14194 ;
  assign y2599 = ~n14195 ;
  assign y2600 = n14201 ;
  assign y2601 = ~1'b0 ;
  assign y2602 = ~n14211 ;
  assign y2603 = n14216 ;
  assign y2604 = n14224 ;
  assign y2605 = ~n14229 ;
  assign y2606 = n14234 ;
  assign y2607 = ~n14236 ;
  assign y2608 = n14241 ;
  assign y2609 = ~n14243 ;
  assign y2610 = ~n14244 ;
  assign y2611 = n14249 ;
  assign y2612 = n14259 ;
  assign y2613 = ~n14264 ;
  assign y2614 = ~n14267 ;
  assign y2615 = n14275 ;
  assign y2616 = ~n14276 ;
  assign y2617 = ~n14284 ;
  assign y2618 = ~n14294 ;
  assign y2619 = n14299 ;
  assign y2620 = n14302 ;
  assign y2621 = n14306 ;
  assign y2622 = n14320 ;
  assign y2623 = n14330 ;
  assign y2624 = ~n14332 ;
  assign y2625 = n14336 ;
  assign y2626 = ~n14344 ;
  assign y2627 = ~n14346 ;
  assign y2628 = ~n14354 ;
  assign y2629 = n14358 ;
  assign y2630 = ~n14362 ;
  assign y2631 = ~n14363 ;
  assign y2632 = ~n14367 ;
  assign y2633 = n14377 ;
  assign y2634 = n14380 ;
  assign y2635 = ~n14391 ;
  assign y2636 = n14392 ;
  assign y2637 = ~1'b0 ;
  assign y2638 = ~1'b0 ;
  assign y2639 = n14400 ;
  assign y2640 = n576 ;
  assign y2641 = n14402 ;
  assign y2642 = n14405 ;
  assign y2643 = n14406 ;
  assign y2644 = n14409 ;
  assign y2645 = n14411 ;
  assign y2646 = ~n14416 ;
  assign y2647 = ~n14425 ;
  assign y2648 = ~n14428 ;
  assign y2649 = ~n14429 ;
  assign y2650 = ~n14432 ;
  assign y2651 = n14434 ;
  assign y2652 = ~n14436 ;
  assign y2653 = n14437 ;
  assign y2654 = ~n14438 ;
  assign y2655 = ~n14441 ;
  assign y2656 = n14446 ;
  assign y2657 = ~n14454 ;
  assign y2658 = ~1'b0 ;
  assign y2659 = ~n14456 ;
  assign y2660 = n14474 ;
  assign y2661 = n14475 ;
  assign y2662 = ~n14476 ;
  assign y2663 = ~n14482 ;
  assign y2664 = ~n14485 ;
  assign y2665 = n14486 ;
  assign y2666 = ~n14489 ;
  assign y2667 = n14505 ;
  assign y2668 = ~1'b0 ;
  assign y2669 = n14521 ;
  assign y2670 = ~n14526 ;
  assign y2671 = ~n14528 ;
  assign y2672 = n14541 ;
  assign y2673 = n14547 ;
  assign y2674 = ~n14553 ;
  assign y2675 = n14559 ;
  assign y2676 = ~n14563 ;
  assign y2677 = ~n14565 ;
  assign y2678 = ~n14575 ;
  assign y2679 = ~n14584 ;
  assign y2680 = ~n14585 ;
  assign y2681 = n14590 ;
  assign y2682 = ~n14598 ;
  assign y2683 = ~n14602 ;
  assign y2684 = n14607 ;
  assign y2685 = ~n14617 ;
  assign y2686 = n14619 ;
  assign y2687 = ~n14627 ;
  assign y2688 = ~n14636 ;
  assign y2689 = ~n14640 ;
  assign y2690 = n14649 ;
  assign y2691 = n14652 ;
  assign y2692 = n14653 ;
  assign y2693 = ~n14657 ;
  assign y2694 = ~n14669 ;
  assign y2695 = ~n14674 ;
  assign y2696 = n14678 ;
  assign y2697 = ~n14684 ;
  assign y2698 = n14690 ;
  assign y2699 = ~1'b0 ;
  assign y2700 = ~n14691 ;
  assign y2701 = n14696 ;
  assign y2702 = n14699 ;
  assign y2703 = ~n14704 ;
  assign y2704 = ~n14708 ;
  assign y2705 = ~1'b0 ;
  assign y2706 = n14711 ;
  assign y2707 = ~n14718 ;
  assign y2708 = ~n14724 ;
  assign y2709 = ~1'b0 ;
  assign y2710 = ~n14725 ;
  assign y2711 = ~n14732 ;
  assign y2712 = n14736 ;
  assign y2713 = ~n14737 ;
  assign y2714 = ~n14741 ;
  assign y2715 = ~n14745 ;
  assign y2716 = ~1'b0 ;
  assign y2717 = n14747 ;
  assign y2718 = ~n14753 ;
  assign y2719 = n14755 ;
  assign y2720 = ~n14760 ;
  assign y2721 = n14774 ;
  assign y2722 = n14783 ;
  assign y2723 = n14786 ;
  assign y2724 = ~n14796 ;
  assign y2725 = ~n14802 ;
  assign y2726 = n14804 ;
  assign y2727 = ~n14808 ;
  assign y2728 = ~n14809 ;
  assign y2729 = ~n14821 ;
  assign y2730 = n14825 ;
  assign y2731 = ~n14826 ;
  assign y2732 = ~n14827 ;
  assign y2733 = ~n14829 ;
  assign y2734 = ~n14835 ;
  assign y2735 = ~n14842 ;
  assign y2736 = ~n14855 ;
  assign y2737 = n14863 ;
  assign y2738 = n14864 ;
  assign y2739 = n14866 ;
  assign y2740 = n14869 ;
  assign y2741 = ~n14871 ;
  assign y2742 = ~n14874 ;
  assign y2743 = n14877 ;
  assign y2744 = n14883 ;
  assign y2745 = n14884 ;
  assign y2746 = ~n14889 ;
  assign y2747 = ~1'b0 ;
  assign y2748 = ~n14890 ;
  assign y2749 = n14898 ;
  assign y2750 = n14900 ;
  assign y2751 = ~n14905 ;
  assign y2752 = n14906 ;
  assign y2753 = ~n14916 ;
  assign y2754 = n14919 ;
  assign y2755 = ~1'b0 ;
  assign y2756 = ~n14929 ;
  assign y2757 = ~n14931 ;
  assign y2758 = ~n14932 ;
  assign y2759 = n14933 ;
  assign y2760 = n14937 ;
  assign y2761 = ~1'b0 ;
  assign y2762 = n14939 ;
  assign y2763 = ~n14940 ;
  assign y2764 = n14944 ;
  assign y2765 = ~n14959 ;
  assign y2766 = ~1'b0 ;
  assign y2767 = ~n14963 ;
  assign y2768 = ~n14971 ;
  assign y2769 = ~n14979 ;
  assign y2770 = n14982 ;
  assign y2771 = ~n14987 ;
  assign y2772 = ~n14990 ;
  assign y2773 = n14991 ;
  assign y2774 = ~n14993 ;
  assign y2775 = n14995 ;
  assign y2776 = n14997 ;
  assign y2777 = n15000 ;
  assign y2778 = n15006 ;
  assign y2779 = ~n15009 ;
  assign y2780 = ~1'b0 ;
  assign y2781 = ~n15012 ;
  assign y2782 = n15014 ;
  assign y2783 = ~n15021 ;
  assign y2784 = ~n15026 ;
  assign y2785 = ~n15027 ;
  assign y2786 = ~n15033 ;
  assign y2787 = n15044 ;
  assign y2788 = n15046 ;
  assign y2789 = ~n15048 ;
  assign y2790 = n15049 ;
  assign y2791 = n15050 ;
  assign y2792 = ~n15053 ;
  assign y2793 = n15063 ;
  assign y2794 = ~n15064 ;
  assign y2795 = ~n15067 ;
  assign y2796 = ~n15069 ;
  assign y2797 = n15071 ;
  assign y2798 = ~1'b0 ;
  assign y2799 = n15073 ;
  assign y2800 = ~n15077 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = ~1'b0 ;
  assign y2803 = ~n15080 ;
  assign y2804 = ~n15083 ;
  assign y2805 = ~n15084 ;
  assign y2806 = ~n15088 ;
  assign y2807 = n15089 ;
  assign y2808 = ~n15090 ;
  assign y2809 = n15091 ;
  assign y2810 = n15095 ;
  assign y2811 = ~n15103 ;
  assign y2812 = n15105 ;
  assign y2813 = n15108 ;
  assign y2814 = ~n15119 ;
  assign y2815 = ~n15130 ;
  assign y2816 = ~n15131 ;
  assign y2817 = n15143 ;
  assign y2818 = ~1'b0 ;
  assign y2819 = ~n15148 ;
  assign y2820 = n15162 ;
  assign y2821 = ~n15165 ;
  assign y2822 = ~n15171 ;
  assign y2823 = n15174 ;
  assign y2824 = n15177 ;
  assign y2825 = n15189 ;
  assign y2826 = ~1'b0 ;
  assign y2827 = ~n15193 ;
  assign y2828 = n15194 ;
  assign y2829 = ~n15201 ;
  assign y2830 = ~n15205 ;
  assign y2831 = ~n15211 ;
  assign y2832 = n15216 ;
  assign y2833 = n15223 ;
  assign y2834 = ~n15234 ;
  assign y2835 = ~n15238 ;
  assign y2836 = ~n15240 ;
  assign y2837 = n15249 ;
  assign y2838 = n15251 ;
  assign y2839 = n15255 ;
  assign y2840 = n15267 ;
  assign y2841 = ~n15268 ;
  assign y2842 = ~n15277 ;
  assign y2843 = ~n15285 ;
  assign y2844 = ~n15289 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = ~n15291 ;
  assign y2847 = n15295 ;
  assign y2848 = n15297 ;
  assign y2849 = ~n15300 ;
  assign y2850 = ~n15308 ;
  assign y2851 = ~n15310 ;
  assign y2852 = ~n15312 ;
  assign y2853 = n15315 ;
  assign y2854 = ~n15317 ;
  assign y2855 = n15321 ;
  assign y2856 = ~n15327 ;
  assign y2857 = n15328 ;
  assign y2858 = ~n15329 ;
  assign y2859 = n15330 ;
  assign y2860 = ~n15332 ;
  assign y2861 = ~n15337 ;
  assign y2862 = ~n15340 ;
  assign y2863 = n15342 ;
  assign y2864 = ~n15352 ;
  assign y2865 = n15359 ;
  assign y2866 = n15363 ;
  assign y2867 = n15367 ;
  assign y2868 = ~n15377 ;
  assign y2869 = ~n15383 ;
  assign y2870 = ~n15384 ;
  assign y2871 = ~1'b0 ;
  assign y2872 = ~1'b0 ;
  assign y2873 = n15389 ;
  assign y2874 = ~n15400 ;
  assign y2875 = ~n15401 ;
  assign y2876 = ~1'b0 ;
  assign y2877 = n15404 ;
  assign y2878 = n15410 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~n15413 ;
  assign y2881 = n15416 ;
  assign y2882 = n15417 ;
  assign y2883 = n15426 ;
  assign y2884 = ~n15428 ;
  assign y2885 = ~n15437 ;
  assign y2886 = ~1'b0 ;
  assign y2887 = ~n15442 ;
  assign y2888 = ~n15447 ;
  assign y2889 = n15449 ;
  assign y2890 = n15452 ;
  assign y2891 = ~n15453 ;
  assign y2892 = n15457 ;
  assign y2893 = ~n15458 ;
  assign y2894 = ~n15465 ;
  assign y2895 = ~1'b0 ;
  assign y2896 = ~n15467 ;
  assign y2897 = n15470 ;
  assign y2898 = n15471 ;
  assign y2899 = n15472 ;
  assign y2900 = n15485 ;
  assign y2901 = n15495 ;
  assign y2902 = ~1'b0 ;
  assign y2903 = n15497 ;
  assign y2904 = ~n15510 ;
  assign y2905 = ~n15513 ;
  assign y2906 = ~1'b0 ;
  assign y2907 = ~n15525 ;
  assign y2908 = ~n15527 ;
  assign y2909 = ~n15529 ;
  assign y2910 = n15537 ;
  assign y2911 = n15539 ;
  assign y2912 = n15544 ;
  assign y2913 = ~n15551 ;
  assign y2914 = n15561 ;
  assign y2915 = ~1'b0 ;
  assign y2916 = ~n15563 ;
  assign y2917 = n15567 ;
  assign y2918 = ~n15573 ;
  assign y2919 = ~n15577 ;
  assign y2920 = n15585 ;
  assign y2921 = n15590 ;
  assign y2922 = n15591 ;
  assign y2923 = ~n15599 ;
  assign y2924 = ~n15603 ;
  assign y2925 = n15616 ;
  assign y2926 = ~n15627 ;
  assign y2927 = n15629 ;
  assign y2928 = n15633 ;
  assign y2929 = n15637 ;
  assign y2930 = ~n15651 ;
  assign y2931 = n15654 ;
  assign y2932 = n15660 ;
  assign y2933 = n15665 ;
  assign y2934 = ~1'b0 ;
  assign y2935 = ~n15670 ;
  assign y2936 = ~n15671 ;
  assign y2937 = ~n15679 ;
  assign y2938 = n15681 ;
  assign y2939 = ~n15683 ;
  assign y2940 = ~n15686 ;
  assign y2941 = ~n15687 ;
  assign y2942 = n15695 ;
  assign y2943 = n15697 ;
  assign y2944 = ~n15698 ;
  assign y2945 = ~n15700 ;
  assign y2946 = ~n15709 ;
  assign y2947 = n15721 ;
  assign y2948 = ~n15728 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = ~n15729 ;
  assign y2951 = n15737 ;
  assign y2952 = ~n15744 ;
  assign y2953 = n15747 ;
  assign y2954 = n15748 ;
  assign y2955 = ~n15751 ;
  assign y2956 = ~n15752 ;
  assign y2957 = ~n15757 ;
  assign y2958 = ~n15767 ;
  assign y2959 = n15783 ;
  assign y2960 = n15786 ;
  assign y2961 = n15791 ;
  assign y2962 = n15798 ;
  assign y2963 = n15808 ;
  assign y2964 = n15820 ;
  assign y2965 = ~n15831 ;
  assign y2966 = ~n15837 ;
  assign y2967 = ~n9347 ;
  assign y2968 = ~n15851 ;
  assign y2969 = ~n15854 ;
  assign y2970 = n15855 ;
  assign y2971 = ~n15856 ;
  assign y2972 = n15859 ;
  assign y2973 = n15869 ;
  assign y2974 = n15870 ;
  assign y2975 = n15872 ;
  assign y2976 = n15877 ;
  assign y2977 = ~n15883 ;
  assign y2978 = ~n15885 ;
  assign y2979 = ~n15890 ;
  assign y2980 = n15894 ;
  assign y2981 = ~n15901 ;
  assign y2982 = n15921 ;
  assign y2983 = n15929 ;
  assign y2984 = ~n15931 ;
  assign y2985 = n15938 ;
  assign y2986 = ~n15950 ;
  assign y2987 = ~n15952 ;
  assign y2988 = n15954 ;
  assign y2989 = ~n15959 ;
  assign y2990 = ~n15966 ;
  assign y2991 = ~n15969 ;
  assign y2992 = n15973 ;
  assign y2993 = ~n15974 ;
  assign y2994 = n15984 ;
  assign y2995 = n15991 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = ~n16001 ;
  assign y2998 = ~n16009 ;
  assign y2999 = ~n16014 ;
  assign y3000 = n16022 ;
  assign y3001 = n16035 ;
  assign y3002 = n16037 ;
  assign y3003 = ~n16041 ;
  assign y3004 = ~n16046 ;
  assign y3005 = ~n16049 ;
  assign y3006 = n16057 ;
  assign y3007 = n16061 ;
  assign y3008 = n16064 ;
  assign y3009 = ~n16067 ;
  assign y3010 = n16075 ;
  assign y3011 = ~n16077 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = n16090 ;
  assign y3014 = ~n16100 ;
  assign y3015 = ~n16104 ;
  assign y3016 = ~n16107 ;
  assign y3017 = ~n16111 ;
  assign y3018 = ~n16112 ;
  assign y3019 = n16119 ;
  assign y3020 = ~1'b0 ;
  assign y3021 = ~n16122 ;
  assign y3022 = n16127 ;
  assign y3023 = n16128 ;
  assign y3024 = ~n16134 ;
  assign y3025 = ~n16135 ;
  assign y3026 = ~n16144 ;
  assign y3027 = ~n16154 ;
  assign y3028 = ~n16156 ;
  assign y3029 = n16162 ;
  assign y3030 = ~n16167 ;
  assign y3031 = ~1'b0 ;
  assign y3032 = n16169 ;
  assign y3033 = n16174 ;
  assign y3034 = ~n16177 ;
  assign y3035 = n16182 ;
  assign y3036 = ~n16183 ;
  assign y3037 = n16186 ;
  assign y3038 = n16200 ;
  assign y3039 = ~1'b0 ;
  assign y3040 = ~n16201 ;
  assign y3041 = n16204 ;
  assign y3042 = n16210 ;
  assign y3043 = n16212 ;
  assign y3044 = ~n16218 ;
  assign y3045 = ~n16223 ;
  assign y3046 = ~n16227 ;
  assign y3047 = n16230 ;
  assign y3048 = ~n16231 ;
  assign y3049 = ~1'b0 ;
  assign y3050 = ~n16232 ;
  assign y3051 = n16234 ;
  assign y3052 = n16241 ;
  assign y3053 = n16243 ;
  assign y3054 = ~n16258 ;
  assign y3055 = ~n16259 ;
  assign y3056 = n16265 ;
  assign y3057 = n16274 ;
  assign y3058 = ~n16275 ;
  assign y3059 = ~n16277 ;
  assign y3060 = n16278 ;
  assign y3061 = n16282 ;
  assign y3062 = n16287 ;
  assign y3063 = n16291 ;
  assign y3064 = ~n16297 ;
  assign y3065 = n16304 ;
  assign y3066 = n16305 ;
  assign y3067 = n16314 ;
  assign y3068 = ~n16319 ;
  assign y3069 = ~n16328 ;
  assign y3070 = n16335 ;
  assign y3071 = n16337 ;
  assign y3072 = ~1'b0 ;
  assign y3073 = n16345 ;
  assign y3074 = n16353 ;
  assign y3075 = ~n16360 ;
  assign y3076 = n16365 ;
  assign y3077 = n16368 ;
  assign y3078 = ~n16371 ;
  assign y3079 = n16372 ;
  assign y3080 = ~n16378 ;
  assign y3081 = ~n16382 ;
  assign y3082 = ~n16385 ;
  assign y3083 = ~n16386 ;
  assign y3084 = ~n16401 ;
  assign y3085 = n16403 ;
  assign y3086 = ~n16410 ;
  assign y3087 = ~n16412 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~n16413 ;
  assign y3090 = ~n16414 ;
  assign y3091 = n16415 ;
  assign y3092 = ~n16417 ;
  assign y3093 = ~1'b0 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = n16424 ;
  assign y3096 = n16428 ;
  assign y3097 = ~n16430 ;
  assign y3098 = n16439 ;
  assign y3099 = ~n16449 ;
  assign y3100 = ~n16452 ;
  assign y3101 = n16462 ;
  assign y3102 = ~n16478 ;
  assign y3103 = ~n16480 ;
  assign y3104 = ~n16481 ;
  assign y3105 = ~n16482 ;
  assign y3106 = n10042 ;
  assign y3107 = ~1'b0 ;
  assign y3108 = ~n16490 ;
  assign y3109 = n16510 ;
  assign y3110 = ~n16515 ;
  assign y3111 = n16519 ;
  assign y3112 = ~n16523 ;
  assign y3113 = ~n16536 ;
  assign y3114 = ~n16539 ;
  assign y3115 = n16550 ;
  assign y3116 = ~n16555 ;
  assign y3117 = ~n16560 ;
  assign y3118 = ~n16563 ;
  assign y3119 = ~n16569 ;
  assign y3120 = ~n16571 ;
  assign y3121 = ~n16583 ;
  assign y3122 = ~1'b0 ;
  assign y3123 = n16586 ;
  assign y3124 = ~n16595 ;
  assign y3125 = n16601 ;
  assign y3126 = ~1'b0 ;
  assign y3127 = ~1'b0 ;
  assign y3128 = n16608 ;
  assign y3129 = n16619 ;
  assign y3130 = ~n16620 ;
  assign y3131 = n16624 ;
  assign y3132 = n16631 ;
  assign y3133 = n16633 ;
  assign y3134 = ~n16638 ;
  assign y3135 = ~n16639 ;
  assign y3136 = ~n16640 ;
  assign y3137 = ~n16645 ;
  assign y3138 = ~n16646 ;
  assign y3139 = n16647 ;
  assign y3140 = n16652 ;
  assign y3141 = ~n16658 ;
  assign y3142 = ~n16659 ;
  assign y3143 = ~n16661 ;
  assign y3144 = n16663 ;
  assign y3145 = ~n16665 ;
  assign y3146 = n16670 ;
  assign y3147 = n16673 ;
  assign y3148 = n16674 ;
  assign y3149 = n16675 ;
  assign y3150 = ~n16678 ;
  assign y3151 = ~n16679 ;
  assign y3152 = ~n16687 ;
  assign y3153 = n16697 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = n16706 ;
  assign y3156 = ~n16712 ;
  assign y3157 = ~n16721 ;
  assign y3158 = ~n16728 ;
  assign y3159 = n16729 ;
  assign y3160 = ~n16730 ;
  assign y3161 = n16736 ;
  assign y3162 = ~n16739 ;
  assign y3163 = n16741 ;
  assign y3164 = n16743 ;
  assign y3165 = n16744 ;
  assign y3166 = ~n16749 ;
  assign y3167 = n16752 ;
  assign y3168 = ~n16761 ;
  assign y3169 = ~n16772 ;
  assign y3170 = n16779 ;
  assign y3171 = ~n16783 ;
  assign y3172 = ~n16786 ;
  assign y3173 = n16803 ;
  assign y3174 = ~n16809 ;
  assign y3175 = n16810 ;
  assign y3176 = n16813 ;
  assign y3177 = ~n16816 ;
  assign y3178 = ~n16821 ;
  assign y3179 = ~n16822 ;
  assign y3180 = ~n16823 ;
  assign y3181 = n16824 ;
  assign y3182 = n16844 ;
  assign y3183 = n16864 ;
  assign y3184 = n16873 ;
  assign y3185 = n16874 ;
  assign y3186 = ~n16875 ;
  assign y3187 = n16876 ;
  assign y3188 = n16885 ;
  assign y3189 = ~n16891 ;
  assign y3190 = n16896 ;
  assign y3191 = n16904 ;
  assign y3192 = n16908 ;
  assign y3193 = ~n16913 ;
  assign y3194 = n16915 ;
  assign y3195 = n16918 ;
  assign y3196 = n16924 ;
  assign y3197 = ~n16929 ;
  assign y3198 = n16930 ;
  assign y3199 = n16931 ;
  assign y3200 = n16938 ;
  assign y3201 = n16939 ;
  assign y3202 = ~n16946 ;
  assign y3203 = n16949 ;
  assign y3204 = n16959 ;
  assign y3205 = n16961 ;
  assign y3206 = n16963 ;
  assign y3207 = n16965 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = n16969 ;
  assign y3210 = n16972 ;
  assign y3211 = n16974 ;
  assign y3212 = n16977 ;
  assign y3213 = ~n16978 ;
  assign y3214 = ~n16983 ;
  assign y3215 = ~n16991 ;
  assign y3216 = ~1'b0 ;
  assign y3217 = ~1'b0 ;
  assign y3218 = ~n16996 ;
  assign y3219 = n17005 ;
  assign y3220 = n17010 ;
  assign y3221 = n17013 ;
  assign y3222 = ~n17017 ;
  assign y3223 = n17024 ;
  assign y3224 = n17026 ;
  assign y3225 = ~n17036 ;
  assign y3226 = ~n17047 ;
  assign y3227 = n17051 ;
  assign y3228 = ~n17057 ;
  assign y3229 = ~n17058 ;
  assign y3230 = n17061 ;
  assign y3231 = n17062 ;
  assign y3232 = ~n17065 ;
  assign y3233 = n17067 ;
  assign y3234 = ~n17068 ;
  assign y3235 = ~n17071 ;
  assign y3236 = n17076 ;
  assign y3237 = ~n17089 ;
  assign y3238 = ~n17090 ;
  assign y3239 = ~n17094 ;
  assign y3240 = n17098 ;
  assign y3241 = n17107 ;
  assign y3242 = ~n17122 ;
  assign y3243 = ~n17127 ;
  assign y3244 = n17129 ;
  assign y3245 = ~n17136 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = ~n17145 ;
  assign y3248 = n17148 ;
  assign y3249 = n17152 ;
  assign y3250 = n17161 ;
  assign y3251 = ~n17169 ;
  assign y3252 = ~n17177 ;
  assign y3253 = ~n17179 ;
  assign y3254 = ~n17182 ;
  assign y3255 = n17189 ;
  assign y3256 = n17194 ;
  assign y3257 = n17197 ;
  assign y3258 = n17200 ;
  assign y3259 = ~n17202 ;
  assign y3260 = ~n17212 ;
  assign y3261 = ~n17216 ;
  assign y3262 = ~n17222 ;
  assign y3263 = n17225 ;
  assign y3264 = n17234 ;
  assign y3265 = ~n17237 ;
  assign y3266 = ~n17238 ;
  assign y3267 = ~n17239 ;
  assign y3268 = n17244 ;
  assign y3269 = n17245 ;
  assign y3270 = ~n17247 ;
  assign y3271 = ~n17250 ;
  assign y3272 = n17254 ;
  assign y3273 = n5222 ;
  assign y3274 = ~n17265 ;
  assign y3275 = n17266 ;
  assign y3276 = n17267 ;
  assign y3277 = ~n17269 ;
  assign y3278 = ~n17277 ;
  assign y3279 = ~n17286 ;
  assign y3280 = n17288 ;
  assign y3281 = ~1'b0 ;
  assign y3282 = n17292 ;
  assign y3283 = ~n17297 ;
  assign y3284 = ~n17300 ;
  assign y3285 = n17310 ;
  assign y3286 = ~n17312 ;
  assign y3287 = ~n17319 ;
  assign y3288 = ~n17321 ;
  assign y3289 = n17323 ;
  assign y3290 = n17325 ;
  assign y3291 = ~n17326 ;
  assign y3292 = ~n17328 ;
  assign y3293 = ~n17333 ;
  assign y3294 = n17343 ;
  assign y3295 = ~n17344 ;
  assign y3296 = ~n17347 ;
  assign y3297 = n17350 ;
  assign y3298 = n17357 ;
  assign y3299 = n17365 ;
  assign y3300 = ~1'b0 ;
  assign y3301 = ~n17370 ;
  assign y3302 = n17373 ;
  assign y3303 = ~1'b0 ;
  assign y3304 = ~n17374 ;
  assign y3305 = n17375 ;
  assign y3306 = n17381 ;
  assign y3307 = n17385 ;
  assign y3308 = n17387 ;
  assign y3309 = ~n17390 ;
  assign y3310 = ~n17395 ;
  assign y3311 = n17410 ;
  assign y3312 = n17414 ;
  assign y3313 = n17417 ;
  assign y3314 = ~1'b0 ;
  assign y3315 = n17419 ;
  assign y3316 = ~n17429 ;
  assign y3317 = n17435 ;
  assign y3318 = ~n17439 ;
  assign y3319 = n17440 ;
  assign y3320 = n17445 ;
  assign y3321 = ~1'b0 ;
  assign y3322 = ~n17447 ;
  assign y3323 = ~n17453 ;
  assign y3324 = n17455 ;
  assign y3325 = n17456 ;
  assign y3326 = ~n17462 ;
  assign y3327 = n17469 ;
  assign y3328 = ~n17473 ;
  assign y3329 = ~n17481 ;
  assign y3330 = ~n17483 ;
  assign y3331 = ~n17490 ;
  assign y3332 = ~n17495 ;
  assign y3333 = ~n17499 ;
  assign y3334 = ~n17506 ;
  assign y3335 = n17509 ;
  assign y3336 = ~n17511 ;
  assign y3337 = n17517 ;
  assign y3338 = ~n17520 ;
  assign y3339 = n17521 ;
  assign y3340 = n17524 ;
  assign y3341 = n17525 ;
  assign y3342 = n17529 ;
  assign y3343 = n17532 ;
  assign y3344 = n17533 ;
  assign y3345 = n17535 ;
  assign y3346 = ~n17539 ;
  assign y3347 = ~n17540 ;
  assign y3348 = ~n17541 ;
  assign y3349 = n17552 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = n17554 ;
  assign y3352 = n17560 ;
  assign y3353 = n17567 ;
  assign y3354 = n17569 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = ~n17572 ;
  assign y3357 = ~n17580 ;
  assign y3358 = n17581 ;
  assign y3359 = ~n17585 ;
  assign y3360 = ~1'b0 ;
  assign y3361 = ~n17587 ;
  assign y3362 = n17590 ;
  assign y3363 = ~n17593 ;
  assign y3364 = ~n17595 ;
  assign y3365 = ~n17599 ;
  assign y3366 = ~n17602 ;
  assign y3367 = n17605 ;
  assign y3368 = n17616 ;
  assign y3369 = ~n17626 ;
  assign y3370 = ~n17628 ;
  assign y3371 = ~n17634 ;
  assign y3372 = ~1'b0 ;
  assign y3373 = ~n17635 ;
  assign y3374 = ~n17644 ;
  assign y3375 = ~n17647 ;
  assign y3376 = ~n17649 ;
  assign y3377 = ~n17657 ;
  assign y3378 = ~n17665 ;
  assign y3379 = ~n17669 ;
  assign y3380 = ~1'b0 ;
  assign y3381 = ~n17670 ;
  assign y3382 = n17679 ;
  assign y3383 = n17688 ;
  assign y3384 = ~n17695 ;
  assign y3385 = n17698 ;
  assign y3386 = ~n17700 ;
  assign y3387 = n17704 ;
  assign y3388 = ~n17711 ;
  assign y3389 = ~n17713 ;
  assign y3390 = n17720 ;
  assign y3391 = n17730 ;
  assign y3392 = n17732 ;
  assign y3393 = n17735 ;
  assign y3394 = n17736 ;
  assign y3395 = ~n17737 ;
  assign y3396 = ~1'b0 ;
  assign y3397 = ~n17739 ;
  assign y3398 = n17740 ;
  assign y3399 = ~n17741 ;
  assign y3400 = n17748 ;
  assign y3401 = n17759 ;
  assign y3402 = n17765 ;
  assign y3403 = n17767 ;
  assign y3404 = n17776 ;
  assign y3405 = n17785 ;
  assign y3406 = ~n17786 ;
  assign y3407 = n17789 ;
  assign y3408 = n17792 ;
  assign y3409 = n17809 ;
  assign y3410 = n17813 ;
  assign y3411 = n17815 ;
  assign y3412 = n17827 ;
  assign y3413 = n17829 ;
  assign y3414 = ~n17837 ;
  assign y3415 = ~n17839 ;
  assign y3416 = n17845 ;
  assign y3417 = ~n17846 ;
  assign y3418 = ~n17848 ;
  assign y3419 = n17850 ;
  assign y3420 = n17852 ;
  assign y3421 = n17855 ;
  assign y3422 = ~n17857 ;
  assign y3423 = ~n17859 ;
  assign y3424 = n17871 ;
  assign y3425 = n17882 ;
  assign y3426 = ~n17888 ;
  assign y3427 = ~n17899 ;
  assign y3428 = ~1'b0 ;
  assign y3429 = ~n17902 ;
  assign y3430 = ~n17921 ;
  assign y3431 = ~n17923 ;
  assign y3432 = ~n17924 ;
  assign y3433 = ~n17937 ;
  assign y3434 = ~1'b0 ;
  assign y3435 = ~n17940 ;
  assign y3436 = n17942 ;
  assign y3437 = ~n17950 ;
  assign y3438 = n17952 ;
  assign y3439 = n17953 ;
  assign y3440 = n17962 ;
  assign y3441 = n17971 ;
  assign y3442 = n17977 ;
  assign y3443 = ~n17996 ;
  assign y3444 = n17998 ;
  assign y3445 = n18002 ;
  assign y3446 = n18009 ;
  assign y3447 = ~n18016 ;
  assign y3448 = n18017 ;
  assign y3449 = n18019 ;
  assign y3450 = ~n18021 ;
  assign y3451 = n18028 ;
  assign y3452 = ~n18032 ;
  assign y3453 = ~n18035 ;
  assign y3454 = ~n18042 ;
  assign y3455 = n18043 ;
  assign y3456 = ~1'b0 ;
  assign y3457 = ~n18047 ;
  assign y3458 = n18049 ;
  assign y3459 = n18050 ;
  assign y3460 = ~n18052 ;
  assign y3461 = n18054 ;
  assign y3462 = ~n18061 ;
  assign y3463 = n18063 ;
  assign y3464 = n18068 ;
  assign y3465 = n18069 ;
  assign y3466 = ~1'b0 ;
  assign y3467 = ~n18077 ;
  assign y3468 = ~n18080 ;
  assign y3469 = ~n18089 ;
  assign y3470 = ~n18090 ;
  assign y3471 = ~1'b0 ;
  assign y3472 = ~1'b0 ;
  assign y3473 = ~n18091 ;
  assign y3474 = n18092 ;
  assign y3475 = ~1'b0 ;
  assign y3476 = ~n18099 ;
  assign y3477 = ~n18106 ;
  assign y3478 = ~n18112 ;
  assign y3479 = n18115 ;
  assign y3480 = ~n18125 ;
  assign y3481 = ~n18126 ;
  assign y3482 = n18130 ;
  assign y3483 = n18137 ;
  assign y3484 = n18139 ;
  assign y3485 = ~n18141 ;
  assign y3486 = ~n18149 ;
  assign y3487 = n18151 ;
  assign y3488 = n18153 ;
  assign y3489 = n18154 ;
  assign y3490 = ~n18159 ;
  assign y3491 = n18162 ;
  assign y3492 = ~n18166 ;
  assign y3493 = ~n18168 ;
  assign y3494 = ~n18170 ;
  assign y3495 = n18183 ;
  assign y3496 = n18186 ;
  assign y3497 = n18188 ;
  assign y3498 = ~n18191 ;
  assign y3499 = ~n18196 ;
  assign y3500 = n18197 ;
  assign y3501 = ~n18201 ;
  assign y3502 = ~n18206 ;
  assign y3503 = ~n18221 ;
  assign y3504 = n18224 ;
  assign y3505 = ~n18227 ;
  assign y3506 = ~n18229 ;
  assign y3507 = ~n18231 ;
  assign y3508 = ~n18232 ;
  assign y3509 = ~n18235 ;
  assign y3510 = ~1'b0 ;
  assign y3511 = ~n18240 ;
  assign y3512 = n18246 ;
  assign y3513 = ~n18247 ;
  assign y3514 = n18249 ;
  assign y3515 = n18252 ;
  assign y3516 = ~n18254 ;
  assign y3517 = ~n18267 ;
  assign y3518 = n18269 ;
  assign y3519 = ~1'b0 ;
  assign y3520 = n8067 ;
  assign y3521 = ~n18272 ;
  assign y3522 = ~n18273 ;
  assign y3523 = ~n18278 ;
  assign y3524 = ~1'b0 ;
  assign y3525 = ~n18294 ;
  assign y3526 = ~n18300 ;
  assign y3527 = ~n18307 ;
  assign y3528 = ~n18309 ;
  assign y3529 = n18323 ;
  assign y3530 = n18335 ;
  assign y3531 = ~1'b0 ;
  assign y3532 = ~n18340 ;
  assign y3533 = ~1'b0 ;
  assign y3534 = ~n18341 ;
  assign y3535 = n18346 ;
  assign y3536 = ~n18348 ;
  assign y3537 = ~n18354 ;
  assign y3538 = n18358 ;
  assign y3539 = n18361 ;
  assign y3540 = ~1'b0 ;
  assign y3541 = ~n18362 ;
  assign y3542 = ~n18368 ;
  assign y3543 = ~n18372 ;
  assign y3544 = n18380 ;
  assign y3545 = n18382 ;
  assign y3546 = ~1'b0 ;
  assign y3547 = n18384 ;
  assign y3548 = n18387 ;
  assign y3549 = ~n18405 ;
  assign y3550 = n18408 ;
  assign y3551 = ~1'b0 ;
  assign y3552 = n18413 ;
  assign y3553 = ~n18414 ;
  assign y3554 = n18421 ;
  assign y3555 = ~n18422 ;
  assign y3556 = n18427 ;
  assign y3557 = n868 ;
  assign y3558 = n18428 ;
  assign y3559 = ~n18432 ;
  assign y3560 = ~n18433 ;
  assign y3561 = ~n18446 ;
  assign y3562 = ~n18448 ;
  assign y3563 = ~n18450 ;
  assign y3564 = ~n18456 ;
  assign y3565 = n18462 ;
  assign y3566 = n18464 ;
  assign y3567 = n18478 ;
  assign y3568 = n18479 ;
  assign y3569 = ~n18481 ;
  assign y3570 = ~n18487 ;
  assign y3571 = ~n18488 ;
  assign y3572 = n18492 ;
  assign y3573 = ~n18501 ;
  assign y3574 = n14888 ;
  assign y3575 = ~n18502 ;
  assign y3576 = n18509 ;
  assign y3577 = ~n18514 ;
  assign y3578 = ~n18519 ;
  assign y3579 = ~n18521 ;
  assign y3580 = n18533 ;
  assign y3581 = n18536 ;
  assign y3582 = ~n18538 ;
  assign y3583 = n18542 ;
  assign y3584 = ~n18548 ;
  assign y3585 = n18549 ;
  assign y3586 = n18554 ;
  assign y3587 = n18555 ;
  assign y3588 = n18561 ;
  assign y3589 = n18566 ;
  assign y3590 = ~n18570 ;
  assign y3591 = ~n18571 ;
  assign y3592 = ~n18573 ;
  assign y3593 = ~n18578 ;
  assign y3594 = ~1'b0 ;
  assign y3595 = ~n18579 ;
  assign y3596 = n18581 ;
  assign y3597 = n18584 ;
  assign y3598 = ~1'b0 ;
  assign y3599 = ~n18591 ;
  assign y3600 = ~n18597 ;
  assign y3601 = ~n18603 ;
  assign y3602 = n18605 ;
  assign y3603 = n18606 ;
  assign y3604 = ~1'b0 ;
  assign y3605 = n18613 ;
  assign y3606 = n18614 ;
  assign y3607 = n18620 ;
  assign y3608 = n18622 ;
  assign y3609 = ~n18623 ;
  assign y3610 = ~n18626 ;
  assign y3611 = n18628 ;
  assign y3612 = ~n18630 ;
  assign y3613 = n18633 ;
  assign y3614 = n18640 ;
  assign y3615 = ~n18642 ;
  assign y3616 = ~n18645 ;
  assign y3617 = ~n18647 ;
  assign y3618 = ~n18653 ;
  assign y3619 = n18663 ;
  assign y3620 = n18665 ;
  assign y3621 = ~n18675 ;
  assign y3622 = n18676 ;
  assign y3623 = n18679 ;
  assign y3624 = ~n18681 ;
  assign y3625 = n18686 ;
  assign y3626 = ~n18687 ;
  assign y3627 = n18691 ;
  assign y3628 = ~n18694 ;
  assign y3629 = n18701 ;
  assign y3630 = ~1'b0 ;
  assign y3631 = n18711 ;
  assign y3632 = ~n18722 ;
  assign y3633 = n18723 ;
  assign y3634 = n18729 ;
  assign y3635 = n18732 ;
  assign y3636 = n18734 ;
  assign y3637 = ~n18737 ;
  assign y3638 = n18750 ;
  assign y3639 = n18755 ;
  assign y3640 = ~n18757 ;
  assign y3641 = n18759 ;
  assign y3642 = n18763 ;
  assign y3643 = ~n18767 ;
  assign y3644 = n18769 ;
  assign y3645 = n18773 ;
  assign y3646 = n18783 ;
  assign y3647 = n18786 ;
  assign y3648 = ~n18793 ;
  assign y3649 = ~n18799 ;
  assign y3650 = ~n18800 ;
  assign y3651 = ~n18804 ;
  assign y3652 = ~n18807 ;
  assign y3653 = ~n18809 ;
  assign y3654 = ~n18810 ;
  assign y3655 = n18815 ;
  assign y3656 = ~n18820 ;
  assign y3657 = ~n18823 ;
  assign y3658 = n18824 ;
  assign y3659 = ~n18826 ;
  assign y3660 = n18827 ;
  assign y3661 = ~n18833 ;
  assign y3662 = n18839 ;
  assign y3663 = n18846 ;
  assign y3664 = n18851 ;
  assign y3665 = n18854 ;
  assign y3666 = ~n18861 ;
  assign y3667 = n18869 ;
  assign y3668 = ~n18872 ;
  assign y3669 = n18876 ;
  assign y3670 = n18880 ;
  assign y3671 = n18884 ;
  assign y3672 = ~n18885 ;
  assign y3673 = ~n18888 ;
  assign y3674 = ~n18899 ;
  assign y3675 = ~n18904 ;
  assign y3676 = n18909 ;
  assign y3677 = ~n18916 ;
  assign y3678 = n18925 ;
  assign y3679 = n18926 ;
  assign y3680 = n18927 ;
  assign y3681 = ~n18929 ;
  assign y3682 = ~1'b0 ;
  assign y3683 = ~n18938 ;
  assign y3684 = ~n18939 ;
  assign y3685 = ~n18944 ;
  assign y3686 = ~1'b0 ;
  assign y3687 = ~n18949 ;
  assign y3688 = n18950 ;
  assign y3689 = n18956 ;
  assign y3690 = n18960 ;
  assign y3691 = ~1'b0 ;
  assign y3692 = ~n18967 ;
  assign y3693 = ~n18970 ;
  assign y3694 = ~n18976 ;
  assign y3695 = ~n18980 ;
  assign y3696 = n18981 ;
  assign y3697 = n18985 ;
  assign y3698 = n18988 ;
  assign y3699 = ~n18992 ;
  assign y3700 = n18998 ;
  assign y3701 = n19001 ;
  assign y3702 = n19004 ;
  assign y3703 = ~n19015 ;
  assign y3704 = n19022 ;
  assign y3705 = n19025 ;
  assign y3706 = ~1'b0 ;
  assign y3707 = ~n19027 ;
  assign y3708 = ~n19028 ;
  assign y3709 = n19032 ;
  assign y3710 = n19042 ;
  assign y3711 = n19044 ;
  assign y3712 = n19049 ;
  assign y3713 = ~n19051 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = n19055 ;
  assign y3716 = ~1'b0 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = n19059 ;
  assign y3719 = ~n19060 ;
  assign y3720 = ~n19063 ;
  assign y3721 = ~n19066 ;
  assign y3722 = n19067 ;
  assign y3723 = n19070 ;
  assign y3724 = ~n19074 ;
  assign y3725 = ~n19076 ;
  assign y3726 = n19079 ;
  assign y3727 = ~n19082 ;
  assign y3728 = ~n19086 ;
  assign y3729 = ~1'b0 ;
  assign y3730 = ~n19091 ;
  assign y3731 = n19092 ;
  assign y3732 = n19096 ;
  assign y3733 = n19099 ;
  assign y3734 = ~n19100 ;
  assign y3735 = n19103 ;
  assign y3736 = n19104 ;
  assign y3737 = ~n19106 ;
  assign y3738 = ~n19113 ;
  assign y3739 = n19116 ;
  assign y3740 = ~n19126 ;
  assign y3741 = ~1'b0 ;
  assign y3742 = n19128 ;
  assign y3743 = ~n19131 ;
  assign y3744 = n19133 ;
  assign y3745 = n19136 ;
  assign y3746 = ~n19137 ;
  assign y3747 = ~n19144 ;
  assign y3748 = n19145 ;
  assign y3749 = ~n19147 ;
  assign y3750 = ~n19154 ;
  assign y3751 = n19162 ;
  assign y3752 = n19163 ;
  assign y3753 = ~n19171 ;
  assign y3754 = ~n19173 ;
  assign y3755 = n19187 ;
  assign y3756 = ~n19197 ;
  assign y3757 = n19202 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = n19210 ;
  assign y3760 = n19212 ;
  assign y3761 = n19217 ;
  assign y3762 = n19231 ;
  assign y3763 = ~n19237 ;
  assign y3764 = n19248 ;
  assign y3765 = ~n19252 ;
  assign y3766 = ~n19254 ;
  assign y3767 = n19260 ;
  assign y3768 = n19278 ;
  assign y3769 = ~n19279 ;
  assign y3770 = n19283 ;
  assign y3771 = ~1'b0 ;
  assign y3772 = ~n19287 ;
  assign y3773 = ~n19292 ;
  assign y3774 = ~n19293 ;
  assign y3775 = ~n19303 ;
  assign y3776 = n19307 ;
  assign y3777 = ~n19309 ;
  assign y3778 = n19312 ;
  assign y3779 = n19319 ;
  assign y3780 = ~1'b0 ;
  assign y3781 = n19329 ;
  assign y3782 = n19335 ;
  assign y3783 = n19345 ;
  assign y3784 = ~n19352 ;
  assign y3785 = n19354 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = ~n19358 ;
  assign y3788 = n19361 ;
  assign y3789 = ~n19364 ;
  assign y3790 = ~1'b0 ;
  assign y3791 = n19374 ;
  assign y3792 = ~n19377 ;
  assign y3793 = ~n19379 ;
  assign y3794 = ~n19389 ;
  assign y3795 = ~n19397 ;
  assign y3796 = n19414 ;
  assign y3797 = ~n19421 ;
  assign y3798 = ~n19422 ;
  assign y3799 = n19427 ;
  assign y3800 = ~n19433 ;
  assign y3801 = n19437 ;
  assign y3802 = n19440 ;
  assign y3803 = ~n19441 ;
  assign y3804 = ~n19443 ;
  assign y3805 = n19445 ;
  assign y3806 = n19447 ;
  assign y3807 = ~1'b0 ;
  assign y3808 = ~n19453 ;
  assign y3809 = ~n19467 ;
  assign y3810 = n19472 ;
  assign y3811 = ~n19474 ;
  assign y3812 = ~n19478 ;
  assign y3813 = n19480 ;
  assign y3814 = ~n10407 ;
  assign y3815 = n19481 ;
  assign y3816 = n19482 ;
  assign y3817 = ~n19489 ;
  assign y3818 = ~n19495 ;
  assign y3819 = n19497 ;
  assign y3820 = n19500 ;
  assign y3821 = n19503 ;
  assign y3822 = n19504 ;
  assign y3823 = ~n19505 ;
  assign y3824 = ~n19508 ;
  assign y3825 = n19509 ;
  assign y3826 = ~n19512 ;
  assign y3827 = n19522 ;
  assign y3828 = ~n19524 ;
  assign y3829 = n19526 ;
  assign y3830 = n19529 ;
  assign y3831 = n19534 ;
  assign y3832 = ~1'b0 ;
  assign y3833 = n19537 ;
  assign y3834 = ~n19540 ;
  assign y3835 = ~n19550 ;
  assign y3836 = ~n19561 ;
  assign y3837 = ~n19565 ;
  assign y3838 = n19569 ;
  assign y3839 = ~n19570 ;
  assign y3840 = ~n19573 ;
  assign y3841 = n19575 ;
  assign y3842 = n19578 ;
  assign y3843 = n19579 ;
  assign y3844 = ~n19583 ;
  assign y3845 = ~n19586 ;
  assign y3846 = ~n19587 ;
  assign y3847 = ~n19589 ;
  assign y3848 = ~1'b0 ;
  assign y3849 = n19590 ;
  assign y3850 = n19597 ;
  assign y3851 = n19601 ;
  assign y3852 = n19608 ;
  assign y3853 = n19610 ;
  assign y3854 = n19618 ;
  assign y3855 = n19621 ;
  assign y3856 = ~1'b0 ;
  assign y3857 = ~n19622 ;
  assign y3858 = ~n19624 ;
  assign y3859 = ~n19629 ;
  assign y3860 = ~n19631 ;
  assign y3861 = ~n19632 ;
  assign y3862 = ~n19637 ;
  assign y3863 = n19638 ;
  assign y3864 = ~n19642 ;
  assign y3865 = n19643 ;
  assign y3866 = n19644 ;
  assign y3867 = n19655 ;
  assign y3868 = n19662 ;
  assign y3869 = n19665 ;
  assign y3870 = ~1'b0 ;
  assign y3871 = ~1'b0 ;
  assign y3872 = n19667 ;
  assign y3873 = ~n19674 ;
  assign y3874 = ~n19676 ;
  assign y3875 = n19680 ;
  assign y3876 = ~n19685 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = ~n19687 ;
  assign y3879 = n19695 ;
  assign y3880 = n19700 ;
  assign y3881 = n19702 ;
  assign y3882 = ~n19703 ;
  assign y3883 = ~n19704 ;
  assign y3884 = n19708 ;
  assign y3885 = ~n19715 ;
  assign y3886 = ~n19723 ;
  assign y3887 = ~n19727 ;
  assign y3888 = n19740 ;
  assign y3889 = ~n19742 ;
  assign y3890 = n19744 ;
  assign y3891 = ~n19749 ;
  assign y3892 = ~n19754 ;
  assign y3893 = n19761 ;
  assign y3894 = n15961 ;
  assign y3895 = ~1'b0 ;
  assign y3896 = ~1'b0 ;
  assign y3897 = n19764 ;
  assign y3898 = ~n19765 ;
  assign y3899 = ~n19770 ;
  assign y3900 = n19772 ;
  assign y3901 = ~n19775 ;
  assign y3902 = ~n19778 ;
  assign y3903 = ~1'b0 ;
  assign y3904 = ~n19780 ;
  assign y3905 = n19787 ;
  assign y3906 = n19789 ;
  assign y3907 = n19793 ;
  assign y3908 = ~n19802 ;
  assign y3909 = ~1'b0 ;
  assign y3910 = n19804 ;
  assign y3911 = ~1'b0 ;
  assign y3912 = n19807 ;
  assign y3913 = n19812 ;
  assign y3914 = n19816 ;
  assign y3915 = ~n19820 ;
  assign y3916 = ~n19827 ;
  assign y3917 = ~1'b0 ;
  assign y3918 = ~n19830 ;
  assign y3919 = n19836 ;
  assign y3920 = ~n19841 ;
  assign y3921 = n19844 ;
  assign y3922 = n19847 ;
  assign y3923 = ~n19850 ;
  assign y3924 = ~n19856 ;
  assign y3925 = ~n19860 ;
  assign y3926 = ~n19868 ;
  assign y3927 = n19870 ;
  assign y3928 = ~n19874 ;
  assign y3929 = n19878 ;
  assign y3930 = ~n19889 ;
  assign y3931 = ~n19890 ;
  assign y3932 = n19892 ;
  assign y3933 = ~n19893 ;
  assign y3934 = n19898 ;
  assign y3935 = n19907 ;
  assign y3936 = ~n19909 ;
  assign y3937 = n19911 ;
  assign y3938 = ~n19912 ;
  assign y3939 = ~1'b0 ;
  assign y3940 = n19916 ;
  assign y3941 = n19920 ;
  assign y3942 = ~n19924 ;
  assign y3943 = ~n19925 ;
  assign y3944 = ~n19926 ;
  assign y3945 = ~n19935 ;
  assign y3946 = ~n19938 ;
  assign y3947 = ~1'b0 ;
  assign y3948 = n19940 ;
  assign y3949 = ~n19944 ;
  assign y3950 = ~n19947 ;
  assign y3951 = ~n19950 ;
  assign y3952 = ~n19954 ;
  assign y3953 = ~n19957 ;
  assign y3954 = ~n19963 ;
  assign y3955 = ~n19969 ;
  assign y3956 = ~n19976 ;
  assign y3957 = ~n19979 ;
  assign y3958 = n19981 ;
  assign y3959 = n19987 ;
  assign y3960 = ~1'b0 ;
  assign y3961 = ~n19989 ;
  assign y3962 = ~n19990 ;
  assign y3963 = n20000 ;
  assign y3964 = ~1'b0 ;
  assign y3965 = n20003 ;
  assign y3966 = ~n20007 ;
  assign y3967 = n20020 ;
  assign y3968 = n20023 ;
  assign y3969 = ~n15773 ;
  assign y3970 = ~n20024 ;
  assign y3971 = n20025 ;
  assign y3972 = ~n20035 ;
  assign y3973 = ~n20046 ;
  assign y3974 = ~n20054 ;
  assign y3975 = ~n20057 ;
  assign y3976 = ~n20060 ;
  assign y3977 = n20064 ;
  assign y3978 = n20071 ;
  assign y3979 = n20076 ;
  assign y3980 = n20083 ;
  assign y3981 = n20088 ;
  assign y3982 = n20093 ;
  assign y3983 = n20098 ;
  assign y3984 = n20103 ;
  assign y3985 = n20107 ;
  assign y3986 = ~n20110 ;
  assign y3987 = ~n20116 ;
  assign y3988 = ~n20117 ;
  assign y3989 = n20125 ;
  assign y3990 = ~n20126 ;
  assign y3991 = n20129 ;
  assign y3992 = ~n20131 ;
  assign y3993 = ~n20135 ;
  assign y3994 = ~n20138 ;
  assign y3995 = n20147 ;
  assign y3996 = ~n20151 ;
  assign y3997 = ~n20157 ;
  assign y3998 = ~n20174 ;
  assign y3999 = ~n20177 ;
  assign y4000 = n20183 ;
  assign y4001 = ~n20187 ;
  assign y4002 = n20191 ;
  assign y4003 = n20193 ;
  assign y4004 = ~n20195 ;
  assign y4005 = n20212 ;
  assign y4006 = ~n20215 ;
  assign y4007 = n20217 ;
  assign y4008 = n20219 ;
  assign y4009 = ~n20221 ;
  assign y4010 = n20225 ;
  assign y4011 = n20228 ;
  assign y4012 = ~n20230 ;
  assign y4013 = ~n20235 ;
  assign y4014 = n20241 ;
  assign y4015 = n20249 ;
  assign y4016 = ~n20256 ;
  assign y4017 = ~n20260 ;
  assign y4018 = n20262 ;
  assign y4019 = ~n20266 ;
  assign y4020 = ~n20271 ;
  assign y4021 = n20273 ;
  assign y4022 = n20281 ;
  assign y4023 = ~n20282 ;
  assign y4024 = n20283 ;
  assign y4025 = ~n20289 ;
  assign y4026 = ~n20293 ;
  assign y4027 = n20299 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = n20301 ;
  assign y4030 = ~n20305 ;
  assign y4031 = ~n20307 ;
  assign y4032 = n20311 ;
  assign y4033 = ~n20312 ;
  assign y4034 = n20314 ;
  assign y4035 = n20320 ;
  assign y4036 = ~n20324 ;
  assign y4037 = n20329 ;
  assign y4038 = ~n20330 ;
  assign y4039 = n20334 ;
  assign y4040 = n20336 ;
  assign y4041 = ~1'b0 ;
  assign y4042 = n20340 ;
  assign y4043 = n20342 ;
  assign y4044 = n20345 ;
  assign y4045 = n20352 ;
  assign y4046 = ~1'b0 ;
  assign y4047 = n20355 ;
  assign y4048 = ~n20358 ;
  assign y4049 = n20363 ;
  assign y4050 = ~n20364 ;
  assign y4051 = n20365 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = n20371 ;
  assign y4054 = ~n20376 ;
  assign y4055 = n20377 ;
  assign y4056 = ~n20381 ;
  assign y4057 = n20388 ;
  assign y4058 = ~n20392 ;
  assign y4059 = n20393 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = n20400 ;
  assign y4062 = n20404 ;
  assign y4063 = n20407 ;
  assign y4064 = ~n20408 ;
  assign y4065 = n20411 ;
  assign y4066 = ~1'b0 ;
  assign y4067 = ~n20423 ;
  assign y4068 = n20425 ;
  assign y4069 = ~n20428 ;
  assign y4070 = n20432 ;
  assign y4071 = ~n20439 ;
  assign y4072 = ~n20444 ;
  assign y4073 = ~n20446 ;
  assign y4074 = ~n20451 ;
  assign y4075 = n20452 ;
  assign y4076 = n20454 ;
  assign y4077 = ~1'b0 ;
  assign y4078 = ~n20456 ;
  assign y4079 = n20461 ;
  assign y4080 = ~n20463 ;
  assign y4081 = n20465 ;
  assign y4082 = ~n20466 ;
  assign y4083 = n20470 ;
  assign y4084 = ~n20472 ;
  assign y4085 = ~n20480 ;
  assign y4086 = ~n20481 ;
  assign y4087 = ~n20483 ;
  assign y4088 = n1967 ;
  assign y4089 = n20486 ;
  assign y4090 = n20494 ;
  assign y4091 = ~n20495 ;
  assign y4092 = n20497 ;
  assign y4093 = ~n20502 ;
  assign y4094 = ~n20503 ;
  assign y4095 = ~n20504 ;
  assign y4096 = ~1'b0 ;
  assign y4097 = n20509 ;
  assign y4098 = n20514 ;
  assign y4099 = ~n20518 ;
  assign y4100 = ~n20521 ;
  assign y4101 = n20525 ;
  assign y4102 = ~n20532 ;
  assign y4103 = ~n20535 ;
  assign y4104 = n20537 ;
  assign y4105 = ~n20541 ;
  assign y4106 = n20543 ;
  assign y4107 = n20553 ;
  assign y4108 = ~n20554 ;
  assign y4109 = ~n20560 ;
  assign y4110 = ~1'b0 ;
  assign y4111 = ~1'b0 ;
  assign y4112 = n20561 ;
  assign y4113 = n20564 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = ~n20566 ;
  assign y4116 = ~n20568 ;
  assign y4117 = n20570 ;
  assign y4118 = ~n20571 ;
  assign y4119 = ~n20578 ;
  assign y4120 = ~1'b0 ;
  assign y4121 = n20579 ;
  assign y4122 = n20584 ;
  assign y4123 = ~n20587 ;
  assign y4124 = n20588 ;
  assign y4125 = n20596 ;
  assign y4126 = n20599 ;
  assign y4127 = ~n20600 ;
  assign y4128 = ~n20604 ;
  assign y4129 = ~n20605 ;
  assign y4130 = ~n20610 ;
  assign y4131 = ~n20612 ;
  assign y4132 = ~n20614 ;
  assign y4133 = ~n20618 ;
  assign y4134 = ~n20627 ;
  assign y4135 = ~n20634 ;
  assign y4136 = ~n20641 ;
  assign y4137 = ~n20646 ;
  assign y4138 = ~n20648 ;
  assign y4139 = n20651 ;
  assign y4140 = ~n20653 ;
  assign y4141 = ~n20656 ;
  assign y4142 = ~n20657 ;
  assign y4143 = n20659 ;
  assign y4144 = n20662 ;
  assign y4145 = ~n20663 ;
  assign y4146 = n20671 ;
  assign y4147 = ~n20673 ;
  assign y4148 = ~n20679 ;
  assign y4149 = ~n20680 ;
  assign y4150 = ~n20681 ;
  assign y4151 = n20686 ;
  assign y4152 = ~n20693 ;
  assign y4153 = ~n20694 ;
  assign y4154 = n20698 ;
  assign y4155 = n20700 ;
  assign y4156 = ~n20701 ;
  assign y4157 = n20709 ;
  assign y4158 = ~n20714 ;
  assign y4159 = ~n20716 ;
  assign y4160 = n20720 ;
  assign y4161 = n20725 ;
  assign y4162 = ~n20734 ;
  assign y4163 = n20740 ;
  assign y4164 = n20745 ;
  assign y4165 = ~n20749 ;
  assign y4166 = ~n20751 ;
  assign y4167 = ~n20760 ;
  assign y4168 = n20766 ;
  assign y4169 = n20770 ;
  assign y4170 = ~n20774 ;
  assign y4171 = ~n20786 ;
  assign y4172 = ~n20792 ;
  assign y4173 = ~n20798 ;
  assign y4174 = n20802 ;
  assign y4175 = ~n20803 ;
  assign y4176 = ~n20804 ;
  assign y4177 = ~n20829 ;
  assign y4178 = ~n20834 ;
  assign y4179 = n20835 ;
  assign y4180 = x134 ;
  assign y4181 = n20837 ;
  assign y4182 = ~n20839 ;
  assign y4183 = ~n20842 ;
  assign y4184 = n20843 ;
  assign y4185 = ~n20846 ;
  assign y4186 = ~n20847 ;
  assign y4187 = ~n20856 ;
  assign y4188 = ~n20866 ;
  assign y4189 = ~n20869 ;
  assign y4190 = n20873 ;
  assign y4191 = n20875 ;
  assign y4192 = n20877 ;
  assign y4193 = ~n20880 ;
  assign y4194 = ~n20881 ;
  assign y4195 = ~n20882 ;
  assign y4196 = n20886 ;
  assign y4197 = ~n20888 ;
  assign y4198 = ~n20891 ;
  assign y4199 = n20895 ;
  assign y4200 = ~n20903 ;
  assign y4201 = ~n20910 ;
  assign y4202 = n20914 ;
  assign y4203 = ~n20918 ;
  assign y4204 = ~n20927 ;
  assign y4205 = n20930 ;
  assign y4206 = ~n20931 ;
  assign y4207 = ~n20938 ;
  assign y4208 = n20939 ;
  assign y4209 = ~n20951 ;
  assign y4210 = ~1'b0 ;
  assign y4211 = ~n20954 ;
  assign y4212 = n20962 ;
  assign y4213 = ~n20966 ;
  assign y4214 = n20974 ;
  assign y4215 = ~1'b0 ;
  assign y4216 = ~n20975 ;
  assign y4217 = n20979 ;
  assign y4218 = n20982 ;
  assign y4219 = n21000 ;
  assign y4220 = ~n21004 ;
  assign y4221 = n21011 ;
  assign y4222 = ~n21013 ;
  assign y4223 = ~n21015 ;
  assign y4224 = ~n8454 ;
  assign y4225 = n21017 ;
  assign y4226 = n21024 ;
  assign y4227 = ~1'b0 ;
  assign y4228 = n21029 ;
  assign y4229 = n21033 ;
  assign y4230 = n21035 ;
  assign y4231 = ~n21046 ;
  assign y4232 = n21048 ;
  assign y4233 = ~n21051 ;
  assign y4234 = n21056 ;
  assign y4235 = n21060 ;
  assign y4236 = ~n21064 ;
  assign y4237 = n21067 ;
  assign y4238 = ~n21069 ;
  assign y4239 = ~n21074 ;
  assign y4240 = n21075 ;
  assign y4241 = n21080 ;
  assign y4242 = ~n21085 ;
  assign y4243 = ~n21088 ;
  assign y4244 = ~1'b0 ;
  assign y4245 = n21089 ;
  assign y4246 = n21093 ;
  assign y4247 = ~n21098 ;
  assign y4248 = ~n21103 ;
  assign y4249 = ~n21104 ;
  assign y4250 = n21105 ;
  assign y4251 = ~n21108 ;
  assign y4252 = ~n21110 ;
  assign y4253 = ~n21114 ;
  assign y4254 = ~n21116 ;
  assign y4255 = n21117 ;
  assign y4256 = n21118 ;
  assign y4257 = ~n21127 ;
  assign y4258 = n21133 ;
  assign y4259 = ~n21135 ;
  assign y4260 = n21137 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = ~n21140 ;
  assign y4263 = n21144 ;
  assign y4264 = ~1'b0 ;
  assign y4265 = n21149 ;
  assign y4266 = ~n21153 ;
  assign y4267 = ~n21156 ;
  assign y4268 = n21159 ;
  assign y4269 = ~n21162 ;
  assign y4270 = ~n21164 ;
  assign y4271 = n21166 ;
  assign y4272 = n21169 ;
  assign y4273 = ~n21171 ;
  assign y4274 = n21174 ;
  assign y4275 = ~n21179 ;
  assign y4276 = n21181 ;
  assign y4277 = n21182 ;
  assign y4278 = ~n21184 ;
  assign y4279 = n21186 ;
  assign y4280 = ~n21196 ;
  assign y4281 = n21197 ;
  assign y4282 = n21198 ;
  assign y4283 = ~n21203 ;
  assign y4284 = ~n21208 ;
  assign y4285 = ~n21214 ;
  assign y4286 = ~n21224 ;
  assign y4287 = ~n21227 ;
  assign y4288 = ~n21228 ;
  assign y4289 = n21230 ;
  assign y4290 = n21231 ;
  assign y4291 = n21249 ;
  assign y4292 = n21264 ;
  assign y4293 = ~n21277 ;
  assign y4294 = ~n21281 ;
  assign y4295 = ~n21283 ;
  assign y4296 = ~n21284 ;
  assign y4297 = n21290 ;
  assign y4298 = ~n21291 ;
  assign y4299 = n21295 ;
  assign y4300 = ~n20246 ;
  assign y4301 = ~1'b0 ;
  assign y4302 = ~n21304 ;
  assign y4303 = n21307 ;
  assign y4304 = ~n13886 ;
  assign y4305 = ~1'b0 ;
  assign y4306 = ~n21310 ;
  assign y4307 = n21313 ;
  assign y4308 = ~n21325 ;
  assign y4309 = n21329 ;
  assign y4310 = ~n21331 ;
  assign y4311 = ~n21333 ;
  assign y4312 = n21336 ;
  assign y4313 = n21338 ;
  assign y4314 = n21342 ;
  assign y4315 = n21347 ;
  assign y4316 = n21351 ;
  assign y4317 = n21354 ;
  assign y4318 = n21356 ;
  assign y4319 = ~n21360 ;
  assign y4320 = ~n21366 ;
  assign y4321 = n21371 ;
  assign y4322 = n21390 ;
  assign y4323 = ~1'b0 ;
  assign y4324 = ~1'b0 ;
  assign y4325 = ~n21395 ;
  assign y4326 = ~n21397 ;
  assign y4327 = ~n21398 ;
  assign y4328 = ~n21401 ;
  assign y4329 = ~1'b0 ;
  assign y4330 = n21403 ;
  assign y4331 = n21404 ;
  assign y4332 = n21411 ;
  assign y4333 = n21414 ;
  assign y4334 = n21415 ;
  assign y4335 = ~n21423 ;
  assign y4336 = ~n21427 ;
  assign y4337 = n21432 ;
  assign y4338 = ~n21434 ;
  assign y4339 = ~n21443 ;
  assign y4340 = ~n21454 ;
  assign y4341 = n21462 ;
  assign y4342 = n21465 ;
  assign y4343 = n21468 ;
  assign y4344 = n21472 ;
  assign y4345 = ~n21474 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = ~n21476 ;
  assign y4348 = ~n21478 ;
  assign y4349 = ~n21489 ;
  assign y4350 = n21498 ;
  assign y4351 = ~n21502 ;
  assign y4352 = ~n21504 ;
  assign y4353 = n21509 ;
  assign y4354 = ~n21513 ;
  assign y4355 = ~n21517 ;
  assign y4356 = n21521 ;
  assign y4357 = n21523 ;
  assign y4358 = ~n21527 ;
  assign y4359 = ~n21530 ;
  assign y4360 = n21531 ;
  assign y4361 = ~n21536 ;
  assign y4362 = ~n21538 ;
  assign y4363 = ~n21540 ;
  assign y4364 = n21546 ;
  assign y4365 = ~n21547 ;
  assign y4366 = n21550 ;
  assign y4367 = n21558 ;
  assign y4368 = n21561 ;
  assign y4369 = n21571 ;
  assign y4370 = n21576 ;
  assign y4371 = n21577 ;
  assign y4372 = ~n21581 ;
  assign y4373 = ~n21596 ;
  assign y4374 = ~n21605 ;
  assign y4375 = ~1'b0 ;
  assign y4376 = n21613 ;
  assign y4377 = n21615 ;
  assign y4378 = ~n21618 ;
  assign y4379 = ~n21619 ;
  assign y4380 = n21620 ;
  assign y4381 = n21621 ;
  assign y4382 = n21625 ;
  assign y4383 = n21627 ;
  assign y4384 = ~n21630 ;
  assign y4385 = ~n21631 ;
  assign y4386 = n21634 ;
  assign y4387 = n21638 ;
  assign y4388 = n21643 ;
  assign y4389 = ~n21646 ;
  assign y4390 = ~n21651 ;
  assign y4391 = ~1'b0 ;
  assign y4392 = n21653 ;
  assign y4393 = n21655 ;
  assign y4394 = ~n21660 ;
  assign y4395 = ~1'b0 ;
  assign y4396 = n21667 ;
  assign y4397 = n21669 ;
  assign y4398 = n21673 ;
  assign y4399 = ~n21688 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = n21693 ;
  assign y4402 = n21694 ;
  assign y4403 = ~n21696 ;
  assign y4404 = n21697 ;
  assign y4405 = ~n21699 ;
  assign y4406 = ~n21703 ;
  assign y4407 = ~n21704 ;
  assign y4408 = n21721 ;
  assign y4409 = ~n21723 ;
  assign y4410 = ~n21729 ;
  assign y4411 = ~n21731 ;
  assign y4412 = ~1'b0 ;
  assign y4413 = ~n21739 ;
  assign y4414 = ~n21740 ;
  assign y4415 = n21744 ;
  assign y4416 = ~n21745 ;
  assign y4417 = ~n21750 ;
  assign y4418 = ~n21751 ;
  assign y4419 = ~1'b0 ;
  assign y4420 = ~n21753 ;
  assign y4421 = n21758 ;
  assign y4422 = ~n21760 ;
  assign y4423 = ~n21771 ;
  assign y4424 = n21775 ;
  assign y4425 = ~1'b0 ;
  assign y4426 = ~n21776 ;
  assign y4427 = n21782 ;
  assign y4428 = n21783 ;
  assign y4429 = n21787 ;
  assign y4430 = n21788 ;
  assign y4431 = n21789 ;
  assign y4432 = ~n21796 ;
  assign y4433 = n21802 ;
  assign y4434 = ~n21807 ;
  assign y4435 = ~n21812 ;
  assign y4436 = n21817 ;
  assign y4437 = n21822 ;
  assign y4438 = ~n21826 ;
  assign y4439 = ~n21837 ;
  assign y4440 = n21838 ;
  assign y4441 = n21844 ;
  assign y4442 = ~n21848 ;
  assign y4443 = ~n21849 ;
  assign y4444 = ~1'b0 ;
  assign y4445 = n21852 ;
  assign y4446 = ~n21853 ;
  assign y4447 = n21859 ;
  assign y4448 = n21866 ;
  assign y4449 = n18091 ;
  assign y4450 = n21873 ;
  assign y4451 = n21874 ;
  assign y4452 = n21875 ;
  assign y4453 = ~n21877 ;
  assign y4454 = n21885 ;
  assign y4455 = n21891 ;
  assign y4456 = n21896 ;
  assign y4457 = ~n21897 ;
  assign y4458 = n21903 ;
  assign y4459 = ~n21906 ;
  assign y4460 = ~n21914 ;
  assign y4461 = ~n21917 ;
  assign y4462 = n21923 ;
  assign y4463 = ~n21924 ;
  assign y4464 = ~n21931 ;
  assign y4465 = ~n21935 ;
  assign y4466 = ~n21938 ;
  assign y4467 = n21946 ;
  assign y4468 = ~n21949 ;
  assign y4469 = ~n21953 ;
  assign y4470 = n21956 ;
  assign y4471 = n21959 ;
  assign y4472 = ~n21962 ;
  assign y4473 = n21975 ;
  assign y4474 = ~n21988 ;
  assign y4475 = ~n21990 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = n21991 ;
  assign y4478 = n21992 ;
  assign y4479 = n21993 ;
  assign y4480 = ~n22000 ;
  assign y4481 = n22001 ;
  assign y4482 = ~n22006 ;
  assign y4483 = ~n22011 ;
  assign y4484 = ~n22017 ;
  assign y4485 = ~n22020 ;
  assign y4486 = ~n22027 ;
  assign y4487 = n22034 ;
  assign y4488 = ~n22042 ;
  assign y4489 = ~n22044 ;
  assign y4490 = ~n22046 ;
  assign y4491 = n22047 ;
  assign y4492 = ~n22050 ;
  assign y4493 = ~n22051 ;
  assign y4494 = ~n22054 ;
  assign y4495 = n22072 ;
  assign y4496 = n22076 ;
  assign y4497 = n22079 ;
  assign y4498 = n22082 ;
  assign y4499 = n22090 ;
  assign y4500 = ~n22091 ;
  assign y4501 = n22092 ;
  assign y4502 = ~n22096 ;
  assign y4503 = ~n22103 ;
  assign y4504 = ~n22104 ;
  assign y4505 = n22105 ;
  assign y4506 = n22106 ;
  assign y4507 = ~n22116 ;
  assign y4508 = ~n22117 ;
  assign y4509 = ~n22123 ;
  assign y4510 = n22127 ;
  assign y4511 = ~n22141 ;
  assign y4512 = n22144 ;
  assign y4513 = n22148 ;
  assign y4514 = ~n22149 ;
  assign y4515 = n22151 ;
  assign y4516 = n22155 ;
  assign y4517 = ~n22156 ;
  assign y4518 = ~n22161 ;
  assign y4519 = n22165 ;
  assign y4520 = n22167 ;
  assign y4521 = n22168 ;
  assign y4522 = n22173 ;
  assign y4523 = ~1'b0 ;
  assign y4524 = ~n22177 ;
  assign y4525 = n22182 ;
  assign y4526 = ~n22186 ;
  assign y4527 = ~n22188 ;
  assign y4528 = n22190 ;
  assign y4529 = ~n22193 ;
  assign y4530 = ~n22195 ;
  assign y4531 = n22198 ;
  assign y4532 = n22203 ;
  assign y4533 = n22205 ;
  assign y4534 = n22207 ;
  assign y4535 = ~n22212 ;
  assign y4536 = n22213 ;
  assign y4537 = ~n22222 ;
  assign y4538 = n22230 ;
  assign y4539 = ~n22234 ;
  assign y4540 = ~n22236 ;
  assign y4541 = ~n22240 ;
  assign y4542 = ~n22241 ;
  assign y4543 = n22248 ;
  assign y4544 = ~n22258 ;
  assign y4545 = n22259 ;
  assign y4546 = n22260 ;
  assign y4547 = ~n22262 ;
  assign y4548 = n22265 ;
  assign y4549 = n22280 ;
  assign y4550 = ~n22286 ;
  assign y4551 = ~n22295 ;
  assign y4552 = ~n22299 ;
  assign y4553 = ~n22304 ;
  assign y4554 = ~n22305 ;
  assign y4555 = n22306 ;
  assign y4556 = n22311 ;
  assign y4557 = n22313 ;
  assign y4558 = n22315 ;
  assign y4559 = ~n22316 ;
  assign y4560 = n22325 ;
  assign y4561 = n22333 ;
  assign y4562 = n22339 ;
  assign y4563 = ~n22342 ;
  assign y4564 = n22349 ;
  assign y4565 = ~n22352 ;
  assign y4566 = n22356 ;
  assign y4567 = n22359 ;
  assign y4568 = ~n22365 ;
  assign y4569 = ~n22366 ;
  assign y4570 = n22368 ;
  assign y4571 = ~n22370 ;
  assign y4572 = ~n22372 ;
  assign y4573 = ~n22375 ;
  assign y4574 = n22378 ;
  assign y4575 = ~n22383 ;
  assign y4576 = n22385 ;
  assign y4577 = n22387 ;
  assign y4578 = ~n22396 ;
  assign y4579 = n22398 ;
  assign y4580 = ~n22399 ;
  assign y4581 = ~1'b0 ;
  assign y4582 = ~n14431 ;
  assign y4583 = ~n22406 ;
  assign y4584 = ~n22409 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = ~n22416 ;
  assign y4587 = n22420 ;
  assign y4588 = n22425 ;
  assign y4589 = ~1'b0 ;
  assign y4590 = n22427 ;
  assign y4591 = ~n22432 ;
  assign y4592 = n22433 ;
  assign y4593 = ~n22435 ;
  assign y4594 = n22439 ;
  assign y4595 = ~n22440 ;
  assign y4596 = ~n22446 ;
  assign y4597 = ~n22452 ;
  assign y4598 = n22454 ;
  assign y4599 = n22458 ;
  assign y4600 = n22460 ;
  assign y4601 = ~n22461 ;
  assign y4602 = n22465 ;
  assign y4603 = n22470 ;
  assign y4604 = ~n22474 ;
  assign y4605 = n22476 ;
  assign y4606 = n22479 ;
  assign y4607 = ~n22480 ;
  assign y4608 = n22483 ;
  assign y4609 = ~n22492 ;
  assign y4610 = n22493 ;
  assign y4611 = n22497 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = n22503 ;
  assign y4614 = n22509 ;
  assign y4615 = n22521 ;
  assign y4616 = ~1'b0 ;
  assign y4617 = n22523 ;
  assign y4618 = ~n22526 ;
  assign y4619 = n22535 ;
  assign y4620 = n22536 ;
  assign y4621 = ~n22544 ;
  assign y4622 = n22545 ;
  assign y4623 = ~n22551 ;
  assign y4624 = ~n22558 ;
  assign y4625 = ~n22562 ;
  assign y4626 = n22573 ;
  assign y4627 = ~n22579 ;
  assign y4628 = n22581 ;
  assign y4629 = ~n22592 ;
  assign y4630 = ~n22598 ;
  assign y4631 = ~n22601 ;
  assign y4632 = n22606 ;
  assign y4633 = ~n22610 ;
  assign y4634 = n22612 ;
  assign y4635 = ~n22614 ;
  assign y4636 = n22618 ;
  assign y4637 = n22624 ;
  assign y4638 = n22625 ;
  assign y4639 = ~n22626 ;
  assign y4640 = ~n22629 ;
  assign y4641 = n22631 ;
  assign y4642 = n22634 ;
  assign y4643 = n22640 ;
  assign y4644 = ~1'b0 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = ~n22644 ;
  assign y4647 = n22645 ;
  assign y4648 = ~n22649 ;
  assign y4649 = ~n22653 ;
  assign y4650 = ~n22659 ;
  assign y4651 = n22661 ;
  assign y4652 = n22668 ;
  assign y4653 = ~1'b0 ;
  assign y4654 = ~1'b0 ;
  assign y4655 = n22669 ;
  assign y4656 = n22673 ;
  assign y4657 = ~1'b0 ;
  assign y4658 = n22674 ;
  assign y4659 = ~n22677 ;
  assign y4660 = ~n22682 ;
  assign y4661 = ~n22689 ;
  assign y4662 = n22693 ;
  assign y4663 = ~n22694 ;
  assign y4664 = ~n22699 ;
  assign y4665 = n22710 ;
  assign y4666 = n22714 ;
  assign y4667 = ~n22716 ;
  assign y4668 = ~n22719 ;
  assign y4669 = n22720 ;
  assign y4670 = n22721 ;
  assign y4671 = ~n22722 ;
  assign y4672 = ~n22731 ;
  assign y4673 = n22737 ;
  assign y4674 = ~n22738 ;
  assign y4675 = ~n22743 ;
  assign y4676 = ~n22746 ;
  assign y4677 = ~n22751 ;
  assign y4678 = n22753 ;
  assign y4679 = ~1'b0 ;
  assign y4680 = n22755 ;
  assign y4681 = n22762 ;
  assign y4682 = ~n22763 ;
  assign y4683 = ~n22767 ;
  assign y4684 = n22769 ;
  assign y4685 = ~n22772 ;
  assign y4686 = ~n22775 ;
  assign y4687 = ~n22785 ;
  assign y4688 = n22786 ;
  assign y4689 = n22792 ;
  assign y4690 = ~n22799 ;
  assign y4691 = ~n22806 ;
  assign y4692 = ~n22810 ;
  assign y4693 = ~n22812 ;
  assign y4694 = ~n22816 ;
  assign y4695 = ~n22818 ;
  assign y4696 = ~n22819 ;
  assign y4697 = n22829 ;
  assign y4698 = ~n22832 ;
  assign y4699 = n22835 ;
  assign y4700 = ~n22837 ;
  assign y4701 = n22838 ;
  assign y4702 = ~n22840 ;
  assign y4703 = ~n22842 ;
  assign y4704 = n22854 ;
  assign y4705 = ~n22860 ;
  assign y4706 = n22863 ;
  assign y4707 = ~1'b0 ;
  assign y4708 = ~n22864 ;
  assign y4709 = n22869 ;
  assign y4710 = ~n22877 ;
  assign y4711 = n22882 ;
  assign y4712 = n22886 ;
  assign y4713 = n22888 ;
  assign y4714 = ~n22890 ;
  assign y4715 = n22900 ;
  assign y4716 = ~n22901 ;
  assign y4717 = ~n22905 ;
  assign y4718 = n22915 ;
  assign y4719 = ~n22916 ;
  assign y4720 = ~n22921 ;
  assign y4721 = n22923 ;
  assign y4722 = ~n22924 ;
  assign y4723 = ~n22929 ;
  assign y4724 = ~n22930 ;
  assign y4725 = ~n22934 ;
  assign y4726 = ~n22937 ;
  assign y4727 = n22940 ;
  assign y4728 = ~n22953 ;
  assign y4729 = n22956 ;
  assign y4730 = ~n22962 ;
  assign y4731 = n22966 ;
  assign y4732 = ~n22967 ;
  assign y4733 = n22970 ;
  assign y4734 = n22973 ;
  assign y4735 = ~n22976 ;
  assign y4736 = n22979 ;
  assign y4737 = n22982 ;
  assign y4738 = ~n22988 ;
  assign y4739 = n22990 ;
  assign y4740 = ~n22992 ;
  assign y4741 = n22993 ;
  assign y4742 = n22994 ;
  assign y4743 = ~n22997 ;
  assign y4744 = ~n22999 ;
  assign y4745 = ~n23005 ;
  assign y4746 = n23006 ;
  assign y4747 = ~n23009 ;
  assign y4748 = n23011 ;
  assign y4749 = n23020 ;
  assign y4750 = ~n23022 ;
  assign y4751 = ~n23035 ;
  assign y4752 = ~n23039 ;
  assign y4753 = ~n23042 ;
  assign y4754 = ~n23045 ;
  assign y4755 = n23046 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = ~n23048 ;
  assign y4758 = ~n23052 ;
  assign y4759 = n23055 ;
  assign y4760 = n23056 ;
  assign y4761 = ~n23068 ;
  assign y4762 = n23070 ;
  assign y4763 = ~n23081 ;
  assign y4764 = ~n23094 ;
  assign y4765 = n23098 ;
  assign y4766 = ~n23106 ;
  assign y4767 = n23108 ;
  assign y4768 = ~n23111 ;
  assign y4769 = n23113 ;
  assign y4770 = n23114 ;
  assign y4771 = n23116 ;
  assign y4772 = ~n23124 ;
  assign y4773 = ~n23125 ;
  assign y4774 = ~n23140 ;
  assign y4775 = ~n23141 ;
  assign y4776 = ~1'b0 ;
  assign y4777 = ~n23148 ;
  assign y4778 = n23155 ;
  assign y4779 = ~n23156 ;
  assign y4780 = n23163 ;
  assign y4781 = n23164 ;
  assign y4782 = n23167 ;
  assign y4783 = ~n23169 ;
  assign y4784 = n23172 ;
  assign y4785 = n23177 ;
  assign y4786 = ~1'b0 ;
  assign y4787 = ~n23179 ;
  assign y4788 = ~n23182 ;
  assign y4789 = ~n23183 ;
  assign y4790 = n23186 ;
  assign y4791 = ~n23188 ;
  assign y4792 = n23195 ;
  assign y4793 = ~n23202 ;
  assign y4794 = ~n23206 ;
  assign y4795 = n23209 ;
  assign y4796 = n23211 ;
  assign y4797 = ~n23212 ;
  assign y4798 = ~n23213 ;
  assign y4799 = n23216 ;
  assign y4800 = ~n23217 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = n23219 ;
  assign y4803 = n23222 ;
  assign y4804 = ~n23223 ;
  assign y4805 = ~n23228 ;
  assign y4806 = n23233 ;
  assign y4807 = ~n23237 ;
  assign y4808 = ~n23242 ;
  assign y4809 = ~n23247 ;
  assign y4810 = n23252 ;
  assign y4811 = ~n23254 ;
  assign y4812 = ~n23255 ;
  assign y4813 = ~1'b0 ;
  assign y4814 = n23263 ;
  assign y4815 = n23264 ;
  assign y4816 = n23267 ;
  assign y4817 = n23269 ;
  assign y4818 = n23270 ;
  assign y4819 = n23271 ;
  assign y4820 = n23273 ;
  assign y4821 = n23274 ;
  assign y4822 = ~1'b0 ;
  assign y4823 = n23282 ;
  assign y4824 = ~n23283 ;
  assign y4825 = ~1'b0 ;
  assign y4826 = n23286 ;
  assign y4827 = ~n23291 ;
  assign y4828 = n23292 ;
  assign y4829 = ~n23297 ;
  assign y4830 = ~n23300 ;
  assign y4831 = n23301 ;
  assign y4832 = n23304 ;
  assign y4833 = n23309 ;
  assign y4834 = n23315 ;
  assign y4835 = n23322 ;
  assign y4836 = ~n23327 ;
  assign y4837 = ~n23330 ;
  assign y4838 = n23337 ;
  assign y4839 = ~n23338 ;
  assign y4840 = ~n23339 ;
  assign y4841 = ~n23341 ;
  assign y4842 = n23342 ;
  assign y4843 = n23345 ;
  assign y4844 = ~n23347 ;
  assign y4845 = ~n23349 ;
  assign y4846 = n23350 ;
  assign y4847 = ~1'b0 ;
  assign y4848 = ~n23357 ;
  assign y4849 = ~n23362 ;
  assign y4850 = ~n23367 ;
  assign y4851 = n23376 ;
  assign y4852 = ~n23381 ;
  assign y4853 = ~n23387 ;
  assign y4854 = ~n23392 ;
  assign y4855 = ~n23396 ;
  assign y4856 = ~n20016 ;
  assign y4857 = ~n23399 ;
  assign y4858 = n23400 ;
  assign y4859 = ~n23405 ;
  assign y4860 = ~1'b0 ;
  assign y4861 = n23407 ;
  assign y4862 = ~n23409 ;
  assign y4863 = n23419 ;
  assign y4864 = n23421 ;
  assign y4865 = ~1'b0 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = ~n23425 ;
  assign y4868 = n23433 ;
  assign y4869 = n23440 ;
  assign y4870 = ~n23441 ;
  assign y4871 = ~n23445 ;
  assign y4872 = n23449 ;
  assign y4873 = n23453 ;
  assign y4874 = n23455 ;
  assign y4875 = ~n23460 ;
  assign y4876 = ~n23467 ;
  assign y4877 = n23469 ;
  assign y4878 = ~1'b0 ;
  assign y4879 = ~n23472 ;
  assign y4880 = ~n23475 ;
  assign y4881 = n23480 ;
  assign y4882 = n23483 ;
  assign y4883 = ~1'b0 ;
  assign y4884 = n23487 ;
  assign y4885 = n23488 ;
  assign y4886 = n23490 ;
  assign y4887 = n23497 ;
  assign y4888 = ~n23499 ;
  assign y4889 = ~n23507 ;
  assign y4890 = ~n23516 ;
  assign y4891 = n23522 ;
  assign y4892 = n23526 ;
  assign y4893 = ~n23527 ;
  assign y4894 = n23528 ;
  assign y4895 = ~n23529 ;
  assign y4896 = n23533 ;
  assign y4897 = n23534 ;
  assign y4898 = n23535 ;
  assign y4899 = ~n23536 ;
  assign y4900 = n23539 ;
  assign y4901 = n23540 ;
  assign y4902 = n23542 ;
  assign y4903 = n23552 ;
  assign y4904 = ~1'b0 ;
  assign y4905 = n23558 ;
  assign y4906 = n23559 ;
  assign y4907 = n23560 ;
  assign y4908 = n6741 ;
  assign y4909 = ~n23562 ;
  assign y4910 = n23564 ;
  assign y4911 = ~n23571 ;
  assign y4912 = n23572 ;
  assign y4913 = ~n23577 ;
  assign y4914 = ~n23581 ;
  assign y4915 = ~1'b0 ;
  assign y4916 = ~n20348 ;
  assign y4917 = n23592 ;
  assign y4918 = ~1'b0 ;
  assign y4919 = ~n23594 ;
  assign y4920 = n23605 ;
  assign y4921 = n23609 ;
  assign y4922 = n23611 ;
  assign y4923 = n23612 ;
  assign y4924 = ~n23614 ;
  assign y4925 = ~n23616 ;
  assign y4926 = ~n23623 ;
  assign y4927 = ~1'b0 ;
  assign y4928 = n23641 ;
  assign y4929 = ~n23642 ;
  assign y4930 = ~n23644 ;
  assign y4931 = n23648 ;
  assign y4932 = ~n23652 ;
  assign y4933 = ~1'b0 ;
  assign y4934 = ~n23653 ;
  assign y4935 = n23654 ;
  assign y4936 = ~n23659 ;
  assign y4937 = ~n23664 ;
  assign y4938 = n23665 ;
  assign y4939 = n23672 ;
  assign y4940 = ~n23675 ;
  assign y4941 = n23681 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = n23683 ;
  assign y4944 = ~n23693 ;
  assign y4945 = n23696 ;
  assign y4946 = ~n23697 ;
  assign y4947 = n23698 ;
  assign y4948 = ~n23700 ;
  assign y4949 = ~n23706 ;
  assign y4950 = n23712 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = ~1'b0 ;
  assign y4953 = n23722 ;
  assign y4954 = ~n23727 ;
  assign y4955 = ~n23731 ;
  assign y4956 = n23739 ;
  assign y4957 = ~n23744 ;
  assign y4958 = n23747 ;
  assign y4959 = ~n23753 ;
  assign y4960 = n23756 ;
  assign y4961 = n23757 ;
  assign y4962 = n23759 ;
  assign y4963 = ~n23769 ;
  assign y4964 = ~n23788 ;
  assign y4965 = ~1'b0 ;
  assign y4966 = ~n23791 ;
  assign y4967 = ~n23795 ;
  assign y4968 = n23797 ;
  assign y4969 = ~n23803 ;
  assign y4970 = ~n23804 ;
  assign y4971 = ~n23810 ;
  assign y4972 = n23811 ;
  assign y4973 = n23817 ;
  assign y4974 = ~n23820 ;
  assign y4975 = n23823 ;
  assign y4976 = n23824 ;
  assign y4977 = n23825 ;
  assign y4978 = ~n23831 ;
  assign y4979 = n23835 ;
  assign y4980 = n23844 ;
  assign y4981 = ~n23845 ;
  assign y4982 = ~n23846 ;
  assign y4983 = ~n23849 ;
  assign y4984 = n23851 ;
  assign y4985 = ~n23852 ;
  assign y4986 = n23855 ;
  assign y4987 = ~n23858 ;
  assign y4988 = n23861 ;
  assign y4989 = ~n23866 ;
  assign y4990 = n23874 ;
  assign y4991 = ~n23878 ;
  assign y4992 = ~1'b0 ;
  assign y4993 = ~n23887 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~n23892 ;
  assign y4996 = n23896 ;
  assign y4997 = n23897 ;
  assign y4998 = n23899 ;
  assign y4999 = n23900 ;
  assign y5000 = ~n23912 ;
  assign y5001 = n23913 ;
  assign y5002 = ~n23914 ;
  assign y5003 = ~1'b0 ;
  assign y5004 = ~1'b0 ;
  assign y5005 = ~n23915 ;
  assign y5006 = n23916 ;
  assign y5007 = n9240 ;
  assign y5008 = ~n23917 ;
  assign y5009 = ~n23925 ;
  assign y5010 = n23930 ;
  assign y5011 = n23932 ;
  assign y5012 = ~n23937 ;
  assign y5013 = ~n23941 ;
  assign y5014 = n23944 ;
  assign y5015 = ~n23947 ;
  assign y5016 = n23952 ;
  assign y5017 = ~n23959 ;
  assign y5018 = ~n23960 ;
  assign y5019 = ~n23965 ;
  assign y5020 = ~n23966 ;
  assign y5021 = n23970 ;
  assign y5022 = ~n23971 ;
  assign y5023 = ~n23976 ;
  assign y5024 = n23983 ;
  assign y5025 = n23984 ;
  assign y5026 = ~n23985 ;
  assign y5027 = ~n23989 ;
  assign y5028 = ~n24003 ;
  assign y5029 = n24005 ;
  assign y5030 = ~n24007 ;
  assign y5031 = n24015 ;
  assign y5032 = n24022 ;
  assign y5033 = n24025 ;
  assign y5034 = ~n24035 ;
  assign y5035 = ~n24041 ;
  assign y5036 = ~n24042 ;
  assign y5037 = ~n24044 ;
  assign y5038 = ~1'b0 ;
  assign y5039 = ~n24045 ;
  assign y5040 = n24050 ;
  assign y5041 = n24051 ;
  assign y5042 = ~n24067 ;
  assign y5043 = n24070 ;
  assign y5044 = ~n24072 ;
  assign y5045 = ~n24073 ;
  assign y5046 = ~n24081 ;
  assign y5047 = n24092 ;
  assign y5048 = ~n24093 ;
  assign y5049 = ~1'b0 ;
  assign y5050 = ~n24097 ;
  assign y5051 = ~1'b0 ;
  assign y5052 = ~n24099 ;
  assign y5053 = ~n6935 ;
  assign y5054 = ~n24104 ;
  assign y5055 = ~n24106 ;
  assign y5056 = ~n24119 ;
  assign y5057 = ~n24121 ;
  assign y5058 = ~n24123 ;
  assign y5059 = ~n24132 ;
  assign y5060 = ~n24133 ;
  assign y5061 = ~n24134 ;
  assign y5062 = n24135 ;
  assign y5063 = ~n24145 ;
  assign y5064 = ~1'b0 ;
  assign y5065 = ~n24151 ;
  assign y5066 = ~n24153 ;
  assign y5067 = n24154 ;
  assign y5068 = n24156 ;
  assign y5069 = ~n24158 ;
  assign y5070 = ~n24161 ;
  assign y5071 = n24166 ;
  assign y5072 = n24176 ;
  assign y5073 = n24188 ;
  assign y5074 = n24190 ;
  assign y5075 = ~n24196 ;
  assign y5076 = ~n24200 ;
  assign y5077 = n24213 ;
  assign y5078 = ~n24216 ;
  assign y5079 = n24222 ;
  assign y5080 = ~n24226 ;
  assign y5081 = n24232 ;
  assign y5082 = n24235 ;
  assign y5083 = ~n24245 ;
  assign y5084 = n24247 ;
  assign y5085 = ~n24250 ;
  assign y5086 = ~n24251 ;
  assign y5087 = n24253 ;
  assign y5088 = ~n24257 ;
  assign y5089 = n24260 ;
  assign y5090 = n24263 ;
  assign y5091 = n24273 ;
  assign y5092 = ~n24275 ;
  assign y5093 = n24277 ;
  assign y5094 = n15728 ;
  assign y5095 = n24281 ;
  assign y5096 = n24283 ;
  assign y5097 = ~n10797 ;
  assign y5098 = ~n24286 ;
  assign y5099 = ~n24290 ;
  assign y5100 = n24292 ;
  assign y5101 = ~n24297 ;
  assign y5102 = ~n24298 ;
  assign y5103 = n24301 ;
  assign y5104 = ~n24305 ;
  assign y5105 = ~n24306 ;
  assign y5106 = ~n24307 ;
  assign y5107 = ~n24309 ;
  assign y5108 = ~n24311 ;
  assign y5109 = n24312 ;
  assign y5110 = ~n24314 ;
  assign y5111 = ~n24320 ;
  assign y5112 = ~n24323 ;
  assign y5113 = ~n24327 ;
  assign y5114 = n24331 ;
  assign y5115 = ~n24334 ;
  assign y5116 = n24336 ;
  assign y5117 = ~1'b0 ;
  assign y5118 = n24341 ;
  assign y5119 = ~n24347 ;
  assign y5120 = n24354 ;
  assign y5121 = n24356 ;
  assign y5122 = ~n24366 ;
  assign y5123 = ~n24368 ;
  assign y5124 = n24378 ;
  assign y5125 = n24379 ;
  assign y5126 = n24381 ;
  assign y5127 = n24382 ;
  assign y5128 = ~n24384 ;
  assign y5129 = ~n24385 ;
  assign y5130 = ~n24389 ;
  assign y5131 = n24390 ;
  assign y5132 = n24399 ;
  assign y5133 = n24404 ;
  assign y5134 = ~n24405 ;
  assign y5135 = ~n24409 ;
  assign y5136 = ~n24412 ;
  assign y5137 = n24413 ;
  assign y5138 = n24415 ;
  assign y5139 = ~n24417 ;
  assign y5140 = ~n24422 ;
  assign y5141 = ~n24424 ;
  assign y5142 = ~n24428 ;
  assign y5143 = ~n24437 ;
  assign y5144 = ~n24438 ;
  assign y5145 = ~n24447 ;
  assign y5146 = n24448 ;
  assign y5147 = ~n24450 ;
  assign y5148 = ~n24451 ;
  assign y5149 = ~n24455 ;
  assign y5150 = n24456 ;
  assign y5151 = ~1'b0 ;
  assign y5152 = ~n24457 ;
  assign y5153 = ~n24458 ;
  assign y5154 = ~n24462 ;
  assign y5155 = n24463 ;
  assign y5156 = n24467 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = ~n24469 ;
  assign y5159 = ~n24470 ;
  assign y5160 = ~n24471 ;
  assign y5161 = ~n24475 ;
  assign y5162 = ~1'b0 ;
  assign y5163 = ~n24477 ;
  assign y5164 = ~n24478 ;
  assign y5165 = ~n24481 ;
  assign y5166 = ~n24483 ;
  assign y5167 = ~n24491 ;
  assign y5168 = n24501 ;
  assign y5169 = n24504 ;
  assign y5170 = ~n24516 ;
  assign y5171 = n24519 ;
  assign y5172 = ~n24527 ;
  assign y5173 = ~n24528 ;
  assign y5174 = ~n24530 ;
  assign y5175 = ~n24536 ;
  assign y5176 = ~n24538 ;
  assign y5177 = ~n24545 ;
  assign y5178 = ~n24549 ;
  assign y5179 = n24553 ;
  assign y5180 = n24554 ;
  assign y5181 = ~n24556 ;
  assign y5182 = ~n24560 ;
  assign y5183 = ~n24563 ;
  assign y5184 = n24567 ;
  assign y5185 = ~n24569 ;
  assign y5186 = ~n24572 ;
  assign y5187 = ~1'b0 ;
  assign y5188 = n24576 ;
  assign y5189 = ~n24577 ;
  assign y5190 = n24583 ;
  assign y5191 = ~1'b0 ;
  assign y5192 = ~n24587 ;
  assign y5193 = ~1'b0 ;
  assign y5194 = n24588 ;
  assign y5195 = n24595 ;
  assign y5196 = n24596 ;
  assign y5197 = ~n24600 ;
  assign y5198 = ~n24601 ;
  assign y5199 = ~n24602 ;
  assign y5200 = n24605 ;
  assign y5201 = ~n24606 ;
  assign y5202 = ~n24608 ;
  assign y5203 = ~n24609 ;
  assign y5204 = ~n24613 ;
  assign y5205 = n24618 ;
  assign y5206 = ~n24624 ;
  assign y5207 = ~n24625 ;
  assign y5208 = n24631 ;
  assign y5209 = ~n24632 ;
  assign y5210 = ~n24635 ;
  assign y5211 = ~n24636 ;
  assign y5212 = ~n24639 ;
  assign y5213 = n24644 ;
  assign y5214 = ~n24655 ;
  assign y5215 = ~n24659 ;
  assign y5216 = n24662 ;
  assign y5217 = n24666 ;
  assign y5218 = ~n24669 ;
  assign y5219 = ~1'b0 ;
  assign y5220 = n24671 ;
  assign y5221 = n24673 ;
  assign y5222 = ~n24676 ;
  assign y5223 = n24683 ;
  assign y5224 = n24688 ;
  assign y5225 = n24692 ;
  assign y5226 = ~1'b0 ;
  assign y5227 = n24693 ;
  assign y5228 = n24697 ;
  assign y5229 = n24706 ;
  assign y5230 = ~n24714 ;
  assign y5231 = ~n24718 ;
  assign y5232 = ~n24720 ;
  assign y5233 = n24724 ;
  assign y5234 = ~n24725 ;
  assign y5235 = ~n24730 ;
  assign y5236 = ~n24732 ;
  assign y5237 = n24736 ;
  assign y5238 = n24738 ;
  assign y5239 = n24743 ;
  assign y5240 = ~n24754 ;
  assign y5241 = ~n24758 ;
  assign y5242 = ~n24760 ;
  assign y5243 = ~n24763 ;
  assign y5244 = n24764 ;
  assign y5245 = n24765 ;
  assign y5246 = ~n24766 ;
  assign y5247 = n24774 ;
  assign y5248 = ~n24779 ;
  assign y5249 = ~n24787 ;
  assign y5250 = ~n24789 ;
  assign y5251 = n24799 ;
  assign y5252 = ~n24803 ;
  assign y5253 = n24813 ;
  assign y5254 = ~1'b0 ;
  assign y5255 = n24816 ;
  assign y5256 = n24821 ;
  assign y5257 = ~n24823 ;
  assign y5258 = ~n24833 ;
  assign y5259 = n24837 ;
  assign y5260 = ~n24840 ;
  assign y5261 = ~n24842 ;
  assign y5262 = ~n24848 ;
  assign y5263 = ~n24856 ;
  assign y5264 = n24859 ;
  assign y5265 = n24863 ;
  assign y5266 = n24864 ;
  assign y5267 = ~n24868 ;
  assign y5268 = n24872 ;
  assign y5269 = n24876 ;
  assign y5270 = n24878 ;
  assign y5271 = n24880 ;
  assign y5272 = n24890 ;
  assign y5273 = ~n24893 ;
  assign y5274 = ~n24894 ;
  assign y5275 = ~n24899 ;
  assign y5276 = n24903 ;
  assign y5277 = ~n24910 ;
  assign y5278 = ~1'b0 ;
  assign y5279 = ~n24911 ;
  assign y5280 = ~n24912 ;
  assign y5281 = ~n24915 ;
  assign y5282 = ~n24917 ;
  assign y5283 = ~n24920 ;
  assign y5284 = ~n24924 ;
  assign y5285 = ~n24926 ;
  assign y5286 = ~n24930 ;
  assign y5287 = ~1'b0 ;
  assign y5288 = n24934 ;
  assign y5289 = ~n24943 ;
  assign y5290 = ~n24944 ;
  assign y5291 = n24953 ;
  assign y5292 = ~n24960 ;
  assign y5293 = n24962 ;
  assign y5294 = ~n24965 ;
  assign y5295 = ~n24971 ;
  assign y5296 = ~n24973 ;
  assign y5297 = n24975 ;
  assign y5298 = n24977 ;
  assign y5299 = ~n24980 ;
  assign y5300 = ~n24987 ;
  assign y5301 = ~n24989 ;
  assign y5302 = ~n24995 ;
  assign y5303 = ~n24997 ;
  assign y5304 = n24999 ;
  assign y5305 = ~n25002 ;
  assign y5306 = n25005 ;
  assign y5307 = n25007 ;
  assign y5308 = n25008 ;
  assign y5309 = ~n25014 ;
  assign y5310 = ~n25017 ;
  assign y5311 = n25018 ;
  assign y5312 = n25024 ;
  assign y5313 = ~n25028 ;
  assign y5314 = ~n25045 ;
  assign y5315 = ~n25046 ;
  assign y5316 = n25048 ;
  assign y5317 = n25054 ;
  assign y5318 = ~n25056 ;
  assign y5319 = ~n25059 ;
  assign y5320 = n25062 ;
  assign y5321 = n25063 ;
  assign y5322 = n25065 ;
  assign y5323 = n25072 ;
  assign y5324 = ~n25077 ;
  assign y5325 = ~1'b0 ;
  assign y5326 = ~n25081 ;
  assign y5327 = ~n25083 ;
  assign y5328 = n25084 ;
  assign y5329 = n25088 ;
  assign y5330 = n25090 ;
  assign y5331 = ~1'b0 ;
  assign y5332 = ~n25092 ;
  assign y5333 = ~n25098 ;
  assign y5334 = ~n25099 ;
  assign y5335 = ~n25106 ;
  assign y5336 = ~1'b0 ;
  assign y5337 = ~1'b0 ;
  assign y5338 = ~n25107 ;
  assign y5339 = n25111 ;
  assign y5340 = n25119 ;
  assign y5341 = ~n25122 ;
  assign y5342 = ~n25123 ;
  assign y5343 = ~n25127 ;
  assign y5344 = n25129 ;
  assign y5345 = ~n25131 ;
  assign y5346 = ~n25138 ;
  assign y5347 = n25144 ;
  assign y5348 = ~n25145 ;
  assign y5349 = n25146 ;
  assign y5350 = n25150 ;
  assign y5351 = ~n25153 ;
  assign y5352 = ~n25161 ;
  assign y5353 = n25163 ;
  assign y5354 = ~n25167 ;
  assign y5355 = ~n25170 ;
  assign y5356 = ~n25174 ;
  assign y5357 = ~n25175 ;
  assign y5358 = ~n25177 ;
  assign y5359 = n25181 ;
  assign y5360 = ~n25182 ;
  assign y5361 = n25184 ;
  assign y5362 = ~n25187 ;
  assign y5363 = ~n25189 ;
  assign y5364 = n25190 ;
  assign y5365 = n25194 ;
  assign y5366 = n25195 ;
  assign y5367 = n25201 ;
  assign y5368 = n25206 ;
  assign y5369 = ~n25212 ;
  assign y5370 = ~n25216 ;
  assign y5371 = ~n25224 ;
  assign y5372 = n25233 ;
  assign y5373 = n25234 ;
  assign y5374 = n25237 ;
  assign y5375 = n25238 ;
  assign y5376 = n25240 ;
  assign y5377 = ~n25245 ;
  assign y5378 = ~n25248 ;
  assign y5379 = n25251 ;
  assign y5380 = ~n25256 ;
  assign y5381 = ~1'b0 ;
  assign y5382 = n25257 ;
  assign y5383 = ~n25258 ;
  assign y5384 = n25268 ;
  assign y5385 = ~n25270 ;
  assign y5386 = ~1'b0 ;
  assign y5387 = ~n25271 ;
  assign y5388 = n25278 ;
  assign y5389 = n25281 ;
  assign y5390 = ~n25284 ;
  assign y5391 = n25288 ;
  assign y5392 = ~n25290 ;
  assign y5393 = n25291 ;
  assign y5394 = ~n25295 ;
  assign y5395 = ~n25302 ;
  assign y5396 = ~n25303 ;
  assign y5397 = n25318 ;
  assign y5398 = ~1'b0 ;
  assign y5399 = ~n25322 ;
  assign y5400 = n25331 ;
  assign y5401 = ~n25333 ;
  assign y5402 = ~n25335 ;
  assign y5403 = ~n25339 ;
  assign y5404 = ~n25351 ;
  assign y5405 = n25359 ;
  assign y5406 = n25361 ;
  assign y5407 = ~n25362 ;
  assign y5408 = ~n25363 ;
  assign y5409 = n25364 ;
  assign y5410 = n25366 ;
  assign y5411 = n25370 ;
  assign y5412 = ~n25372 ;
  assign y5413 = ~n25374 ;
  assign y5414 = n25382 ;
  assign y5415 = ~n25383 ;
  assign y5416 = n25385 ;
  assign y5417 = n25386 ;
  assign y5418 = ~n25387 ;
  assign y5419 = ~n25392 ;
  assign y5420 = ~n25397 ;
  assign y5421 = n25398 ;
  assign y5422 = n25404 ;
  assign y5423 = n25409 ;
  assign y5424 = ~n25410 ;
  assign y5425 = n25418 ;
  assign y5426 = ~n25424 ;
  assign y5427 = n25427 ;
  assign y5428 = ~n25430 ;
  assign y5429 = ~n25434 ;
  assign y5430 = ~n25436 ;
  assign y5431 = ~n25440 ;
  assign y5432 = ~n25444 ;
  assign y5433 = n25449 ;
  assign y5434 = n25457 ;
  assign y5435 = n25460 ;
  assign y5436 = n25470 ;
  assign y5437 = n25476 ;
  assign y5438 = ~n25480 ;
  assign y5439 = ~n25482 ;
  assign y5440 = ~n25483 ;
  assign y5441 = ~n25484 ;
  assign y5442 = ~n25488 ;
  assign y5443 = n25489 ;
  assign y5444 = ~n25492 ;
  assign y5445 = n25494 ;
  assign y5446 = n25497 ;
  assign y5447 = n25502 ;
  assign y5448 = ~1'b0 ;
  assign y5449 = n25503 ;
  assign y5450 = n25505 ;
  assign y5451 = ~n25513 ;
  assign y5452 = ~n25517 ;
  assign y5453 = n25519 ;
  assign y5454 = n25520 ;
  assign y5455 = n25523 ;
  assign y5456 = ~n25526 ;
  assign y5457 = n25535 ;
  assign y5458 = n25536 ;
  assign y5459 = n25539 ;
  assign y5460 = n25544 ;
  assign y5461 = n25554 ;
  assign y5462 = ~n25558 ;
  assign y5463 = ~1'b0 ;
  assign y5464 = n25568 ;
  assign y5465 = ~n25570 ;
  assign y5466 = n25583 ;
  assign y5467 = ~n25584 ;
  assign y5468 = ~n25589 ;
  assign y5469 = n25593 ;
  assign y5470 = n25594 ;
  assign y5471 = n25598 ;
  assign y5472 = n25602 ;
  assign y5473 = n25605 ;
  assign y5474 = ~n25607 ;
  assign y5475 = ~n25610 ;
  assign y5476 = ~n25615 ;
  assign y5477 = ~n25620 ;
  assign y5478 = ~1'b0 ;
  assign y5479 = n25621 ;
  assign y5480 = n25629 ;
  assign y5481 = ~n25631 ;
  assign y5482 = n25634 ;
  assign y5483 = ~n25636 ;
  assign y5484 = ~n25638 ;
  assign y5485 = n25640 ;
  assign y5486 = ~n25641 ;
  assign y5487 = n25645 ;
  assign y5488 = ~n25653 ;
  assign y5489 = ~n25656 ;
  assign y5490 = ~n25658 ;
  assign y5491 = ~n25659 ;
  assign y5492 = ~n25663 ;
  assign y5493 = n25668 ;
  assign y5494 = ~n25675 ;
  assign y5495 = n25677 ;
  assign y5496 = ~n25678 ;
  assign y5497 = ~n25687 ;
  assign y5498 = ~n25689 ;
  assign y5499 = n25692 ;
  assign y5500 = ~n25695 ;
  assign y5501 = n25697 ;
  assign y5502 = ~n25706 ;
  assign y5503 = ~n25710 ;
  assign y5504 = ~n25722 ;
  assign y5505 = ~1'b0 ;
  assign y5506 = n25723 ;
  assign y5507 = ~n25728 ;
  assign y5508 = ~n25731 ;
  assign y5509 = n25733 ;
  assign y5510 = n25736 ;
  assign y5511 = ~n25741 ;
  assign y5512 = ~n25742 ;
  assign y5513 = ~n25743 ;
  assign y5514 = n25748 ;
  assign y5515 = ~n25752 ;
  assign y5516 = n25753 ;
  assign y5517 = n25754 ;
  assign y5518 = n25758 ;
  assign y5519 = ~1'b0 ;
  assign y5520 = ~n25763 ;
  assign y5521 = n25767 ;
  assign y5522 = ~n25775 ;
  assign y5523 = n25776 ;
  assign y5524 = ~n25780 ;
  assign y5525 = ~n25790 ;
  assign y5526 = n25802 ;
  assign y5527 = ~n25806 ;
  assign y5528 = n25812 ;
  assign y5529 = n25816 ;
  assign y5530 = n25819 ;
  assign y5531 = n25822 ;
  assign y5532 = ~n25824 ;
  assign y5533 = ~n25825 ;
  assign y5534 = ~n25832 ;
  assign y5535 = n25834 ;
  assign y5536 = ~n25836 ;
  assign y5537 = ~n25838 ;
  assign y5538 = ~n25839 ;
  assign y5539 = ~n25849 ;
  assign y5540 = n25852 ;
  assign y5541 = n25853 ;
  assign y5542 = n25854 ;
  assign y5543 = ~n25857 ;
  assign y5544 = ~n25859 ;
  assign y5545 = n25863 ;
  assign y5546 = n25866 ;
  assign y5547 = ~n25869 ;
  assign y5548 = n25873 ;
  assign y5549 = n25874 ;
  assign y5550 = n25878 ;
  assign y5551 = ~n25881 ;
  assign y5552 = ~n25883 ;
  assign y5553 = n25885 ;
  assign y5554 = ~n25886 ;
  assign y5555 = n25890 ;
  assign y5556 = n25898 ;
  assign y5557 = n25904 ;
  assign y5558 = ~n25906 ;
  assign y5559 = n25911 ;
  assign y5560 = n25913 ;
  assign y5561 = ~n25914 ;
  assign y5562 = n25916 ;
  assign y5563 = ~n25920 ;
  assign y5564 = n25922 ;
  assign y5565 = n25923 ;
  assign y5566 = ~n25926 ;
  assign y5567 = ~n25927 ;
  assign y5568 = ~n25928 ;
  assign y5569 = ~1'b0 ;
  assign y5570 = n25930 ;
  assign y5571 = ~n25934 ;
  assign y5572 = ~n25945 ;
  assign y5573 = ~n25949 ;
  assign y5574 = n25956 ;
  assign y5575 = n25957 ;
  assign y5576 = ~n25960 ;
  assign y5577 = n25972 ;
  assign y5578 = ~n25974 ;
  assign y5579 = ~n25978 ;
  assign y5580 = n25979 ;
  assign y5581 = ~n25981 ;
  assign y5582 = ~n25982 ;
  assign y5583 = n25986 ;
  assign y5584 = n25992 ;
  assign y5585 = ~n25996 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = n25998 ;
  assign y5588 = ~n26007 ;
  assign y5589 = n26014 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = ~n26019 ;
  assign y5592 = ~n26024 ;
  assign y5593 = n26026 ;
  assign y5594 = ~n26036 ;
  assign y5595 = n26040 ;
  assign y5596 = ~n26045 ;
  assign y5597 = ~n26049 ;
  assign y5598 = ~n26060 ;
  assign y5599 = ~n26067 ;
  assign y5600 = n26070 ;
  assign y5601 = n26076 ;
  assign y5602 = n26079 ;
  assign y5603 = ~1'b0 ;
  assign y5604 = n26080 ;
  assign y5605 = n26083 ;
  assign y5606 = n26088 ;
  assign y5607 = n26091 ;
  assign y5608 = ~1'b0 ;
  assign y5609 = ~1'b0 ;
  assign y5610 = n26095 ;
  assign y5611 = ~n26098 ;
  assign y5612 = ~n26102 ;
  assign y5613 = ~1'b0 ;
  assign y5614 = ~n26104 ;
  assign y5615 = ~n26108 ;
  assign y5616 = n26109 ;
  assign y5617 = ~n26110 ;
  assign y5618 = n26115 ;
  assign y5619 = ~1'b0 ;
  assign y5620 = n26117 ;
  assign y5621 = n26119 ;
  assign y5622 = ~n26120 ;
  assign y5623 = n26126 ;
  assign y5624 = n26133 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = n26138 ;
  assign y5627 = n26139 ;
  assign y5628 = n26143 ;
  assign y5629 = n26144 ;
  assign y5630 = ~1'b0 ;
  assign y5631 = ~n26145 ;
  assign y5632 = ~n26150 ;
  assign y5633 = ~n26159 ;
  assign y5634 = n26161 ;
  assign y5635 = ~n26165 ;
  assign y5636 = ~n26170 ;
  assign y5637 = n26171 ;
  assign y5638 = ~1'b0 ;
  assign y5639 = ~n26172 ;
  assign y5640 = ~n26174 ;
  assign y5641 = n26175 ;
  assign y5642 = ~n26179 ;
  assign y5643 = ~n26181 ;
  assign y5644 = n26185 ;
  assign y5645 = n26188 ;
  assign y5646 = ~n26195 ;
  assign y5647 = n26196 ;
  assign y5648 = ~n26201 ;
  assign y5649 = n26211 ;
  assign y5650 = ~n26215 ;
  assign y5651 = ~n26219 ;
  assign y5652 = ~n26225 ;
  assign y5653 = n26228 ;
  assign y5654 = ~n26232 ;
  assign y5655 = ~n26233 ;
  assign y5656 = ~n26236 ;
  assign y5657 = n26240 ;
  assign y5658 = n26248 ;
  assign y5659 = n26253 ;
  assign y5660 = ~n26254 ;
  assign y5661 = ~n26258 ;
  assign y5662 = ~n26260 ;
  assign y5663 = n26261 ;
  assign y5664 = ~n26262 ;
  assign y5665 = n26268 ;
  assign y5666 = ~1'b0 ;
  assign y5667 = ~n26276 ;
  assign y5668 = n26277 ;
  assign y5669 = n26285 ;
  assign y5670 = ~n26288 ;
  assign y5671 = n26289 ;
  assign y5672 = ~n26292 ;
  assign y5673 = n26297 ;
  assign y5674 = ~n26301 ;
  assign y5675 = ~1'b0 ;
  assign y5676 = n26305 ;
  assign y5677 = ~1'b0 ;
  assign y5678 = ~n26309 ;
  assign y5679 = ~n26310 ;
  assign y5680 = ~1'b0 ;
  assign y5681 = ~n26314 ;
  assign y5682 = n26322 ;
  assign y5683 = n26325 ;
  assign y5684 = ~n26329 ;
  assign y5685 = ~n26331 ;
  assign y5686 = n26332 ;
  assign y5687 = ~n26334 ;
  assign y5688 = ~n26337 ;
  assign y5689 = ~n26342 ;
  assign y5690 = n26347 ;
  assign y5691 = ~n26348 ;
  assign y5692 = ~n26350 ;
  assign y5693 = n826 ;
  assign y5694 = n26355 ;
  assign y5695 = n26357 ;
  assign y5696 = n26363 ;
  assign y5697 = n26367 ;
  assign y5698 = ~n26369 ;
  assign y5699 = n26371 ;
  assign y5700 = n26375 ;
  assign y5701 = ~n26379 ;
  assign y5702 = n26382 ;
  assign y5703 = n26385 ;
  assign y5704 = ~n26387 ;
  assign y5705 = ~n26393 ;
  assign y5706 = ~1'b0 ;
  assign y5707 = ~n26398 ;
  assign y5708 = n26401 ;
  assign y5709 = n26405 ;
  assign y5710 = ~n26408 ;
  assign y5711 = n26412 ;
  assign y5712 = n26413 ;
  assign y5713 = ~n26415 ;
  assign y5714 = ~n26417 ;
  assign y5715 = ~n26418 ;
  assign y5716 = n26424 ;
  assign y5717 = n26427 ;
  assign y5718 = ~n26430 ;
  assign y5719 = ~n26431 ;
  assign y5720 = ~n26436 ;
  assign y5721 = n26438 ;
  assign y5722 = n26440 ;
  assign y5723 = ~n26443 ;
  assign y5724 = ~n26444 ;
  assign y5725 = n26446 ;
  assign y5726 = ~1'b0 ;
  assign y5727 = ~1'b0 ;
  assign y5728 = ~n26453 ;
  assign y5729 = ~n26454 ;
  assign y5730 = ~n26456 ;
  assign y5731 = ~1'b0 ;
  assign y5732 = n26458 ;
  assign y5733 = n26461 ;
  assign y5734 = n26463 ;
  assign y5735 = ~n26471 ;
  assign y5736 = ~n26481 ;
  assign y5737 = n26482 ;
  assign y5738 = n26486 ;
  assign y5739 = ~1'b0 ;
  assign y5740 = ~n26487 ;
  assign y5741 = n26488 ;
  assign y5742 = n26491 ;
  assign y5743 = n26493 ;
  assign y5744 = n17432 ;
  assign y5745 = ~n26495 ;
  assign y5746 = ~1'b0 ;
  assign y5747 = ~n26496 ;
  assign y5748 = n26497 ;
  assign y5749 = n26501 ;
  assign y5750 = n26502 ;
  assign y5751 = ~n26505 ;
  assign y5752 = n26506 ;
  assign y5753 = ~n26507 ;
  assign y5754 = ~n26515 ;
  assign y5755 = n26518 ;
  assign y5756 = ~n26523 ;
  assign y5757 = ~n26524 ;
  assign y5758 = n26530 ;
  assign y5759 = ~n26537 ;
  assign y5760 = n26538 ;
  assign y5761 = n26540 ;
  assign y5762 = n26543 ;
  assign y5763 = ~n26547 ;
  assign y5764 = ~n26550 ;
  assign y5765 = ~n26551 ;
  assign y5766 = ~n26553 ;
  assign y5767 = ~n26555 ;
  assign y5768 = n26558 ;
  assign y5769 = ~n26559 ;
  assign y5770 = ~1'b0 ;
  assign y5771 = ~n26560 ;
  assign y5772 = n26563 ;
  assign y5773 = ~n26565 ;
  assign y5774 = n26568 ;
  assign y5775 = ~n26572 ;
  assign y5776 = n26574 ;
  assign y5777 = n26580 ;
  assign y5778 = ~n26581 ;
  assign y5779 = ~n26582 ;
  assign y5780 = n26584 ;
  assign y5781 = n26585 ;
  assign y5782 = n26589 ;
  assign y5783 = ~n26592 ;
  assign y5784 = n26599 ;
  assign y5785 = ~n26601 ;
  assign y5786 = ~n26603 ;
  assign y5787 = ~n26605 ;
  assign y5788 = ~n26609 ;
  assign y5789 = ~n26614 ;
  assign y5790 = ~n26616 ;
  assign y5791 = n26621 ;
  assign y5792 = ~n26624 ;
  assign y5793 = n26629 ;
  assign y5794 = ~n26630 ;
  assign y5795 = ~n26635 ;
  assign y5796 = ~n26644 ;
  assign y5797 = ~1'b0 ;
  assign y5798 = n26650 ;
  assign y5799 = ~n26657 ;
  assign y5800 = n26660 ;
  assign y5801 = n26665 ;
  assign y5802 = n26666 ;
  assign y5803 = ~n26668 ;
  assign y5804 = n26675 ;
  assign y5805 = ~n26677 ;
  assign y5806 = n26679 ;
  assign y5807 = n26680 ;
  assign y5808 = ~1'b0 ;
  assign y5809 = n26692 ;
  assign y5810 = ~n26696 ;
  assign y5811 = n26704 ;
  assign y5812 = n26705 ;
  assign y5813 = ~n26706 ;
  assign y5814 = n26714 ;
  assign y5815 = ~n26726 ;
  assign y5816 = n26727 ;
  assign y5817 = n26728 ;
  assign y5818 = ~n26733 ;
  assign y5819 = n17498 ;
  assign y5820 = n26736 ;
  assign y5821 = ~n2662 ;
  assign y5822 = n26746 ;
  assign y5823 = n26747 ;
  assign y5824 = ~n26750 ;
  assign y5825 = ~n26753 ;
  assign y5826 = ~n26754 ;
  assign y5827 = n26756 ;
  assign y5828 = ~n26761 ;
  assign y5829 = n26767 ;
  assign y5830 = ~n26768 ;
  assign y5831 = ~1'b0 ;
  assign y5832 = ~n26769 ;
  assign y5833 = ~n26770 ;
  assign y5834 = n26771 ;
  assign y5835 = n26775 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = n26776 ;
  assign y5838 = ~n26780 ;
  assign y5839 = ~n26787 ;
  assign y5840 = ~n26788 ;
  assign y5841 = ~n26790 ;
  assign y5842 = n26792 ;
  assign y5843 = ~n26796 ;
  assign y5844 = ~1'b0 ;
  assign y5845 = ~n26797 ;
  assign y5846 = n26807 ;
  assign y5847 = ~n26809 ;
  assign y5848 = ~n26810 ;
  assign y5849 = n26816 ;
  assign y5850 = n26817 ;
  assign y5851 = ~n26819 ;
  assign y5852 = n26821 ;
  assign y5853 = ~n26822 ;
  assign y5854 = n26830 ;
  assign y5855 = ~n26834 ;
  assign y5856 = ~n26835 ;
  assign y5857 = ~n26837 ;
  assign y5858 = ~n26839 ;
  assign y5859 = ~n26841 ;
  assign y5860 = ~n26851 ;
  assign y5861 = ~n26854 ;
  assign y5862 = n26864 ;
  assign y5863 = n26866 ;
  assign y5864 = ~n26868 ;
  assign y5865 = ~n26871 ;
  assign y5866 = ~n26874 ;
  assign y5867 = ~n26875 ;
  assign y5868 = ~n26887 ;
  assign y5869 = ~n26892 ;
  assign y5870 = n26894 ;
  assign y5871 = ~n26902 ;
  assign y5872 = ~n26904 ;
  assign y5873 = ~n26905 ;
  assign y5874 = n26911 ;
  assign y5875 = ~n26914 ;
  assign y5876 = n26923 ;
  assign y5877 = n26933 ;
  assign y5878 = ~n26935 ;
  assign y5879 = n26937 ;
  assign y5880 = n26941 ;
  assign y5881 = n26949 ;
  assign y5882 = ~n26952 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~n26954 ;
  assign y5885 = ~n26962 ;
  assign y5886 = ~n26963 ;
  assign y5887 = n26966 ;
  assign y5888 = ~n20845 ;
  assign y5889 = ~n26969 ;
  assign y5890 = n26973 ;
  assign y5891 = n26981 ;
  assign y5892 = ~n26982 ;
  assign y5893 = ~n26984 ;
  assign y5894 = n26989 ;
  assign y5895 = n26990 ;
  assign y5896 = n26993 ;
  assign y5897 = ~n26996 ;
  assign y5898 = ~n26997 ;
  assign y5899 = ~n27004 ;
  assign y5900 = ~n27006 ;
  assign y5901 = n27008 ;
  assign y5902 = n27009 ;
  assign y5903 = ~n27015 ;
  assign y5904 = n27018 ;
  assign y5905 = n27021 ;
  assign y5906 = n27024 ;
  assign y5907 = n27029 ;
  assign y5908 = ~n27033 ;
  assign y5909 = ~n27038 ;
  assign y5910 = n27047 ;
  assign y5911 = n27048 ;
  assign y5912 = ~n27049 ;
  assign y5913 = n27052 ;
  assign y5914 = n27061 ;
  assign y5915 = n27064 ;
  assign y5916 = n27066 ;
  assign y5917 = ~1'b0 ;
  assign y5918 = ~1'b0 ;
  assign y5919 = n27067 ;
  assign y5920 = n27071 ;
  assign y5921 = n27073 ;
  assign y5922 = ~n27075 ;
  assign y5923 = ~n27076 ;
  assign y5924 = n27083 ;
  assign y5925 = n27094 ;
  assign y5926 = n27095 ;
  assign y5927 = n27096 ;
  assign y5928 = ~n27097 ;
  assign y5929 = ~n27098 ;
  assign y5930 = n27100 ;
  assign y5931 = n27104 ;
  assign y5932 = ~1'b0 ;
  assign y5933 = n27107 ;
  assign y5934 = n27108 ;
  assign y5935 = ~n27109 ;
  assign y5936 = n27113 ;
  assign y5937 = ~n27114 ;
  assign y5938 = ~n27121 ;
  assign y5939 = ~1'b0 ;
  assign y5940 = ~n27124 ;
  assign y5941 = ~n27131 ;
  assign y5942 = ~n27132 ;
  assign y5943 = n27138 ;
  assign y5944 = ~n27140 ;
  assign y5945 = ~n27143 ;
  assign y5946 = ~n27146 ;
  assign y5947 = ~n27148 ;
  assign y5948 = ~1'b0 ;
  assign y5949 = ~n27155 ;
  assign y5950 = ~n27164 ;
  assign y5951 = ~n27170 ;
  assign y5952 = n27171 ;
  assign y5953 = ~n27173 ;
  assign y5954 = n27174 ;
  assign y5955 = n27182 ;
  assign y5956 = ~n27183 ;
  assign y5957 = ~n27185 ;
  assign y5958 = ~n27194 ;
  assign y5959 = ~n27196 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = ~n27199 ;
  assign y5962 = ~n27210 ;
  assign y5963 = ~n27212 ;
  assign y5964 = n27217 ;
  assign y5965 = ~n27227 ;
  assign y5966 = ~1'b0 ;
  assign y5967 = ~n27235 ;
  assign y5968 = n27245 ;
  assign y5969 = n27249 ;
  assign y5970 = ~n27253 ;
  assign y5971 = n27254 ;
  assign y5972 = n27266 ;
  assign y5973 = n27270 ;
  assign y5974 = n27276 ;
  assign y5975 = ~n27278 ;
  assign y5976 = ~n27288 ;
  assign y5977 = n27290 ;
  assign y5978 = n27291 ;
  assign y5979 = ~n27301 ;
  assign y5980 = n27302 ;
  assign y5981 = ~n27304 ;
  assign y5982 = n27307 ;
  assign y5983 = ~n27309 ;
  assign y5984 = ~n27312 ;
  assign y5985 = n27314 ;
  assign y5986 = ~n27315 ;
  assign y5987 = ~n27316 ;
  assign y5988 = ~1'b0 ;
  assign y5989 = n27317 ;
  assign y5990 = ~n27321 ;
  assign y5991 = ~n27329 ;
  assign y5992 = ~n27332 ;
  assign y5993 = ~n27333 ;
  assign y5994 = ~n27334 ;
  assign y5995 = n27336 ;
  assign y5996 = ~n27339 ;
  assign y5997 = ~n27344 ;
  assign y5998 = n27348 ;
  assign y5999 = n27351 ;
  assign y6000 = ~1'b0 ;
  assign y6001 = ~n27356 ;
  assign y6002 = ~n27358 ;
  assign y6003 = n27361 ;
  assign y6004 = n4773 ;
  assign y6005 = n27362 ;
  assign y6006 = n27366 ;
  assign y6007 = n27379 ;
  assign y6008 = n27382 ;
  assign y6009 = n27390 ;
  assign y6010 = n27395 ;
  assign y6011 = ~n27396 ;
  assign y6012 = n27398 ;
  assign y6013 = ~n27399 ;
  assign y6014 = n27401 ;
  assign y6015 = n27405 ;
  assign y6016 = n27407 ;
  assign y6017 = ~n27412 ;
  assign y6018 = n27422 ;
  assign y6019 = n27425 ;
  assign y6020 = ~n27429 ;
  assign y6021 = ~n27441 ;
  assign y6022 = n27442 ;
  assign y6023 = ~n27445 ;
  assign y6024 = n27450 ;
  assign y6025 = n27452 ;
  assign y6026 = n27453 ;
  assign y6027 = ~n27454 ;
  assign y6028 = n27465 ;
  assign y6029 = ~n27466 ;
  assign y6030 = ~n27480 ;
  assign y6031 = n27483 ;
  assign y6032 = n27486 ;
  assign y6033 = ~n27488 ;
  assign y6034 = ~n27489 ;
  assign y6035 = ~n27496 ;
  assign y6036 = ~n27498 ;
  assign y6037 = ~n27499 ;
  assign y6038 = n27501 ;
  assign y6039 = ~n27505 ;
  assign y6040 = ~n27511 ;
  assign y6041 = n27515 ;
  assign y6042 = n27517 ;
  assign y6043 = ~n27525 ;
  assign y6044 = n27527 ;
  assign y6045 = n27529 ;
  assign y6046 = ~n27532 ;
  assign y6047 = ~n27537 ;
  assign y6048 = ~n27541 ;
  assign y6049 = n27546 ;
  assign y6050 = n27550 ;
  assign y6051 = ~n27558 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = ~n27559 ;
  assign y6054 = n27561 ;
  assign y6055 = ~n27565 ;
  assign y6056 = ~1'b0 ;
  assign y6057 = ~n27567 ;
  assign y6058 = n27576 ;
  assign y6059 = ~n27577 ;
  assign y6060 = n27584 ;
  assign y6061 = ~n27593 ;
  assign y6062 = ~n27594 ;
  assign y6063 = ~n27598 ;
  assign y6064 = ~n27605 ;
  assign y6065 = ~n27610 ;
  assign y6066 = ~1'b0 ;
  assign y6067 = ~n27615 ;
  assign y6068 = ~n27629 ;
  assign y6069 = n27630 ;
  assign y6070 = n27637 ;
  assign y6071 = n27642 ;
  assign y6072 = n27644 ;
  assign y6073 = n27645 ;
  assign y6074 = ~n27646 ;
  assign y6075 = ~n27652 ;
  assign y6076 = n27653 ;
  assign y6077 = n27658 ;
  assign y6078 = n27660 ;
  assign y6079 = ~n27661 ;
  assign y6080 = ~n27667 ;
  assign y6081 = ~n27668 ;
  assign y6082 = ~n27671 ;
  assign y6083 = n27672 ;
  assign y6084 = ~n27673 ;
  assign y6085 = n27676 ;
  assign y6086 = n27686 ;
  assign y6087 = ~n27691 ;
  assign y6088 = n27694 ;
  assign y6089 = n27699 ;
  assign y6090 = ~n27701 ;
  assign y6091 = n27704 ;
  assign y6092 = ~n27709 ;
  assign y6093 = ~n27715 ;
  assign y6094 = n27718 ;
  assign y6095 = ~n27721 ;
  assign y6096 = ~n27730 ;
  assign y6097 = n27732 ;
  assign y6098 = n27734 ;
  assign y6099 = n27735 ;
  assign y6100 = n27737 ;
  assign y6101 = n27741 ;
  assign y6102 = ~n27747 ;
  assign y6103 = ~n27760 ;
  assign y6104 = n27761 ;
  assign y6105 = n27764 ;
  assign y6106 = n27770 ;
  assign y6107 = ~n27775 ;
  assign y6108 = ~n27776 ;
  assign y6109 = ~n27779 ;
  assign y6110 = n27780 ;
  assign y6111 = n27784 ;
  assign y6112 = n27786 ;
  assign y6113 = n27799 ;
  assign y6114 = n27803 ;
  assign y6115 = n27806 ;
  assign y6116 = n27811 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = n27812 ;
  assign y6119 = ~n27813 ;
  assign y6120 = ~n27825 ;
  assign y6121 = n27829 ;
  assign y6122 = ~n27831 ;
  assign y6123 = n27840 ;
  assign y6124 = ~n27846 ;
  assign y6125 = n27847 ;
  assign y6126 = ~n27848 ;
  assign y6127 = ~n27850 ;
  assign y6128 = n27852 ;
  assign y6129 = n27853 ;
  assign y6130 = n27866 ;
  assign y6131 = n27868 ;
  assign y6132 = ~n27872 ;
  assign y6133 = n27873 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = n27874 ;
  assign y6136 = ~n27877 ;
  assign y6137 = n27880 ;
  assign y6138 = ~n27884 ;
  assign y6139 = ~n27887 ;
  assign y6140 = ~n27891 ;
  assign y6141 = ~1'b0 ;
  assign y6142 = ~n27895 ;
  assign y6143 = n27896 ;
  assign y6144 = n27897 ;
  assign y6145 = n27899 ;
  assign y6146 = ~n27902 ;
  assign y6147 = ~n27903 ;
  assign y6148 = ~n27906 ;
  assign y6149 = n27913 ;
  assign y6150 = ~n27915 ;
  assign y6151 = n27917 ;
  assign y6152 = n27920 ;
  assign y6153 = ~n27923 ;
  assign y6154 = n27926 ;
  assign y6155 = ~n27927 ;
  assign y6156 = n27930 ;
  assign y6157 = ~n27931 ;
  assign y6158 = ~n27939 ;
  assign y6159 = ~n27942 ;
  assign y6160 = ~n27944 ;
  assign y6161 = n27952 ;
  assign y6162 = n27959 ;
  assign y6163 = n27963 ;
  assign y6164 = ~n27965 ;
  assign y6165 = ~n27967 ;
  assign y6166 = n27969 ;
  assign y6167 = ~n27970 ;
  assign y6168 = n27972 ;
  assign y6169 = ~n27974 ;
  assign y6170 = ~n27975 ;
  assign y6171 = n27993 ;
  assign y6172 = n27994 ;
  assign y6173 = n27999 ;
  assign y6174 = n28001 ;
  assign y6175 = ~n28003 ;
  assign y6176 = n28005 ;
  assign y6177 = n28008 ;
  assign y6178 = ~n28010 ;
  assign y6179 = n28024 ;
  assign y6180 = n28027 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = n28029 ;
  assign y6183 = ~n28030 ;
  assign y6184 = ~n28032 ;
  assign y6185 = n28045 ;
  assign y6186 = n28046 ;
  assign y6187 = n28049 ;
  assign y6188 = n28052 ;
  assign y6189 = n28074 ;
  assign y6190 = ~1'b0 ;
  assign y6191 = n28075 ;
  assign y6192 = n28080 ;
  assign y6193 = ~1'b0 ;
  assign y6194 = n28086 ;
  assign y6195 = n28089 ;
  assign y6196 = ~n28093 ;
  assign y6197 = ~n28095 ;
  assign y6198 = n28096 ;
  assign y6199 = n28100 ;
  assign y6200 = n28102 ;
  assign y6201 = n28104 ;
  assign y6202 = ~n28109 ;
  assign y6203 = n28111 ;
  assign y6204 = ~n28115 ;
  assign y6205 = n28118 ;
  assign y6206 = n28121 ;
  assign y6207 = n28127 ;
  assign y6208 = ~n28129 ;
  assign y6209 = n28137 ;
  assign y6210 = ~n28141 ;
  assign y6211 = ~n28145 ;
  assign y6212 = ~n28153 ;
  assign y6213 = n28156 ;
  assign y6214 = n28157 ;
  assign y6215 = n28159 ;
  assign y6216 = ~n28160 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = ~1'b0 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = ~n28163 ;
  assign y6221 = ~n28167 ;
  assign y6222 = ~n28168 ;
  assign y6223 = ~n28169 ;
  assign y6224 = ~n28172 ;
  assign y6225 = n28182 ;
  assign y6226 = ~n28187 ;
  assign y6227 = n28190 ;
  assign y6228 = ~n28201 ;
  assign y6229 = ~n28204 ;
  assign y6230 = n28214 ;
  assign y6231 = n28216 ;
  assign y6232 = ~n28217 ;
  assign y6233 = n28218 ;
  assign y6234 = n28221 ;
  assign y6235 = n28225 ;
  assign y6236 = ~n28235 ;
  assign y6237 = n28245 ;
  assign y6238 = n28246 ;
  assign y6239 = ~n28251 ;
  assign y6240 = n28252 ;
  assign y6241 = n28257 ;
  assign y6242 = ~n28258 ;
  assign y6243 = ~n28264 ;
  assign y6244 = n28267 ;
  assign y6245 = ~1'b0 ;
  assign y6246 = n28273 ;
  assign y6247 = ~n28275 ;
  assign y6248 = n28279 ;
  assign y6249 = ~n28281 ;
  assign y6250 = ~n28282 ;
  assign y6251 = ~n28287 ;
  assign y6252 = ~n28289 ;
  assign y6253 = ~n28294 ;
  assign y6254 = n28297 ;
  assign y6255 = ~n28298 ;
  assign y6256 = n28301 ;
  assign y6257 = ~n28302 ;
  assign y6258 = n28307 ;
  assign y6259 = ~1'b0 ;
  assign y6260 = ~n28309 ;
  assign y6261 = ~n28311 ;
  assign y6262 = ~1'b0 ;
  assign y6263 = n28314 ;
  assign y6264 = n28317 ;
  assign y6265 = ~n28319 ;
  assign y6266 = n28323 ;
  assign y6267 = n28330 ;
  assign y6268 = n28332 ;
  assign y6269 = n28338 ;
  assign y6270 = ~n28348 ;
  assign y6271 = n28370 ;
  assign y6272 = ~n28373 ;
  assign y6273 = ~n28375 ;
  assign y6274 = n13071 ;
  assign y6275 = n28378 ;
  assign y6276 = ~1'b0 ;
  assign y6277 = n28381 ;
  assign y6278 = ~n28387 ;
  assign y6279 = n28389 ;
  assign y6280 = n28390 ;
  assign y6281 = ~n28393 ;
  assign y6282 = ~n28395 ;
  assign y6283 = n28396 ;
  assign y6284 = n28400 ;
  assign y6285 = ~n28407 ;
  assign y6286 = ~1'b0 ;
  assign y6287 = ~n28413 ;
  assign y6288 = n28416 ;
  assign y6289 = n28419 ;
  assign y6290 = n28420 ;
  assign y6291 = ~n28423 ;
  assign y6292 = ~n28434 ;
  assign y6293 = n28437 ;
  assign y6294 = ~n28444 ;
  assign y6295 = ~n28446 ;
  assign y6296 = n28447 ;
  assign y6297 = n28449 ;
  assign y6298 = n28450 ;
  assign y6299 = ~n28451 ;
  assign y6300 = ~n28452 ;
  assign y6301 = n28453 ;
  assign y6302 = n28458 ;
  assign y6303 = n28461 ;
  assign y6304 = n28463 ;
  assign y6305 = n28464 ;
  assign y6306 = n28466 ;
  assign y6307 = ~n28467 ;
  assign y6308 = ~n28469 ;
  assign y6309 = ~1'b0 ;
  assign y6310 = ~n28482 ;
  assign y6311 = n28483 ;
  assign y6312 = ~n28485 ;
  assign y6313 = ~1'b0 ;
  assign y6314 = ~n28491 ;
  assign y6315 = ~n28495 ;
  assign y6316 = n28499 ;
  assign y6317 = ~n28501 ;
  assign y6318 = ~n28510 ;
  assign y6319 = ~n28512 ;
  assign y6320 = ~n28514 ;
  assign y6321 = n28515 ;
  assign y6322 = n28519 ;
  assign y6323 = ~1'b0 ;
  assign y6324 = ~n28526 ;
  assign y6325 = n28529 ;
  assign y6326 = ~n28535 ;
  assign y6327 = n28539 ;
  assign y6328 = n15659 ;
  assign y6329 = ~n28543 ;
  assign y6330 = ~1'b0 ;
  assign y6331 = n28545 ;
  assign y6332 = ~n28550 ;
  assign y6333 = ~n28555 ;
  assign y6334 = n28559 ;
  assign y6335 = ~1'b0 ;
  assign y6336 = ~n28560 ;
  assign y6337 = ~n28563 ;
  assign y6338 = ~n28570 ;
  assign y6339 = n28571 ;
  assign y6340 = ~n28579 ;
  assign y6341 = ~n28590 ;
  assign y6342 = n28600 ;
  assign y6343 = ~1'b0 ;
  assign y6344 = n28605 ;
  assign y6345 = ~n28607 ;
  assign y6346 = ~n28609 ;
  assign y6347 = n28610 ;
  assign y6348 = n28612 ;
  assign y6349 = n28613 ;
  assign y6350 = n28614 ;
  assign y6351 = n28618 ;
  assign y6352 = ~n28619 ;
  assign y6353 = ~n28620 ;
  assign y6354 = n28623 ;
  assign y6355 = ~n28626 ;
  assign y6356 = n28628 ;
  assign y6357 = ~n28633 ;
  assign y6358 = n28639 ;
  assign y6359 = n28640 ;
  assign y6360 = n28644 ;
  assign y6361 = n28646 ;
  assign y6362 = n28657 ;
  assign y6363 = ~n28671 ;
  assign y6364 = n28674 ;
  assign y6365 = n28676 ;
  assign y6366 = ~n28678 ;
  assign y6367 = n28684 ;
  assign y6368 = ~n28686 ;
  assign y6369 = n28690 ;
  assign y6370 = ~n28691 ;
  assign y6371 = ~n28695 ;
  assign y6372 = n28696 ;
  assign y6373 = ~n28698 ;
  assign y6374 = ~1'b0 ;
  assign y6375 = n28701 ;
  assign y6376 = ~n28704 ;
  assign y6377 = n28708 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = ~n28710 ;
  assign y6380 = ~n28711 ;
  assign y6381 = n28713 ;
  assign y6382 = n28715 ;
  assign y6383 = n28718 ;
  assign y6384 = ~n28723 ;
  assign y6385 = ~n28725 ;
  assign y6386 = n28732 ;
  assign y6387 = ~n28738 ;
  assign y6388 = n28740 ;
  assign y6389 = ~n28741 ;
  assign y6390 = n28745 ;
  assign y6391 = ~n28747 ;
  assign y6392 = n28749 ;
  assign y6393 = ~n28750 ;
  assign y6394 = ~n28753 ;
  assign y6395 = n28758 ;
  assign y6396 = ~1'b0 ;
  assign y6397 = n12789 ;
  assign y6398 = n28759 ;
  assign y6399 = n28765 ;
  assign y6400 = ~n28767 ;
  assign y6401 = n28773 ;
  assign y6402 = ~n28774 ;
  assign y6403 = ~n28778 ;
  assign y6404 = ~1'b0 ;
  assign y6405 = ~n28783 ;
  assign y6406 = n28786 ;
  assign y6407 = n28787 ;
  assign y6408 = ~n28793 ;
  assign y6409 = n28795 ;
  assign y6410 = ~n28796 ;
  assign y6411 = n28801 ;
  assign y6412 = ~n28802 ;
  assign y6413 = ~n28803 ;
  assign y6414 = ~n28809 ;
  assign y6415 = ~n28811 ;
  assign y6416 = n28813 ;
  assign y6417 = n28815 ;
  assign y6418 = n28816 ;
  assign y6419 = n28817 ;
  assign y6420 = ~n28819 ;
  assign y6421 = ~n28821 ;
  assign y6422 = n28822 ;
  assign y6423 = n28824 ;
  assign y6424 = ~n28826 ;
  assign y6425 = ~n28834 ;
  assign y6426 = ~n28837 ;
  assign y6427 = ~n28838 ;
  assign y6428 = ~1'b0 ;
  assign y6429 = n28842 ;
  assign y6430 = n28846 ;
  assign y6431 = ~n28851 ;
  assign y6432 = n28859 ;
  assign y6433 = ~n28862 ;
  assign y6434 = n28867 ;
  assign y6435 = ~1'b0 ;
  assign y6436 = ~n28875 ;
  assign y6437 = n28882 ;
  assign y6438 = n28886 ;
  assign y6439 = ~n28887 ;
  assign y6440 = ~n28889 ;
  assign y6441 = ~n28894 ;
  assign y6442 = n28897 ;
  assign y6443 = ~1'b0 ;
  assign y6444 = ~n28901 ;
  assign y6445 = ~n28904 ;
  assign y6446 = n28907 ;
  assign y6447 = ~n28909 ;
  assign y6448 = ~n28919 ;
  assign y6449 = n28924 ;
  assign y6450 = n28925 ;
  assign y6451 = ~n28926 ;
  assign y6452 = ~n28927 ;
  assign y6453 = n28928 ;
  assign y6454 = ~n28933 ;
  assign y6455 = ~n28936 ;
  assign y6456 = ~n28937 ;
  assign y6457 = ~n28940 ;
  assign y6458 = ~1'b0 ;
  assign y6459 = n28941 ;
  assign y6460 = n28947 ;
  assign y6461 = n28950 ;
  assign y6462 = n28954 ;
  assign y6463 = n28957 ;
  assign y6464 = ~n28965 ;
  assign y6465 = ~n28966 ;
  assign y6466 = ~n28971 ;
  assign y6467 = n28972 ;
  assign y6468 = ~n28977 ;
  assign y6469 = n28979 ;
  assign y6470 = n28986 ;
  assign y6471 = ~n28988 ;
  assign y6472 = ~n28995 ;
  assign y6473 = n29000 ;
  assign y6474 = n29003 ;
  assign y6475 = n29009 ;
  assign y6476 = ~n29013 ;
  assign y6477 = ~n29015 ;
  assign y6478 = n29017 ;
  assign y6479 = n29018 ;
  assign y6480 = n29019 ;
  assign y6481 = ~n29021 ;
  assign y6482 = ~n29026 ;
  assign y6483 = ~n29029 ;
  assign y6484 = n29034 ;
  assign y6485 = ~n29037 ;
  assign y6486 = ~n29039 ;
  assign y6487 = ~n29041 ;
  assign y6488 = ~n29043 ;
  assign y6489 = ~n29047 ;
  assign y6490 = ~n29053 ;
  assign y6491 = ~1'b0 ;
  assign y6492 = ~n29056 ;
  assign y6493 = n29061 ;
  assign y6494 = ~n29074 ;
  assign y6495 = ~n29076 ;
  assign y6496 = ~n29081 ;
  assign y6497 = n29086 ;
  assign y6498 = ~n29091 ;
  assign y6499 = ~n29092 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~1'b0 ;
  assign y6502 = ~n29095 ;
  assign y6503 = n29096 ;
  assign y6504 = n29098 ;
  assign y6505 = n29109 ;
  assign y6506 = n29112 ;
  assign y6507 = n29113 ;
  assign y6508 = n29120 ;
  assign y6509 = n29124 ;
  assign y6510 = ~n29131 ;
  assign y6511 = n29134 ;
  assign y6512 = ~n29139 ;
  assign y6513 = ~1'b0 ;
  assign y6514 = ~n29145 ;
  assign y6515 = n29149 ;
  assign y6516 = ~n29159 ;
  assign y6517 = n29161 ;
  assign y6518 = ~1'b0 ;
  assign y6519 = n29163 ;
  assign y6520 = ~n29164 ;
  assign y6521 = n29165 ;
  assign y6522 = ~n29169 ;
  assign y6523 = n29171 ;
  assign y6524 = ~n29173 ;
  assign y6525 = n29176 ;
  assign y6526 = ~n29179 ;
  assign y6527 = ~n29182 ;
  assign y6528 = ~n29184 ;
  assign y6529 = ~n29185 ;
  assign y6530 = n29186 ;
  assign y6531 = n29187 ;
  assign y6532 = n29188 ;
  assign y6533 = ~n29192 ;
  assign y6534 = ~n29194 ;
  assign y6535 = n29196 ;
  assign y6536 = ~n29199 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = n29201 ;
  assign y6540 = n29207 ;
  assign y6541 = n29211 ;
  assign y6542 = ~n29212 ;
  assign y6543 = ~n29215 ;
  assign y6544 = ~n29217 ;
  assign y6545 = ~n29219 ;
  assign y6546 = n29220 ;
  assign y6547 = n29221 ;
  assign y6548 = n29223 ;
  assign y6549 = ~n29226 ;
  assign y6550 = n29227 ;
  assign y6551 = n29229 ;
  assign y6552 = n29232 ;
  assign y6553 = ~n29236 ;
  assign y6554 = n29241 ;
  assign y6555 = n29249 ;
  assign y6556 = n29252 ;
  assign y6557 = n29262 ;
  assign y6558 = ~n29263 ;
  assign y6559 = ~n29265 ;
  assign y6560 = ~1'b0 ;
  assign y6561 = n29266 ;
  assign y6562 = ~n29271 ;
  assign y6563 = ~n29287 ;
  assign y6564 = ~n29298 ;
  assign y6565 = ~n29304 ;
  assign y6566 = ~1'b0 ;
  assign y6567 = ~1'b0 ;
  assign y6568 = n29317 ;
  assign y6569 = n29323 ;
  assign y6570 = ~n29325 ;
  assign y6571 = ~n29330 ;
  assign y6572 = ~1'b0 ;
  assign y6573 = ~1'b0 ;
  assign y6574 = n29335 ;
  assign y6575 = ~n29338 ;
  assign y6576 = ~n29342 ;
  assign y6577 = ~n29346 ;
  assign y6578 = ~1'b0 ;
  assign y6579 = n29350 ;
  assign y6580 = ~n29356 ;
  assign y6581 = ~n29358 ;
  assign y6582 = n29359 ;
  assign y6583 = ~n29362 ;
  assign y6584 = ~n29368 ;
  assign y6585 = n29375 ;
  assign y6586 = ~n29376 ;
  assign y6587 = ~n29378 ;
  assign y6588 = ~n29380 ;
  assign y6589 = ~n29384 ;
  assign y6590 = ~n29385 ;
  assign y6591 = ~n29386 ;
  assign y6592 = n29389 ;
  assign y6593 = n29391 ;
  assign y6594 = ~n29393 ;
  assign y6595 = ~n29394 ;
  assign y6596 = n29395 ;
  assign y6597 = n29406 ;
  assign y6598 = ~n29418 ;
  assign y6599 = ~n29422 ;
  assign y6600 = n29424 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = ~n29425 ;
  assign y6603 = n29430 ;
  assign y6604 = ~n29431 ;
  assign y6605 = ~n29434 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = n29440 ;
  assign y6608 = n29442 ;
  assign y6609 = n29447 ;
  assign y6610 = n29448 ;
  assign y6611 = n29451 ;
  assign y6612 = n29453 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = n29458 ;
  assign y6615 = ~n29462 ;
  assign y6616 = ~n29465 ;
  assign y6617 = n29470 ;
  assign y6618 = ~n29475 ;
  assign y6619 = ~n29477 ;
  assign y6620 = n29484 ;
  assign y6621 = n29486 ;
  assign y6622 = ~n29497 ;
  assign y6623 = ~n29503 ;
  assign y6624 = ~n29507 ;
  assign y6625 = ~n29508 ;
  assign y6626 = ~n29511 ;
  assign y6627 = n29512 ;
  assign y6628 = n29515 ;
  assign y6629 = n29523 ;
  assign y6630 = n29524 ;
  assign y6631 = n29526 ;
  assign y6632 = ~n29527 ;
  assign y6633 = n29528 ;
  assign y6634 = ~n29530 ;
  assign y6635 = n29533 ;
  assign y6636 = ~1'b0 ;
  assign y6637 = ~1'b0 ;
  assign y6638 = n29538 ;
  assign y6639 = n29539 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = ~n29541 ;
  assign y6642 = ~n29544 ;
  assign y6643 = n29546 ;
  assign y6644 = n29550 ;
  assign y6645 = n29552 ;
  assign y6646 = n29562 ;
  assign y6647 = ~n29564 ;
  assign y6648 = n29567 ;
  assign y6649 = ~n29568 ;
  assign y6650 = n29571 ;
  assign y6651 = ~n29576 ;
  assign y6652 = n29591 ;
  assign y6653 = n29595 ;
  assign y6654 = ~n29600 ;
  assign y6655 = ~n29601 ;
  assign y6656 = n29605 ;
  assign y6657 = ~n29611 ;
  assign y6658 = n29615 ;
  assign y6659 = n29617 ;
  assign y6660 = ~1'b0 ;
  assign y6661 = ~1'b0 ;
  assign y6662 = n29620 ;
  assign y6663 = n29621 ;
  assign y6664 = n29625 ;
  assign y6665 = n29632 ;
  assign y6666 = n29633 ;
  assign y6667 = n29634 ;
  assign y6668 = ~1'b0 ;
  assign y6669 = ~1'b0 ;
  assign y6670 = ~n29636 ;
  assign y6671 = ~n29640 ;
  assign y6672 = ~n29644 ;
  assign y6673 = n29645 ;
  assign y6674 = n29647 ;
  assign y6675 = n29652 ;
  assign y6676 = n29653 ;
  assign y6677 = ~n29654 ;
  assign y6678 = n29656 ;
  assign y6679 = ~n29659 ;
  assign y6680 = n29660 ;
  assign y6681 = ~1'b0 ;
  assign y6682 = n29662 ;
  assign y6683 = ~n29665 ;
  assign y6684 = ~n29667 ;
  assign y6685 = ~n29672 ;
  assign y6686 = n29678 ;
  assign y6687 = ~n29679 ;
  assign y6688 = ~n29680 ;
  assign y6689 = n29686 ;
  assign y6690 = n29689 ;
  assign y6691 = n29697 ;
  assign y6692 = ~n29701 ;
  assign y6693 = ~n29704 ;
  assign y6694 = n29709 ;
  assign y6695 = ~n29710 ;
  assign y6696 = ~n29711 ;
  assign y6697 = n29718 ;
  assign y6698 = ~1'b0 ;
  assign y6699 = n29722 ;
  assign y6700 = ~n29723 ;
  assign y6701 = n29725 ;
  assign y6702 = n29727 ;
  assign y6703 = ~n29730 ;
  assign y6704 = ~n29737 ;
  assign y6705 = ~n29739 ;
  assign y6706 = n29744 ;
  assign y6707 = ~n29747 ;
  assign y6708 = n29748 ;
  assign y6709 = n29750 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = n29753 ;
  assign y6712 = n29755 ;
  assign y6713 = ~n23965 ;
  assign y6714 = ~n29760 ;
  assign y6715 = n29761 ;
  assign y6716 = ~n29762 ;
  assign y6717 = n29765 ;
  assign y6718 = ~n29771 ;
  assign y6719 = n29775 ;
  assign y6720 = n29782 ;
  assign y6721 = ~n29783 ;
  assign y6722 = n29784 ;
  assign y6723 = n29788 ;
  assign y6724 = ~n29793 ;
  assign y6725 = n29794 ;
  assign y6726 = n29795 ;
  assign y6727 = ~n29800 ;
  assign y6728 = ~n29802 ;
  assign y6729 = n29805 ;
  assign y6730 = ~n29808 ;
  assign y6731 = n29819 ;
  assign y6732 = n29822 ;
  assign y6733 = n29826 ;
  assign y6734 = ~n29834 ;
  assign y6735 = ~n29836 ;
  assign y6736 = n29845 ;
  assign y6737 = ~n29850 ;
  assign y6738 = n29851 ;
  assign y6739 = n29857 ;
  assign y6740 = n29861 ;
  assign y6741 = n29866 ;
  assign y6742 = ~n29872 ;
  assign y6743 = ~1'b0 ;
  assign y6744 = ~n29874 ;
  assign y6745 = ~n29876 ;
  assign y6746 = n29883 ;
  assign y6747 = ~n29885 ;
  assign y6748 = n29897 ;
  assign y6749 = n29899 ;
  assign y6750 = n29903 ;
  assign y6751 = ~n29906 ;
  assign y6752 = ~n29911 ;
  assign y6753 = ~n29913 ;
  assign y6754 = ~n29917 ;
  assign y6755 = ~n29920 ;
  assign y6756 = ~n29921 ;
  assign y6757 = n29932 ;
  assign y6758 = n29941 ;
  assign y6759 = ~n29943 ;
  assign y6760 = n29944 ;
  assign y6761 = ~n29950 ;
  assign y6762 = ~n29955 ;
  assign y6763 = n29960 ;
  assign y6764 = ~n29961 ;
  assign y6765 = n29965 ;
  assign y6766 = ~n29966 ;
  assign y6767 = n29968 ;
  assign y6768 = ~n29969 ;
  assign y6769 = ~n29973 ;
  assign y6770 = ~n29978 ;
  assign y6771 = n29981 ;
  assign y6772 = n29983 ;
  assign y6773 = ~n29986 ;
  assign y6774 = n29991 ;
  assign y6775 = ~n29998 ;
  assign y6776 = n30003 ;
  assign y6777 = ~n30009 ;
  assign y6778 = n30010 ;
  assign y6779 = ~1'b0 ;
  assign y6780 = ~n30011 ;
  assign y6781 = ~n30013 ;
  assign y6782 = n30019 ;
  assign y6783 = n30022 ;
  assign y6784 = ~n30023 ;
  assign y6785 = n30028 ;
  assign y6786 = n30032 ;
  assign y6787 = n30037 ;
  assign y6788 = ~1'b0 ;
  assign y6789 = ~n30042 ;
  assign y6790 = n30044 ;
  assign y6791 = n30047 ;
  assign y6792 = n30051 ;
  assign y6793 = n30054 ;
  assign y6794 = ~n30061 ;
  assign y6795 = n30066 ;
  assign y6796 = n30067 ;
  assign y6797 = n30069 ;
  assign y6798 = n30072 ;
  assign y6799 = ~n30074 ;
  assign y6800 = ~1'b0 ;
  assign y6801 = n30075 ;
  assign y6802 = n30076 ;
  assign y6803 = n30082 ;
  assign y6804 = ~n30084 ;
  assign y6805 = n30089 ;
  assign y6806 = ~n30092 ;
  assign y6807 = n30096 ;
  assign y6808 = ~n30098 ;
  assign y6809 = ~n30100 ;
  assign y6810 = n30101 ;
  assign y6811 = n30103 ;
  assign y6812 = n30104 ;
  assign y6813 = n30106 ;
  assign y6814 = ~n30112 ;
  assign y6815 = n30123 ;
  assign y6816 = n30126 ;
  assign y6817 = ~n30127 ;
  assign y6818 = ~n30130 ;
  assign y6819 = ~n30132 ;
  assign y6820 = n30134 ;
  assign y6821 = n30136 ;
  assign y6822 = n30137 ;
  assign y6823 = n30138 ;
  assign y6824 = n30146 ;
  assign y6825 = ~n30147 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = n30149 ;
  assign y6828 = n30151 ;
  assign y6829 = ~n30153 ;
  assign y6830 = ~1'b0 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = n30154 ;
  assign y6833 = ~n30156 ;
  assign y6834 = ~n30159 ;
  assign y6835 = n30160 ;
  assign y6836 = ~n30166 ;
  assign y6837 = n30168 ;
  assign y6838 = ~1'b0 ;
  assign y6839 = ~n30174 ;
  assign y6840 = ~n30176 ;
  assign y6841 = ~1'b0 ;
  assign y6842 = ~1'b0 ;
  assign y6843 = ~n30179 ;
  assign y6844 = n30181 ;
  assign y6845 = ~n30184 ;
  assign y6846 = n30188 ;
  assign y6847 = n30189 ;
  assign y6848 = n30193 ;
  assign y6849 = ~n30199 ;
  assign y6850 = ~n30204 ;
  assign y6851 = ~n30206 ;
  assign y6852 = n30208 ;
  assign y6853 = n30212 ;
  assign y6854 = n30219 ;
  assign y6855 = ~n30225 ;
  assign y6856 = ~1'b0 ;
  assign y6857 = n30228 ;
  assign y6858 = ~n30231 ;
  assign y6859 = ~n30233 ;
  assign y6860 = ~n30234 ;
  assign y6861 = n30241 ;
  assign y6862 = ~n30242 ;
  assign y6863 = n30244 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = n30245 ;
  assign y6866 = n30246 ;
  assign y6867 = ~n30249 ;
  assign y6868 = n30251 ;
  assign y6869 = ~n30253 ;
  assign y6870 = n30257 ;
  assign y6871 = ~n30259 ;
  assign y6872 = ~n30264 ;
  assign y6873 = ~n30266 ;
  assign y6874 = ~n30269 ;
  assign y6875 = ~n30270 ;
  assign y6876 = ~n30271 ;
  assign y6877 = ~n30272 ;
  assign y6878 = ~n30273 ;
  assign y6879 = ~1'b0 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = n30275 ;
  assign y6882 = n30281 ;
  assign y6883 = ~n30282 ;
  assign y6884 = ~n30283 ;
  assign y6885 = n30287 ;
  assign y6886 = n30289 ;
  assign y6887 = n30291 ;
  assign y6888 = ~n30295 ;
  assign y6889 = ~n30297 ;
  assign y6890 = n30301 ;
  assign y6891 = ~n30304 ;
  assign y6892 = n30306 ;
  assign y6893 = n30307 ;
  assign y6894 = n30309 ;
  assign y6895 = ~n30313 ;
  assign y6896 = ~n30317 ;
  assign y6897 = ~n30319 ;
  assign y6898 = ~n30320 ;
  assign y6899 = n30327 ;
  assign y6900 = ~n30328 ;
  assign y6901 = ~n30330 ;
  assign y6902 = ~n30336 ;
  assign y6903 = ~n30343 ;
  assign y6904 = ~n30344 ;
  assign y6905 = ~n30347 ;
  assign y6906 = ~1'b0 ;
  assign y6907 = ~n30349 ;
  assign y6908 = ~n30357 ;
  assign y6909 = ~n30360 ;
  assign y6910 = n30363 ;
  assign y6911 = n30365 ;
  assign y6912 = ~n30367 ;
  assign y6913 = ~n30374 ;
  assign y6914 = n30375 ;
  assign y6915 = ~n30382 ;
  assign y6916 = ~1'b0 ;
  assign y6917 = ~n30389 ;
  assign y6918 = ~n30395 ;
  assign y6919 = n30396 ;
  assign y6920 = ~n30397 ;
  assign y6921 = ~n30399 ;
  assign y6922 = ~n30404 ;
  assign y6923 = n30406 ;
  assign y6924 = ~1'b0 ;
  assign y6925 = ~n30413 ;
  assign y6926 = n30416 ;
  assign y6927 = n30420 ;
  assign y6928 = ~n30427 ;
  assign y6929 = ~n30430 ;
  assign y6930 = ~1'b0 ;
  assign y6931 = ~1'b0 ;
  assign y6932 = ~n30439 ;
  assign y6933 = ~n30440 ;
  assign y6934 = ~n30447 ;
  assign y6935 = n30448 ;
  assign y6936 = n30452 ;
  assign y6937 = n30456 ;
  assign y6938 = ~n30458 ;
  assign y6939 = ~n30461 ;
  assign y6940 = n30466 ;
  assign y6941 = n30470 ;
  assign y6942 = ~n30475 ;
  assign y6943 = ~n30479 ;
  assign y6944 = ~n30480 ;
  assign y6945 = ~1'b0 ;
  assign y6946 = n30481 ;
  assign y6947 = n30484 ;
  assign y6948 = n30488 ;
  assign y6949 = ~n30489 ;
  assign y6950 = ~n30494 ;
  assign y6951 = n30497 ;
  assign y6952 = ~n30502 ;
  assign y6953 = ~n30504 ;
  assign y6954 = ~n30506 ;
  assign y6955 = n30509 ;
  assign y6956 = ~n30512 ;
  assign y6957 = n30514 ;
  assign y6958 = ~1'b0 ;
  assign y6959 = ~n30516 ;
  assign y6960 = n30518 ;
  assign y6961 = n30520 ;
  assign y6962 = n30527 ;
  assign y6963 = n30529 ;
  assign y6964 = ~n30530 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = ~n30532 ;
  assign y6967 = n30535 ;
  assign y6968 = ~n30537 ;
  assign y6969 = ~n30538 ;
  assign y6970 = ~n30540 ;
  assign y6971 = ~n30542 ;
  assign y6972 = n30543 ;
  assign y6973 = ~1'b0 ;
  assign y6974 = ~n30545 ;
  assign y6975 = n30549 ;
  assign y6976 = n30551 ;
  assign y6977 = n30553 ;
  assign y6978 = ~n30555 ;
  assign y6979 = n30558 ;
  assign y6980 = ~n30560 ;
  assign y6981 = n30566 ;
  assign y6982 = n30570 ;
  assign y6983 = n30572 ;
  assign y6984 = ~n30576 ;
  assign y6985 = n30579 ;
  assign y6986 = n30580 ;
  assign y6987 = ~n30581 ;
  assign y6988 = n30583 ;
  assign y6989 = ~n30585 ;
  assign y6990 = n30590 ;
  assign y6991 = n30592 ;
  assign y6992 = ~n30598 ;
  assign y6993 = n30600 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = ~n30603 ;
  assign y6996 = n30605 ;
  assign y6997 = n30610 ;
  assign y6998 = ~n30611 ;
  assign y6999 = ~n30614 ;
  assign y7000 = n30620 ;
  assign y7001 = ~n30633 ;
  assign y7002 = ~n30635 ;
  assign y7003 = ~n30636 ;
  assign y7004 = n30641 ;
  assign y7005 = ~n30646 ;
  assign y7006 = ~1'b0 ;
  assign y7007 = n30647 ;
  assign y7008 = ~n30653 ;
  assign y7009 = n30656 ;
  assign y7010 = n30657 ;
  assign y7011 = n30661 ;
  assign y7012 = ~1'b0 ;
  assign y7013 = ~n30663 ;
  assign y7014 = ~n30666 ;
  assign y7015 = ~n30668 ;
  assign y7016 = n30671 ;
  assign y7017 = ~n30675 ;
  assign y7018 = ~n30679 ;
  assign y7019 = ~1'b0 ;
  assign y7020 = n30682 ;
  assign y7021 = ~n30683 ;
  assign y7022 = n30688 ;
  assign y7023 = n30695 ;
  assign y7024 = n30701 ;
  assign y7025 = n30702 ;
  assign y7026 = ~n30706 ;
  assign y7027 = ~n30709 ;
  assign y7028 = n30710 ;
  assign y7029 = n30711 ;
  assign y7030 = ~n30713 ;
  assign y7031 = ~n30715 ;
  assign y7032 = n30716 ;
  assign y7033 = n30719 ;
  assign y7034 = ~n30723 ;
  assign y7035 = ~n30726 ;
  assign y7036 = ~n30743 ;
  assign y7037 = ~1'b0 ;
  assign y7038 = ~n30749 ;
  assign y7039 = ~n30751 ;
  assign y7040 = n30754 ;
  assign y7041 = n30756 ;
  assign y7042 = ~n30759 ;
  assign y7043 = n30760 ;
  assign y7044 = n30762 ;
  assign y7045 = ~n30763 ;
  assign y7046 = ~n30766 ;
  assign y7047 = ~n30767 ;
  assign y7048 = ~n30768 ;
  assign y7049 = n30769 ;
  assign y7050 = n30771 ;
  assign y7051 = ~n30773 ;
  assign y7052 = ~n30778 ;
  assign y7053 = ~n30780 ;
  assign y7054 = n30784 ;
  assign y7055 = n30786 ;
  assign y7056 = n30787 ;
  assign y7057 = n30788 ;
  assign y7058 = ~n30790 ;
  assign y7059 = n30791 ;
  assign y7060 = ~n30795 ;
  assign y7061 = ~1'b0 ;
  assign y7062 = ~n30798 ;
  assign y7063 = ~n30800 ;
  assign y7064 = n30803 ;
  assign y7065 = n30804 ;
  assign y7066 = n30805 ;
  assign y7067 = ~n30814 ;
  assign y7068 = n30816 ;
  assign y7069 = n30822 ;
  assign y7070 = n30828 ;
  assign y7071 = ~n30829 ;
  assign y7072 = n30832 ;
  assign y7073 = n30837 ;
  assign y7074 = ~n30841 ;
  assign y7075 = ~n30844 ;
  assign y7076 = n3109 ;
  assign y7077 = n30847 ;
  assign y7078 = n30853 ;
  assign y7079 = n30860 ;
  assign y7080 = ~n30864 ;
  assign y7081 = ~n30871 ;
  assign y7082 = n30875 ;
  assign y7083 = ~1'b0 ;
  assign y7084 = n30884 ;
  assign y7085 = n30885 ;
  assign y7086 = n30891 ;
  assign y7087 = n30898 ;
  assign y7088 = ~n30899 ;
  assign y7089 = ~n30904 ;
  assign y7090 = ~n30907 ;
  assign y7091 = n30909 ;
  assign y7092 = n30923 ;
  assign y7093 = n30924 ;
  assign y7094 = n30926 ;
  assign y7095 = ~n30930 ;
  assign y7096 = n30933 ;
  assign y7097 = ~1'b0 ;
  assign y7098 = n30937 ;
  assign y7099 = ~n30941 ;
  assign y7100 = n30944 ;
  assign y7101 = n30945 ;
  assign y7102 = n30950 ;
  assign y7103 = n30951 ;
  assign y7104 = ~n30954 ;
  assign y7105 = n30959 ;
  assign y7106 = ~n30961 ;
  assign y7107 = ~n30967 ;
  assign y7108 = n30969 ;
  assign y7109 = n30971 ;
  assign y7110 = ~n30972 ;
  assign y7111 = ~n30976 ;
  assign y7112 = ~n30977 ;
  assign y7113 = ~n30981 ;
  assign y7114 = ~n30982 ;
  assign y7115 = ~n30988 ;
  assign y7116 = ~n30991 ;
  assign y7117 = n30992 ;
  assign y7118 = n30999 ;
  assign y7119 = ~n31005 ;
  assign y7120 = ~n31007 ;
  assign y7121 = ~n31008 ;
  assign y7122 = ~n31009 ;
  assign y7123 = ~n31012 ;
  assign y7124 = ~n31015 ;
  assign y7125 = n31019 ;
  assign y7126 = n31024 ;
  assign y7127 = ~n31027 ;
  assign y7128 = ~n31030 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = n31033 ;
  assign y7131 = n31040 ;
  assign y7132 = ~n31046 ;
  assign y7133 = n31049 ;
  assign y7134 = ~n31053 ;
  assign y7135 = ~n31059 ;
  assign y7136 = n31064 ;
  assign y7137 = n31066 ;
  assign y7138 = ~n31069 ;
  assign y7139 = ~n31073 ;
  assign y7140 = ~n31082 ;
  assign y7141 = n31086 ;
  assign y7142 = ~n31088 ;
  assign y7143 = ~n31097 ;
  assign y7144 = n31099 ;
  assign y7145 = n31100 ;
  assign y7146 = ~n31103 ;
  assign y7147 = n31110 ;
  assign y7148 = n31113 ;
  assign y7149 = n31116 ;
  assign y7150 = n31124 ;
  assign y7151 = n31130 ;
  assign y7152 = ~n31131 ;
  assign y7153 = n31132 ;
  assign y7154 = ~n31135 ;
  assign y7155 = ~1'b0 ;
  assign y7156 = n31140 ;
  assign y7157 = n31145 ;
  assign y7158 = ~n31148 ;
  assign y7159 = ~n31152 ;
  assign y7160 = ~n31155 ;
  assign y7161 = ~n31160 ;
  assign y7162 = ~n31163 ;
  assign y7163 = ~n31171 ;
  assign y7164 = ~n31176 ;
  assign y7165 = n31183 ;
  assign y7166 = ~n31185 ;
  assign y7167 = n31186 ;
  assign y7168 = n31192 ;
  assign y7169 = n31209 ;
  assign y7170 = ~n31212 ;
  assign y7171 = ~n31215 ;
  assign y7172 = ~n31217 ;
  assign y7173 = n31229 ;
  assign y7174 = ~n31235 ;
  assign y7175 = ~n31236 ;
  assign y7176 = ~n31239 ;
  assign y7177 = ~n31242 ;
  assign y7178 = ~n31244 ;
  assign y7179 = n31249 ;
  assign y7180 = n31251 ;
  assign y7181 = n31252 ;
  assign y7182 = ~n31255 ;
  assign y7183 = n31256 ;
  assign y7184 = ~n31258 ;
  assign y7185 = ~n31259 ;
  assign y7186 = ~n31262 ;
  assign y7187 = n31267 ;
  assign y7188 = n31269 ;
  assign y7189 = ~n31271 ;
  assign y7190 = n31274 ;
  assign y7191 = ~n31278 ;
  assign y7192 = ~1'b0 ;
  assign y7193 = n31280 ;
  assign y7194 = ~n31294 ;
  assign y7195 = ~n31300 ;
  assign y7196 = n31305 ;
  assign y7197 = ~1'b0 ;
  assign y7198 = n31309 ;
  assign y7199 = n31312 ;
  assign y7200 = ~n31316 ;
  assign y7201 = n31323 ;
  assign y7202 = n31327 ;
  assign y7203 = ~n31331 ;
  assign y7204 = n31332 ;
  assign y7205 = n31334 ;
  assign y7206 = n31337 ;
  assign y7207 = n31338 ;
  assign y7208 = ~n31341 ;
  assign y7209 = ~n31342 ;
  assign y7210 = n31346 ;
  assign y7211 = ~n31348 ;
  assign y7212 = ~n31351 ;
  assign y7213 = ~n31352 ;
  assign y7214 = ~n31358 ;
  assign y7215 = ~n31360 ;
  assign y7216 = n31361 ;
  assign y7217 = ~n31366 ;
  assign y7218 = n31368 ;
  assign y7219 = ~n31372 ;
  assign y7220 = n31373 ;
  assign y7221 = ~n31378 ;
  assign y7222 = n31386 ;
  assign y7223 = ~n31389 ;
  assign y7224 = ~1'b0 ;
  assign y7225 = n31393 ;
  assign y7226 = n31395 ;
  assign y7227 = n31398 ;
  assign y7228 = n31407 ;
  assign y7229 = ~n31408 ;
  assign y7230 = ~n31410 ;
  assign y7231 = n31414 ;
  assign y7232 = n31415 ;
  assign y7233 = n31417 ;
  assign y7234 = n31419 ;
  assign y7235 = n31421 ;
  assign y7236 = ~n31425 ;
  assign y7237 = n31431 ;
  assign y7238 = ~n31432 ;
  assign y7239 = ~n31433 ;
  assign y7240 = n31434 ;
  assign y7241 = ~n31436 ;
  assign y7242 = ~n31440 ;
  assign y7243 = ~n31450 ;
  assign y7244 = ~n31453 ;
  assign y7245 = ~n31457 ;
  assign y7246 = ~n31458 ;
  assign y7247 = n31459 ;
  assign y7248 = n31461 ;
  assign y7249 = ~n31464 ;
  assign y7250 = ~n31466 ;
  assign y7251 = ~n31477 ;
  assign y7252 = n31478 ;
  assign y7253 = n31479 ;
  assign y7254 = ~n31490 ;
  assign y7255 = n31501 ;
  assign y7256 = ~n31506 ;
  assign y7257 = ~n31507 ;
  assign y7258 = ~n31510 ;
  assign y7259 = n31515 ;
  assign y7260 = n31516 ;
  assign y7261 = ~1'b0 ;
  assign y7262 = n31519 ;
  assign y7263 = n31521 ;
  assign y7264 = ~n31523 ;
  assign y7265 = ~n31527 ;
  assign y7266 = n31537 ;
  assign y7267 = n31541 ;
  assign y7268 = n31542 ;
  assign y7269 = n31546 ;
  assign y7270 = n31549 ;
  assign y7271 = ~n31550 ;
  assign y7272 = ~n31551 ;
  assign y7273 = ~n31553 ;
  assign y7274 = ~1'b0 ;
  assign y7275 = n31556 ;
  assign y7276 = ~n31565 ;
  assign y7277 = n31566 ;
  assign y7278 = n31567 ;
  assign y7279 = ~n31572 ;
  assign y7280 = ~n31573 ;
  assign y7281 = n31578 ;
  assign y7282 = n31581 ;
  assign y7283 = ~n31582 ;
  assign y7284 = ~1'b0 ;
  assign y7285 = ~n31587 ;
  assign y7286 = ~n31588 ;
  assign y7287 = n31590 ;
  assign y7288 = n31591 ;
  assign y7289 = ~n31595 ;
  assign y7290 = n31597 ;
  assign y7291 = n31598 ;
  assign y7292 = ~n31599 ;
  assign y7293 = ~n31600 ;
  assign y7294 = ~n31604 ;
  assign y7295 = ~n31606 ;
  assign y7296 = n31616 ;
  assign y7297 = n31618 ;
  assign y7298 = ~n31629 ;
  assign y7299 = ~n31632 ;
  assign y7300 = ~1'b0 ;
  assign y7301 = ~n31639 ;
  assign y7302 = n31640 ;
  assign y7303 = ~n31644 ;
  assign y7304 = ~n31648 ;
  assign y7305 = ~1'b0 ;
  assign y7306 = n31651 ;
  assign y7307 = ~n31655 ;
  assign y7308 = n31656 ;
  assign y7309 = ~n31657 ;
  assign y7310 = n31658 ;
  assign y7311 = ~n31662 ;
  assign y7312 = ~n31669 ;
  assign y7313 = ~n31672 ;
  assign y7314 = n31674 ;
  assign y7315 = ~n31677 ;
  assign y7316 = n31681 ;
  assign y7317 = n31683 ;
  assign y7318 = ~n31688 ;
  assign y7319 = n31691 ;
  assign y7320 = ~n31693 ;
  assign y7321 = ~n31701 ;
  assign y7322 = ~n31707 ;
  assign y7323 = n31710 ;
  assign y7324 = n31717 ;
  assign y7325 = ~n31718 ;
  assign y7326 = ~n31726 ;
  assign y7327 = n31728 ;
  assign y7328 = n31734 ;
  assign y7329 = n31735 ;
  assign y7330 = ~n31744 ;
  assign y7331 = ~n31748 ;
  assign y7332 = ~n31751 ;
  assign y7333 = n31753 ;
  assign y7334 = ~n31754 ;
  assign y7335 = ~n31757 ;
  assign y7336 = ~n31759 ;
  assign y7337 = n31760 ;
  assign y7338 = ~n31764 ;
  assign y7339 = n31771 ;
  assign y7340 = ~n31781 ;
  assign y7341 = n31785 ;
  assign y7342 = ~1'b0 ;
  assign y7343 = ~n31786 ;
  assign y7344 = ~n31788 ;
  assign y7345 = ~n31789 ;
  assign y7346 = ~n31794 ;
  assign y7347 = ~n31797 ;
  assign y7348 = ~n31800 ;
  assign y7349 = n31803 ;
  assign y7350 = n31804 ;
  assign y7351 = ~n31808 ;
  assign y7352 = 1'b0 ;
  assign y7353 = n31809 ;
  assign y7354 = ~n31810 ;
  assign y7355 = ~n31813 ;
  assign y7356 = n31824 ;
  assign y7357 = ~n31831 ;
  assign y7358 = ~n31835 ;
  assign y7359 = ~n31837 ;
  assign y7360 = ~n31838 ;
  assign y7361 = ~n31839 ;
  assign y7362 = n31843 ;
  assign y7363 = ~n31845 ;
  assign y7364 = n31849 ;
  assign y7365 = n31850 ;
  assign y7366 = ~n31851 ;
  assign y7367 = n31852 ;
  assign y7368 = n31854 ;
  assign y7369 = ~1'b0 ;
  assign y7370 = n31859 ;
  assign y7371 = n31862 ;
  assign y7372 = n31867 ;
  assign y7373 = n31873 ;
  assign y7374 = n31874 ;
  assign y7375 = n31878 ;
  assign y7376 = ~n31886 ;
  assign y7377 = n31891 ;
  assign y7378 = ~n31892 ;
  assign y7379 = n31896 ;
  assign y7380 = ~1'b0 ;
  assign y7381 = ~n31899 ;
  assign y7382 = n31905 ;
  assign y7383 = n31908 ;
  assign y7384 = n31920 ;
  assign y7385 = ~n31925 ;
  assign y7386 = ~n31927 ;
  assign y7387 = ~n31928 ;
  assign y7388 = n31933 ;
  assign y7389 = ~n31934 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = n31940 ;
  assign y7392 = n31944 ;
  assign y7393 = ~n31945 ;
  assign y7394 = ~n31950 ;
  assign y7395 = ~n31952 ;
  assign y7396 = ~n31956 ;
  assign y7397 = ~n31957 ;
  assign y7398 = ~n31958 ;
  assign y7399 = ~n31960 ;
  assign y7400 = ~1'b0 ;
  assign y7401 = n31962 ;
  assign y7402 = n31966 ;
  assign y7403 = n31969 ;
  assign y7404 = ~n31972 ;
  assign y7405 = ~1'b0 ;
  assign y7406 = ~n31974 ;
  assign y7407 = n31976 ;
  assign y7408 = ~n31978 ;
  assign y7409 = ~n31986 ;
  assign y7410 = ~n23112 ;
  assign y7411 = ~n31988 ;
  assign y7412 = n31990 ;
  assign y7413 = n31994 ;
  assign y7414 = n31996 ;
  assign y7415 = n32001 ;
  assign y7416 = n32011 ;
  assign y7417 = n32018 ;
  assign y7418 = ~1'b0 ;
  assign y7419 = ~n32020 ;
  assign y7420 = n32024 ;
  assign y7421 = n32028 ;
  assign y7422 = n32029 ;
  assign y7423 = ~n32034 ;
  assign y7424 = n32039 ;
  assign y7425 = n32043 ;
  assign y7426 = ~n32049 ;
  assign y7427 = n32052 ;
  assign y7428 = ~n32053 ;
  assign y7429 = ~n32058 ;
  assign y7430 = n32061 ;
  assign y7431 = ~1'b0 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = n32069 ;
  assign y7434 = n32070 ;
  assign y7435 = ~n32081 ;
  assign y7436 = ~n32085 ;
  assign y7437 = ~n32092 ;
  assign y7438 = n32093 ;
  assign y7439 = n32097 ;
  assign y7440 = n32099 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = n32100 ;
  assign y7443 = ~n32101 ;
  assign y7444 = ~n32104 ;
  assign y7445 = ~1'b0 ;
  assign y7446 = ~n32109 ;
  assign y7447 = ~n32117 ;
  assign y7448 = n32119 ;
  assign y7449 = n32126 ;
  assign y7450 = ~n32127 ;
  assign y7451 = ~n32130 ;
  assign y7452 = n32132 ;
  assign y7453 = ~n32136 ;
  assign y7454 = ~n32141 ;
  assign y7455 = n32142 ;
  assign y7456 = n32144 ;
  assign y7457 = n32148 ;
  assign y7458 = n32154 ;
  assign y7459 = n32157 ;
  assign y7460 = ~n32166 ;
  assign y7461 = n32167 ;
  assign y7462 = n32170 ;
  assign y7463 = n32175 ;
  assign y7464 = ~1'b0 ;
  assign y7465 = ~n32176 ;
  assign y7466 = ~n32183 ;
  assign y7467 = n32188 ;
  assign y7468 = n32191 ;
  assign y7469 = ~n32193 ;
  assign y7470 = n32199 ;
  assign y7471 = n32200 ;
  assign y7472 = n32202 ;
  assign y7473 = ~n32205 ;
  assign y7474 = n32207 ;
  assign y7475 = n32208 ;
  assign y7476 = ~n32215 ;
  assign y7477 = n32219 ;
  assign y7478 = n32221 ;
  assign y7479 = ~1'b0 ;
  assign y7480 = ~n32228 ;
  assign y7481 = n32230 ;
  assign y7482 = n32231 ;
  assign y7483 = n32234 ;
  assign y7484 = ~n32237 ;
  assign y7485 = ~1'b0 ;
  assign y7486 = n32238 ;
  assign y7487 = n32239 ;
  assign y7488 = n32240 ;
  assign y7489 = ~n32247 ;
  assign y7490 = ~n32250 ;
  assign y7491 = ~n32251 ;
  assign y7492 = n32255 ;
  assign y7493 = ~n32257 ;
  assign y7494 = n32263 ;
  assign y7495 = ~n32265 ;
  assign y7496 = n32267 ;
  assign y7497 = n32269 ;
  assign y7498 = ~n32271 ;
  assign y7499 = ~n32272 ;
  assign y7500 = ~n32274 ;
  assign y7501 = n32276 ;
  assign y7502 = ~n32277 ;
  assign y7503 = ~n32278 ;
  assign y7504 = ~n32281 ;
  assign y7505 = ~n32283 ;
  assign y7506 = n32285 ;
  assign y7507 = ~n32290 ;
  assign y7508 = n32291 ;
  assign y7509 = n32298 ;
  assign y7510 = n32306 ;
  assign y7511 = ~n32314 ;
  assign y7512 = ~n32317 ;
  assign y7513 = n32320 ;
  assign y7514 = ~n32323 ;
  assign y7515 = n32327 ;
  assign y7516 = n32330 ;
  assign y7517 = ~n32331 ;
  assign y7518 = ~n32336 ;
  assign y7519 = n32342 ;
  assign y7520 = ~n32345 ;
  assign y7521 = ~n32348 ;
  assign y7522 = ~n32351 ;
  assign y7523 = n32355 ;
  assign y7524 = ~n32360 ;
  assign y7525 = n32371 ;
  assign y7526 = n13173 ;
  assign y7527 = ~n32374 ;
  assign y7528 = ~n32383 ;
  assign y7529 = ~n32390 ;
  assign y7530 = ~n32393 ;
  assign y7531 = ~n32397 ;
  assign y7532 = n32399 ;
  assign y7533 = ~n32404 ;
  assign y7534 = ~n32405 ;
  assign y7535 = n32407 ;
  assign y7536 = n32409 ;
  assign y7537 = n32410 ;
  assign y7538 = ~n32411 ;
  assign y7539 = n32420 ;
  assign y7540 = ~n32424 ;
  assign y7541 = n32425 ;
  assign y7542 = ~n32426 ;
  assign y7543 = n32427 ;
  assign y7544 = ~n32428 ;
  assign y7545 = ~n32429 ;
  assign y7546 = n32433 ;
  assign y7547 = ~n32440 ;
  assign y7548 = n32442 ;
  assign y7549 = n32445 ;
  assign y7550 = ~n32446 ;
  assign y7551 = n32451 ;
  assign y7552 = n32453 ;
  assign y7553 = ~n32454 ;
  assign y7554 = ~n32461 ;
  assign y7555 = ~n32463 ;
  assign y7556 = n32465 ;
  assign y7557 = n32467 ;
  assign y7558 = ~1'b0 ;
  assign y7559 = n32470 ;
  assign y7560 = n32475 ;
  assign y7561 = n32478 ;
  assign y7562 = ~n32483 ;
  assign y7563 = ~n32485 ;
  assign y7564 = n32488 ;
  assign y7565 = n32490 ;
  assign y7566 = ~n32492 ;
  assign y7567 = n32496 ;
  assign y7568 = ~n32499 ;
  assign y7569 = n32502 ;
  assign y7570 = ~n3053 ;
  assign y7571 = n32503 ;
  assign y7572 = ~n32505 ;
  assign y7573 = ~1'b0 ;
  assign y7574 = ~n32509 ;
  assign y7575 = ~n32511 ;
  assign y7576 = n32513 ;
  assign y7577 = ~n32514 ;
  assign y7578 = ~n32515 ;
  assign y7579 = n32516 ;
  assign y7580 = n32521 ;
  assign y7581 = ~1'b0 ;
  assign y7582 = n32523 ;
  assign y7583 = n32527 ;
  assign y7584 = ~n32529 ;
  assign y7585 = n32531 ;
  assign y7586 = n32535 ;
  assign y7587 = n32538 ;
  assign y7588 = ~n32541 ;
  assign y7589 = ~n32549 ;
  assign y7590 = n32551 ;
  assign y7591 = ~n32554 ;
  assign y7592 = ~n32559 ;
  assign y7593 = n32560 ;
  assign y7594 = n32561 ;
  assign y7595 = n32562 ;
  assign y7596 = ~n32572 ;
  assign y7597 = ~n32574 ;
  assign y7598 = n32575 ;
  assign y7599 = ~n32580 ;
  assign y7600 = ~1'b0 ;
  assign y7601 = ~n32585 ;
  assign y7602 = ~n32593 ;
  assign y7603 = n32594 ;
  assign y7604 = n32597 ;
  assign y7605 = ~n32601 ;
  assign y7606 = ~n32602 ;
  assign y7607 = n32604 ;
  assign y7608 = n32607 ;
  assign y7609 = n32610 ;
  assign y7610 = ~n32613 ;
  assign y7611 = n32614 ;
  assign y7612 = ~n32616 ;
  assign y7613 = n32618 ;
  assign y7614 = ~n32627 ;
  assign y7615 = n32629 ;
  assign y7616 = ~n32632 ;
  assign y7617 = n32635 ;
  assign y7618 = ~n32637 ;
  assign y7619 = n32638 ;
  assign y7620 = n32639 ;
  assign y7621 = ~n32640 ;
  assign y7622 = ~n32645 ;
  assign y7623 = n32652 ;
  assign y7624 = ~n32655 ;
  assign y7625 = n32658 ;
  assign y7626 = ~n32662 ;
  assign y7627 = n32667 ;
  assign y7628 = ~1'b0 ;
  assign y7629 = n32670 ;
  assign y7630 = ~n32673 ;
  assign y7631 = ~1'b0 ;
  assign y7632 = n32680 ;
  assign y7633 = ~n32681 ;
  assign y7634 = ~n32683 ;
  assign y7635 = n32692 ;
  assign y7636 = n32693 ;
  assign y7637 = ~n32695 ;
  assign y7638 = n32698 ;
  assign y7639 = ~n32699 ;
  assign y7640 = n32706 ;
  assign y7641 = ~n32707 ;
  assign y7642 = n32711 ;
  assign y7643 = ~n32714 ;
  assign y7644 = n32723 ;
  assign y7645 = ~n32725 ;
  assign y7646 = ~n32727 ;
  assign y7647 = n32728 ;
  assign y7648 = ~n32735 ;
  assign y7649 = n32736 ;
  assign y7650 = ~n32738 ;
  assign y7651 = n32746 ;
  assign y7652 = n32749 ;
  assign y7653 = ~1'b0 ;
  assign y7654 = n32753 ;
  assign y7655 = n32754 ;
  assign y7656 = n32756 ;
  assign y7657 = ~n32757 ;
  assign y7658 = ~n32766 ;
  assign y7659 = ~n32770 ;
  assign y7660 = n32771 ;
  assign y7661 = ~n32773 ;
  assign y7662 = ~n32776 ;
  assign y7663 = ~n32780 ;
  assign y7664 = ~n32784 ;
  assign y7665 = n32786 ;
  assign y7666 = n32788 ;
  assign y7667 = n32789 ;
  assign y7668 = n32791 ;
  assign y7669 = n32793 ;
  assign y7670 = ~n32796 ;
  assign y7671 = n32800 ;
  assign y7672 = ~1'b0 ;
  assign y7673 = ~n32802 ;
  assign y7674 = ~n32803 ;
  assign y7675 = n32805 ;
  assign y7676 = ~n32813 ;
  assign y7677 = ~n32815 ;
  assign y7678 = ~n32822 ;
  assign y7679 = ~n32823 ;
  assign y7680 = n32826 ;
  assign y7681 = ~1'b0 ;
  assign y7682 = n32831 ;
  assign y7683 = n32837 ;
  assign y7684 = ~n32838 ;
  assign y7685 = n32844 ;
  assign y7686 = n32847 ;
  assign y7687 = n32848 ;
  assign y7688 = ~n32850 ;
  assign y7689 = ~n32851 ;
  assign y7690 = n32853 ;
  assign y7691 = n32857 ;
  assign y7692 = n32859 ;
  assign y7693 = ~n32868 ;
  assign y7694 = ~n32870 ;
  assign y7695 = ~n32875 ;
  assign y7696 = n32877 ;
  assign y7697 = ~n32880 ;
  assign y7698 = ~n32881 ;
  assign y7699 = ~n32882 ;
  assign y7700 = ~n32885 ;
  assign y7701 = ~1'b0 ;
  assign y7702 = ~n32889 ;
  assign y7703 = n32891 ;
  assign y7704 = ~n32894 ;
  assign y7705 = n32899 ;
  assign y7706 = ~1'b0 ;
  assign y7707 = ~n32903 ;
  assign y7708 = ~n32906 ;
  assign y7709 = n32907 ;
  assign y7710 = n32909 ;
  assign y7711 = ~n32912 ;
  assign y7712 = n32915 ;
  assign y7713 = ~n32917 ;
  assign y7714 = n32918 ;
  assign y7715 = n32927 ;
  assign y7716 = ~n32931 ;
  assign y7717 = ~n32937 ;
  assign y7718 = ~n32939 ;
  assign y7719 = n32940 ;
  assign y7720 = ~n32949 ;
  assign y7721 = ~n32950 ;
  assign y7722 = ~n32952 ;
  assign y7723 = n32959 ;
  assign y7724 = ~n32962 ;
  assign y7725 = ~n32963 ;
  assign y7726 = ~n32971 ;
  assign y7727 = ~n32977 ;
  assign y7728 = n32981 ;
  assign y7729 = ~n32984 ;
  assign y7730 = ~n32989 ;
  assign y7731 = ~n32997 ;
  assign y7732 = ~1'b0 ;
  assign y7733 = ~n33012 ;
  assign y7734 = ~n33019 ;
  assign y7735 = ~n33022 ;
  assign y7736 = ~n33025 ;
  assign y7737 = ~n33026 ;
  assign y7738 = ~n33028 ;
  assign y7739 = n33031 ;
  assign y7740 = ~1'b0 ;
  assign y7741 = ~n33034 ;
  assign y7742 = ~n33042 ;
  assign y7743 = ~n33043 ;
  assign y7744 = ~n33044 ;
  assign y7745 = ~n33045 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = n33046 ;
  assign y7748 = n33047 ;
  assign y7749 = n33048 ;
  assign y7750 = n33051 ;
  assign y7751 = ~n33053 ;
  assign y7752 = ~n33054 ;
  assign y7753 = n33055 ;
  assign y7754 = n33057 ;
  assign y7755 = ~n33059 ;
  assign y7756 = n33072 ;
  assign y7757 = ~n33074 ;
  assign y7758 = n33079 ;
  assign y7759 = n33080 ;
  assign y7760 = ~n33082 ;
  assign y7761 = ~1'b0 ;
  assign y7762 = ~n33084 ;
  assign y7763 = ~n33087 ;
  assign y7764 = ~n33089 ;
  assign y7765 = n33097 ;
  assign y7766 = n33110 ;
  assign y7767 = ~1'b0 ;
  assign y7768 = n33114 ;
  assign y7769 = n33116 ;
  assign y7770 = ~n33119 ;
  assign y7771 = ~n33120 ;
  assign y7772 = n33121 ;
  assign y7773 = ~n33123 ;
  assign y7774 = n33128 ;
  assign y7775 = n33133 ;
  assign y7776 = ~n33135 ;
  assign y7777 = n33136 ;
  assign y7778 = n33138 ;
  assign y7779 = n33143 ;
  assign y7780 = ~n33149 ;
  assign y7781 = ~n33151 ;
  assign y7782 = ~n33153 ;
  assign y7783 = ~n33155 ;
  assign y7784 = n33156 ;
  assign y7785 = ~n33162 ;
  assign y7786 = n33164 ;
  assign y7787 = n33170 ;
  assign y7788 = n33177 ;
  assign y7789 = ~n33179 ;
  assign y7790 = n33182 ;
  assign y7791 = n33183 ;
  assign y7792 = ~n33187 ;
  assign y7793 = n33195 ;
  assign y7794 = ~n33204 ;
  assign y7795 = n33209 ;
  assign y7796 = ~1'b0 ;
  assign y7797 = ~n33210 ;
  assign y7798 = n33211 ;
  assign y7799 = ~n33215 ;
  assign y7800 = n33217 ;
  assign y7801 = n33219 ;
  assign y7802 = n33220 ;
  assign y7803 = ~n33225 ;
  assign y7804 = n33229 ;
  assign y7805 = n33231 ;
  assign y7806 = n33234 ;
  assign y7807 = n33237 ;
  assign y7808 = n33247 ;
  assign y7809 = ~n33248 ;
  assign y7810 = ~n33249 ;
  assign y7811 = n33250 ;
  assign y7812 = ~n33251 ;
  assign y7813 = ~n33252 ;
  assign y7814 = ~n33254 ;
  assign y7815 = ~n33257 ;
  assign y7816 = ~n33260 ;
  assign y7817 = n33262 ;
  assign y7818 = ~n33265 ;
  assign y7819 = ~n33266 ;
  assign y7820 = ~n33268 ;
  assign y7821 = ~n33275 ;
  assign y7822 = n33276 ;
  assign y7823 = ~n33277 ;
  assign y7824 = n33280 ;
  assign y7825 = ~n33285 ;
  assign y7826 = ~n33293 ;
  assign y7827 = n33295 ;
  assign y7828 = ~n33297 ;
  assign y7829 = ~n33298 ;
  assign y7830 = n33300 ;
  assign y7831 = ~n33301 ;
  assign y7832 = ~n33302 ;
  assign y7833 = n33308 ;
  assign y7834 = n33311 ;
  assign y7835 = ~n33313 ;
  assign y7836 = ~n33314 ;
  assign y7837 = n33317 ;
  assign y7838 = n33320 ;
  assign y7839 = ~n33321 ;
  assign y7840 = n33322 ;
  assign y7841 = n33328 ;
  assign y7842 = ~n33329 ;
  assign y7843 = ~n33334 ;
  assign y7844 = n33342 ;
  assign y7845 = n33344 ;
  assign y7846 = ~n33345 ;
  assign y7847 = ~n33347 ;
  assign y7848 = ~n33349 ;
  assign y7849 = n33350 ;
  assign y7850 = ~n33365 ;
  assign y7851 = ~n33369 ;
  assign y7852 = n33370 ;
  assign y7853 = n33371 ;
  assign y7854 = n33373 ;
  assign y7855 = n33377 ;
  assign y7856 = n33380 ;
  assign y7857 = ~1'b0 ;
  assign y7858 = n33382 ;
  assign y7859 = ~n33383 ;
  assign y7860 = n33387 ;
  assign y7861 = ~1'b0 ;
  assign y7862 = ~n33402 ;
  assign y7863 = n33405 ;
  assign y7864 = ~n33408 ;
  assign y7865 = ~n33411 ;
  assign y7866 = ~n33414 ;
  assign y7867 = ~n33417 ;
  assign y7868 = ~n33418 ;
  assign y7869 = n33420 ;
  assign y7870 = ~n33424 ;
  assign y7871 = n33425 ;
  assign y7872 = n33428 ;
  assign y7873 = n33430 ;
  assign y7874 = ~n33434 ;
  assign y7875 = n33439 ;
  assign y7876 = ~n33446 ;
  assign y7877 = ~n33453 ;
  assign y7878 = ~n33456 ;
  assign y7879 = ~1'b0 ;
  assign y7880 = ~n33457 ;
  assign y7881 = ~n33459 ;
  assign y7882 = n33462 ;
  assign y7883 = ~n33466 ;
  assign y7884 = ~1'b0 ;
  assign y7885 = n33468 ;
  assign y7886 = n33469 ;
  assign y7887 = n33473 ;
  assign y7888 = n33475 ;
  assign y7889 = n33477 ;
  assign y7890 = ~n33481 ;
  assign y7891 = n33482 ;
  assign y7892 = ~n33483 ;
  assign y7893 = n33489 ;
  assign y7894 = ~n33490 ;
  assign y7895 = n33492 ;
  assign y7896 = n33495 ;
  assign y7897 = n33502 ;
  assign y7898 = n33509 ;
  assign y7899 = ~1'b0 ;
  assign y7900 = n33512 ;
  assign y7901 = n33513 ;
  assign y7902 = n33514 ;
  assign y7903 = ~n33516 ;
  assign y7904 = ~n33518 ;
  assign y7905 = ~n33519 ;
  assign y7906 = n33521 ;
  assign y7907 = n33524 ;
  assign y7908 = ~n33529 ;
  assign y7909 = ~n33535 ;
  assign y7910 = ~n33537 ;
  assign y7911 = ~n33539 ;
  assign y7912 = ~n33540 ;
  assign y7913 = ~n33544 ;
  assign y7914 = ~n33546 ;
  assign y7915 = ~n33547 ;
  assign y7916 = ~n33549 ;
  assign y7917 = ~n33553 ;
  assign y7918 = ~n33558 ;
  assign y7919 = ~n33560 ;
  assign y7920 = n33561 ;
  assign y7921 = n33565 ;
  assign y7922 = ~n33567 ;
  assign y7923 = ~1'b0 ;
  assign y7924 = n33569 ;
  assign y7925 = n33572 ;
  assign y7926 = n33575 ;
  assign y7927 = ~n33578 ;
  assign y7928 = ~n33582 ;
  assign y7929 = n33586 ;
  assign y7930 = ~n33590 ;
  assign y7931 = n33600 ;
  assign y7932 = ~n33602 ;
  assign y7933 = ~n33611 ;
  assign y7934 = n33613 ;
  assign y7935 = n33616 ;
  assign y7936 = ~1'b0 ;
  assign y7937 = n33618 ;
  assign y7938 = ~n33619 ;
  assign y7939 = n33622 ;
  assign y7940 = ~n33631 ;
  assign y7941 = n33640 ;
  assign y7942 = n33643 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = ~n33649 ;
  assign y7945 = n33657 ;
  assign y7946 = ~n33660 ;
  assign y7947 = ~n33663 ;
  assign y7948 = ~n33669 ;
  assign y7949 = n33675 ;
  assign y7950 = ~n33681 ;
  assign y7951 = n33684 ;
  assign y7952 = n33685 ;
  assign y7953 = n33686 ;
  assign y7954 = ~n33687 ;
  assign y7955 = ~n33690 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = ~n33691 ;
  assign y7958 = n33696 ;
  assign y7959 = ~n33699 ;
  assign y7960 = n33706 ;
  assign y7961 = ~n33709 ;
  assign y7962 = n33710 ;
  assign y7963 = n33716 ;
  assign y7964 = n33717 ;
  assign y7965 = ~n33721 ;
  assign y7966 = ~n33725 ;
  assign y7967 = ~1'b0 ;
  assign y7968 = ~n33727 ;
  assign y7969 = n33730 ;
  assign y7970 = ~n33731 ;
  assign y7971 = n33733 ;
  assign y7972 = n33734 ;
  assign y7973 = n33739 ;
  assign y7974 = n33745 ;
  assign y7975 = n33746 ;
  assign y7976 = ~n33752 ;
  assign y7977 = ~n33755 ;
  assign y7978 = ~n33761 ;
  assign y7979 = n33762 ;
  assign y7980 = ~1'b0 ;
  assign y7981 = ~n33770 ;
  assign y7982 = n33774 ;
  assign y7983 = n33776 ;
  assign y7984 = ~n33783 ;
  assign y7985 = ~n33786 ;
  assign y7986 = n33787 ;
  assign y7987 = n33789 ;
  assign y7988 = ~n33796 ;
  assign y7989 = ~n33800 ;
  assign y7990 = ~n33803 ;
  assign y7991 = n16453 ;
  assign y7992 = n33805 ;
  assign y7993 = ~n33806 ;
  assign y7994 = ~1'b0 ;
  assign y7995 = n33807 ;
  assign y7996 = ~n33810 ;
  assign y7997 = ~n33816 ;
  assign y7998 = n33820 ;
  assign y7999 = n33823 ;
  assign y8000 = ~n33828 ;
  assign y8001 = ~n33830 ;
  assign y8002 = ~n33834 ;
  assign y8003 = n33838 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = n33839 ;
  assign y8006 = n33840 ;
  assign y8007 = ~n33844 ;
  assign y8008 = n33846 ;
  assign y8009 = n33847 ;
  assign y8010 = n33851 ;
  assign y8011 = ~n33854 ;
  assign y8012 = n33859 ;
  assign y8013 = ~n33863 ;
  assign y8014 = ~n33865 ;
  assign y8015 = ~n33868 ;
  assign y8016 = ~n33871 ;
  assign y8017 = n33873 ;
  assign y8018 = ~n33875 ;
  assign y8019 = n33879 ;
  assign y8020 = n33894 ;
  assign y8021 = n33895 ;
  assign y8022 = ~n33901 ;
  assign y8023 = n33902 ;
  assign y8024 = n33906 ;
  assign y8025 = ~n33909 ;
  assign y8026 = ~n33915 ;
  assign y8027 = n33916 ;
  assign y8028 = ~n33919 ;
  assign y8029 = n33923 ;
  assign y8030 = n12082 ;
  assign y8031 = ~n33929 ;
  assign y8032 = ~n33930 ;
  assign y8033 = ~n33931 ;
  assign y8034 = ~n33935 ;
  assign y8035 = ~n33938 ;
  assign y8036 = ~n33945 ;
  assign y8037 = ~n33946 ;
  assign y8038 = n33948 ;
  assign y8039 = ~n33950 ;
  assign y8040 = n33953 ;
  assign y8041 = ~n33958 ;
  assign y8042 = n33960 ;
  assign y8043 = ~n12426 ;
  assign y8044 = ~n33968 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = ~1'b0 ;
  assign y8047 = n33975 ;
  assign y8048 = ~n33980 ;
  assign y8049 = ~n33984 ;
  assign y8050 = ~n33985 ;
  assign y8051 = n33990 ;
  assign y8052 = ~n33994 ;
  assign y8053 = n33999 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = n34000 ;
  assign y8056 = n34002 ;
  assign y8057 = ~n34011 ;
  assign y8058 = ~n34019 ;
  assign y8059 = n34025 ;
  assign y8060 = ~n34026 ;
  assign y8061 = ~n34027 ;
  assign y8062 = ~n34028 ;
  assign y8063 = ~n34030 ;
  assign y8064 = n34034 ;
  assign y8065 = ~n34036 ;
  assign y8066 = n34037 ;
  assign y8067 = n34038 ;
  assign y8068 = ~n34039 ;
  assign y8069 = n34041 ;
  assign y8070 = n34044 ;
  assign y8071 = n34049 ;
  assign y8072 = n34052 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = ~n34053 ;
  assign y8075 = ~n34064 ;
  assign y8076 = n34065 ;
  assign y8077 = ~1'b0 ;
  assign y8078 = n34067 ;
  assign y8079 = n34069 ;
  assign y8080 = ~n34070 ;
  assign y8081 = ~n34075 ;
  assign y8082 = n34077 ;
  assign y8083 = ~n34078 ;
  assign y8084 = n34082 ;
  assign y8085 = ~n34091 ;
  assign y8086 = n34093 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~n34096 ;
  assign y8089 = n34098 ;
  assign y8090 = n34100 ;
  assign y8091 = ~n34102 ;
  assign y8092 = ~1'b0 ;
  assign y8093 = ~1'b0 ;
  assign y8094 = n34104 ;
  assign y8095 = ~n34105 ;
  assign y8096 = ~n34108 ;
  assign y8097 = n34109 ;
  assign y8098 = ~n34114 ;
  assign y8099 = ~n34122 ;
  assign y8100 = ~n34124 ;
  assign y8101 = ~n34125 ;
  assign y8102 = ~n34126 ;
  assign y8103 = n34128 ;
  assign y8104 = n34130 ;
  assign y8105 = n34136 ;
  assign y8106 = n34140 ;
  assign y8107 = ~n34147 ;
  assign y8108 = n34150 ;
  assign y8109 = n34152 ;
  assign y8110 = n34158 ;
  assign y8111 = ~n34161 ;
  assign y8112 = ~n34164 ;
  assign y8113 = n34168 ;
  assign y8114 = n34169 ;
  assign y8115 = n34171 ;
  assign y8116 = n34172 ;
  assign y8117 = n34173 ;
  assign y8118 = n34177 ;
  assign y8119 = n34179 ;
  assign y8120 = ~n34180 ;
  assign y8121 = n34187 ;
  assign y8122 = n34188 ;
  assign y8123 = n34189 ;
  assign y8124 = ~n34197 ;
  assign y8125 = ~n34199 ;
  assign y8126 = ~n34200 ;
  assign y8127 = ~n34201 ;
  assign y8128 = ~n34204 ;
  assign y8129 = ~n34210 ;
  assign y8130 = n34211 ;
  assign y8131 = ~n34212 ;
  assign y8132 = ~n34215 ;
  assign y8133 = n34219 ;
  assign y8134 = ~n34223 ;
  assign y8135 = ~n34226 ;
  assign y8136 = ~n34227 ;
  assign y8137 = ~n34228 ;
  assign y8138 = ~n34245 ;
  assign y8139 = ~n34251 ;
  assign y8140 = ~n34253 ;
  assign y8141 = ~1'b0 ;
  assign y8142 = n34264 ;
  assign y8143 = ~n34267 ;
  assign y8144 = n34268 ;
  assign y8145 = n34279 ;
  assign y8146 = n34288 ;
  assign y8147 = ~n34289 ;
  assign y8148 = n34290 ;
  assign y8149 = n34292 ;
  assign y8150 = n34297 ;
  assign y8151 = n34300 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = n34303 ;
  assign y8154 = n34305 ;
  assign y8155 = n34309 ;
  assign y8156 = n34311 ;
  assign y8157 = ~n34312 ;
  assign y8158 = ~n34313 ;
  assign y8159 = n34316 ;
  assign y8160 = n34318 ;
  assign y8161 = ~n34319 ;
  assign y8162 = ~1'b0 ;
  assign y8163 = n34324 ;
  assign y8164 = ~1'b0 ;
  assign y8165 = ~n34325 ;
  assign y8166 = ~n34328 ;
  assign y8167 = ~n34330 ;
  assign y8168 = n34333 ;
  assign y8169 = ~1'b0 ;
  assign y8170 = ~1'b0 ;
  assign y8171 = ~1'b0 ;
  assign y8172 = ~n34336 ;
  assign y8173 = n34338 ;
  assign y8174 = n34340 ;
  assign y8175 = ~n34342 ;
  assign y8176 = ~n34343 ;
  assign y8177 = n34344 ;
  assign y8178 = ~n34349 ;
  assign y8179 = n34354 ;
  assign y8180 = n34356 ;
  assign y8181 = n34357 ;
  assign y8182 = ~n34360 ;
  assign y8183 = ~1'b0 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~n34363 ;
  assign y8186 = ~n34364 ;
  assign y8187 = ~n34366 ;
  assign y8188 = n34368 ;
  assign y8189 = ~n34370 ;
  assign y8190 = ~n34374 ;
  assign y8191 = ~n34376 ;
  assign y8192 = ~n34379 ;
  assign y8193 = ~n34385 ;
  assign y8194 = n34387 ;
  assign y8195 = ~1'b0 ;
  assign y8196 = n34396 ;
  assign y8197 = ~n34403 ;
  assign y8198 = ~n34406 ;
  assign y8199 = n34408 ;
  assign y8200 = n34411 ;
  assign y8201 = ~n34414 ;
  assign y8202 = n34416 ;
  assign y8203 = n34422 ;
  assign y8204 = ~n34424 ;
  assign y8205 = ~n34428 ;
  assign y8206 = n34429 ;
  assign y8207 = ~n34430 ;
  assign y8208 = ~n34434 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = ~n34435 ;
  assign y8211 = ~n34437 ;
  assign y8212 = ~n34440 ;
  assign y8213 = n34446 ;
  assign y8214 = ~n34450 ;
  assign y8215 = n34452 ;
  assign y8216 = ~n34455 ;
  assign y8217 = n34457 ;
  assign y8218 = ~n34460 ;
  assign y8219 = n34461 ;
  assign y8220 = ~n34465 ;
  assign y8221 = ~1'b0 ;
  assign y8222 = n34466 ;
  assign y8223 = ~n34468 ;
  assign y8224 = n34473 ;
  assign y8225 = n34477 ;
  assign y8226 = n34478 ;
  assign y8227 = n34480 ;
  assign y8228 = ~n34484 ;
  assign y8229 = ~n34494 ;
  assign y8230 = ~n34496 ;
  assign y8231 = n34497 ;
  assign y8232 = n34501 ;
  assign y8233 = n34502 ;
  assign y8234 = ~n34505 ;
  assign y8235 = ~1'b0 ;
  assign y8236 = n34510 ;
  assign y8237 = n34513 ;
  assign y8238 = ~n34514 ;
  assign y8239 = n34516 ;
  assign y8240 = n34518 ;
  assign y8241 = ~1'b0 ;
  assign y8242 = n34520 ;
  assign y8243 = ~n34522 ;
  assign y8244 = ~n34525 ;
  assign y8245 = ~n34534 ;
  assign y8246 = ~n34536 ;
  assign y8247 = n34540 ;
  assign y8248 = ~1'b0 ;
  assign y8249 = ~n34544 ;
  assign y8250 = ~n34545 ;
  assign y8251 = ~n34549 ;
  assign y8252 = n34552 ;
  assign y8253 = n34553 ;
  assign y8254 = ~1'b0 ;
  assign y8255 = ~n34554 ;
  assign y8256 = n34555 ;
  assign y8257 = ~n34556 ;
  assign y8258 = ~n34560 ;
  assign y8259 = ~n34561 ;
  assign y8260 = n34562 ;
  assign y8261 = ~n34569 ;
  assign y8262 = n34570 ;
  assign y8263 = ~n34573 ;
  assign y8264 = ~n34575 ;
  assign y8265 = n34586 ;
  assign y8266 = n34595 ;
  assign y8267 = n34599 ;
  assign y8268 = n34600 ;
  assign y8269 = n34603 ;
  assign y8270 = ~1'b0 ;
  assign y8271 = ~n34605 ;
  assign y8272 = ~n34606 ;
  assign y8273 = n34609 ;
  assign y8274 = ~n34616 ;
  assign y8275 = ~n34619 ;
  assign y8276 = ~1'b0 ;
  assign y8277 = n34621 ;
  assign y8278 = ~n34623 ;
  assign y8279 = ~n34628 ;
  assign y8280 = n34632 ;
  assign y8281 = ~n34638 ;
  assign y8282 = n34643 ;
  assign y8283 = n34646 ;
  assign y8284 = ~1'b0 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = ~n34648 ;
  assign y8287 = n34652 ;
  assign y8288 = n34655 ;
  assign y8289 = ~n34657 ;
  assign y8290 = ~n34660 ;
  assign y8291 = n34662 ;
  assign y8292 = n34664 ;
  assign y8293 = n34666 ;
  assign y8294 = n34668 ;
  assign y8295 = n34680 ;
  assign y8296 = n34681 ;
  assign y8297 = ~n34683 ;
  assign y8298 = n34687 ;
  assign y8299 = ~n34689 ;
  assign y8300 = n34690 ;
  assign y8301 = ~n34692 ;
  assign y8302 = n34698 ;
  assign y8303 = n34699 ;
  assign y8304 = n34702 ;
  assign y8305 = ~n34707 ;
  assign y8306 = ~n34708 ;
  assign y8307 = ~1'b0 ;
  assign y8308 = ~1'b0 ;
  assign y8309 = ~n34712 ;
  assign y8310 = ~n34713 ;
  assign y8311 = ~n34714 ;
  assign y8312 = ~n34717 ;
  assign y8313 = ~n34718 ;
  assign y8314 = ~n34723 ;
  assign y8315 = ~n34724 ;
  assign y8316 = n34729 ;
  assign y8317 = ~n34730 ;
  assign y8318 = ~n34734 ;
  assign y8319 = ~n34740 ;
  assign y8320 = n34741 ;
  assign y8321 = n34742 ;
  assign y8322 = n34743 ;
  assign y8323 = n34744 ;
  assign y8324 = ~n34747 ;
  assign y8325 = ~n34748 ;
  assign y8326 = ~n34749 ;
  assign y8327 = n34750 ;
  assign y8328 = ~n34751 ;
  assign y8329 = n34752 ;
  assign y8330 = n34755 ;
  assign y8331 = ~n34757 ;
  assign y8332 = ~1'b0 ;
  assign y8333 = n34758 ;
  assign y8334 = ~n34761 ;
  assign y8335 = n34770 ;
  assign y8336 = n34771 ;
  assign y8337 = ~n34776 ;
  assign y8338 = ~n34779 ;
  assign y8339 = ~n34781 ;
  assign y8340 = ~n34784 ;
  assign y8341 = ~n34785 ;
  assign y8342 = n34786 ;
  assign y8343 = n34788 ;
  assign y8344 = n34792 ;
  assign y8345 = ~n34797 ;
  assign y8346 = ~n34799 ;
  assign y8347 = n34803 ;
  assign y8348 = ~n34804 ;
  assign y8349 = n34805 ;
  assign y8350 = n34809 ;
  assign y8351 = ~n34811 ;
  assign y8352 = ~n34813 ;
  assign y8353 = ~n34815 ;
  assign y8354 = n34816 ;
  assign y8355 = n34819 ;
  assign y8356 = ~n34826 ;
  assign y8357 = n34827 ;
  assign y8358 = ~n34831 ;
  assign y8359 = ~n34834 ;
  assign y8360 = n34837 ;
  assign y8361 = n34838 ;
  assign y8362 = ~n34841 ;
  assign y8363 = n34843 ;
  assign y8364 = ~n34847 ;
  assign y8365 = ~n34849 ;
  assign y8366 = ~n34850 ;
  assign y8367 = ~n34851 ;
  assign y8368 = ~n34852 ;
  assign y8369 = n34853 ;
  assign y8370 = ~n34854 ;
  assign y8371 = ~1'b0 ;
  assign y8372 = ~n34857 ;
  assign y8373 = ~n34861 ;
  assign y8374 = n34867 ;
  assign y8375 = n34868 ;
  assign y8376 = n34869 ;
  assign y8377 = n34871 ;
  assign y8378 = ~n34873 ;
  assign y8379 = n34875 ;
  assign y8380 = ~n2952 ;
  assign y8381 = n34879 ;
  assign y8382 = ~n34880 ;
  assign y8383 = n34888 ;
  assign y8384 = n34891 ;
  assign y8385 = ~n34897 ;
  assign y8386 = n34905 ;
  assign y8387 = ~n34906 ;
  assign y8388 = ~n34911 ;
  assign y8389 = ~1'b0 ;
  assign y8390 = ~1'b0 ;
  assign y8391 = ~1'b0 ;
  assign y8392 = ~n34914 ;
  assign y8393 = ~1'b0 ;
  assign y8394 = ~n34918 ;
  assign y8395 = n34919 ;
  assign y8396 = ~n34920 ;
  assign y8397 = n34921 ;
  assign y8398 = n34925 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = n34946 ;
  assign y8401 = n34955 ;
  assign y8402 = ~n34958 ;
  assign y8403 = ~n34963 ;
  assign y8404 = ~n34967 ;
  assign y8405 = ~1'b0 ;
  assign y8406 = ~1'b0 ;
  assign y8407 = ~1'b0 ;
  assign y8408 = n34968 ;
  assign y8409 = n34969 ;
  assign y8410 = n34971 ;
  assign y8411 = n34972 ;
  assign y8412 = ~n34974 ;
  assign y8413 = ~n34977 ;
  assign y8414 = ~n34982 ;
  assign y8415 = n34983 ;
  assign y8416 = ~n34984 ;
  assign y8417 = ~n34985 ;
  assign y8418 = ~n34986 ;
  assign y8419 = n34988 ;
  assign y8420 = ~1'b0 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = ~n34989 ;
  assign y8423 = n34996 ;
  assign y8424 = ~n34997 ;
  assign y8425 = n35002 ;
  assign y8426 = n35004 ;
  assign y8427 = ~n35012 ;
  assign y8428 = ~n35015 ;
  assign y8429 = n35019 ;
  assign y8430 = n35021 ;
  assign y8431 = ~n35027 ;
  assign y8432 = n35031 ;
  assign y8433 = ~n35032 ;
  assign y8434 = ~n35039 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~n35040 ;
  assign y8437 = n35043 ;
  assign y8438 = n35047 ;
  assign y8439 = n35049 ;
  assign y8440 = n35050 ;
  assign y8441 = n35053 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = ~n35056 ;
  assign y8444 = ~n35059 ;
  assign y8445 = ~n35062 ;
  assign y8446 = n35068 ;
  assign y8447 = ~n35071 ;
  assign y8448 = ~n35075 ;
  assign y8449 = n35078 ;
  assign y8450 = ~1'b0 ;
  assign y8451 = ~n35081 ;
  assign y8452 = n35083 ;
  assign y8453 = ~n35084 ;
  assign y8454 = n35086 ;
  assign y8455 = n35087 ;
  assign y8456 = ~n35089 ;
  assign y8457 = ~n35091 ;
  assign y8458 = ~n35094 ;
  assign y8459 = n35096 ;
  assign y8460 = n35099 ;
  assign y8461 = n35101 ;
  assign y8462 = ~n35103 ;
  assign y8463 = ~n35104 ;
  assign y8464 = n35108 ;
  assign y8465 = ~n35116 ;
  assign y8466 = n35122 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = n35124 ;
  assign y8469 = n35135 ;
  assign y8470 = ~n35136 ;
  assign y8471 = n6464 ;
  assign y8472 = ~n35141 ;
  assign y8473 = n35143 ;
  assign y8474 = n35147 ;
  assign y8475 = n35150 ;
  assign y8476 = ~n35152 ;
  assign y8477 = ~1'b0 ;
  assign y8478 = n35154 ;
  assign y8479 = ~n35160 ;
  assign y8480 = n35161 ;
  assign y8481 = ~n35162 ;
  assign y8482 = ~n35167 ;
  assign y8483 = ~n35169 ;
  assign y8484 = n35172 ;
  assign y8485 = n35177 ;
  assign y8486 = ~n35186 ;
  assign y8487 = ~n35187 ;
  assign y8488 = ~n35189 ;
  assign y8489 = ~n35193 ;
  assign y8490 = ~n35199 ;
  assign y8491 = n35203 ;
  assign y8492 = n35204 ;
  assign y8493 = ~1'b0 ;
  assign y8494 = ~n35206 ;
  assign y8495 = ~n35208 ;
  assign y8496 = ~n35212 ;
  assign y8497 = n35215 ;
  assign y8498 = ~n35216 ;
  assign y8499 = n35217 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = n35219 ;
  assign y8502 = n35220 ;
  assign y8503 = n35221 ;
  assign y8504 = n35222 ;
  assign y8505 = ~n35225 ;
  assign y8506 = n35239 ;
  assign y8507 = ~n35241 ;
  assign y8508 = ~n35242 ;
  assign y8509 = n35245 ;
  assign y8510 = ~n35246 ;
  assign y8511 = ~n35249 ;
  assign y8512 = n35251 ;
  assign y8513 = n35252 ;
  assign y8514 = ~1'b0 ;
  assign y8515 = ~1'b0 ;
  assign y8516 = ~n35255 ;
  assign y8517 = n35258 ;
  assign y8518 = ~n35259 ;
  assign y8519 = ~n35263 ;
  assign y8520 = ~n35264 ;
  assign y8521 = ~1'b0 ;
  assign y8522 = n35265 ;
  assign y8523 = n35267 ;
  assign y8524 = ~n25122 ;
  assign y8525 = n35268 ;
  assign y8526 = ~n35271 ;
  assign y8527 = ~n35274 ;
  assign y8528 = n35276 ;
  assign y8529 = ~n35277 ;
  assign y8530 = ~n35279 ;
  assign y8531 = ~1'b0 ;
  assign y8532 = n35280 ;
  assign y8533 = n35281 ;
  assign y8534 = ~n35284 ;
  assign y8535 = n35285 ;
  assign y8536 = ~n35288 ;
  assign y8537 = n35290 ;
  assign y8538 = ~n35295 ;
  assign y8539 = n35297 ;
  assign y8540 = ~n35298 ;
  assign y8541 = ~n35302 ;
  assign y8542 = ~n35304 ;
  assign y8543 = n35306 ;
  assign y8544 = n35309 ;
  assign y8545 = n35313 ;
  assign y8546 = ~n35315 ;
  assign y8547 = ~n35319 ;
  assign y8548 = n35323 ;
  assign y8549 = ~n35324 ;
  assign y8550 = ~n35325 ;
  assign y8551 = n35326 ;
  assign y8552 = n35331 ;
  assign y8553 = ~n35336 ;
  assign y8554 = ~1'b0 ;
  assign y8555 = ~1'b0 ;
  assign y8556 = n35339 ;
  assign y8557 = n35340 ;
  assign y8558 = n35343 ;
  assign y8559 = ~n35344 ;
  assign y8560 = n35346 ;
  assign y8561 = n35348 ;
  assign y8562 = n35351 ;
  assign y8563 = ~n35357 ;
  assign y8564 = n35360 ;
  assign y8565 = ~n35363 ;
  assign y8566 = n35364 ;
  assign y8567 = n35366 ;
  assign y8568 = n35367 ;
  assign y8569 = ~n35374 ;
  assign y8570 = ~n35377 ;
  assign y8571 = ~n35383 ;
  assign y8572 = ~n35394 ;
  assign y8573 = ~n35396 ;
  assign y8574 = ~n35400 ;
  assign y8575 = n35401 ;
  assign y8576 = ~n35402 ;
  assign y8577 = n35403 ;
  assign y8578 = ~n35406 ;
  assign y8579 = n35410 ;
  assign y8580 = ~n35414 ;
  assign y8581 = ~n35422 ;
  assign y8582 = n35423 ;
  assign y8583 = ~n35425 ;
  assign y8584 = ~n35429 ;
  assign y8585 = ~n35431 ;
  assign y8586 = ~n35433 ;
  assign y8587 = ~1'b0 ;
  assign y8588 = ~1'b0 ;
  assign y8589 = ~n35434 ;
  assign y8590 = n35440 ;
  assign y8591 = ~n35441 ;
  assign y8592 = ~1'b0 ;
  assign y8593 = ~n35442 ;
  assign y8594 = ~n35443 ;
  assign y8595 = n35445 ;
  assign y8596 = n35446 ;
  assign y8597 = ~n35447 ;
  assign y8598 = ~n35449 ;
  assign y8599 = ~n35463 ;
  assign y8600 = n35466 ;
  assign y8601 = ~n35467 ;
  assign y8602 = ~n35468 ;
  assign y8603 = ~n35469 ;
  assign y8604 = ~n35471 ;
  assign y8605 = n35472 ;
  assign y8606 = ~n35477 ;
  assign y8607 = n35478 ;
  assign y8608 = n35479 ;
  assign y8609 = n35480 ;
  assign y8610 = ~n35483 ;
  assign y8611 = n35487 ;
  assign y8612 = n35488 ;
  assign y8613 = n35489 ;
  assign y8614 = n35491 ;
  assign y8615 = ~n35499 ;
  assign y8616 = n35500 ;
  assign y8617 = ~n35506 ;
  assign y8618 = n35509 ;
  assign y8619 = n35510 ;
  assign y8620 = n35512 ;
  assign y8621 = ~n35514 ;
  assign y8622 = n35515 ;
  assign y8623 = ~n35521 ;
  assign y8624 = ~1'b0 ;
  assign y8625 = n35522 ;
  assign y8626 = ~n35525 ;
  assign y8627 = n35526 ;
  assign y8628 = ~n35528 ;
  assign y8629 = n35536 ;
  assign y8630 = ~n35539 ;
  assign y8631 = n35541 ;
  assign y8632 = n35542 ;
  assign y8633 = n35545 ;
  assign y8634 = ~n35547 ;
  assign y8635 = n35548 ;
  assign y8636 = n35550 ;
  assign y8637 = ~n35552 ;
  assign y8638 = n35553 ;
  assign y8639 = ~n35554 ;
  assign y8640 = ~n35557 ;
  assign y8641 = n35558 ;
  assign y8642 = n35560 ;
  assign y8643 = n35561 ;
  assign y8644 = n35564 ;
  assign y8645 = ~n35573 ;
  assign y8646 = ~n35576 ;
  assign y8647 = n35579 ;
  assign y8648 = n35580 ;
  assign y8649 = n6171 ;
  assign y8650 = ~1'b0 ;
  assign y8651 = ~n35581 ;
  assign y8652 = n35584 ;
  assign y8653 = n35586 ;
  assign y8654 = n35591 ;
  assign y8655 = ~n35595 ;
  assign y8656 = ~n35607 ;
  assign y8657 = ~1'b0 ;
  assign y8658 = ~n35609 ;
  assign y8659 = n35611 ;
  assign y8660 = n35612 ;
  assign y8661 = ~n35616 ;
  assign y8662 = n35617 ;
  assign y8663 = ~n35621 ;
  assign y8664 = ~n35623 ;
  assign y8665 = n35624 ;
  assign y8666 = ~n35627 ;
  assign y8667 = n35631 ;
  assign y8668 = n35636 ;
  assign y8669 = ~n35639 ;
  assign y8670 = ~n35645 ;
  assign y8671 = ~1'b0 ;
  assign y8672 = n35646 ;
  assign y8673 = ~n35647 ;
  assign y8674 = ~n35652 ;
  assign y8675 = ~n35659 ;
  assign y8676 = ~n35661 ;
  assign y8677 = ~1'b0 ;
  assign y8678 = ~n35662 ;
  assign y8679 = ~n35664 ;
  assign y8680 = n35667 ;
  assign y8681 = n35669 ;
  assign y8682 = ~n35671 ;
  assign y8683 = ~n35673 ;
  assign y8684 = n35674 ;
  assign y8685 = ~n35679 ;
  assign y8686 = ~n35682 ;
  assign y8687 = n35685 ;
  assign y8688 = n35690 ;
  assign y8689 = ~n35692 ;
  assign y8690 = n35698 ;
  assign y8691 = ~n35699 ;
  assign y8692 = ~n35703 ;
  assign y8693 = ~n35707 ;
  assign y8694 = ~n35713 ;
  assign y8695 = ~n35717 ;
  assign y8696 = n35723 ;
  assign y8697 = n35725 ;
  assign y8698 = ~n35726 ;
  assign y8699 = ~n35727 ;
  assign y8700 = ~n35728 ;
  assign y8701 = n35730 ;
  assign y8702 = ~n35731 ;
  assign y8703 = n35732 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = n35741 ;
  assign y8707 = n35743 ;
  assign y8708 = n35744 ;
  assign y8709 = n35748 ;
  assign y8710 = n35750 ;
  assign y8711 = ~n35752 ;
  assign y8712 = n35753 ;
  assign y8713 = n35756 ;
  assign y8714 = ~n35759 ;
  assign y8715 = n35763 ;
  assign y8716 = n35767 ;
  assign y8717 = ~n35770 ;
  assign y8718 = n35775 ;
  assign y8719 = ~n35776 ;
  assign y8720 = n35781 ;
  assign y8721 = n35785 ;
  assign y8722 = ~1'b0 ;
  assign y8723 = n35786 ;
  assign y8724 = ~n35788 ;
  assign y8725 = n35790 ;
  assign y8726 = ~n12507 ;
  assign y8727 = ~n35794 ;
  assign y8728 = n35797 ;
  assign y8729 = ~n35802 ;
  assign y8730 = ~n35803 ;
  assign y8731 = ~n35808 ;
  assign y8732 = n35812 ;
  assign y8733 = ~n35814 ;
  assign y8734 = n35815 ;
  assign y8735 = ~1'b0 ;
  assign y8736 = ~n35817 ;
  assign y8737 = n35823 ;
  assign y8738 = n35825 ;
  assign y8739 = n35828 ;
  assign y8740 = ~n35829 ;
  assign y8741 = n35837 ;
  assign y8742 = ~n35839 ;
  assign y8743 = n35841 ;
  assign y8744 = ~n35842 ;
  assign y8745 = ~n35853 ;
  assign y8746 = ~n35854 ;
  assign y8747 = ~n35856 ;
  assign y8748 = n35862 ;
  assign y8749 = ~n35863 ;
  assign y8750 = n35864 ;
  assign y8751 = ~n35867 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = n35870 ;
  assign y8754 = n35879 ;
  assign y8755 = n35880 ;
  assign y8756 = ~n35884 ;
  assign y8757 = n35885 ;
  assign y8758 = ~n35887 ;
  assign y8759 = n35889 ;
  assign y8760 = ~n35891 ;
  assign y8761 = ~n35897 ;
  assign y8762 = ~n35903 ;
  assign y8763 = n35908 ;
  assign y8764 = ~n35912 ;
  assign y8765 = ~n35913 ;
  assign y8766 = n35914 ;
  assign y8767 = ~n35915 ;
  assign y8768 = ~n35920 ;
  assign y8769 = n35926 ;
  assign y8770 = ~1'b0 ;
  assign y8771 = ~n35937 ;
  assign y8772 = n35942 ;
  assign y8773 = n35944 ;
  assign y8774 = ~n35949 ;
  assign y8775 = n35950 ;
  assign y8776 = n35955 ;
  assign y8777 = ~n35959 ;
  assign y8778 = ~n35961 ;
  assign y8779 = n35962 ;
  assign y8780 = n35965 ;
  assign y8781 = n35966 ;
  assign y8782 = ~n35971 ;
  assign y8783 = ~1'b0 ;
  assign y8784 = n35972 ;
  assign y8785 = ~n35975 ;
  assign y8786 = ~n35983 ;
  assign y8787 = ~n35988 ;
  assign y8788 = n35992 ;
  assign y8789 = n35993 ;
  assign y8790 = n35996 ;
  assign y8791 = ~1'b0 ;
  assign y8792 = ~n35997 ;
  assign y8793 = ~n36000 ;
  assign y8794 = ~n36006 ;
  assign y8795 = ~n36007 ;
  assign y8796 = ~n36010 ;
  assign y8797 = ~n36019 ;
  assign y8798 = n36020 ;
  assign y8799 = ~n36023 ;
  assign y8800 = ~n36025 ;
  assign y8801 = n36026 ;
  assign y8802 = n36027 ;
  assign y8803 = n36029 ;
  assign y8804 = ~1'b0 ;
  assign y8805 = ~n36032 ;
  assign y8806 = ~n36033 ;
  assign y8807 = ~n36035 ;
  assign y8808 = n36038 ;
  assign y8809 = ~n36039 ;
  assign y8810 = n36049 ;
  assign y8811 = n36051 ;
  assign y8812 = ~n36053 ;
  assign y8813 = n36065 ;
  assign y8814 = n36066 ;
  assign y8815 = ~n36067 ;
  assign y8816 = ~n36072 ;
  assign y8817 = n36073 ;
  assign y8818 = ~n36080 ;
  assign y8819 = ~1'b0 ;
  assign y8820 = n36082 ;
  assign y8821 = ~n36085 ;
  assign y8822 = n36093 ;
  assign y8823 = ~n36097 ;
  assign y8824 = n36098 ;
  assign y8825 = ~n36102 ;
  assign y8826 = ~1'b0 ;
  assign y8827 = n36105 ;
  assign y8828 = n36106 ;
  assign y8829 = n36109 ;
  assign y8830 = ~n36110 ;
  assign y8831 = n36113 ;
  assign y8832 = ~n36114 ;
  assign y8833 = ~n36119 ;
  assign y8834 = ~n36121 ;
  assign y8835 = n36122 ;
  assign y8836 = ~n36124 ;
  assign y8837 = ~n36126 ;
  assign y8838 = ~n36130 ;
  assign y8839 = ~1'b0 ;
  assign y8840 = n36132 ;
  assign y8841 = ~1'b0 ;
  assign y8842 = ~n36135 ;
  assign y8843 = n36137 ;
  assign y8844 = n36140 ;
  assign y8845 = ~n36147 ;
  assign y8846 = ~n36153 ;
  assign y8847 = ~n36159 ;
  assign y8848 = n36168 ;
  assign y8849 = n36179 ;
  assign y8850 = n36182 ;
  assign y8851 = ~n36183 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = n36186 ;
  assign y8854 = ~n36187 ;
  assign y8855 = n36194 ;
  assign y8856 = n36197 ;
  assign y8857 = n36201 ;
  assign y8858 = ~n36207 ;
  assign y8859 = ~n36208 ;
  assign y8860 = n36214 ;
  assign y8861 = n36216 ;
  assign y8862 = ~n36219 ;
  assign y8863 = ~n36223 ;
  assign y8864 = ~n36225 ;
  assign y8865 = ~n36226 ;
  assign y8866 = n36233 ;
  assign y8867 = n36240 ;
  assign y8868 = ~n36241 ;
  assign y8869 = n36245 ;
  assign y8870 = ~n36249 ;
  assign y8871 = n36251 ;
  assign y8872 = ~n36252 ;
  assign y8873 = ~n36263 ;
  assign y8874 = n36268 ;
  assign y8875 = ~n36270 ;
  assign y8876 = n36271 ;
  assign y8877 = ~1'b0 ;
  assign y8878 = n36274 ;
  assign y8879 = ~n36276 ;
  assign y8880 = n36282 ;
  assign y8881 = n36285 ;
  assign y8882 = n36290 ;
  assign y8883 = ~n36295 ;
  assign y8884 = n36297 ;
  assign y8885 = n36299 ;
  assign y8886 = ~n36301 ;
  assign y8887 = ~n36303 ;
  assign y8888 = ~n36305 ;
  assign y8889 = ~n36306 ;
  assign y8890 = ~n36308 ;
  assign y8891 = n36310 ;
  assign y8892 = n36313 ;
  assign y8893 = ~n36314 ;
  assign y8894 = ~n36319 ;
  assign y8895 = ~1'b0 ;
  assign y8896 = ~n36321 ;
  assign y8897 = ~n36322 ;
  assign y8898 = ~n36329 ;
  assign y8899 = n36334 ;
  assign y8900 = n36336 ;
  assign y8901 = ~n36338 ;
  assign y8902 = n36345 ;
  assign y8903 = ~n36348 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = n36349 ;
  assign y8906 = ~n36352 ;
  assign y8907 = n36353 ;
  assign y8908 = n36355 ;
  assign y8909 = n36361 ;
  assign y8910 = ~n36366 ;
  assign y8911 = n36369 ;
  assign y8912 = ~n36373 ;
  assign y8913 = n36375 ;
  assign y8914 = n36376 ;
  assign y8915 = n36381 ;
  assign y8916 = ~n36383 ;
  assign y8917 = ~n36385 ;
  assign y8918 = ~n36386 ;
  assign y8919 = ~1'b0 ;
  assign y8920 = n36389 ;
  assign y8921 = ~n36391 ;
  assign y8922 = n36392 ;
  assign y8923 = ~n36396 ;
  assign y8924 = n36397 ;
  assign y8925 = ~n36411 ;
  assign y8926 = ~n36418 ;
  assign y8927 = ~n36419 ;
  assign y8928 = n36422 ;
  assign y8929 = n36427 ;
  assign y8930 = n36429 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = n36433 ;
  assign y8933 = n36434 ;
  assign y8934 = n36435 ;
  assign y8935 = ~n36437 ;
  assign y8936 = n36438 ;
  assign y8937 = ~n36442 ;
  assign y8938 = n36446 ;
  assign y8939 = n36449 ;
  assign y8940 = ~n36451 ;
  assign y8941 = ~n36458 ;
  assign y8942 = n36459 ;
  assign y8943 = ~n36463 ;
  assign y8944 = ~n36465 ;
  assign y8945 = ~n36468 ;
  assign y8946 = ~n36470 ;
  assign y8947 = n36471 ;
  assign y8948 = ~n36476 ;
  assign y8949 = ~n36478 ;
  assign y8950 = ~n36482 ;
  assign y8951 = ~n36483 ;
  assign y8952 = ~n36484 ;
  assign y8953 = ~n36488 ;
  assign y8954 = ~n36489 ;
  assign y8955 = ~n36491 ;
  assign y8956 = n36492 ;
  assign y8957 = n36494 ;
  assign y8958 = ~1'b0 ;
  assign y8959 = n36496 ;
  assign y8960 = n36498 ;
  assign y8961 = n36501 ;
  assign y8962 = n36506 ;
  assign y8963 = ~1'b0 ;
  assign y8964 = ~1'b0 ;
  assign y8965 = n36509 ;
  assign y8966 = ~n36517 ;
  assign y8967 = n36518 ;
  assign y8968 = n36519 ;
  assign y8969 = n36524 ;
  assign y8970 = ~n36526 ;
  assign y8971 = ~1'b0 ;
  assign y8972 = ~n36534 ;
  assign y8973 = ~n36535 ;
  assign y8974 = n36538 ;
  assign y8975 = n36539 ;
  assign y8976 = ~1'b0 ;
  assign y8977 = ~1'b0 ;
  assign y8978 = ~n36542 ;
  assign y8979 = ~n36543 ;
  assign y8980 = ~n36544 ;
  assign y8981 = ~n36546 ;
  assign y8982 = ~n36547 ;
  assign y8983 = n36549 ;
  assign y8984 = ~n36550 ;
  assign y8985 = ~n36554 ;
  assign y8986 = n36555 ;
  assign y8987 = n36563 ;
  assign y8988 = ~n36566 ;
  assign y8989 = ~n36570 ;
  assign y8990 = ~1'b0 ;
  assign y8991 = ~n36572 ;
  assign y8992 = ~n36573 ;
  assign y8993 = n36574 ;
  assign y8994 = n36575 ;
  assign y8995 = ~n36578 ;
  assign y8996 = n36579 ;
  assign y8997 = n36581 ;
  assign y8998 = n36586 ;
  assign y8999 = n36587 ;
  assign y9000 = n36588 ;
  assign y9001 = ~n36592 ;
  assign y9002 = ~n36598 ;
  assign y9003 = ~1'b0 ;
  assign y9004 = ~1'b0 ;
  assign y9005 = ~n36602 ;
  assign y9006 = n36605 ;
  assign y9007 = ~n36610 ;
  assign y9008 = ~n36612 ;
  assign y9009 = n36615 ;
  assign y9010 = n36618 ;
  assign y9011 = n36621 ;
  assign y9012 = n36626 ;
  assign y9013 = ~n36627 ;
  assign y9014 = ~n4699 ;
  assign y9015 = n36631 ;
  assign y9016 = ~n36634 ;
  assign y9017 = n36639 ;
  assign y9018 = n36642 ;
  assign y9019 = ~n36645 ;
  assign y9020 = n36651 ;
  assign y9021 = n36652 ;
  assign y9022 = ~n36654 ;
  assign y9023 = n36659 ;
  assign y9024 = n36660 ;
  assign y9025 = ~n36663 ;
  assign y9026 = n36666 ;
  assign y9027 = ~n36667 ;
  assign y9028 = ~n36670 ;
  assign y9029 = ~n36673 ;
  assign y9030 = ~n36678 ;
  assign y9031 = ~n36680 ;
  assign y9032 = n36682 ;
  assign y9033 = ~n36684 ;
  assign y9034 = ~n36685 ;
  assign y9035 = n8382 ;
  assign y9036 = ~n36691 ;
  assign y9037 = ~n36693 ;
  assign y9038 = n36699 ;
  assign y9039 = n36701 ;
  assign y9040 = ~n36703 ;
  assign y9041 = ~n36704 ;
  assign y9042 = ~n36712 ;
  assign y9043 = ~n36716 ;
  assign y9044 = ~n36718 ;
  assign y9045 = ~1'b0 ;
  assign y9046 = n36720 ;
  assign y9047 = ~n36721 ;
  assign y9048 = n22486 ;
  assign y9049 = ~n36722 ;
  assign y9050 = n36724 ;
  assign y9051 = ~n36725 ;
  assign y9052 = n36726 ;
  assign y9053 = ~1'b0 ;
  assign y9054 = n36729 ;
  assign y9055 = ~n36736 ;
  assign y9056 = n36740 ;
  assign y9057 = ~n36742 ;
  assign y9058 = n36744 ;
  assign y9059 = ~n36747 ;
  assign y9060 = n36752 ;
  assign y9061 = ~n36753 ;
  assign y9062 = ~n36756 ;
  assign y9063 = n36757 ;
  assign y9064 = ~n36761 ;
  assign y9065 = n36768 ;
  assign y9066 = ~n36769 ;
  assign y9067 = ~n36772 ;
  assign y9068 = n36774 ;
  assign y9069 = n36776 ;
  assign y9070 = ~n36779 ;
  assign y9071 = n36780 ;
  assign y9072 = ~n36784 ;
  assign y9073 = ~n36786 ;
  assign y9074 = ~1'b0 ;
  assign y9075 = ~n36787 ;
  assign y9076 = ~n36788 ;
  assign y9077 = n36793 ;
  assign y9078 = ~n36794 ;
  assign y9079 = n36797 ;
  assign y9080 = ~n36799 ;
  assign y9081 = n36802 ;
  assign y9082 = ~n36805 ;
  assign y9083 = ~n36806 ;
  assign y9084 = n36810 ;
  assign y9085 = ~n36813 ;
  assign y9086 = n36817 ;
  assign y9087 = n36818 ;
  assign y9088 = n36825 ;
  assign y9089 = n36827 ;
  assign y9090 = n36828 ;
  assign y9091 = ~n36829 ;
  assign y9092 = n36832 ;
  assign y9093 = n36836 ;
  assign y9094 = n36839 ;
  assign y9095 = n36841 ;
  assign y9096 = ~1'b0 ;
  assign y9097 = ~n36843 ;
  assign y9098 = n36844 ;
  assign y9099 = ~n36847 ;
  assign y9100 = n36850 ;
  assign y9101 = n36857 ;
  assign y9102 = n36858 ;
  assign y9103 = ~1'b0 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = n36860 ;
  assign y9106 = ~n36861 ;
  assign y9107 = ~n36864 ;
  assign y9108 = n36866 ;
  assign y9109 = ~n36868 ;
  assign y9110 = n36871 ;
  assign y9111 = ~n36875 ;
  assign y9112 = ~1'b0 ;
  assign y9113 = ~n36879 ;
  assign y9114 = n36880 ;
  assign y9115 = n36881 ;
  assign y9116 = n36882 ;
  assign y9117 = n36898 ;
  assign y9118 = n36899 ;
  assign y9119 = ~n36904 ;
  assign y9120 = ~n36906 ;
  assign y9121 = ~n36911 ;
  assign y9122 = ~n36912 ;
  assign y9123 = ~n36913 ;
  assign y9124 = ~n36914 ;
  assign y9125 = ~n36915 ;
  assign y9126 = ~n36917 ;
  assign y9127 = ~n36920 ;
  assign y9128 = n36922 ;
  assign y9129 = n36925 ;
  assign y9130 = ~n36928 ;
  assign y9131 = n36929 ;
  assign y9132 = n36932 ;
  assign y9133 = ~n36936 ;
  assign y9134 = ~n36941 ;
  assign y9135 = ~n36947 ;
  assign y9136 = n36949 ;
  assign y9137 = n36951 ;
  assign y9138 = ~n36956 ;
  assign y9139 = ~n36961 ;
  assign y9140 = ~n36967 ;
  assign y9141 = ~n36973 ;
  assign y9142 = ~n36977 ;
  assign y9143 = n36980 ;
  assign y9144 = n36985 ;
  assign y9145 = n36986 ;
  assign y9146 = n36988 ;
  assign y9147 = n36993 ;
  assign y9148 = n37002 ;
  assign y9149 = n37008 ;
  assign y9150 = ~n37010 ;
  assign y9151 = ~n37012 ;
  assign y9152 = n37016 ;
  assign y9153 = n37021 ;
  assign y9154 = ~1'b0 ;
  assign y9155 = n37023 ;
  assign y9156 = ~n37030 ;
  assign y9157 = n37032 ;
  assign y9158 = ~n37036 ;
  assign y9159 = ~n37045 ;
  assign y9160 = ~n37049 ;
  assign y9161 = n37054 ;
  assign y9162 = ~n37057 ;
  assign y9163 = n37061 ;
  assign y9164 = n37062 ;
  assign y9165 = ~n37064 ;
  assign y9166 = n37065 ;
  assign y9167 = ~n37072 ;
  assign y9168 = ~n37074 ;
  assign y9169 = n37078 ;
  assign y9170 = n37080 ;
  assign y9171 = n37083 ;
  assign y9172 = ~n37087 ;
  assign y9173 = ~n37091 ;
  assign y9174 = n37092 ;
  assign y9175 = ~n37094 ;
  assign y9176 = n37096 ;
  assign y9177 = n37097 ;
  assign y9178 = ~n37099 ;
  assign y9179 = ~1'b0 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = n37109 ;
  assign y9182 = ~n37111 ;
  assign y9183 = ~n37116 ;
  assign y9184 = n37120 ;
  assign y9185 = ~n37121 ;
  assign y9186 = ~n37124 ;
  assign y9187 = ~1'b0 ;
  assign y9188 = n37125 ;
  assign y9189 = n37127 ;
  assign y9190 = ~n37128 ;
  assign y9191 = n37136 ;
  assign y9192 = ~n37139 ;
  assign y9193 = n37147 ;
  assign y9194 = n37150 ;
  assign y9195 = n37152 ;
  assign y9196 = n37158 ;
  assign y9197 = ~1'b0 ;
  assign y9198 = ~n37161 ;
  assign y9199 = ~n37163 ;
  assign y9200 = ~n37166 ;
  assign y9201 = n37170 ;
  assign y9202 = n37180 ;
  assign y9203 = ~n37182 ;
  assign y9204 = ~n37183 ;
  assign y9205 = ~n37187 ;
  assign y9206 = ~n37191 ;
  assign y9207 = n37192 ;
  assign y9208 = ~n37193 ;
  assign y9209 = n37194 ;
  assign y9210 = ~n37196 ;
  assign y9211 = n37198 ;
  assign y9212 = n37200 ;
  assign y9213 = n37209 ;
  assign y9214 = ~n37210 ;
  assign y9215 = ~n37213 ;
  assign y9216 = ~n37214 ;
  assign y9217 = ~1'b0 ;
  assign y9218 = ~n37220 ;
  assign y9219 = ~n37224 ;
  assign y9220 = ~n37228 ;
  assign y9221 = n37230 ;
  assign y9222 = n37232 ;
  assign y9223 = ~n37248 ;
  assign y9224 = ~n37255 ;
  assign y9225 = n37257 ;
  assign y9226 = ~n37258 ;
  assign y9227 = ~n37259 ;
  assign y9228 = n37261 ;
  assign y9229 = ~n37266 ;
  assign y9230 = n37271 ;
  assign y9231 = n37272 ;
  assign y9232 = ~n37277 ;
  assign y9233 = n37278 ;
  assign y9234 = n37279 ;
  assign y9235 = ~n37280 ;
  assign y9236 = ~n37284 ;
  assign y9237 = n37285 ;
  assign y9238 = ~n37286 ;
  assign y9239 = n37287 ;
  assign y9240 = n37289 ;
  assign y9241 = ~n37291 ;
  assign y9242 = ~n37294 ;
  assign y9243 = ~n37295 ;
  assign y9244 = n37296 ;
  assign y9245 = n37299 ;
  assign y9246 = n37304 ;
  assign y9247 = n37310 ;
  assign y9248 = ~n37312 ;
  assign y9249 = n37313 ;
  assign y9250 = n37314 ;
  assign y9251 = ~1'b0 ;
  assign y9252 = ~1'b0 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = n37316 ;
  assign y9255 = ~n37322 ;
  assign y9256 = n37327 ;
  assign y9257 = ~n37330 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = n37332 ;
  assign y9260 = ~n37339 ;
  assign y9261 = n37342 ;
  assign y9262 = n37344 ;
  assign y9263 = n37345 ;
  assign y9264 = ~n37347 ;
  assign y9265 = n37348 ;
  assign y9266 = ~n37359 ;
  assign y9267 = ~n37363 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = n37365 ;
  assign y9270 = ~n37366 ;
  assign y9271 = n37370 ;
  assign y9272 = ~n37373 ;
  assign y9273 = ~n37376 ;
  assign y9274 = n37377 ;
  assign y9275 = ~1'b0 ;
  assign y9276 = n37379 ;
  assign y9277 = n37383 ;
  assign y9278 = ~n37385 ;
  assign y9279 = n37387 ;
  assign y9280 = ~1'b0 ;
  assign y9281 = ~n37392 ;
  assign y9282 = n37394 ;
  assign y9283 = n37398 ;
  assign y9284 = n37399 ;
  assign y9285 = ~n37404 ;
  assign y9286 = ~n37409 ;
  assign y9287 = ~n37410 ;
  assign y9288 = n37412 ;
  assign y9289 = n37414 ;
  assign y9290 = n37417 ;
  assign y9291 = n37424 ;
  assign y9292 = ~n37426 ;
  assign y9293 = ~n37434 ;
  assign y9294 = n37436 ;
  assign y9295 = n37445 ;
  assign y9296 = ~n37447 ;
  assign y9297 = n37448 ;
  assign y9298 = ~n37452 ;
  assign y9299 = ~n37457 ;
  assign y9300 = n37464 ;
  assign y9301 = ~n37469 ;
  assign y9302 = n37471 ;
  assign y9303 = ~n37475 ;
  assign y9304 = n37476 ;
  assign y9305 = ~n37479 ;
  assign y9306 = n37481 ;
  assign y9307 = ~n37482 ;
  assign y9308 = ~n37486 ;
  assign y9309 = n37488 ;
  assign y9310 = n37492 ;
  assign y9311 = ~1'b0 ;
  assign y9312 = n37495 ;
  assign y9313 = n37501 ;
  assign y9314 = ~n37505 ;
  assign y9315 = n37507 ;
  assign y9316 = ~n37509 ;
  assign y9317 = ~n37510 ;
  assign y9318 = n37514 ;
  assign y9319 = n37516 ;
  assign y9320 = ~n37517 ;
  assign y9321 = n37525 ;
  assign y9322 = ~n37526 ;
  assign y9323 = ~n37530 ;
  assign y9324 = ~n37534 ;
  assign y9325 = ~n37540 ;
  assign y9326 = n37544 ;
  assign y9327 = n37551 ;
  assign y9328 = n37554 ;
  assign y9329 = ~n37560 ;
  assign y9330 = ~n37564 ;
  assign y9331 = n37571 ;
  assign y9332 = ~n37572 ;
  assign y9333 = n37579 ;
  assign y9334 = n37582 ;
  assign y9335 = ~1'b0 ;
  assign y9336 = ~n37583 ;
  assign y9337 = n37585 ;
  assign y9338 = n37590 ;
  assign y9339 = n37591 ;
  assign y9340 = ~n37593 ;
  assign y9341 = n37598 ;
  assign y9342 = ~n37599 ;
  assign y9343 = n37602 ;
  assign y9344 = ~n37604 ;
  assign y9345 = ~n37605 ;
  assign y9346 = n37607 ;
  assign y9347 = ~1'b0 ;
  assign y9348 = ~n37613 ;
  assign y9349 = ~n37614 ;
  assign y9350 = ~n37618 ;
  assign y9351 = n37620 ;
  assign y9352 = ~n37623 ;
  assign y9353 = n37629 ;
  assign y9354 = ~n37632 ;
  assign y9355 = n37633 ;
  assign y9356 = n37634 ;
  assign y9357 = ~n37641 ;
  assign y9358 = ~n37644 ;
  assign y9359 = ~n37645 ;
  assign y9360 = n37649 ;
  assign y9361 = ~n37650 ;
  assign y9362 = n37651 ;
  assign y9363 = ~n37652 ;
  assign y9364 = ~n37654 ;
  assign y9365 = ~n37655 ;
  assign y9366 = n37656 ;
  assign y9367 = ~n37663 ;
  assign y9368 = ~n37664 ;
  assign y9369 = n37671 ;
  assign y9370 = ~n37673 ;
  assign y9371 = n37676 ;
  assign y9372 = ~n37680 ;
  assign y9373 = ~n37682 ;
  assign y9374 = ~n37685 ;
  assign y9375 = n37688 ;
  assign y9376 = n37695 ;
  assign y9377 = n37696 ;
  assign y9378 = ~n37699 ;
  assign y9379 = ~1'b0 ;
  assign y9380 = ~n37701 ;
  assign y9381 = ~n37702 ;
  assign y9382 = n37703 ;
  assign y9383 = ~n37706 ;
  assign y9384 = n37708 ;
  assign y9385 = n37711 ;
  assign y9386 = ~n37712 ;
  assign y9387 = n37719 ;
  assign y9388 = ~1'b0 ;
  assign y9389 = n37724 ;
  assign y9390 = ~n37728 ;
  assign y9391 = ~n37730 ;
  assign y9392 = n37731 ;
  assign y9393 = n37733 ;
  assign y9394 = n37735 ;
  assign y9395 = ~n37738 ;
  assign y9396 = n37739 ;
  assign y9397 = n37740 ;
  assign y9398 = ~n37741 ;
  assign y9399 = ~n37742 ;
  assign y9400 = n37743 ;
  assign y9401 = n37745 ;
  assign y9402 = n37750 ;
  assign y9403 = ~1'b0 ;
  assign y9404 = ~1'b0 ;
  assign y9405 = ~n37751 ;
  assign y9406 = ~n37758 ;
  assign y9407 = ~n37765 ;
  assign y9408 = n37771 ;
  assign y9409 = ~n37775 ;
  assign y9410 = n37777 ;
  assign y9411 = n37779 ;
  assign y9412 = ~n37785 ;
  assign y9413 = n37786 ;
  assign y9414 = ~n37789 ;
  assign y9415 = n37791 ;
  assign y9416 = n37799 ;
  assign y9417 = ~n37803 ;
  assign y9418 = n37805 ;
  assign y9419 = ~1'b0 ;
  assign y9420 = ~n37807 ;
  assign y9421 = ~n37811 ;
  assign y9422 = n37813 ;
  assign y9423 = ~n37815 ;
  assign y9424 = ~n37819 ;
  assign y9425 = ~n37822 ;
  assign y9426 = ~n37825 ;
  assign y9427 = ~n37826 ;
  assign y9428 = n37828 ;
  assign y9429 = ~n37831 ;
  assign y9430 = n37834 ;
  assign y9431 = n37835 ;
  assign y9432 = n37837 ;
  assign y9433 = n37839 ;
  assign y9434 = ~1'b0 ;
  assign y9435 = ~1'b0 ;
  assign y9436 = ~n37841 ;
  assign y9437 = ~n37842 ;
  assign y9438 = n37844 ;
  assign y9439 = ~n37849 ;
  assign y9440 = ~n37852 ;
  assign y9441 = ~n37853 ;
  assign y9442 = n37857 ;
  assign y9443 = n37860 ;
  assign y9444 = n37866 ;
  assign y9445 = ~1'b0 ;
  assign y9446 = n37868 ;
  assign y9447 = n37874 ;
  assign y9448 = n37879 ;
  assign y9449 = ~n37881 ;
  assign y9450 = n37884 ;
  assign y9451 = ~1'b0 ;
  assign y9452 = ~n37887 ;
  assign y9453 = ~n37893 ;
  assign y9454 = n37896 ;
  assign y9455 = n37897 ;
  assign y9456 = ~n37902 ;
  assign y9457 = ~n37906 ;
  assign y9458 = n37909 ;
  assign y9459 = n37916 ;
  assign y9460 = ~n37919 ;
  assign y9461 = n37921 ;
  assign y9462 = ~n37927 ;
  assign y9463 = ~n37929 ;
  assign y9464 = ~n37932 ;
  assign y9465 = ~n37935 ;
  assign y9466 = ~n37943 ;
  assign y9467 = n37944 ;
  assign y9468 = ~n37945 ;
  assign y9469 = ~n37946 ;
  assign y9470 = ~1'b0 ;
  assign y9471 = ~n37949 ;
  assign y9472 = n37954 ;
  assign y9473 = ~n37959 ;
  assign y9474 = ~n37960 ;
  assign y9475 = ~n37963 ;
  assign y9476 = ~n37966 ;
  assign y9477 = ~n37968 ;
  assign y9478 = ~n37974 ;
  assign y9479 = n37980 ;
  assign y9480 = ~n37981 ;
  assign y9481 = n37984 ;
  assign y9482 = ~n37989 ;
  assign y9483 = n37995 ;
  assign y9484 = n37996 ;
  assign y9485 = n38004 ;
  assign y9486 = ~n38006 ;
  assign y9487 = n38009 ;
  assign y9488 = ~n38010 ;
  assign y9489 = ~n38012 ;
  assign y9490 = ~n38015 ;
  assign y9491 = n38018 ;
  assign y9492 = ~n38019 ;
  assign y9493 = n38021 ;
  assign y9494 = n38026 ;
  assign y9495 = n38027 ;
  assign y9496 = n38029 ;
  assign y9497 = ~n38030 ;
  assign y9498 = ~n38034 ;
  assign y9499 = ~n38035 ;
  assign y9500 = n38041 ;
  assign y9501 = ~n38043 ;
  assign y9502 = n38044 ;
  assign y9503 = ~n38045 ;
  assign y9504 = n38047 ;
  assign y9505 = n38051 ;
  assign y9506 = ~1'b0 ;
  assign y9507 = n38057 ;
  assign y9508 = n38059 ;
  assign y9509 = ~n38060 ;
  assign y9510 = n38061 ;
  assign y9511 = ~n38062 ;
  assign y9512 = ~1'b0 ;
  assign y9513 = ~n38064 ;
  assign y9514 = n38065 ;
  assign y9515 = ~n38066 ;
  assign y9516 = ~n38069 ;
  assign y9517 = n38073 ;
  assign y9518 = n38075 ;
  assign y9519 = n38080 ;
  assign y9520 = ~n1865 ;
  assign y9521 = n38083 ;
  assign y9522 = ~n38085 ;
  assign y9523 = ~n38086 ;
  assign y9524 = ~n38091 ;
  assign y9525 = ~n38094 ;
  assign y9526 = n38095 ;
  assign y9527 = ~n38096 ;
  assign y9528 = ~n38098 ;
  assign y9529 = n38100 ;
  assign y9530 = ~n38102 ;
  assign y9531 = n38103 ;
  assign y9532 = ~n38104 ;
  assign y9533 = ~n38108 ;
  assign y9534 = ~n38115 ;
  assign y9535 = ~1'b0 ;
  assign y9536 = ~n38116 ;
  assign y9537 = ~n38118 ;
  assign y9538 = ~n38121 ;
  assign y9539 = n38126 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = n38128 ;
  assign y9542 = ~n38133 ;
  assign y9543 = n38135 ;
  assign y9544 = n38136 ;
  assign y9545 = n38137 ;
  assign y9546 = ~1'b0 ;
  assign y9547 = n38140 ;
  assign y9548 = n38142 ;
  assign y9549 = ~n38144 ;
  assign y9550 = ~n38146 ;
  assign y9551 = ~n38149 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = ~1'b0 ;
  assign y9554 = ~n38151 ;
  assign y9555 = ~n38154 ;
  assign y9556 = n38155 ;
  assign y9557 = ~n38158 ;
  assign y9558 = ~n38163 ;
  assign y9559 = ~n38165 ;
  assign y9560 = ~1'b0 ;
  assign y9561 = n38167 ;
  assign y9562 = n38168 ;
  assign y9563 = ~n38171 ;
  assign y9564 = ~n38172 ;
  assign y9565 = ~n38174 ;
  assign y9566 = ~n38180 ;
  assign y9567 = n38184 ;
  assign y9568 = n38187 ;
  assign y9569 = n38189 ;
  assign y9570 = n38190 ;
  assign y9571 = n38193 ;
  assign y9572 = n38194 ;
  assign y9573 = ~n38196 ;
  assign y9574 = n38200 ;
  assign y9575 = n38201 ;
  assign y9576 = n38202 ;
  assign y9577 = n38203 ;
  assign y9578 = n38206 ;
  assign y9579 = n38207 ;
  assign y9580 = ~n37089 ;
  assign y9581 = ~n38209 ;
  assign y9582 = n38217 ;
  assign y9583 = ~1'b0 ;
  assign y9584 = ~1'b0 ;
  assign y9585 = ~n607 ;
  assign y9586 = ~n38220 ;
  assign y9587 = n38221 ;
  assign y9588 = n38222 ;
  assign y9589 = ~1'b0 ;
  assign y9590 = n38228 ;
  assign y9591 = n38232 ;
  assign y9592 = n38234 ;
  assign y9593 = ~n38235 ;
  assign y9594 = ~n38241 ;
  assign y9595 = ~n38244 ;
  assign y9596 = 1'b0 ;
  assign y9597 = ~n38249 ;
  assign y9598 = ~1'b0 ;
  assign y9599 = ~n38250 ;
  assign y9600 = ~n38251 ;
  assign y9601 = n38255 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = ~n38257 ;
  assign y9604 = ~n38262 ;
  assign y9605 = n38265 ;
  assign y9606 = ~n38271 ;
  assign y9607 = ~n38272 ;
  assign y9608 = n38275 ;
  assign y9609 = n38276 ;
  assign y9610 = ~n38282 ;
  assign y9611 = n38284 ;
  assign y9612 = n38286 ;
  assign y9613 = n38290 ;
  assign y9614 = ~n38291 ;
  assign y9615 = n38293 ;
  assign y9616 = n38297 ;
  assign y9617 = n38302 ;
  assign y9618 = ~n38303 ;
  assign y9619 = ~n38304 ;
  assign y9620 = n38310 ;
  assign y9621 = ~n38315 ;
  assign y9622 = n38317 ;
  assign y9623 = n38322 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = ~n38325 ;
  assign y9626 = ~n38326 ;
  assign y9627 = ~n38328 ;
  assign y9628 = n38330 ;
  assign y9629 = n38332 ;
  assign y9630 = n38335 ;
  assign y9631 = ~n38337 ;
  assign y9632 = n38339 ;
  assign y9633 = ~n38340 ;
  assign y9634 = n38347 ;
  assign y9635 = ~n38348 ;
  assign y9636 = ~n38353 ;
  assign y9637 = n38354 ;
  assign y9638 = ~n38357 ;
  assign y9639 = n38359 ;
  assign y9640 = n38362 ;
  assign y9641 = ~n38364 ;
  assign y9642 = ~n38368 ;
  assign y9643 = ~n38373 ;
  assign y9644 = n38376 ;
  assign y9645 = n38379 ;
  assign y9646 = ~n38381 ;
  assign y9647 = n38384 ;
  assign y9648 = ~1'b0 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = n38388 ;
  assign y9651 = n38389 ;
  assign y9652 = n38392 ;
  assign y9653 = ~n38395 ;
  assign y9654 = n38399 ;
  assign y9655 = n38406 ;
  assign y9656 = n38408 ;
  assign y9657 = n38409 ;
  assign y9658 = ~n38419 ;
  assign y9659 = ~n38421 ;
  assign y9660 = n38425 ;
  assign y9661 = ~n38428 ;
  assign y9662 = ~1'b0 ;
  assign y9663 = ~n38433 ;
  assign y9664 = n38435 ;
  assign y9665 = ~n38440 ;
  assign y9666 = ~n38441 ;
  assign y9667 = n38446 ;
  assign y9668 = n38447 ;
  assign y9669 = ~n38448 ;
  assign y9670 = ~n38449 ;
  assign y9671 = n38452 ;
  assign y9672 = ~n38454 ;
  assign y9673 = ~n38456 ;
  assign y9674 = ~n38459 ;
  assign y9675 = n38464 ;
  assign y9676 = n38467 ;
  assign y9677 = n38475 ;
  assign y9678 = ~n38476 ;
  assign y9679 = ~n38478 ;
  assign y9680 = n38480 ;
  assign y9681 = ~n38482 ;
  assign y9682 = ~n38485 ;
  assign y9683 = n38486 ;
  assign y9684 = n38487 ;
  assign y9685 = n38489 ;
  assign y9686 = ~n38491 ;
  assign y9687 = ~1'b0 ;
  assign y9688 = n38493 ;
  assign y9689 = ~n38496 ;
  assign y9690 = ~n38498 ;
  assign y9691 = ~n38501 ;
  assign y9692 = n38504 ;
  assign y9693 = ~n38507 ;
  assign y9694 = ~n38508 ;
  assign y9695 = n38509 ;
  assign y9696 = n38515 ;
  assign y9697 = ~n38521 ;
  assign y9698 = n38523 ;
  assign y9699 = n38529 ;
  assign y9700 = n38532 ;
  assign y9701 = ~n38536 ;
  assign y9702 = ~n38540 ;
  assign y9703 = ~n38548 ;
  assign y9704 = n38551 ;
  assign y9705 = n38556 ;
  assign y9706 = n38567 ;
  assign y9707 = n38569 ;
  assign y9708 = n38570 ;
  assign y9709 = n38571 ;
  assign y9710 = n38573 ;
  assign y9711 = ~n38574 ;
  assign y9712 = ~n38575 ;
  assign y9713 = n38576 ;
  assign y9714 = n38577 ;
  assign y9715 = ~n38582 ;
  assign y9716 = n38585 ;
  assign y9717 = n38587 ;
  assign y9718 = ~n38592 ;
  assign y9719 = ~n38596 ;
  assign y9720 = ~n38605 ;
  assign y9721 = ~n38607 ;
  assign y9722 = ~n38609 ;
  assign y9723 = n38610 ;
  assign y9724 = n38617 ;
  assign y9725 = n38618 ;
  assign y9726 = ~n38620 ;
  assign y9727 = ~1'b0 ;
  assign y9728 = n38621 ;
  assign y9729 = n38623 ;
  assign y9730 = n38628 ;
  assign y9731 = ~n38629 ;
  assign y9732 = n38635 ;
  assign y9733 = n38638 ;
  assign y9734 = ~n38646 ;
  assign y9735 = ~n38648 ;
  assign y9736 = n38652 ;
  assign y9737 = ~n38661 ;
  assign y9738 = ~n38662 ;
  assign y9739 = n38664 ;
  assign y9740 = n38665 ;
  assign y9741 = ~n38675 ;
  assign y9742 = ~n38677 ;
  assign y9743 = n38682 ;
  assign y9744 = ~n38683 ;
  assign y9745 = ~n38684 ;
  assign y9746 = ~n38685 ;
  assign y9747 = ~n38688 ;
  assign y9748 = ~1'b0 ;
  assign y9749 = n38690 ;
  assign y9750 = n38693 ;
  assign y9751 = n38695 ;
  assign y9752 = ~n38697 ;
  assign y9753 = ~n38698 ;
  assign y9754 = n38700 ;
  assign y9755 = ~n38702 ;
  assign y9756 = n38704 ;
  assign y9757 = ~n38710 ;
  assign y9758 = n38712 ;
  assign y9759 = ~n38714 ;
  assign y9760 = ~n38721 ;
  assign y9761 = n38726 ;
  assign y9762 = n38727 ;
  assign y9763 = n38728 ;
  assign y9764 = ~n38733 ;
  assign y9765 = n38739 ;
  assign y9766 = n38741 ;
  assign y9767 = n38746 ;
  assign y9768 = n38747 ;
  assign y9769 = ~1'b0 ;
  assign y9770 = ~n38751 ;
  assign y9771 = n38755 ;
  assign y9772 = ~n38761 ;
  assign y9773 = n38765 ;
  assign y9774 = n38768 ;
  assign y9775 = ~n38774 ;
  assign y9776 = n38776 ;
  assign y9777 = ~n38780 ;
  assign y9778 = n38781 ;
  assign y9779 = n38783 ;
  assign y9780 = ~n38784 ;
  assign y9781 = ~n38785 ;
  assign y9782 = ~n38790 ;
  assign y9783 = n38792 ;
  assign y9784 = ~n38799 ;
  assign y9785 = n38804 ;
  assign y9786 = n38807 ;
  assign y9787 = ~n38812 ;
  assign y9788 = ~n38816 ;
  assign y9789 = n38817 ;
  assign y9790 = n38818 ;
  assign y9791 = n38820 ;
  assign y9792 = n38821 ;
  assign y9793 = ~n11925 ;
  assign y9794 = n38825 ;
  assign y9795 = n38826 ;
  assign y9796 = n38827 ;
  assign y9797 = ~n38829 ;
  assign y9798 = n38830 ;
  assign y9799 = n12760 ;
  assign y9800 = n38833 ;
  assign y9801 = ~n38835 ;
  assign y9802 = ~1'b0 ;
  assign y9803 = ~n38837 ;
  assign y9804 = n38838 ;
  assign y9805 = ~n38842 ;
  assign y9806 = ~n38845 ;
  assign y9807 = n38846 ;
  assign y9808 = n38849 ;
  assign y9809 = n38851 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~n38856 ;
  assign y9812 = n38858 ;
  assign y9813 = n38859 ;
  assign y9814 = ~n38863 ;
  assign y9815 = ~n38864 ;
  assign y9816 = n38866 ;
  assign y9817 = n38868 ;
  assign y9818 = ~n38869 ;
  assign y9819 = ~n38870 ;
  assign y9820 = n38885 ;
  assign y9821 = ~n38889 ;
  assign y9822 = n38891 ;
  assign y9823 = ~n38892 ;
  assign y9824 = n38895 ;
  assign y9825 = ~n38896 ;
  assign y9826 = ~n38900 ;
  assign y9827 = ~n38911 ;
  assign y9828 = ~1'b0 ;
  assign y9829 = ~n38912 ;
  assign y9830 = n38915 ;
  assign y9831 = ~n38919 ;
  assign y9832 = ~n38920 ;
  assign y9833 = ~1'b0 ;
  assign y9834 = ~1'b0 ;
  assign y9835 = n38922 ;
  assign y9836 = n38924 ;
  assign y9837 = ~n38925 ;
  assign y9838 = ~n38926 ;
  assign y9839 = ~n38927 ;
  assign y9840 = n38934 ;
  assign y9841 = n38936 ;
  assign y9842 = ~1'b0 ;
  assign y9843 = ~1'b0 ;
  assign y9844 = ~n38939 ;
  assign y9845 = ~n38940 ;
  assign y9846 = ~n38941 ;
  assign y9847 = ~n38949 ;
  assign y9848 = n38950 ;
  assign y9849 = ~n38953 ;
  assign y9850 = ~n38956 ;
  assign y9851 = ~n38959 ;
  assign y9852 = n38961 ;
  assign y9853 = n38963 ;
  assign y9854 = n38969 ;
  assign y9855 = n38976 ;
  assign y9856 = ~n38977 ;
  assign y9857 = ~n38980 ;
  assign y9858 = n38984 ;
  assign y9859 = n38988 ;
  assign y9860 = ~n38989 ;
  assign y9861 = ~n38992 ;
  assign y9862 = ~n38996 ;
  assign y9863 = n38997 ;
  assign y9864 = ~n38999 ;
  assign y9865 = n39000 ;
  assign y9866 = ~n39001 ;
  assign y9867 = ~n39004 ;
  assign y9868 = n39007 ;
  assign y9869 = ~n39009 ;
  assign y9870 = ~n39011 ;
  assign y9871 = ~n39013 ;
  assign y9872 = ~n39014 ;
  assign y9873 = n39019 ;
  assign y9874 = n39020 ;
  assign y9875 = ~n39026 ;
  assign y9876 = ~1'b0 ;
  assign y9877 = ~n39030 ;
  assign y9878 = n39034 ;
  assign y9879 = ~n39040 ;
  assign y9880 = ~n39044 ;
  assign y9881 = n39045 ;
  assign y9882 = ~n39047 ;
  assign y9883 = ~n39049 ;
  assign y9884 = n39056 ;
  assign y9885 = n39058 ;
  assign y9886 = n39061 ;
  assign y9887 = n39065 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = ~n39069 ;
  assign y9890 = n39078 ;
  assign y9891 = ~n39087 ;
  assign y9892 = ~n39088 ;
  assign y9893 = n39090 ;
  assign y9894 = ~n39093 ;
  assign y9895 = ~n39096 ;
  assign y9896 = n39105 ;
  assign y9897 = n39106 ;
  assign y9898 = ~n39108 ;
  assign y9899 = ~n39114 ;
  assign y9900 = ~n39118 ;
  assign y9901 = ~n39126 ;
  assign y9902 = ~n39127 ;
  assign y9903 = n39128 ;
  assign y9904 = ~n39132 ;
  assign y9905 = ~n39134 ;
  assign y9906 = n39139 ;
  assign y9907 = n39140 ;
  assign y9908 = n39142 ;
  assign y9909 = n39143 ;
  assign y9910 = ~n39146 ;
  assign y9911 = ~n39150 ;
  assign y9912 = n39152 ;
  assign y9913 = ~n39156 ;
  assign y9914 = ~n39158 ;
  assign y9915 = n39159 ;
  assign y9916 = n39169 ;
  assign y9917 = ~n39172 ;
  assign y9918 = n39174 ;
  assign y9919 = n39175 ;
  assign y9920 = ~n39178 ;
  assign y9921 = ~n39182 ;
  assign y9922 = n39184 ;
  assign y9923 = ~n39188 ;
  assign y9924 = n39197 ;
  assign y9925 = ~1'b0 ;
  assign y9926 = ~n39203 ;
  assign y9927 = ~n39204 ;
  assign y9928 = ~n39205 ;
  assign y9929 = n39206 ;
  assign y9930 = ~n39208 ;
  assign y9931 = n39217 ;
  assign y9932 = ~n39220 ;
  assign y9933 = ~n39221 ;
  assign y9934 = n39222 ;
  assign y9935 = n39230 ;
  assign y9936 = n39233 ;
  assign y9937 = ~n39236 ;
  assign y9938 = n39243 ;
  assign y9939 = n39244 ;
  assign y9940 = ~n39251 ;
  assign y9941 = ~n39252 ;
  assign y9942 = ~1'b0 ;
  assign y9943 = n39256 ;
  assign y9944 = n8065 ;
  assign y9945 = ~n39257 ;
  assign y9946 = n39258 ;
  assign y9947 = n39263 ;
  assign y9948 = n39268 ;
  assign y9949 = n39269 ;
  assign y9950 = n39274 ;
  assign y9951 = n39276 ;
  assign y9952 = ~1'b0 ;
  assign y9953 = ~1'b0 ;
  assign y9954 = ~n39277 ;
  assign y9955 = ~n39280 ;
  assign y9956 = n39283 ;
  assign y9957 = ~n39292 ;
  assign y9958 = n39298 ;
  assign y9959 = ~n39300 ;
  assign y9960 = n39302 ;
  assign y9961 = ~n39305 ;
  assign y9962 = ~n39310 ;
  assign y9963 = n39312 ;
  assign y9964 = n39316 ;
  assign y9965 = n39318 ;
  assign y9966 = ~n39321 ;
  assign y9967 = ~1'b0 ;
  assign y9968 = n39326 ;
  assign y9969 = n39329 ;
  assign y9970 = n39330 ;
  assign y9971 = n39331 ;
  assign y9972 = ~n39332 ;
  assign y9973 = n39339 ;
  assign y9974 = ~n39342 ;
  assign y9975 = n39345 ;
  assign y9976 = n39347 ;
  assign y9977 = ~n39351 ;
  assign y9978 = ~1'b0 ;
  assign y9979 = ~n39352 ;
  assign y9980 = n39361 ;
  assign y9981 = n39363 ;
  assign y9982 = ~n39365 ;
  assign y9983 = n39367 ;
  assign y9984 = n39369 ;
  assign y9985 = ~n39372 ;
  assign y9986 = n39378 ;
  assign y9987 = ~n39380 ;
  assign y9988 = ~n39384 ;
  assign y9989 = n39390 ;
  assign y9990 = ~n39395 ;
  assign y9991 = ~n39396 ;
  assign y9992 = ~n39398 ;
  assign y9993 = n39399 ;
  assign y9994 = ~n39400 ;
  assign y9995 = ~n39401 ;
  assign y9996 = ~1'b0 ;
  assign y9997 = n39402 ;
  assign y9998 = ~n39407 ;
  assign y9999 = n39409 ;
  assign y10000 = ~n39412 ;
  assign y10001 = n39415 ;
  assign y10002 = ~n39419 ;
  assign y10003 = n39420 ;
  assign y10004 = n39424 ;
  assign y10005 = ~n39433 ;
  assign y10006 = n39434 ;
  assign y10007 = n39435 ;
  assign y10008 = n39437 ;
  assign y10009 = ~n39439 ;
  assign y10010 = n39440 ;
  assign y10011 = n39443 ;
  assign y10012 = n39444 ;
  assign y10013 = ~n39445 ;
  assign y10014 = ~n39450 ;
  assign y10015 = n39452 ;
  assign y10016 = ~n39453 ;
  assign y10017 = ~n39456 ;
  assign y10018 = n39462 ;
  assign y10019 = ~n39469 ;
  assign y10020 = ~n39470 ;
  assign y10021 = n39474 ;
  assign y10022 = n35344 ;
  assign y10023 = ~1'b0 ;
  assign y10024 = ~n39475 ;
  assign y10025 = n39480 ;
  assign y10026 = ~n39481 ;
  assign y10027 = ~n39484 ;
  assign y10028 = n39485 ;
  assign y10029 = ~n39495 ;
  assign y10030 = ~n39497 ;
  assign y10031 = n39499 ;
  assign y10032 = n39500 ;
  assign y10033 = ~n39503 ;
  assign y10034 = n39507 ;
  assign y10035 = ~n39509 ;
  assign y10036 = ~1'b0 ;
  assign y10037 = n39512 ;
  assign y10038 = ~n39515 ;
  assign y10039 = ~n39516 ;
  assign y10040 = ~n39517 ;
  assign y10041 = ~n39518 ;
  assign y10042 = n39521 ;
  assign y10043 = ~n39523 ;
  assign y10044 = n39525 ;
  assign y10045 = n39529 ;
  assign y10046 = ~n39534 ;
  assign y10047 = n39535 ;
  assign y10048 = n39537 ;
  assign y10049 = ~n39539 ;
  assign y10050 = ~n39542 ;
  assign y10051 = n39546 ;
  assign y10052 = n39547 ;
  assign y10053 = n39548 ;
  assign y10054 = ~n39554 ;
  assign y10055 = ~n39557 ;
  assign y10056 = ~n39558 ;
  assign y10057 = ~n39559 ;
  assign y10058 = ~1'b0 ;
  assign y10059 = ~n39564 ;
  assign y10060 = n39568 ;
  assign y10061 = ~n39572 ;
  assign y10062 = n39574 ;
  assign y10063 = n39575 ;
  assign y10064 = n39576 ;
  assign y10065 = ~n39579 ;
  assign y10066 = n39585 ;
  assign y10067 = n39591 ;
  assign y10068 = ~n39595 ;
  assign y10069 = ~n39596 ;
  assign y10070 = ~n39599 ;
  assign y10071 = n39601 ;
  assign y10072 = ~n39603 ;
  assign y10073 = ~n39606 ;
  assign y10074 = n39607 ;
  assign y10075 = n39611 ;
  assign y10076 = ~n39612 ;
  assign y10077 = n39617 ;
  assign y10078 = ~n39619 ;
  assign y10079 = ~n39621 ;
  assign y10080 = n39622 ;
  assign y10081 = n39627 ;
  assign y10082 = ~n39632 ;
  assign y10083 = ~n39634 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = ~n39637 ;
  assign y10086 = ~n39639 ;
  assign y10087 = ~n39640 ;
  assign y10088 = ~n39646 ;
  assign y10089 = ~n39647 ;
  assign y10090 = n39651 ;
  assign y10091 = ~n39657 ;
  assign y10092 = ~n39658 ;
  assign y10093 = n39660 ;
  assign y10094 = n39662 ;
  assign y10095 = n39663 ;
  assign y10096 = n39667 ;
  assign y10097 = ~n39668 ;
  assign y10098 = ~n39671 ;
  assign y10099 = ~1'b0 ;
  assign y10100 = n39678 ;
  assign y10101 = ~n39680 ;
  assign y10102 = n39681 ;
  assign y10103 = ~1'b0 ;
  assign y10104 = n39682 ;
  assign y10105 = ~n39686 ;
  assign y10106 = ~n39689 ;
  assign y10107 = ~n39693 ;
  assign y10108 = n39694 ;
  assign y10109 = n39695 ;
  assign y10110 = n39697 ;
  assign y10111 = ~n39698 ;
  assign y10112 = n39702 ;
  assign y10113 = ~n39703 ;
  assign y10114 = n39706 ;
  assign y10115 = n39712 ;
  assign y10116 = ~n39717 ;
  assign y10117 = ~n39719 ;
  assign y10118 = n39721 ;
  assign y10119 = n39722 ;
  assign y10120 = ~n39724 ;
  assign y10121 = ~n39725 ;
  assign y10122 = n39729 ;
  assign y10123 = n39730 ;
  assign y10124 = ~n39732 ;
  assign y10125 = ~n39739 ;
  assign y10126 = n39741 ;
  assign y10127 = n39744 ;
  assign y10128 = n39748 ;
  assign y10129 = n39749 ;
  assign y10130 = ~n39751 ;
  assign y10131 = n39754 ;
  assign y10132 = n39760 ;
  assign y10133 = ~n39766 ;
  assign y10134 = n39767 ;
  assign y10135 = ~n39768 ;
  assign y10136 = n39769 ;
  assign y10137 = n39774 ;
  assign y10138 = n39777 ;
  assign y10139 = n39779 ;
  assign y10140 = n39783 ;
  assign y10141 = n39785 ;
  assign y10142 = n39791 ;
  assign y10143 = ~n39795 ;
  assign y10144 = ~n39797 ;
  assign y10145 = ~n39798 ;
  assign y10146 = ~n39803 ;
  assign y10147 = n39807 ;
  assign y10148 = ~1'b0 ;
  assign y10149 = ~1'b0 ;
  assign y10150 = ~n39808 ;
  assign y10151 = n39811 ;
  assign y10152 = ~n39814 ;
  assign y10153 = ~n39815 ;
  assign y10154 = n39817 ;
  assign y10155 = ~n39822 ;
  assign y10156 = ~n39828 ;
  assign y10157 = ~1'b0 ;
  assign y10158 = ~n39830 ;
  assign y10159 = ~n39832 ;
  assign y10160 = n39835 ;
  assign y10161 = ~n39836 ;
  assign y10162 = n39839 ;
  assign y10163 = ~n39840 ;
  assign y10164 = ~1'b0 ;
  assign y10165 = ~1'b0 ;
  assign y10166 = ~n39844 ;
  assign y10167 = n39849 ;
  assign y10168 = n39857 ;
  assign y10169 = ~n39861 ;
  assign y10170 = ~n39869 ;
  assign y10171 = n39872 ;
  assign y10172 = n39874 ;
  assign y10173 = ~n39875 ;
  assign y10174 = ~n39880 ;
  assign y10175 = n39883 ;
  assign y10176 = n39884 ;
  assign y10177 = ~n39888 ;
  assign y10178 = n39889 ;
  assign y10179 = ~n39892 ;
  assign y10180 = n39899 ;
  assign y10181 = ~n39900 ;
  assign y10182 = n39905 ;
  assign y10183 = n39906 ;
  assign y10184 = n39909 ;
  assign y10185 = ~n39911 ;
  assign y10186 = n39912 ;
  assign y10187 = ~n39918 ;
  assign y10188 = ~n39923 ;
  assign y10189 = ~n39933 ;
  assign y10190 = n39942 ;
  assign y10191 = n39946 ;
  assign y10192 = ~n39949 ;
  assign y10193 = ~n39952 ;
  assign y10194 = ~n39954 ;
  assign y10195 = ~n39955 ;
  assign y10196 = ~n39956 ;
  assign y10197 = n39958 ;
  assign y10198 = n39961 ;
  assign y10199 = ~n39962 ;
  assign y10200 = ~n39965 ;
  assign y10201 = n39966 ;
  assign y10202 = ~1'b0 ;
  assign y10203 = ~n39969 ;
  assign y10204 = ~n39970 ;
  assign y10205 = ~n39977 ;
  assign y10206 = n39978 ;
  assign y10207 = ~n39979 ;
  assign y10208 = ~n39980 ;
  assign y10209 = ~1'b0 ;
  assign y10210 = n39984 ;
  assign y10211 = ~n39989 ;
  assign y10212 = ~n39990 ;
  assign y10213 = n39991 ;
  assign y10214 = n39999 ;
  assign y10215 = ~n40003 ;
  assign y10216 = ~n40005 ;
  assign y10217 = n40006 ;
  assign y10218 = n40007 ;
  assign y10219 = ~n40008 ;
  assign y10220 = n40011 ;
  assign y10221 = ~n40012 ;
  assign y10222 = n40020 ;
  assign y10223 = n40026 ;
  assign y10224 = ~n40029 ;
  assign y10225 = ~n40032 ;
  assign y10226 = ~n40033 ;
  assign y10227 = ~n40034 ;
  assign y10228 = ~n40037 ;
  assign y10229 = n40038 ;
  assign y10230 = n40039 ;
  assign y10231 = n40040 ;
  assign y10232 = ~n40047 ;
  assign y10233 = ~n40049 ;
  assign y10234 = ~n40050 ;
  assign y10235 = n40055 ;
  assign y10236 = ~n40057 ;
  assign y10237 = ~n40058 ;
  assign y10238 = ~n40059 ;
  assign y10239 = ~1'b0 ;
  assign y10240 = n40063 ;
  assign y10241 = ~n40071 ;
  assign y10242 = ~n40072 ;
  assign y10243 = n40074 ;
  assign y10244 = ~n40075 ;
  assign y10245 = ~n40077 ;
  assign y10246 = ~n40080 ;
  assign y10247 = ~1'b0 ;
  assign y10248 = ~n40082 ;
  assign y10249 = ~n40084 ;
  assign y10250 = ~n40085 ;
  assign y10251 = ~n40087 ;
  assign y10252 = ~n40094 ;
  assign y10253 = ~n40095 ;
  assign y10254 = n40099 ;
  assign y10255 = n40104 ;
  assign y10256 = ~n40106 ;
  assign y10257 = ~n40108 ;
  assign y10258 = ~n40110 ;
  assign y10259 = ~n40111 ;
  assign y10260 = ~n40114 ;
  assign y10261 = ~1'b0 ;
  assign y10262 = ~n40117 ;
  assign y10263 = ~n40121 ;
  assign y10264 = n40122 ;
  assign y10265 = n40125 ;
  assign y10266 = ~n40127 ;
  assign y10267 = n40130 ;
  assign y10268 = ~n40131 ;
  assign y10269 = ~n40135 ;
  assign y10270 = n40138 ;
  assign y10271 = ~n40140 ;
  assign y10272 = n40142 ;
  assign y10273 = n40146 ;
  assign y10274 = ~n40147 ;
  assign y10275 = n40150 ;
  assign y10276 = ~n40152 ;
  assign y10277 = ~n40155 ;
  assign y10278 = ~n40159 ;
  assign y10279 = ~1'b0 ;
  assign y10280 = ~n40161 ;
  assign y10281 = n40164 ;
  assign y10282 = ~n40165 ;
  assign y10283 = ~n40168 ;
  assign y10284 = n40171 ;
  assign y10285 = n40172 ;
  assign y10286 = ~n40173 ;
  assign y10287 = ~n40175 ;
  assign y10288 = n40176 ;
  assign y10289 = n40179 ;
  assign y10290 = ~n40182 ;
  assign y10291 = ~n40188 ;
  assign y10292 = ~n40191 ;
  assign y10293 = ~1'b0 ;
  assign y10294 = ~n40192 ;
  assign y10295 = ~n40193 ;
  assign y10296 = ~1'b0 ;
  assign y10297 = n40194 ;
  assign y10298 = n40199 ;
  assign y10299 = n40202 ;
  assign y10300 = ~n40207 ;
  assign y10301 = ~n40211 ;
  assign y10302 = n40212 ;
  assign y10303 = ~1'b0 ;
  assign y10304 = n40217 ;
  assign y10305 = n40218 ;
  assign y10306 = n40223 ;
  assign y10307 = n40224 ;
  assign y10308 = n40231 ;
  assign y10309 = ~n40232 ;
  assign y10310 = ~n40236 ;
  assign y10311 = n40238 ;
  assign y10312 = ~n40242 ;
  assign y10313 = n40247 ;
  assign y10314 = ~n40251 ;
  assign y10315 = ~n40253 ;
  assign y10316 = ~n40259 ;
  assign y10317 = n40262 ;
  assign y10318 = ~n40264 ;
  assign y10319 = n40267 ;
  assign y10320 = n40269 ;
  assign y10321 = ~n40270 ;
  assign y10322 = n40275 ;
  assign y10323 = ~n40276 ;
  assign y10324 = n40277 ;
  assign y10325 = ~n40278 ;
  assign y10326 = ~n40280 ;
  assign y10327 = ~n40283 ;
  assign y10328 = n40286 ;
  assign y10329 = n40287 ;
  assign y10330 = n40288 ;
  assign y10331 = ~n40291 ;
  assign y10332 = n40295 ;
  assign y10333 = n40299 ;
  assign y10334 = ~n40308 ;
  assign y10335 = n40312 ;
  assign y10336 = n40315 ;
  assign y10337 = n40316 ;
  assign y10338 = n40319 ;
  assign y10339 = n40326 ;
  assign y10340 = n40329 ;
  assign y10341 = n40330 ;
  assign y10342 = ~n40332 ;
  assign y10343 = n40336 ;
  assign y10344 = ~n40338 ;
  assign y10345 = n40339 ;
  assign y10346 = n40340 ;
  assign y10347 = n40342 ;
  assign y10348 = n40345 ;
  assign y10349 = n40347 ;
  assign y10350 = n40351 ;
  assign y10351 = ~n40352 ;
  assign y10352 = ~n40355 ;
  assign y10353 = ~n40359 ;
  assign y10354 = n40367 ;
  assign y10355 = ~n40371 ;
  assign y10356 = ~1'b0 ;
  assign y10357 = ~n40372 ;
  assign y10358 = ~n40376 ;
  assign y10359 = n40377 ;
  assign y10360 = ~n40379 ;
  assign y10361 = ~1'b0 ;
  assign y10362 = n40384 ;
  assign y10363 = n40385 ;
  assign y10364 = ~n40386 ;
  assign y10365 = n40387 ;
  assign y10366 = ~n40388 ;
  assign y10367 = ~n40393 ;
  assign y10368 = n40398 ;
  assign y10369 = ~n40403 ;
  assign y10370 = n40404 ;
  assign y10371 = ~n40405 ;
  assign y10372 = ~n40408 ;
  assign y10373 = n40410 ;
  assign y10374 = ~n40412 ;
  assign y10375 = ~n40413 ;
  assign y10376 = ~1'b0 ;
  assign y10377 = n40415 ;
  assign y10378 = n40418 ;
  assign y10379 = n40420 ;
  assign y10380 = ~n40422 ;
  assign y10381 = n40423 ;
  assign y10382 = ~n40425 ;
  assign y10383 = n40427 ;
  assign y10384 = ~n40431 ;
  assign y10385 = n40434 ;
  assign y10386 = n40437 ;
  assign y10387 = ~1'b0 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = ~n40438 ;
  assign y10390 = ~n40444 ;
  assign y10391 = n40446 ;
  assign y10392 = n40448 ;
  assign y10393 = ~n40452 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = n40454 ;
  assign y10396 = ~n40456 ;
  assign y10397 = ~n40459 ;
  assign y10398 = ~n40460 ;
  assign y10399 = ~n40465 ;
  assign y10400 = ~n40472 ;
  assign y10401 = n40474 ;
  assign y10402 = ~n40478 ;
  assign y10403 = n40482 ;
  assign y10404 = n40484 ;
  assign y10405 = ~n40486 ;
  assign y10406 = n40487 ;
  assign y10407 = ~n40489 ;
  assign y10408 = ~n40491 ;
  assign y10409 = n40492 ;
  assign y10410 = n40493 ;
  assign y10411 = n40498 ;
  assign y10412 = ~1'b0 ;
  assign y10413 = ~n40505 ;
  assign y10414 = ~n40514 ;
  assign y10415 = ~n40515 ;
  assign y10416 = n40518 ;
  assign y10417 = ~n40521 ;
  assign y10418 = ~1'b0 ;
  assign y10419 = ~n40524 ;
  assign y10420 = ~n40525 ;
  assign y10421 = n40526 ;
  assign y10422 = ~1'b0 ;
  assign y10423 = ~n40528 ;
  assign y10424 = n40530 ;
  assign y10425 = ~n40535 ;
  assign y10426 = ~n40538 ;
  assign y10427 = ~n40542 ;
  assign y10428 = n40543 ;
  assign y10429 = n40545 ;
  assign y10430 = ~1'b0 ;
  assign y10431 = n40546 ;
  assign y10432 = n40547 ;
  assign y10433 = n40548 ;
  assign y10434 = ~n40552 ;
  assign y10435 = ~n40554 ;
  assign y10436 = ~n40559 ;
  assign y10437 = ~1'b0 ;
  assign y10438 = ~1'b0 ;
  assign y10439 = n40563 ;
  assign y10440 = n40569 ;
  assign y10441 = n40572 ;
  assign y10442 = n40573 ;
  assign y10443 = ~n40575 ;
  assign y10444 = ~1'b0 ;
  assign y10445 = ~1'b0 ;
  assign y10446 = ~1'b0 ;
  assign y10447 = n40576 ;
  assign y10448 = ~n40583 ;
  assign y10449 = ~n40586 ;
  assign y10450 = n40588 ;
  assign y10451 = ~n40595 ;
  assign y10452 = n40604 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = n40610 ;
  assign y10455 = ~n40612 ;
  assign y10456 = ~n40613 ;
  assign y10457 = n40616 ;
  assign y10458 = ~n40617 ;
  assign y10459 = n40619 ;
  assign y10460 = ~n40624 ;
  assign y10461 = ~1'b0 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = ~n40628 ;
  assign y10464 = ~n40630 ;
  assign y10465 = ~n40631 ;
  assign y10466 = n40637 ;
  assign y10467 = n40639 ;
  assign y10468 = ~n40642 ;
  assign y10469 = ~n40643 ;
  assign y10470 = ~n40644 ;
  assign y10471 = n40647 ;
  assign y10472 = ~n40648 ;
  assign y10473 = n40652 ;
  assign y10474 = ~n40657 ;
  assign y10475 = n40663 ;
  assign y10476 = n40668 ;
  assign y10477 = n40669 ;
  assign y10478 = n40670 ;
  assign y10479 = ~n40672 ;
  assign y10480 = n40673 ;
  assign y10481 = n40675 ;
  assign y10482 = n40678 ;
  assign y10483 = ~1'b0 ;
  assign y10484 = n40686 ;
  assign y10485 = n40688 ;
  assign y10486 = n40690 ;
  assign y10487 = n40691 ;
  assign y10488 = n40697 ;
  assign y10489 = ~n40699 ;
  assign y10490 = ~1'b0 ;
  assign y10491 = n40707 ;
  assign y10492 = n40709 ;
  assign y10493 = ~n40714 ;
  assign y10494 = n40716 ;
  assign y10495 = n40720 ;
  assign y10496 = n40721 ;
  assign y10497 = n40728 ;
  assign y10498 = n40731 ;
  assign y10499 = ~n40734 ;
  assign y10500 = ~n40736 ;
  assign y10501 = ~n40737 ;
  assign y10502 = ~n40741 ;
  assign y10503 = ~n40745 ;
  assign y10504 = n40746 ;
  assign y10505 = n40747 ;
  assign y10506 = n40751 ;
  assign y10507 = n40755 ;
  assign y10508 = ~1'b0 ;
  assign y10509 = n40756 ;
  assign y10510 = ~n40757 ;
  assign y10511 = n40758 ;
  assign y10512 = n40762 ;
  assign y10513 = n40763 ;
  assign y10514 = n40764 ;
  assign y10515 = n40765 ;
  assign y10516 = n40766 ;
  assign y10517 = n40770 ;
  assign y10518 = n40773 ;
  assign y10519 = n40777 ;
  assign y10520 = ~n40779 ;
  assign y10521 = ~1'b0 ;
  assign y10522 = ~1'b0 ;
  assign y10523 = ~1'b0 ;
  assign y10524 = n40781 ;
  assign y10525 = ~n40783 ;
  assign y10526 = ~n40784 ;
  assign y10527 = n40786 ;
  assign y10528 = ~1'b0 ;
  assign y10529 = n40798 ;
  assign y10530 = n40799 ;
  assign y10531 = n40800 ;
  assign y10532 = n40803 ;
  assign y10533 = ~1'b0 ;
  assign y10534 = ~n40805 ;
  assign y10535 = n40811 ;
  assign y10536 = ~n40812 ;
  assign y10537 = ~n40814 ;
  assign y10538 = n40817 ;
  assign y10539 = ~n40823 ;
  assign y10540 = n40826 ;
  assign y10541 = ~n40830 ;
  assign y10542 = ~n40834 ;
  assign y10543 = n40837 ;
  assign y10544 = ~n40840 ;
  assign y10545 = n40842 ;
  assign y10546 = ~n40843 ;
  assign y10547 = n40844 ;
  assign y10548 = ~1'b0 ;
  assign y10549 = n40849 ;
  assign y10550 = ~n40851 ;
  assign y10551 = ~n40855 ;
  assign y10552 = n40857 ;
  assign y10553 = ~n40859 ;
  assign y10554 = ~n40863 ;
  assign y10555 = ~n40867 ;
  assign y10556 = ~n40869 ;
  assign y10557 = n40871 ;
  assign y10558 = ~n40880 ;
  assign y10559 = n40882 ;
  assign y10560 = ~n40884 ;
  assign y10561 = ~n40891 ;
  assign y10562 = n40892 ;
  assign y10563 = ~n40894 ;
  assign y10564 = n40895 ;
  assign y10565 = n40896 ;
  assign y10566 = ~n40905 ;
  assign y10567 = n40907 ;
  assign y10568 = ~n40908 ;
  assign y10569 = n40917 ;
  assign y10570 = n40920 ;
  assign y10571 = ~1'b0 ;
  assign y10572 = ~n40922 ;
  assign y10573 = ~n40927 ;
  assign y10574 = ~n40928 ;
  assign y10575 = n40933 ;
  assign y10576 = ~n40935 ;
  assign y10577 = n40936 ;
  assign y10578 = ~n40940 ;
  assign y10579 = n40942 ;
  assign y10580 = ~n40943 ;
  assign y10581 = ~n40944 ;
  assign y10582 = ~n40945 ;
  assign y10583 = n40946 ;
  assign y10584 = n40948 ;
  assign y10585 = n40951 ;
  assign y10586 = ~n40953 ;
  assign y10587 = ~n40954 ;
  assign y10588 = n40957 ;
  assign y10589 = n40958 ;
  assign y10590 = n40961 ;
  assign y10591 = ~n40963 ;
  assign y10592 = n40964 ;
  assign y10593 = ~n40965 ;
  assign y10594 = ~n40968 ;
  assign y10595 = ~n40970 ;
  assign y10596 = ~1'b0 ;
  assign y10597 = ~n40977 ;
  assign y10598 = n40984 ;
  assign y10599 = n40986 ;
  assign y10600 = ~n40987 ;
  assign y10601 = n40988 ;
  assign y10602 = ~n40996 ;
  assign y10603 = n40998 ;
  assign y10604 = ~n41001 ;
  assign y10605 = n41004 ;
  assign y10606 = ~n41012 ;
  assign y10607 = ~n41015 ;
  assign y10608 = ~n41020 ;
  assign y10609 = n41025 ;
  assign y10610 = n41029 ;
  assign y10611 = n41034 ;
  assign y10612 = ~n41037 ;
  assign y10613 = ~n41038 ;
  assign y10614 = n41045 ;
  assign y10615 = n41048 ;
  assign y10616 = ~1'b0 ;
  assign y10617 = ~n41049 ;
  assign y10618 = n41050 ;
  assign y10619 = ~n41055 ;
  assign y10620 = n41057 ;
  assign y10621 = ~n41059 ;
  assign y10622 = n41063 ;
  assign y10623 = ~1'b0 ;
  assign y10624 = ~1'b0 ;
  assign y10625 = ~n41065 ;
  assign y10626 = n41070 ;
  assign y10627 = ~n41074 ;
  assign y10628 = n41079 ;
  assign y10629 = n41081 ;
  assign y10630 = n41086 ;
  assign y10631 = ~n41093 ;
  assign y10632 = ~n41096 ;
  assign y10633 = n41104 ;
  assign y10634 = ~n41105 ;
  assign y10635 = ~n41108 ;
  assign y10636 = n41110 ;
  assign y10637 = n41113 ;
  assign y10638 = n41116 ;
  assign y10639 = ~n41117 ;
  assign y10640 = n41120 ;
  assign y10641 = ~n41122 ;
  assign y10642 = ~n41123 ;
  assign y10643 = ~n41128 ;
  assign y10644 = n41131 ;
  assign y10645 = ~1'b0 ;
  assign y10646 = n41133 ;
  assign y10647 = ~n41135 ;
  assign y10648 = n41142 ;
  assign y10649 = ~n41143 ;
  assign y10650 = ~n41144 ;
  assign y10651 = n41145 ;
  assign y10652 = ~n41150 ;
  assign y10653 = ~n41151 ;
  assign y10654 = ~n41152 ;
  assign y10655 = n41158 ;
  assign y10656 = ~n41159 ;
  assign y10657 = ~n41162 ;
  assign y10658 = n41163 ;
  assign y10659 = n41175 ;
  assign y10660 = n41177 ;
  assign y10661 = ~n41179 ;
  assign y10662 = n41188 ;
  assign y10663 = ~n41193 ;
  assign y10664 = n41198 ;
  assign y10665 = ~n41209 ;
  assign y10666 = n27822 ;
  assign y10667 = n41212 ;
  assign y10668 = n15783 ;
  assign y10669 = ~n41215 ;
  assign y10670 = n41217 ;
  assign y10671 = ~n41221 ;
  assign y10672 = n41227 ;
  assign y10673 = ~n41228 ;
  assign y10674 = n41229 ;
  assign y10675 = n41230 ;
  assign y10676 = ~n41235 ;
  assign y10677 = n41239 ;
  assign y10678 = n41244 ;
  assign y10679 = n41251 ;
  assign y10680 = ~n41253 ;
  assign y10681 = n41255 ;
  assign y10682 = ~n41257 ;
  assign y10683 = n41259 ;
  assign y10684 = n41264 ;
  assign y10685 = ~n41269 ;
  assign y10686 = ~n41273 ;
  assign y10687 = n41277 ;
  assign y10688 = ~n41280 ;
  assign y10689 = n41284 ;
  assign y10690 = ~n41292 ;
  assign y10691 = ~n41297 ;
  assign y10692 = ~1'b0 ;
  assign y10693 = n41302 ;
  assign y10694 = n41303 ;
  assign y10695 = n41304 ;
  assign y10696 = n41305 ;
  assign y10697 = n41306 ;
  assign y10698 = n41308 ;
  assign y10699 = ~1'b0 ;
  assign y10700 = ~n41311 ;
  assign y10701 = ~n41313 ;
  assign y10702 = ~n41315 ;
  assign y10703 = ~n41316 ;
  assign y10704 = n41317 ;
  assign y10705 = ~n41319 ;
  assign y10706 = ~n41321 ;
  assign y10707 = ~1'b0 ;
  assign y10708 = ~1'b0 ;
  assign y10709 = n41323 ;
  assign y10710 = n41327 ;
  assign y10711 = ~n41330 ;
  assign y10712 = ~n41332 ;
  assign y10713 = n41338 ;
  assign y10714 = ~n6138 ;
  assign y10715 = ~n41339 ;
  assign y10716 = ~n41340 ;
  assign y10717 = n41341 ;
  assign y10718 = n41346 ;
  assign y10719 = ~n41350 ;
  assign y10720 = ~n41360 ;
  assign y10721 = n41361 ;
  assign y10722 = n41363 ;
  assign y10723 = ~1'b0 ;
  assign y10724 = n41367 ;
  assign y10725 = ~1'b0 ;
  assign y10726 = n41369 ;
  assign y10727 = n41371 ;
  assign y10728 = n41373 ;
  assign y10729 = ~n41378 ;
  assign y10730 = ~n41381 ;
  assign y10731 = ~n41383 ;
  assign y10732 = ~1'b0 ;
  assign y10733 = n41387 ;
  assign y10734 = ~n41389 ;
  assign y10735 = n41395 ;
  assign y10736 = ~n41399 ;
  assign y10737 = ~n41400 ;
  assign y10738 = ~n41413 ;
  assign y10739 = n41415 ;
  assign y10740 = n41417 ;
  assign y10741 = ~n41419 ;
  assign y10742 = n41422 ;
  assign y10743 = n41426 ;
  assign y10744 = n41428 ;
  assign y10745 = n41430 ;
  assign y10746 = ~n41432 ;
  assign y10747 = n41433 ;
  assign y10748 = ~n41434 ;
  assign y10749 = ~n41438 ;
  assign y10750 = ~n41447 ;
  assign y10751 = n41448 ;
  assign y10752 = n41449 ;
  assign y10753 = ~n41454 ;
  assign y10754 = ~n41455 ;
  assign y10755 = n41460 ;
  assign y10756 = n41467 ;
  assign y10757 = ~n41472 ;
  assign y10758 = n41473 ;
  assign y10759 = ~n41474 ;
  assign y10760 = ~1'b0 ;
  assign y10761 = ~n41476 ;
  assign y10762 = n41478 ;
  assign y10763 = ~n41479 ;
  assign y10764 = n41480 ;
  assign y10765 = ~n41486 ;
  assign y10766 = n41488 ;
  assign y10767 = ~n41492 ;
  assign y10768 = ~n41496 ;
  assign y10769 = ~n41499 ;
  assign y10770 = ~n41500 ;
  assign y10771 = ~n41502 ;
  assign y10772 = ~n41503 ;
  assign y10773 = n41508 ;
  assign y10774 = ~n41511 ;
  assign y10775 = ~n41513 ;
  assign y10776 = ~n41514 ;
  assign y10777 = n41520 ;
  assign y10778 = ~n41523 ;
  assign y10779 = ~n41526 ;
  assign y10780 = ~n41530 ;
  assign y10781 = n41535 ;
  assign y10782 = n41536 ;
  assign y10783 = n41537 ;
  assign y10784 = ~n41542 ;
  assign y10785 = n41545 ;
  assign y10786 = ~1'b0 ;
  assign y10787 = ~n41546 ;
  assign y10788 = ~1'b0 ;
  assign y10789 = ~n41551 ;
  assign y10790 = ~n41554 ;
  assign y10791 = n41558 ;
  assign y10792 = n41560 ;
  assign y10793 = ~n41027 ;
  assign y10794 = n41562 ;
  assign y10795 = ~n41564 ;
  assign y10796 = n41569 ;
  assign y10797 = ~n41570 ;
  assign y10798 = n41572 ;
  assign y10799 = ~n41579 ;
  assign y10800 = ~n41580 ;
  assign y10801 = ~n41582 ;
  assign y10802 = n41592 ;
  assign y10803 = n41596 ;
  assign y10804 = ~n41598 ;
  assign y10805 = n41599 ;
  assign y10806 = n41602 ;
  assign y10807 = ~n41604 ;
  assign y10808 = ~n41606 ;
  assign y10809 = n41607 ;
  assign y10810 = n41609 ;
  assign y10811 = ~1'b0 ;
  assign y10812 = ~n41610 ;
  assign y10813 = n41614 ;
  assign y10814 = n41615 ;
  assign y10815 = n41617 ;
  assign y10816 = n41622 ;
  assign y10817 = n41625 ;
  assign y10818 = ~n41627 ;
  assign y10819 = ~n41630 ;
  assign y10820 = n41634 ;
  assign y10821 = ~n41635 ;
  assign y10822 = ~n41636 ;
  assign y10823 = ~n41639 ;
  assign y10824 = ~n41640 ;
  assign y10825 = ~n41646 ;
  assign y10826 = ~n41648 ;
  assign y10827 = n41650 ;
  assign y10828 = ~n41655 ;
  assign y10829 = ~n41659 ;
  assign y10830 = n41660 ;
  assign y10831 = ~n41663 ;
  assign y10832 = ~n41665 ;
  assign y10833 = ~n41666 ;
  assign y10834 = n41667 ;
  assign y10835 = n41668 ;
  assign y10836 = n41670 ;
  assign y10837 = n41671 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = ~n41679 ;
  assign y10840 = n41680 ;
  assign y10841 = n41681 ;
  assign y10842 = ~n41682 ;
  assign y10843 = n41686 ;
  assign y10844 = ~n41688 ;
  assign y10845 = ~n41692 ;
  assign y10846 = ~1'b0 ;
  assign y10847 = n41697 ;
  assign y10848 = n41701 ;
  assign y10849 = ~n41705 ;
  assign y10850 = ~n41707 ;
  assign y10851 = ~n41708 ;
  assign y10852 = n41710 ;
  assign y10853 = ~n41714 ;
  assign y10854 = ~1'b0 ;
  assign y10855 = ~n41716 ;
  assign y10856 = n41719 ;
  assign y10857 = n41721 ;
  assign y10858 = n41722 ;
  assign y10859 = n41726 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = n41727 ;
  assign y10862 = ~n41731 ;
  assign y10863 = n41738 ;
  assign y10864 = n41739 ;
  assign y10865 = n41741 ;
  assign y10866 = n41743 ;
  assign y10867 = ~n41744 ;
  assign y10868 = n41751 ;
  assign y10869 = n41753 ;
  assign y10870 = n41758 ;
  assign y10871 = ~n41760 ;
  assign y10872 = n41763 ;
  assign y10873 = ~n41767 ;
  assign y10874 = ~n41770 ;
  assign y10875 = n41772 ;
  assign y10876 = ~n41776 ;
  assign y10877 = ~n41780 ;
  assign y10878 = ~1'b0 ;
  assign y10879 = ~n41788 ;
  assign y10880 = ~n41789 ;
  assign y10881 = n41793 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = ~n41795 ;
  assign y10884 = n41798 ;
  assign y10885 = ~n41801 ;
  assign y10886 = ~n41802 ;
  assign y10887 = ~1'b0 ;
  assign y10888 = ~n41805 ;
  assign y10889 = ~n41809 ;
  assign y10890 = n41812 ;
  assign y10891 = ~n41815 ;
  assign y10892 = ~n41816 ;
  assign y10893 = n41819 ;
  assign y10894 = ~n41821 ;
  assign y10895 = n41823 ;
  assign y10896 = ~n41826 ;
  assign y10897 = n41827 ;
  assign y10898 = n41828 ;
  assign y10899 = n41829 ;
  assign y10900 = ~1'b0 ;
  assign y10901 = ~1'b0 ;
  assign y10902 = ~1'b0 ;
  assign y10903 = ~n41831 ;
  assign y10904 = n41833 ;
  assign y10905 = n41836 ;
  assign y10906 = ~n41844 ;
  assign y10907 = n41846 ;
  assign y10908 = n41847 ;
  assign y10909 = n41850 ;
  assign y10910 = n41854 ;
  assign y10911 = n41857 ;
  assign y10912 = ~n41860 ;
  assign y10913 = ~n41865 ;
  assign y10914 = ~n41866 ;
  assign y10915 = n41868 ;
  assign y10916 = ~n41872 ;
  assign y10917 = ~n41873 ;
  assign y10918 = ~n41876 ;
  assign y10919 = ~n41885 ;
  assign y10920 = ~n41889 ;
  assign y10921 = n41891 ;
  assign y10922 = n41893 ;
  assign y10923 = n41895 ;
  assign y10924 = n41900 ;
  assign y10925 = n41904 ;
  assign y10926 = ~n41910 ;
  assign y10927 = ~n41915 ;
  assign y10928 = ~n41916 ;
  assign y10929 = ~n41918 ;
  assign y10930 = n41922 ;
  assign y10931 = ~1'b0 ;
  assign y10932 = n41924 ;
  assign y10933 = n41928 ;
  assign y10934 = ~n41931 ;
  assign y10935 = ~n41934 ;
  assign y10936 = n41936 ;
  assign y10937 = ~n41939 ;
  assign y10938 = n41944 ;
  assign y10939 = n41950 ;
  assign y10940 = ~n41952 ;
  assign y10941 = n41958 ;
  assign y10942 = ~n41959 ;
  assign y10943 = ~n41961 ;
  assign y10944 = n41962 ;
  assign y10945 = ~n41963 ;
  assign y10946 = ~1'b0 ;
  assign y10947 = ~n41964 ;
  assign y10948 = ~n41965 ;
  assign y10949 = ~n41966 ;
  assign y10950 = n41968 ;
  assign y10951 = ~n41971 ;
  assign y10952 = n41972 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~n41974 ;
  assign y10955 = ~n41977 ;
  assign y10956 = ~n41979 ;
  assign y10957 = ~n41980 ;
  assign y10958 = n41981 ;
  assign y10959 = n41983 ;
  assign y10960 = ~n41984 ;
  assign y10961 = n41988 ;
  assign y10962 = n41991 ;
  assign y10963 = ~n41994 ;
  assign y10964 = ~n41998 ;
  assign y10965 = ~n41999 ;
  assign y10966 = ~n42001 ;
  assign y10967 = ~n42005 ;
  assign y10968 = n42006 ;
  assign y10969 = n42010 ;
  assign y10970 = ~n42012 ;
  assign y10971 = ~n42014 ;
  assign y10972 = n42016 ;
  assign y10973 = ~n42018 ;
  assign y10974 = n42020 ;
  assign y10975 = n42021 ;
  assign y10976 = n42022 ;
  assign y10977 = ~n42025 ;
  assign y10978 = ~n42030 ;
  assign y10979 = ~n42034 ;
  assign y10980 = ~n42036 ;
  assign y10981 = n42037 ;
  assign y10982 = n42038 ;
  assign y10983 = ~n42042 ;
  assign y10984 = n42044 ;
  assign y10985 = ~n42045 ;
  assign y10986 = n42046 ;
  assign y10987 = n42048 ;
  assign y10988 = ~n42051 ;
  assign y10989 = ~n42057 ;
  assign y10990 = n42062 ;
  assign y10991 = n42065 ;
  assign y10992 = n42066 ;
  assign y10993 = n42068 ;
  assign y10994 = ~1'b0 ;
  assign y10995 = ~n42072 ;
  assign y10996 = ~n42079 ;
  assign y10997 = n42082 ;
  assign y10998 = ~n42084 ;
  assign y10999 = n42088 ;
  assign y11000 = n42089 ;
  assign y11001 = n42094 ;
  assign y11002 = n42098 ;
  assign y11003 = n42100 ;
  assign y11004 = ~n42101 ;
  assign y11005 = ~n42102 ;
  assign y11006 = n42104 ;
  assign y11007 = ~n42105 ;
  assign y11008 = ~n42108 ;
  assign y11009 = ~n42112 ;
  assign y11010 = ~n42116 ;
  assign y11011 = n42118 ;
  assign y11012 = n42121 ;
  assign y11013 = ~n42127 ;
  assign y11014 = n42131 ;
  assign y11015 = n42133 ;
  assign y11016 = n42137 ;
  assign y11017 = ~n42138 ;
  assign y11018 = n42142 ;
  assign y11019 = n42143 ;
  assign y11020 = ~n42145 ;
  assign y11021 = n42149 ;
  assign y11022 = ~n42152 ;
  assign y11023 = ~n42156 ;
  assign y11024 = ~n42161 ;
  assign y11025 = ~n42166 ;
  assign y11026 = ~n42167 ;
  assign y11027 = n42172 ;
  assign y11028 = n42177 ;
  assign y11029 = ~n42179 ;
  assign y11030 = ~n42183 ;
  assign y11031 = n42184 ;
  assign y11032 = ~n42189 ;
  assign y11033 = n42194 ;
  assign y11034 = ~n42199 ;
  assign y11035 = n42204 ;
  assign y11036 = ~n42208 ;
  assign y11037 = ~n42212 ;
  assign y11038 = n42213 ;
  assign y11039 = n42217 ;
  assign y11040 = ~n42219 ;
  assign y11041 = ~n42224 ;
  assign y11042 = ~n42226 ;
  assign y11043 = n42229 ;
  assign y11044 = n42230 ;
  assign y11045 = ~n42232 ;
  assign y11046 = n42233 ;
  assign y11047 = ~1'b0 ;
  assign y11048 = ~n42236 ;
  assign y11049 = ~n42240 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = ~1'b0 ;
  assign y11052 = ~n42245 ;
  assign y11053 = ~n42248 ;
  assign y11054 = n42255 ;
  assign y11055 = ~n42257 ;
  assign y11056 = n42258 ;
  assign y11057 = ~n42259 ;
  assign y11058 = n42260 ;
  assign y11059 = ~1'b0 ;
  assign y11060 = ~n42261 ;
  assign y11061 = ~n42263 ;
  assign y11062 = n42266 ;
  assign y11063 = ~n42267 ;
  assign y11064 = n42273 ;
  assign y11065 = ~n42274 ;
  assign y11066 = ~n42275 ;
  assign y11067 = ~n42276 ;
  assign y11068 = ~n18255 ;
  assign y11069 = n42279 ;
  assign y11070 = n42283 ;
  assign y11071 = n42285 ;
  assign y11072 = n42287 ;
  assign y11073 = ~n42290 ;
  assign y11074 = n42294 ;
  assign y11075 = ~n42298 ;
  assign y11076 = ~1'b0 ;
  assign y11077 = n42300 ;
  assign y11078 = n42302 ;
  assign y11079 = ~n42308 ;
  assign y11080 = ~n42310 ;
  assign y11081 = ~n42313 ;
  assign y11082 = ~n29823 ;
  assign y11083 = n42315 ;
  assign y11084 = ~1'b0 ;
  assign y11085 = ~n42319 ;
  assign y11086 = n42323 ;
  assign y11087 = ~n42326 ;
  assign y11088 = ~n42328 ;
  assign y11089 = ~n42329 ;
  assign y11090 = n42331 ;
  assign y11091 = ~n42334 ;
  assign y11092 = ~1'b0 ;
  assign y11093 = n42338 ;
  assign y11094 = n42341 ;
  assign y11095 = ~n42344 ;
  assign y11096 = ~n42349 ;
  assign y11097 = ~n42350 ;
  assign y11098 = ~n42354 ;
  assign y11099 = ~n42355 ;
  assign y11100 = ~1'b0 ;
  assign y11101 = ~n42357 ;
  assign y11102 = n42360 ;
  assign y11103 = n42361 ;
  assign y11104 = n42362 ;
  assign y11105 = n42364 ;
  assign y11106 = ~n42368 ;
  assign y11107 = n42370 ;
  assign y11108 = ~n42371 ;
  assign y11109 = n42373 ;
  assign y11110 = n42378 ;
  assign y11111 = ~n42380 ;
  assign y11112 = ~n42382 ;
  assign y11113 = ~n42384 ;
  assign y11114 = n42386 ;
  assign y11115 = ~n42388 ;
  assign y11116 = n42389 ;
  assign y11117 = ~n42394 ;
  assign y11118 = n42399 ;
  assign y11119 = n42400 ;
  assign y11120 = n42402 ;
  assign y11121 = n42406 ;
  assign y11122 = n42407 ;
  assign y11123 = n42409 ;
  assign y11124 = ~n42411 ;
  assign y11125 = ~n42413 ;
  assign y11126 = n42416 ;
  assign y11127 = n42420 ;
  assign y11128 = ~n42423 ;
  assign y11129 = n42428 ;
  assign y11130 = ~n42430 ;
  assign y11131 = ~n42435 ;
  assign y11132 = ~n42436 ;
  assign y11133 = ~n42437 ;
  assign y11134 = n42438 ;
  assign y11135 = n42442 ;
  assign y11136 = n42446 ;
  assign y11137 = ~1'b0 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = ~n42448 ;
  assign y11140 = n42449 ;
  assign y11141 = n42450 ;
  assign y11142 = n42455 ;
  assign y11143 = ~n42459 ;
  assign y11144 = ~n42462 ;
  assign y11145 = ~1'b0 ;
  assign y11146 = ~n42465 ;
  assign y11147 = n42467 ;
  assign y11148 = n42468 ;
  assign y11149 = n42469 ;
  assign y11150 = ~n42470 ;
  assign y11151 = n42480 ;
  assign y11152 = n42482 ;
  assign y11153 = ~1'b0 ;
  assign y11154 = n42483 ;
  assign y11155 = ~n42485 ;
  assign y11156 = n42491 ;
  assign y11157 = ~n42492 ;
  assign y11158 = ~n42496 ;
  assign y11159 = n42501 ;
  assign y11160 = n42503 ;
  assign y11161 = ~n42506 ;
  assign y11162 = n42511 ;
  assign y11163 = n42512 ;
  assign y11164 = n42514 ;
  assign y11165 = n42516 ;
  assign y11166 = ~n42519 ;
  assign y11167 = ~n42521 ;
  assign y11168 = n42522 ;
  assign y11169 = n42523 ;
  assign y11170 = n42524 ;
  assign y11171 = n42527 ;
  assign y11172 = ~n42531 ;
  assign y11173 = ~n42533 ;
  assign y11174 = ~n42535 ;
  assign y11175 = n42536 ;
  assign y11176 = ~n42537 ;
  assign y11177 = ~n42540 ;
  assign y11178 = n42542 ;
  assign y11179 = n42544 ;
  assign y11180 = ~n42549 ;
  assign y11181 = ~n42557 ;
  assign y11182 = ~n42561 ;
  assign y11183 = ~n42565 ;
  assign y11184 = n42566 ;
  assign y11185 = ~n42568 ;
  assign y11186 = n42571 ;
  assign y11187 = n42576 ;
  assign y11188 = n42578 ;
  assign y11189 = ~n42581 ;
  assign y11190 = ~1'b0 ;
  assign y11191 = n42583 ;
  assign y11192 = n42584 ;
  assign y11193 = n42585 ;
  assign y11194 = n42590 ;
  assign y11195 = ~n42592 ;
  assign y11196 = ~n42593 ;
  assign y11197 = n42595 ;
  assign y11198 = n42596 ;
  assign y11199 = ~n42600 ;
  assign y11200 = n42605 ;
  assign y11201 = n42609 ;
  assign y11202 = n42610 ;
  assign y11203 = ~n42617 ;
  assign y11204 = ~n373 ;
  assign y11205 = ~n42620 ;
  assign y11206 = n42625 ;
  assign y11207 = n42632 ;
  assign y11208 = ~1'b0 ;
  assign y11209 = ~1'b0 ;
  assign y11210 = ~n42635 ;
  assign y11211 = n42636 ;
  assign y11212 = n42637 ;
  assign y11213 = n42638 ;
  assign y11214 = n42643 ;
  assign y11215 = n42646 ;
  assign y11216 = n42648 ;
  assign y11217 = ~n42650 ;
  assign y11218 = ~n42653 ;
  assign y11219 = n42657 ;
  assign y11220 = n42659 ;
  assign y11221 = ~n42660 ;
  assign y11222 = n42663 ;
  assign y11223 = ~n42671 ;
  assign y11224 = ~n42674 ;
  assign y11225 = ~n42677 ;
  assign y11226 = n42678 ;
  assign y11227 = n42680 ;
  assign y11228 = n42681 ;
  assign y11229 = n42685 ;
  assign y11230 = n42686 ;
  assign y11231 = ~n42688 ;
  assign y11232 = ~n42691 ;
  assign y11233 = ~n42695 ;
  assign y11234 = n42696 ;
  assign y11235 = n42698 ;
  assign y11236 = n42700 ;
  assign y11237 = ~n42701 ;
  assign y11238 = ~n42704 ;
  assign y11239 = ~1'b0 ;
  assign y11240 = n42707 ;
  assign y11241 = n42708 ;
  assign y11242 = ~n42709 ;
  assign y11243 = ~n42710 ;
  assign y11244 = ~n42712 ;
  assign y11245 = ~n42715 ;
  assign y11246 = ~1'b0 ;
  assign y11247 = ~n42718 ;
  assign y11248 = n42720 ;
  assign y11249 = n42722 ;
  assign y11250 = n42725 ;
  assign y11251 = ~n42726 ;
  assign y11252 = ~1'b0 ;
  assign y11253 = ~n42728 ;
  assign y11254 = n42731 ;
  assign y11255 = n42733 ;
  assign y11256 = n42734 ;
  assign y11257 = n42738 ;
  assign y11258 = n42739 ;
  assign y11259 = ~n42741 ;
  assign y11260 = ~n42744 ;
  assign y11261 = ~1'b0 ;
  assign y11262 = ~n42745 ;
  assign y11263 = n42747 ;
  assign y11264 = ~n42752 ;
  assign y11265 = n42755 ;
  assign y11266 = ~n42756 ;
  assign y11267 = ~n42758 ;
  assign y11268 = n42761 ;
  assign y11269 = n42765 ;
  assign y11270 = n42766 ;
  assign y11271 = ~n42767 ;
  assign y11272 = ~n42768 ;
  assign y11273 = ~n42772 ;
  assign y11274 = ~n42775 ;
  assign y11275 = n42776 ;
  assign y11276 = n42779 ;
  assign y11277 = n42780 ;
  assign y11278 = n42782 ;
  assign y11279 = ~1'b0 ;
  assign y11280 = n42784 ;
  assign y11281 = ~n42785 ;
  assign y11282 = n42787 ;
  assign y11283 = ~n42793 ;
  assign y11284 = n42794 ;
  assign y11285 = ~n42803 ;
  assign y11286 = n42807 ;
  assign y11287 = n42810 ;
  assign y11288 = ~n42811 ;
  assign y11289 = n42812 ;
  assign y11290 = n42813 ;
  assign y11291 = n42814 ;
  assign y11292 = ~n42815 ;
  assign y11293 = ~n42817 ;
  assign y11294 = n42824 ;
  assign y11295 = n42826 ;
  assign y11296 = ~n42827 ;
  assign y11297 = n42831 ;
  assign y11298 = n42833 ;
  assign y11299 = n42834 ;
  assign y11300 = ~n42838 ;
  assign y11301 = n42841 ;
  assign y11302 = ~n42848 ;
  assign y11303 = n42853 ;
  assign y11304 = n42859 ;
  assign y11305 = ~n42860 ;
  assign y11306 = n42862 ;
  assign y11307 = ~n42864 ;
  assign y11308 = n42866 ;
  assign y11309 = n42869 ;
  assign y11310 = ~n42873 ;
  assign y11311 = ~n42874 ;
  assign y11312 = n42876 ;
  assign y11313 = n42879 ;
  assign y11314 = ~n42880 ;
  assign y11315 = n42885 ;
  assign y11316 = ~n42886 ;
  assign y11317 = ~n42889 ;
  assign y11318 = n42896 ;
  assign y11319 = n42899 ;
  assign y11320 = n42903 ;
  assign y11321 = ~n42904 ;
  assign y11322 = n42906 ;
  assign y11323 = ~n42909 ;
  assign y11324 = ~n42915 ;
  assign y11325 = ~n42916 ;
  assign y11326 = ~n42917 ;
  assign y11327 = n42919 ;
  assign y11328 = n42920 ;
  assign y11329 = ~n15697 ;
  assign y11330 = n42921 ;
  assign y11331 = n42924 ;
  assign y11332 = ~n42926 ;
  assign y11333 = ~n42930 ;
  assign y11334 = ~1'b0 ;
  assign y11335 = ~1'b0 ;
  assign y11336 = ~n42933 ;
  assign y11337 = ~n42936 ;
  assign y11338 = n42940 ;
  assign y11339 = n42941 ;
  assign y11340 = ~n42949 ;
  assign y11341 = n42955 ;
  assign y11342 = ~n42957 ;
  assign y11343 = n42959 ;
  assign y11344 = ~1'b0 ;
  assign y11345 = ~n42960 ;
  assign y11346 = n42973 ;
  assign y11347 = ~n42976 ;
  assign y11348 = n42977 ;
  assign y11349 = ~n42980 ;
  assign y11350 = n42982 ;
  assign y11351 = ~n42993 ;
  assign y11352 = ~n42997 ;
  assign y11353 = ~n43000 ;
  assign y11354 = ~1'b0 ;
  assign y11355 = n43004 ;
  assign y11356 = n43005 ;
  assign y11357 = n43006 ;
  assign y11358 = n43007 ;
  assign y11359 = n43010 ;
  assign y11360 = ~n43011 ;
  assign y11361 = n43013 ;
  assign y11362 = n43021 ;
  assign y11363 = ~1'b0 ;
  assign y11364 = ~n43025 ;
  assign y11365 = n43033 ;
  assign y11366 = n43037 ;
  assign y11367 = n43041 ;
  assign y11368 = n43044 ;
  assign y11369 = ~n43047 ;
  assign y11370 = n43049 ;
  assign y11371 = ~n43054 ;
  assign y11372 = ~n43056 ;
  assign y11373 = n43057 ;
  assign y11374 = n43059 ;
  assign y11375 = ~n43061 ;
  assign y11376 = ~n43063 ;
  assign y11377 = n43064 ;
  assign y11378 = ~1'b0 ;
  assign y11379 = n43067 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = n43070 ;
  assign y11382 = ~n43083 ;
  assign y11383 = n43085 ;
  assign y11384 = n43087 ;
  assign y11385 = ~n43091 ;
  assign y11386 = ~n43093 ;
  assign y11387 = ~n43098 ;
  assign y11388 = n43100 ;
  assign y11389 = n43101 ;
  assign y11390 = n43102 ;
  assign y11391 = ~n43109 ;
  assign y11392 = n43110 ;
  assign y11393 = n43118 ;
  assign y11394 = n43123 ;
  assign y11395 = ~n43125 ;
  assign y11396 = ~n43129 ;
  assign y11397 = n43133 ;
  assign y11398 = ~n43135 ;
  assign y11399 = ~n43137 ;
  assign y11400 = n43139 ;
  assign y11401 = n43143 ;
  assign y11402 = ~n43146 ;
  assign y11403 = ~n43151 ;
  assign y11404 = ~n43154 ;
  assign y11405 = n43156 ;
  assign y11406 = ~n43157 ;
  assign y11407 = n43162 ;
  assign y11408 = ~n43165 ;
  assign y11409 = n43167 ;
  assign y11410 = ~n43168 ;
  assign y11411 = ~n43169 ;
  assign y11412 = n43170 ;
  assign y11413 = ~n43172 ;
  assign y11414 = n43178 ;
  assign y11415 = n43182 ;
  assign y11416 = ~n43184 ;
  assign y11417 = ~n43186 ;
  assign y11418 = n43187 ;
  assign y11419 = ~n43191 ;
  assign y11420 = ~n43195 ;
  assign y11421 = ~n43196 ;
  assign y11422 = ~1'b0 ;
  assign y11423 = n43201 ;
  assign y11424 = ~n43203 ;
  assign y11425 = n43208 ;
  assign y11426 = ~n43210 ;
  assign y11427 = ~n43211 ;
  assign y11428 = n43214 ;
  assign y11429 = n43215 ;
  assign y11430 = ~n17675 ;
  assign y11431 = ~1'b0 ;
  assign y11432 = ~1'b0 ;
  assign y11433 = n43221 ;
  assign y11434 = ~n43223 ;
  assign y11435 = n43224 ;
  assign y11436 = ~n43225 ;
  assign y11437 = n43234 ;
  assign y11438 = n43236 ;
  assign y11439 = ~n43237 ;
  assign y11440 = n43243 ;
  assign y11441 = ~n43245 ;
  assign y11442 = n43246 ;
  assign y11443 = ~1'b0 ;
  assign y11444 = n43248 ;
  assign y11445 = ~n43251 ;
  assign y11446 = ~n43253 ;
  assign y11447 = ~n43254 ;
  assign y11448 = ~n43258 ;
  assign y11449 = n43265 ;
  assign y11450 = ~n43267 ;
  assign y11451 = ~1'b0 ;
  assign y11452 = ~n43278 ;
  assign y11453 = n43280 ;
  assign y11454 = n43283 ;
  assign y11455 = ~n43286 ;
  assign y11456 = n43291 ;
  assign y11457 = n43300 ;
  assign y11458 = n43303 ;
  assign y11459 = n43304 ;
  assign y11460 = ~n43306 ;
  assign y11461 = ~1'b0 ;
  assign y11462 = ~n43307 ;
  assign y11463 = ~n43308 ;
  assign y11464 = n43313 ;
  assign y11465 = ~n43314 ;
  assign y11466 = ~n43316 ;
  assign y11467 = n43317 ;
  assign y11468 = ~n43319 ;
  assign y11469 = n43323 ;
  assign y11470 = ~n43324 ;
  assign y11471 = ~n43326 ;
  assign y11472 = ~n43330 ;
  assign y11473 = n43333 ;
  assign y11474 = ~n43336 ;
  assign y11475 = ~n43337 ;
  assign y11476 = ~n43338 ;
  assign y11477 = ~1'b0 ;
  assign y11478 = n43340 ;
  assign y11479 = ~n43341 ;
  assign y11480 = ~n43342 ;
  assign y11481 = n43344 ;
  assign y11482 = n43345 ;
  assign y11483 = ~n43346 ;
  assign y11484 = ~n43351 ;
  assign y11485 = ~n43355 ;
  assign y11486 = n43358 ;
  assign y11487 = n43362 ;
  assign y11488 = ~n43369 ;
  assign y11489 = n43370 ;
  assign y11490 = ~n43373 ;
  assign y11491 = ~n43374 ;
  assign y11492 = n43382 ;
  assign y11493 = ~n43384 ;
  assign y11494 = n43392 ;
  assign y11495 = n43397 ;
  assign y11496 = n43399 ;
  assign y11497 = n43400 ;
  assign y11498 = ~n43402 ;
  assign y11499 = n43407 ;
  assign y11500 = n43414 ;
  assign y11501 = n43419 ;
  assign y11502 = ~1'b0 ;
  assign y11503 = n43421 ;
  assign y11504 = n43422 ;
  assign y11505 = n43423 ;
  assign y11506 = ~n43431 ;
  assign y11507 = n43434 ;
  assign y11508 = n43435 ;
  assign y11509 = n43437 ;
  assign y11510 = ~n43440 ;
  assign y11511 = ~n43447 ;
  assign y11512 = n43451 ;
  assign y11513 = ~n43455 ;
  assign y11514 = ~n43456 ;
  assign y11515 = n43460 ;
  assign y11516 = ~n43461 ;
  assign y11517 = n43462 ;
  assign y11518 = ~n43467 ;
  assign y11519 = n43469 ;
  assign y11520 = n43472 ;
  assign y11521 = n43479 ;
  assign y11522 = n43481 ;
  assign y11523 = ~n43482 ;
  assign y11524 = n43491 ;
  assign y11525 = n43494 ;
  assign y11526 = ~1'b0 ;
  assign y11527 = n43495 ;
  assign y11528 = n43497 ;
  assign y11529 = ~n43501 ;
  assign y11530 = ~n43504 ;
  assign y11531 = ~n43506 ;
  assign y11532 = n43508 ;
  assign y11533 = n43509 ;
  assign y11534 = ~n43512 ;
  assign y11535 = n43514 ;
  assign y11536 = ~n43516 ;
  assign y11537 = n43519 ;
  assign y11538 = n43521 ;
  assign y11539 = n43522 ;
  assign y11540 = ~n43524 ;
  assign y11541 = ~n43525 ;
  assign y11542 = ~n43528 ;
  assign y11543 = n43535 ;
  assign y11544 = n43537 ;
  assign y11545 = n43540 ;
  assign y11546 = ~1'b0 ;
  assign y11547 = ~n43541 ;
  assign y11548 = n43542 ;
  assign y11549 = ~n43548 ;
  assign y11550 = ~1'b0 ;
  assign y11551 = n43553 ;
  assign y11552 = n43554 ;
  assign y11553 = n43555 ;
  assign y11554 = ~n43556 ;
  assign y11555 = n43557 ;
  assign y11556 = n43565 ;
  assign y11557 = n43567 ;
  assign y11558 = n43570 ;
  assign y11559 = ~n43572 ;
  assign y11560 = n43573 ;
  assign y11561 = n43576 ;
  assign y11562 = ~n43579 ;
  assign y11563 = n25524 ;
  assign y11564 = ~n43582 ;
  assign y11565 = ~n43594 ;
  assign y11566 = ~n43596 ;
  assign y11567 = ~n43597 ;
  assign y11568 = ~n43600 ;
  assign y11569 = n43601 ;
  assign y11570 = n43602 ;
  assign y11571 = ~n43603 ;
  assign y11572 = n43605 ;
  assign y11573 = ~n43606 ;
  assign y11574 = ~n43609 ;
  assign y11575 = ~n43614 ;
  assign y11576 = ~n43615 ;
  assign y11577 = ~n43619 ;
  assign y11578 = ~n43623 ;
  assign y11579 = n43629 ;
  assign y11580 = n43630 ;
  assign y11581 = n43632 ;
  assign y11582 = n43634 ;
  assign y11583 = ~1'b0 ;
  assign y11584 = ~n43635 ;
  assign y11585 = ~n43636 ;
  assign y11586 = n43640 ;
  assign y11587 = n43648 ;
  assign y11588 = ~1'b0 ;
  assign y11589 = n43651 ;
  assign y11590 = ~1'b0 ;
  assign y11591 = ~n43655 ;
  assign y11592 = ~n43658 ;
  assign y11593 = ~n43660 ;
  assign y11594 = ~n43663 ;
  assign y11595 = ~n43666 ;
  assign y11596 = n43669 ;
  assign y11597 = ~n43678 ;
  assign y11598 = n43680 ;
  assign y11599 = ~1'b0 ;
  assign y11600 = n43683 ;
  assign y11601 = n43684 ;
  assign y11602 = ~n43689 ;
  assign y11603 = ~n43690 ;
  assign y11604 = n43695 ;
  assign y11605 = n43697 ;
  assign y11606 = ~n43698 ;
  assign y11607 = ~n43701 ;
  assign y11608 = n43702 ;
  assign y11609 = n43703 ;
  assign y11610 = ~n43710 ;
  assign y11611 = n43713 ;
  assign y11612 = n43714 ;
  assign y11613 = n43717 ;
  assign y11614 = ~n43725 ;
  assign y11615 = n43730 ;
  assign y11616 = n43733 ;
  assign y11617 = ~n43734 ;
  assign y11618 = n43735 ;
  assign y11619 = n43740 ;
  assign y11620 = ~n43741 ;
  assign y11621 = ~n43745 ;
  assign y11622 = ~n43748 ;
  assign y11623 = n43751 ;
  assign y11624 = ~n43753 ;
  assign y11625 = ~n43760 ;
  assign y11626 = n43762 ;
  assign y11627 = ~n43766 ;
  assign y11628 = n43768 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = ~n43771 ;
  assign y11631 = n43773 ;
  assign y11632 = n43782 ;
  assign y11633 = ~n43784 ;
  assign y11634 = n43786 ;
  assign y11635 = ~n43788 ;
  assign y11636 = n43789 ;
  assign y11637 = ~n43790 ;
  assign y11638 = ~n43792 ;
  assign y11639 = ~1'b0 ;
  assign y11640 = ~n43794 ;
  assign y11641 = n43797 ;
  assign y11642 = ~n43799 ;
  assign y11643 = n43801 ;
  assign y11644 = n43805 ;
  assign y11645 = ~n43810 ;
  assign y11646 = n43811 ;
  assign y11647 = ~n43815 ;
  assign y11648 = ~n43817 ;
  assign y11649 = ~n43822 ;
  assign y11650 = n43825 ;
  assign y11651 = n43827 ;
  assign y11652 = n43830 ;
  assign y11653 = n43837 ;
  assign y11654 = ~n10801 ;
  assign y11655 = ~n43843 ;
  assign y11656 = ~n43846 ;
  assign y11657 = ~n43848 ;
  assign y11658 = n43849 ;
  assign y11659 = n43850 ;
  assign y11660 = ~n43852 ;
  assign y11661 = n43859 ;
  assign y11662 = n43863 ;
  assign y11663 = ~n43864 ;
  assign y11664 = ~n43865 ;
  assign y11665 = ~n43866 ;
  assign y11666 = ~n43870 ;
  assign y11667 = ~n43872 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = n43874 ;
  assign y11670 = n43877 ;
  assign y11671 = ~n43883 ;
  assign y11672 = n43884 ;
  assign y11673 = n43886 ;
  assign y11674 = n43887 ;
  assign y11675 = ~n43889 ;
  assign y11676 = n43890 ;
  assign y11677 = n43892 ;
  assign y11678 = ~n43894 ;
  assign y11679 = ~n43895 ;
  assign y11680 = n43896 ;
  assign y11681 = ~n43897 ;
  assign y11682 = ~n43898 ;
  assign y11683 = ~n43906 ;
  assign y11684 = ~n43909 ;
  assign y11685 = ~n43912 ;
  assign y11686 = n43913 ;
  assign y11687 = ~n43917 ;
  assign y11688 = ~n43920 ;
  assign y11689 = ~n43926 ;
  assign y11690 = n43928 ;
  assign y11691 = n43930 ;
  assign y11692 = n43931 ;
  assign y11693 = n43932 ;
  assign y11694 = n43934 ;
  assign y11695 = ~n43936 ;
  assign y11696 = ~n43940 ;
  assign y11697 = ~n43941 ;
  assign y11698 = n43945 ;
  assign y11699 = ~n43949 ;
  assign y11700 = n43950 ;
  assign y11701 = n43951 ;
  assign y11702 = ~n43953 ;
  assign y11703 = ~n43955 ;
  assign y11704 = n43956 ;
  assign y11705 = ~n43957 ;
  assign y11706 = n43958 ;
  assign y11707 = ~n43961 ;
  assign y11708 = ~n43962 ;
  assign y11709 = n43963 ;
  assign y11710 = ~n43964 ;
  assign y11711 = n43967 ;
  assign y11712 = n43968 ;
  assign y11713 = ~n43969 ;
  assign y11714 = ~n43978 ;
  assign y11715 = ~n43979 ;
  assign y11716 = ~n43982 ;
  assign y11717 = ~n43984 ;
  assign y11718 = ~n43986 ;
  assign y11719 = n43989 ;
  assign y11720 = ~n43993 ;
  assign y11721 = ~n43995 ;
  assign y11722 = n43997 ;
  assign y11723 = ~n43999 ;
  assign y11724 = ~n44000 ;
  assign y11725 = n44003 ;
  assign y11726 = n44004 ;
  assign y11727 = n44007 ;
  assign y11728 = n44008 ;
  assign y11729 = n44011 ;
  assign y11730 = ~n44017 ;
  assign y11731 = n44026 ;
  assign y11732 = n44028 ;
  assign y11733 = ~n44030 ;
  assign y11734 = n44032 ;
  assign y11735 = ~n44034 ;
  assign y11736 = ~n44036 ;
  assign y11737 = ~n44039 ;
  assign y11738 = n44040 ;
  assign y11739 = ~n44041 ;
  assign y11740 = n44043 ;
  assign y11741 = ~1'b0 ;
  assign y11742 = n44046 ;
  assign y11743 = ~n44047 ;
  assign y11744 = ~n44052 ;
  assign y11745 = n44054 ;
  assign y11746 = n44058 ;
  assign y11747 = ~n44062 ;
  assign y11748 = n44065 ;
  assign y11749 = ~n44067 ;
  assign y11750 = n44069 ;
  assign y11751 = ~1'b0 ;
  assign y11752 = ~n44072 ;
  assign y11753 = ~n44081 ;
  assign y11754 = ~n44083 ;
  assign y11755 = ~n44085 ;
  assign y11756 = n44091 ;
  assign y11757 = ~n44097 ;
  assign y11758 = ~n44098 ;
  assign y11759 = ~n44100 ;
  assign y11760 = ~n44102 ;
  assign y11761 = n44103 ;
  assign y11762 = n44104 ;
  assign y11763 = ~n44105 ;
  assign y11764 = ~n44107 ;
  assign y11765 = n44110 ;
  assign y11766 = n44112 ;
  assign y11767 = ~n44114 ;
  assign y11768 = ~n44115 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = n44117 ;
  assign y11771 = ~n44118 ;
  assign y11772 = ~n44120 ;
  assign y11773 = ~n44123 ;
  assign y11774 = ~n44125 ;
  assign y11775 = n44128 ;
  assign y11776 = n44130 ;
  assign y11777 = ~1'b0 ;
  assign y11778 = n44134 ;
  assign y11779 = n44136 ;
  assign y11780 = ~n44138 ;
  assign y11781 = ~n44140 ;
  assign y11782 = n44144 ;
  assign y11783 = ~n44145 ;
  assign y11784 = ~n44147 ;
  assign y11785 = ~n44152 ;
  assign y11786 = n44154 ;
  assign y11787 = ~1'b0 ;
  assign y11788 = ~n44156 ;
  assign y11789 = ~n44158 ;
  assign y11790 = ~n44159 ;
  assign y11791 = n44160 ;
  assign y11792 = n44161 ;
  assign y11793 = ~1'b0 ;
  assign y11794 = ~n44163 ;
  assign y11795 = ~n44165 ;
  assign y11796 = ~n44168 ;
  assign y11797 = n44172 ;
  assign y11798 = ~n44174 ;
  assign y11799 = ~n44178 ;
  assign y11800 = ~n44182 ;
  assign y11801 = ~n44183 ;
  assign y11802 = n44186 ;
  assign y11803 = ~1'b0 ;
  assign y11804 = ~1'b0 ;
  assign y11805 = ~n44187 ;
  assign y11806 = ~n44191 ;
  assign y11807 = ~n44192 ;
  assign y11808 = n44194 ;
  assign y11809 = n44204 ;
  assign y11810 = ~n44209 ;
  assign y11811 = n44210 ;
  assign y11812 = ~1'b0 ;
  assign y11813 = ~1'b0 ;
  assign y11814 = ~n44212 ;
  assign y11815 = n44215 ;
  assign y11816 = ~n44216 ;
  assign y11817 = ~n44218 ;
  assign y11818 = ~n44219 ;
  assign y11819 = n44224 ;
  assign y11820 = ~n44226 ;
  assign y11821 = n44235 ;
  assign y11822 = ~n44237 ;
  assign y11823 = n44242 ;
  assign y11824 = ~n44245 ;
  assign y11825 = ~n44246 ;
  assign y11826 = n44247 ;
  assign y11827 = ~1'b0 ;
  assign y11828 = ~n44249 ;
  assign y11829 = n44251 ;
  assign y11830 = n16322 ;
  assign y11831 = ~n44254 ;
  assign y11832 = ~n44255 ;
  assign y11833 = ~n44256 ;
  assign y11834 = n44259 ;
  assign y11835 = ~n44261 ;
  assign y11836 = ~n44264 ;
  assign y11837 = ~n44265 ;
  assign y11838 = ~n44266 ;
  assign y11839 = n44269 ;
  assign y11840 = n44272 ;
  assign y11841 = n44274 ;
  assign y11842 = n44275 ;
  assign y11843 = ~n44277 ;
  assign y11844 = ~n44279 ;
  assign y11845 = ~n44283 ;
  assign y11846 = n44291 ;
  assign y11847 = n44292 ;
  assign y11848 = ~n44300 ;
  assign y11849 = n44302 ;
  assign y11850 = n44303 ;
  assign y11851 = n44304 ;
  assign y11852 = n44305 ;
  assign y11853 = n44308 ;
  assign y11854 = ~n44311 ;
  assign y11855 = ~n44313 ;
  assign y11856 = n44315 ;
  assign y11857 = n44316 ;
  assign y11858 = ~n44322 ;
  assign y11859 = ~n44324 ;
  assign y11860 = n44327 ;
  assign y11861 = n44328 ;
  assign y11862 = n44332 ;
  assign y11863 = n44334 ;
  assign y11864 = ~n44338 ;
  assign y11865 = n44340 ;
  assign y11866 = ~1'b0 ;
  assign y11867 = ~n44341 ;
  assign y11868 = n44344 ;
  assign y11869 = n44348 ;
  assign y11870 = ~n44349 ;
  assign y11871 = n44353 ;
  assign y11872 = ~1'b0 ;
  assign y11873 = n44356 ;
  assign y11874 = ~n44360 ;
  assign y11875 = n44362 ;
  assign y11876 = ~n44363 ;
  assign y11877 = ~n44365 ;
  assign y11878 = n44373 ;
  assign y11879 = n44374 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = ~n44377 ;
  assign y11882 = n44378 ;
  assign y11883 = n44385 ;
  assign y11884 = n44394 ;
  assign y11885 = ~n44395 ;
  assign y11886 = n44396 ;
  assign y11887 = n44400 ;
  assign y11888 = n44403 ;
  assign y11889 = n44404 ;
  assign y11890 = ~n44407 ;
  assign y11891 = n44409 ;
  assign y11892 = ~n44411 ;
  assign y11893 = n44412 ;
  assign y11894 = n44417 ;
  assign y11895 = n44418 ;
  assign y11896 = ~n44420 ;
  assign y11897 = ~n44421 ;
  assign y11898 = n44427 ;
  assign y11899 = ~n44432 ;
  assign y11900 = ~n44434 ;
  assign y11901 = ~n44437 ;
  assign y11902 = n44439 ;
  assign y11903 = n44440 ;
  assign y11904 = n44442 ;
  assign y11905 = n44443 ;
  assign y11906 = n44450 ;
  assign y11907 = ~n44452 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = n44457 ;
  assign y11910 = ~n44458 ;
  assign y11911 = n44460 ;
  assign y11912 = ~n31245 ;
  assign y11913 = ~n44462 ;
  assign y11914 = ~n44464 ;
  assign y11915 = ~n44465 ;
  assign y11916 = n44467 ;
  assign y11917 = n44474 ;
  assign y11918 = ~n44477 ;
  assign y11919 = n44478 ;
  assign y11920 = ~n44479 ;
  assign y11921 = n44480 ;
  assign y11922 = n44481 ;
  assign y11923 = ~n44486 ;
  assign y11924 = ~n44488 ;
  assign y11925 = n44489 ;
  assign y11926 = n44493 ;
  assign y11927 = ~n44498 ;
  assign y11928 = ~n44500 ;
  assign y11929 = ~n44501 ;
  assign y11930 = n44503 ;
  assign y11931 = n44504 ;
  assign y11932 = n44505 ;
  assign y11933 = ~n44508 ;
  assign y11934 = n44510 ;
  assign y11935 = n44514 ;
  assign y11936 = ~n5219 ;
  assign y11937 = ~n44522 ;
  assign y11938 = n44532 ;
  assign y11939 = n44538 ;
  assign y11940 = n44542 ;
  assign y11941 = ~n44555 ;
  assign y11942 = ~n44556 ;
  assign y11943 = n44559 ;
  assign y11944 = n44564 ;
  assign y11945 = n44568 ;
  assign y11946 = ~n44569 ;
  assign y11947 = ~n44570 ;
  assign y11948 = n44580 ;
  assign y11949 = ~n44581 ;
  assign y11950 = n44585 ;
  assign y11951 = ~n44589 ;
  assign y11952 = ~n44592 ;
  assign y11953 = n44594 ;
  assign y11954 = n44601 ;
  assign y11955 = n44602 ;
  assign y11956 = n44604 ;
  assign y11957 = ~n44607 ;
  assign y11958 = n44613 ;
  assign y11959 = ~n44616 ;
  assign y11960 = n44618 ;
  assign y11961 = n44620 ;
  assign y11962 = n44622 ;
  assign y11963 = n44623 ;
  assign y11964 = n44626 ;
  assign y11965 = n44628 ;
  assign y11966 = ~n44630 ;
  assign y11967 = ~n44633 ;
  assign y11968 = ~n44634 ;
  assign y11969 = ~n44640 ;
  assign y11970 = ~n44647 ;
  assign y11971 = ~n44654 ;
  assign y11972 = ~n44656 ;
  assign y11973 = ~n44659 ;
  assign y11974 = n44660 ;
  assign y11975 = ~n44663 ;
  assign y11976 = ~n44669 ;
  assign y11977 = n44674 ;
  assign y11978 = ~1'b0 ;
  assign y11979 = ~n44677 ;
  assign y11980 = ~n44679 ;
  assign y11981 = n44680 ;
  assign y11982 = ~n44681 ;
  assign y11983 = n44682 ;
  assign y11984 = ~n44684 ;
  assign y11985 = ~n44685 ;
  assign y11986 = ~1'b0 ;
  assign y11987 = ~1'b0 ;
  assign y11988 = ~n44689 ;
  assign y11989 = ~n44690 ;
  assign y11990 = ~n44692 ;
  assign y11991 = ~n44695 ;
  assign y11992 = n44696 ;
  assign y11993 = n44697 ;
  assign y11994 = ~n44698 ;
  assign y11995 = ~n44699 ;
  assign y11996 = n44702 ;
  assign y11997 = n44712 ;
  assign y11998 = ~n44714 ;
  assign y11999 = ~n44717 ;
  assign y12000 = ~n44719 ;
  assign y12001 = ~n44722 ;
  assign y12002 = ~n44726 ;
  assign y12003 = ~n44727 ;
  assign y12004 = n44729 ;
  assign y12005 = n44730 ;
  assign y12006 = n44733 ;
  assign y12007 = n44734 ;
  assign y12008 = n44736 ;
  assign y12009 = ~n44737 ;
  assign y12010 = ~n44738 ;
  assign y12011 = n44741 ;
  assign y12012 = n44742 ;
  assign y12013 = n44744 ;
  assign y12014 = n20396 ;
  assign y12015 = ~n44745 ;
  assign y12016 = ~n44746 ;
  assign y12017 = ~n44748 ;
  assign y12018 = ~n44754 ;
  assign y12019 = n44758 ;
  assign y12020 = n44760 ;
  assign y12021 = ~n44763 ;
  assign y12022 = n44765 ;
  assign y12023 = ~n44772 ;
  assign y12024 = n44773 ;
  assign y12025 = n44775 ;
  assign y12026 = n44776 ;
  assign y12027 = n44782 ;
  assign y12028 = n44783 ;
  assign y12029 = n44785 ;
  assign y12030 = ~n44789 ;
  assign y12031 = ~n44794 ;
  assign y12032 = ~n44797 ;
  assign y12033 = n44798 ;
  assign y12034 = ~n44799 ;
  assign y12035 = ~n44801 ;
  assign y12036 = n44804 ;
  assign y12037 = ~n44806 ;
  assign y12038 = ~n44808 ;
  assign y12039 = n44809 ;
  assign y12040 = ~n44810 ;
  assign y12041 = ~n44811 ;
  assign y12042 = n44812 ;
  assign y12043 = n44816 ;
  assign y12044 = ~n44817 ;
  assign y12045 = ~n44821 ;
  assign y12046 = ~n44822 ;
  assign y12047 = n44827 ;
  assign y12048 = ~n44829 ;
  assign y12049 = ~n44833 ;
  assign y12050 = n44836 ;
  assign y12051 = n44837 ;
  assign y12052 = ~n44838 ;
  assign y12053 = n44839 ;
  assign y12054 = ~1'b0 ;
  assign y12055 = n44841 ;
  assign y12056 = ~n44843 ;
  assign y12057 = n44845 ;
  assign y12058 = n44846 ;
  assign y12059 = n27209 ;
  assign y12060 = ~n44847 ;
  assign y12061 = ~n44848 ;
  assign y12062 = ~n44849 ;
  assign y12063 = ~1'b0 ;
  assign y12064 = ~n44851 ;
  assign y12065 = ~n44852 ;
  assign y12066 = ~n44853 ;
  assign y12067 = n44854 ;
  assign y12068 = ~n44856 ;
  assign y12069 = ~n44859 ;
  assign y12070 = ~n44861 ;
  assign y12071 = n44863 ;
  assign y12072 = n44865 ;
  assign y12073 = n44869 ;
  assign y12074 = ~n44870 ;
  assign y12075 = ~n44871 ;
  assign y12076 = n44873 ;
  assign y12077 = ~n44875 ;
  assign y12078 = n44877 ;
  assign y12079 = ~n44879 ;
  assign y12080 = ~1'b0 ;
  assign y12081 = ~n44882 ;
  assign y12082 = ~n44886 ;
  assign y12083 = ~n44890 ;
  assign y12084 = ~n44893 ;
  assign y12085 = n44895 ;
  assign y12086 = n44899 ;
  assign y12087 = n44900 ;
  assign y12088 = ~n44906 ;
  assign y12089 = ~n44909 ;
  assign y12090 = ~n44910 ;
  assign y12091 = ~1'b0 ;
  assign y12092 = n44911 ;
  assign y12093 = n44913 ;
  assign y12094 = ~n44914 ;
  assign y12095 = n44916 ;
  assign y12096 = n44918 ;
  assign y12097 = n44920 ;
  assign y12098 = n44924 ;
  assign y12099 = ~1'b0 ;
  assign y12100 = ~1'b0 ;
  assign y12101 = ~n44926 ;
  assign y12102 = n44927 ;
  assign y12103 = ~n44928 ;
  assign y12104 = ~n44931 ;
  assign y12105 = n44932 ;
  assign y12106 = n44935 ;
  assign y12107 = ~n44937 ;
  assign y12108 = ~n44938 ;
  assign y12109 = ~n44939 ;
  assign y12110 = n44940 ;
  assign y12111 = ~n44945 ;
  assign y12112 = n44947 ;
  assign y12113 = ~n44948 ;
  assign y12114 = ~n44949 ;
  assign y12115 = n44953 ;
  assign y12116 = n44956 ;
  assign y12117 = n44957 ;
  assign y12118 = ~n44959 ;
  assign y12119 = ~1'b0 ;
  assign y12120 = n44961 ;
  assign y12121 = ~n44963 ;
  assign y12122 = n44973 ;
  assign y12123 = n44979 ;
  assign y12124 = n44982 ;
  assign y12125 = ~n44983 ;
  assign y12126 = ~n44989 ;
  assign y12127 = ~n44991 ;
  assign y12128 = ~n44997 ;
  assign y12129 = ~n44999 ;
  assign y12130 = n45000 ;
  assign y12131 = n45003 ;
  assign y12132 = n45004 ;
  assign y12133 = ~n45006 ;
  assign y12134 = ~1'b0 ;
  assign y12135 = n45008 ;
  assign y12136 = n45011 ;
  assign y12137 = ~n45014 ;
  assign y12138 = ~n45015 ;
  assign y12139 = ~n45016 ;
  assign y12140 = ~n45020 ;
  assign y12141 = ~n45025 ;
  assign y12142 = n45028 ;
  assign y12143 = n45029 ;
  assign y12144 = n45032 ;
  assign y12145 = ~n45037 ;
  assign y12146 = n45039 ;
  assign y12147 = ~1'b0 ;
  assign y12148 = ~n45046 ;
  assign y12149 = n45047 ;
  assign y12150 = ~n45050 ;
  assign y12151 = n45052 ;
  assign y12152 = n45053 ;
  assign y12153 = ~n45054 ;
  assign y12154 = ~1'b0 ;
  assign y12155 = n45055 ;
  assign y12156 = ~n45057 ;
  assign y12157 = n45058 ;
  assign y12158 = n45063 ;
  assign y12159 = ~n45065 ;
  assign y12160 = n45067 ;
  assign y12161 = n45068 ;
  assign y12162 = ~n45071 ;
  assign y12163 = n45073 ;
  assign y12164 = ~n45077 ;
  assign y12165 = n45078 ;
  assign y12166 = ~1'b0 ;
  assign y12167 = ~n45081 ;
  assign y12168 = n45086 ;
  assign y12169 = n45087 ;
  assign y12170 = n45088 ;
  assign y12171 = ~n45089 ;
  assign y12172 = ~n45092 ;
  assign y12173 = ~n45093 ;
  assign y12174 = n45096 ;
  assign y12175 = n45100 ;
  assign y12176 = ~n45103 ;
  assign y12177 = n45110 ;
  assign y12178 = ~n45111 ;
  assign y12179 = n45118 ;
  assign y12180 = n45121 ;
  assign y12181 = n45124 ;
  assign y12182 = ~n45127 ;
  assign y12183 = n45128 ;
  assign y12184 = ~n45131 ;
  assign y12185 = ~n45132 ;
  assign y12186 = n45135 ;
  assign y12187 = ~n45138 ;
  assign y12188 = ~n45146 ;
  assign y12189 = ~n45150 ;
  assign y12190 = n45158 ;
  assign y12191 = n45159 ;
  assign y12192 = n45162 ;
  assign y12193 = ~n45164 ;
  assign y12194 = ~n45166 ;
  assign y12195 = ~n45169 ;
  assign y12196 = n45171 ;
  assign y12197 = n45172 ;
  assign y12198 = ~n45173 ;
  assign y12199 = ~n45174 ;
  assign y12200 = ~n45175 ;
  assign y12201 = ~n45182 ;
  assign y12202 = n45184 ;
  assign y12203 = ~1'b0 ;
  assign y12204 = ~n45190 ;
  assign y12205 = ~n45191 ;
  assign y12206 = n45192 ;
  assign y12207 = n45193 ;
  assign y12208 = ~n45194 ;
  assign y12209 = ~n45195 ;
  assign y12210 = ~n45203 ;
  assign y12211 = ~n45204 ;
  assign y12212 = n45206 ;
  assign y12213 = ~n45212 ;
  assign y12214 = n45213 ;
  assign y12215 = ~1'b0 ;
  assign y12216 = ~1'b0 ;
  assign y12217 = ~1'b0 ;
  assign y12218 = n45219 ;
  assign y12219 = ~n45221 ;
  assign y12220 = ~n45222 ;
  assign y12221 = n45224 ;
  assign y12222 = n45230 ;
  assign y12223 = n45231 ;
  assign y12224 = n45233 ;
  assign y12225 = ~n45237 ;
  assign y12226 = ~n45247 ;
  assign y12227 = n45250 ;
  assign y12228 = n45253 ;
  assign y12229 = n45254 ;
  assign y12230 = ~n45256 ;
  assign y12231 = n45258 ;
  assign y12232 = ~n45260 ;
  assign y12233 = n45268 ;
  assign y12234 = ~n45272 ;
  assign y12235 = ~n45273 ;
  assign y12236 = ~n45278 ;
  assign y12237 = ~n45280 ;
  assign y12238 = ~1'b0 ;
  assign y12239 = n45282 ;
  assign y12240 = ~n45283 ;
  assign y12241 = ~n45284 ;
  assign y12242 = ~n45285 ;
  assign y12243 = ~n45287 ;
  assign y12244 = ~n45290 ;
  assign y12245 = n45295 ;
  assign y12246 = ~n45296 ;
  assign y12247 = ~n45300 ;
  assign y12248 = ~1'b0 ;
  assign y12249 = ~1'b0 ;
  assign y12250 = n45311 ;
  assign y12251 = ~n45313 ;
  assign y12252 = ~n45316 ;
  assign y12253 = n45318 ;
  assign y12254 = ~n45323 ;
  assign y12255 = ~1'b0 ;
  assign y12256 = ~n45325 ;
  assign y12257 = n45328 ;
  assign y12258 = n45330 ;
  assign y12259 = ~n45332 ;
  assign y12260 = ~n45333 ;
  assign y12261 = ~n45338 ;
  assign y12262 = ~1'b0 ;
  assign y12263 = ~n45341 ;
  assign y12264 = n45343 ;
  assign y12265 = ~n45346 ;
  assign y12266 = ~n45348 ;
  assign y12267 = n45355 ;
  assign y12268 = ~n45358 ;
  assign y12269 = n45359 ;
  assign y12270 = ~n45365 ;
  assign y12271 = ~1'b0 ;
  assign y12272 = n45370 ;
  assign y12273 = n45381 ;
  assign y12274 = n45382 ;
  assign y12275 = n45385 ;
  assign y12276 = ~n45386 ;
  assign y12277 = ~n45389 ;
  assign y12278 = n45392 ;
  assign y12279 = ~n45395 ;
  assign y12280 = ~n45397 ;
  assign y12281 = ~n45398 ;
  assign y12282 = n45401 ;
  assign y12283 = n45402 ;
  assign y12284 = n45405 ;
  assign y12285 = ~n45408 ;
  assign y12286 = ~n45412 ;
  assign y12287 = ~n45413 ;
  assign y12288 = n45415 ;
  assign y12289 = n45417 ;
  assign y12290 = n45420 ;
  assign y12291 = n45421 ;
  assign y12292 = ~n45422 ;
  assign y12293 = ~n45426 ;
  assign y12294 = ~n45427 ;
  assign y12295 = n45430 ;
  assign y12296 = ~n45431 ;
  assign y12297 = n45438 ;
  assign y12298 = n45441 ;
  assign y12299 = ~n45444 ;
  assign y12300 = n45445 ;
  assign y12301 = ~n45446 ;
  assign y12302 = n45453 ;
  assign y12303 = ~n45454 ;
  assign y12304 = n45455 ;
  assign y12305 = ~n45458 ;
  assign y12306 = ~1'b0 ;
  assign y12307 = ~n45460 ;
  assign y12308 = ~n45463 ;
  assign y12309 = ~n45464 ;
  assign y12310 = ~n45466 ;
  assign y12311 = n45469 ;
  assign y12312 = n45476 ;
  assign y12313 = ~n45478 ;
  assign y12314 = ~n45481 ;
  assign y12315 = n45484 ;
  assign y12316 = n45486 ;
  assign y12317 = n45488 ;
  assign y12318 = ~n45490 ;
  assign y12319 = ~1'b0 ;
  assign y12320 = ~n45492 ;
  assign y12321 = ~n45493 ;
  assign y12322 = n45494 ;
  assign y12323 = n45496 ;
  assign y12324 = n45502 ;
  assign y12325 = ~n45505 ;
  assign y12326 = n45506 ;
  assign y12327 = n45511 ;
  assign y12328 = ~n45514 ;
  assign y12329 = n45515 ;
  assign y12330 = ~n45516 ;
  assign y12331 = n45520 ;
  assign y12332 = n45521 ;
  assign y12333 = ~n45529 ;
  assign y12334 = n45530 ;
  assign y12335 = ~n45532 ;
  assign y12336 = n45535 ;
  assign y12337 = ~n45536 ;
  assign y12338 = n45537 ;
  assign y12339 = ~n45540 ;
  assign y12340 = n45545 ;
  assign y12341 = ~n45548 ;
  assign y12342 = ~n45550 ;
  assign y12343 = ~n45557 ;
  assign y12344 = n45561 ;
  assign y12345 = ~n45565 ;
  assign y12346 = ~n45566 ;
  assign y12347 = n45569 ;
  assign y12348 = n45573 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = ~n45575 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = ~n45578 ;
  assign y12353 = n45582 ;
  assign y12354 = n45585 ;
  assign y12355 = ~n45586 ;
  assign y12356 = ~n45587 ;
  assign y12357 = n45589 ;
  assign y12358 = ~n45591 ;
  assign y12359 = n45593 ;
  assign y12360 = n45594 ;
  assign y12361 = n45598 ;
  assign y12362 = ~n45601 ;
  assign y12363 = n45602 ;
  assign y12364 = n45604 ;
  assign y12365 = ~n45607 ;
  assign y12366 = n45609 ;
  assign y12367 = ~1'b0 ;
  assign y12368 = n45613 ;
  assign y12369 = ~n45614 ;
  assign y12370 = n45617 ;
  assign y12371 = ~n45620 ;
  assign y12372 = ~n45622 ;
  assign y12373 = n45623 ;
  assign y12374 = n45624 ;
  assign y12375 = n45625 ;
  assign y12376 = ~n45626 ;
  assign y12377 = ~1'b0 ;
  assign y12378 = n45627 ;
  assign y12379 = n45631 ;
  assign y12380 = n45633 ;
  assign y12381 = ~n45636 ;
  assign y12382 = ~n45639 ;
  assign y12383 = n45641 ;
  assign y12384 = ~n45646 ;
  assign y12385 = ~n45647 ;
  assign y12386 = ~n45650 ;
  assign y12387 = ~n45654 ;
  assign y12388 = ~n45655 ;
  assign y12389 = ~n45658 ;
  assign y12390 = n45661 ;
  assign y12391 = n45665 ;
  assign y12392 = ~n45669 ;
  assign y12393 = n45670 ;
  assign y12394 = n45671 ;
  assign y12395 = n45680 ;
  assign y12396 = ~n45681 ;
  assign y12397 = ~n45682 ;
  assign y12398 = ~n45684 ;
  assign y12399 = n45688 ;
  assign y12400 = ~n45690 ;
  assign y12401 = ~n45692 ;
  assign y12402 = ~n45695 ;
  assign y12403 = ~n45696 ;
  assign y12404 = n45697 ;
  assign y12405 = ~n45699 ;
  assign y12406 = ~n45702 ;
  assign y12407 = ~n45704 ;
  assign y12408 = n45705 ;
  assign y12409 = n45709 ;
  assign y12410 = ~n45713 ;
  assign y12411 = n45715 ;
  assign y12412 = ~n45721 ;
  assign y12413 = n45724 ;
  assign y12414 = ~n45726 ;
  assign y12415 = ~n45727 ;
  assign y12416 = ~1'b0 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = ~n45730 ;
  assign y12419 = ~n45732 ;
  assign y12420 = ~n45735 ;
  assign y12421 = n45736 ;
  assign y12422 = n45738 ;
  assign y12423 = n45740 ;
  assign y12424 = ~n45742 ;
  assign y12425 = n45744 ;
  assign y12426 = ~1'b0 ;
  assign y12427 = n45745 ;
  assign y12428 = n45746 ;
  assign y12429 = n45756 ;
  assign y12430 = ~n45757 ;
  assign y12431 = ~n45759 ;
  assign y12432 = ~n45760 ;
  assign y12433 = n45762 ;
  assign y12434 = ~1'b0 ;
  assign y12435 = n45764 ;
  assign y12436 = ~n45765 ;
  assign y12437 = n45770 ;
  assign y12438 = ~n45777 ;
  assign y12439 = n45778 ;
  assign y12440 = n45780 ;
  assign y12441 = ~n45782 ;
  assign y12442 = ~n45783 ;
  assign y12443 = n45787 ;
  assign y12444 = ~n45791 ;
  assign y12445 = ~n45792 ;
  assign y12446 = n45793 ;
  assign y12447 = n45794 ;
  assign y12448 = n45795 ;
  assign y12449 = ~n45797 ;
  assign y12450 = ~n45799 ;
  assign y12451 = ~n45801 ;
  assign y12452 = n45803 ;
  assign y12453 = ~n45804 ;
  assign y12454 = n45809 ;
  assign y12455 = ~n45811 ;
  assign y12456 = ~n45818 ;
  assign y12457 = n45821 ;
  assign y12458 = n45823 ;
  assign y12459 = ~1'b0 ;
  assign y12460 = ~n45824 ;
  assign y12461 = ~n45827 ;
  assign y12462 = n45830 ;
  assign y12463 = ~n45832 ;
  assign y12464 = ~n45834 ;
  assign y12465 = n45836 ;
  assign y12466 = n45838 ;
  assign y12467 = n45840 ;
  assign y12468 = ~n45844 ;
  assign y12469 = n45845 ;
  assign y12470 = n45848 ;
  assign y12471 = n45849 ;
  assign y12472 = n45850 ;
  assign y12473 = ~n45853 ;
  assign y12474 = ~n45856 ;
  assign y12475 = n45859 ;
  assign y12476 = ~n45861 ;
  assign y12477 = ~n45862 ;
  assign y12478 = n45865 ;
  assign y12479 = n45869 ;
  assign y12480 = n45874 ;
  assign y12481 = n45875 ;
  assign y12482 = ~n45881 ;
  assign y12483 = ~n45883 ;
  assign y12484 = ~1'b0 ;
  assign y12485 = ~n45885 ;
  assign y12486 = ~n45886 ;
  assign y12487 = n45890 ;
  assign y12488 = n45891 ;
  assign y12489 = n45893 ;
  assign y12490 = ~n45895 ;
  assign y12491 = n45899 ;
  assign y12492 = ~1'b0 ;
  assign y12493 = n45904 ;
  assign y12494 = n45906 ;
  assign y12495 = ~n45907 ;
  assign y12496 = n45912 ;
  assign y12497 = n45917 ;
  assign y12498 = ~n45920 ;
  assign y12499 = ~1'b0 ;
  assign y12500 = n45922 ;
  assign y12501 = n45924 ;
  assign y12502 = n45926 ;
  assign y12503 = n45928 ;
  assign y12504 = ~n45929 ;
  assign y12505 = ~n45931 ;
  assign y12506 = n45935 ;
  assign y12507 = n45939 ;
  assign y12508 = n45941 ;
  assign y12509 = ~1'b0 ;
  assign y12510 = ~1'b0 ;
  assign y12511 = n45942 ;
  assign y12512 = n45943 ;
  assign y12513 = ~n45948 ;
  assign y12514 = ~n45949 ;
  assign y12515 = n45954 ;
  assign y12516 = n45957 ;
  assign y12517 = ~n45963 ;
  assign y12518 = n45966 ;
  assign y12519 = ~n45969 ;
  assign y12520 = n45970 ;
  assign y12521 = ~n45971 ;
  assign y12522 = ~n45972 ;
  assign y12523 = n45974 ;
  assign y12524 = ~n45979 ;
  assign y12525 = n45981 ;
  assign y12526 = ~n45983 ;
  assign y12527 = ~n45985 ;
  assign y12528 = ~n45995 ;
  assign y12529 = ~n45996 ;
  assign y12530 = n45997 ;
  assign y12531 = ~n46002 ;
  assign y12532 = n46007 ;
  assign y12533 = n46012 ;
  assign y12534 = n46016 ;
  assign y12535 = ~n46021 ;
  assign y12536 = n46023 ;
  assign y12537 = ~n46024 ;
  assign y12538 = n46028 ;
  assign y12539 = ~n46030 ;
  assign y12540 = ~n46035 ;
  assign y12541 = n46036 ;
  assign y12542 = ~n46040 ;
  assign y12543 = ~n46041 ;
  assign y12544 = ~n46046 ;
  assign y12545 = n46053 ;
  assign y12546 = ~n46055 ;
  assign y12547 = ~n46057 ;
  assign y12548 = n46058 ;
  assign y12549 = ~n46059 ;
  assign y12550 = ~n46061 ;
  assign y12551 = ~n46064 ;
  assign y12552 = ~n46070 ;
  assign y12553 = n46073 ;
  assign y12554 = n46074 ;
  assign y12555 = ~n46079 ;
  assign y12556 = ~n46080 ;
  assign y12557 = n46082 ;
  assign y12558 = n46084 ;
  assign y12559 = n46086 ;
  assign y12560 = n46088 ;
  assign y12561 = ~n46092 ;
  assign y12562 = n46093 ;
  assign y12563 = n46094 ;
  assign y12564 = ~n46095 ;
  assign y12565 = ~n46096 ;
  assign y12566 = n46098 ;
  assign y12567 = ~n46099 ;
  assign y12568 = n46100 ;
  assign y12569 = ~n46105 ;
  assign y12570 = n46109 ;
  assign y12571 = ~1'b0 ;
  assign y12572 = ~n46111 ;
  assign y12573 = ~n46114 ;
  assign y12574 = ~n46116 ;
  assign y12575 = ~n46119 ;
  assign y12576 = ~n46120 ;
  assign y12577 = ~n46123 ;
  assign y12578 = ~n46124 ;
  assign y12579 = ~1'b0 ;
  assign y12580 = ~1'b0 ;
  assign y12581 = n46126 ;
  assign y12582 = n15742 ;
  assign y12583 = ~n46130 ;
  assign y12584 = n46132 ;
  assign y12585 = ~n46133 ;
  assign y12586 = ~n46134 ;
  assign y12587 = n46139 ;
  assign y12588 = ~n46141 ;
  assign y12589 = ~n46144 ;
  assign y12590 = n46145 ;
  assign y12591 = n46146 ;
  assign y12592 = ~n46147 ;
  assign y12593 = n46148 ;
  assign y12594 = ~n46149 ;
  assign y12595 = n46150 ;
  assign y12596 = ~n46151 ;
  assign y12597 = ~1'b0 ;
  assign y12598 = ~n46155 ;
  assign y12599 = ~n46157 ;
  assign y12600 = ~n46160 ;
  assign y12601 = ~n46165 ;
  assign y12602 = ~n46166 ;
  assign y12603 = n46170 ;
  assign y12604 = ~n46171 ;
  assign y12605 = n46172 ;
  assign y12606 = n46173 ;
  assign y12607 = ~1'b0 ;
  assign y12608 = ~n46177 ;
  assign y12609 = ~1'b0 ;
  assign y12610 = ~n46179 ;
  assign y12611 = n46182 ;
  assign y12612 = n46184 ;
  assign y12613 = ~1'b0 ;
  assign y12614 = ~n46186 ;
  assign y12615 = n46189 ;
  assign y12616 = n46191 ;
  assign y12617 = ~n46193 ;
  assign y12618 = n46195 ;
  assign y12619 = n46196 ;
  assign y12620 = ~n46199 ;
  assign y12621 = n46200 ;
  assign y12622 = n46201 ;
  assign y12623 = n46203 ;
  assign y12624 = ~n46205 ;
  assign y12625 = n46208 ;
  assign y12626 = ~1'b0 ;
  assign y12627 = ~n46212 ;
  assign y12628 = n46214 ;
  assign y12629 = n46217 ;
  assign y12630 = n46219 ;
  assign y12631 = ~n46228 ;
  assign y12632 = n46230 ;
  assign y12633 = ~n46232 ;
  assign y12634 = ~1'b0 ;
  assign y12635 = ~n46234 ;
  assign y12636 = ~n46238 ;
  assign y12637 = n46241 ;
  assign y12638 = n46245 ;
  assign y12639 = n46250 ;
  assign y12640 = ~n46251 ;
  assign y12641 = ~n46252 ;
  assign y12642 = ~n46254 ;
  assign y12643 = ~1'b0 ;
  assign y12644 = ~n46255 ;
  assign y12645 = ~n46256 ;
  assign y12646 = ~n46261 ;
  assign y12647 = ~n46262 ;
  assign y12648 = ~n46263 ;
  assign y12649 = ~n46270 ;
  assign y12650 = n46271 ;
  assign y12651 = ~1'b0 ;
  assign y12652 = ~n46272 ;
  assign y12653 = ~n46276 ;
  assign y12654 = ~n46277 ;
  assign y12655 = n46282 ;
  assign y12656 = n46283 ;
  assign y12657 = n46285 ;
  assign y12658 = ~n46288 ;
  assign y12659 = ~n46291 ;
  assign y12660 = ~n46293 ;
  assign y12661 = ~n46295 ;
  assign y12662 = ~1'b0 ;
  assign y12663 = ~1'b0 ;
  assign y12664 = n46297 ;
  assign y12665 = ~n46300 ;
  assign y12666 = ~n46301 ;
  assign y12667 = n46304 ;
  assign y12668 = n46312 ;
  assign y12669 = n46313 ;
  assign y12670 = n46315 ;
  assign y12671 = n46316 ;
  assign y12672 = ~1'b0 ;
  assign y12673 = ~n46319 ;
  assign y12674 = ~n46322 ;
  assign y12675 = ~n46324 ;
  assign y12676 = n46327 ;
  assign y12677 = ~n46328 ;
  assign y12678 = ~n46330 ;
  assign y12679 = ~n46332 ;
  assign y12680 = ~n46334 ;
  assign y12681 = ~n46337 ;
  assign y12682 = ~n46339 ;
  assign y12683 = ~n46340 ;
  assign y12684 = n46342 ;
  assign y12685 = n46344 ;
  assign y12686 = n46346 ;
  assign y12687 = n46347 ;
  assign y12688 = ~n46348 ;
  assign y12689 = ~1'b0 ;
  assign y12690 = ~n46349 ;
  assign y12691 = n46353 ;
  assign y12692 = n46354 ;
  assign y12693 = n46358 ;
  assign y12694 = ~n46359 ;
  assign y12695 = ~n46360 ;
  assign y12696 = ~n46362 ;
  assign y12697 = ~n46364 ;
  assign y12698 = ~1'b0 ;
  assign y12699 = ~1'b0 ;
  assign y12700 = n46365 ;
  assign y12701 = ~n46367 ;
  assign y12702 = ~n46369 ;
  assign y12703 = n46370 ;
  assign y12704 = ~n46372 ;
  assign y12705 = n46373 ;
  assign y12706 = ~n46375 ;
  assign y12707 = ~1'b0 ;
  assign y12708 = n46376 ;
  assign y12709 = ~n46377 ;
  assign y12710 = ~n46382 ;
  assign y12711 = ~n46384 ;
  assign y12712 = n46385 ;
  assign y12713 = ~n46388 ;
  assign y12714 = n46391 ;
  assign y12715 = ~n46392 ;
  assign y12716 = ~n46393 ;
  assign y12717 = ~n46399 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = ~n46401 ;
  assign y12720 = n46404 ;
  assign y12721 = n46406 ;
  assign y12722 = ~n46411 ;
  assign y12723 = n46412 ;
  assign y12724 = ~n46417 ;
  assign y12725 = ~1'b0 ;
  assign y12726 = n46419 ;
  assign y12727 = n46421 ;
  assign y12728 = n46423 ;
  assign y12729 = n46425 ;
  assign y12730 = n46428 ;
  assign y12731 = n46429 ;
  assign y12732 = n46433 ;
  assign y12733 = ~n46437 ;
  assign y12734 = ~n46439 ;
  assign y12735 = n46441 ;
  assign y12736 = ~n46442 ;
  assign y12737 = ~n46443 ;
  assign y12738 = n46448 ;
  assign y12739 = ~n46451 ;
  assign y12740 = ~n46452 ;
  assign y12741 = ~n46454 ;
  assign y12742 = ~n46455 ;
  assign y12743 = ~1'b0 ;
  assign y12744 = n46458 ;
  assign y12745 = n46466 ;
  assign y12746 = ~n46467 ;
  assign y12747 = n46469 ;
  assign y12748 = ~n46470 ;
  assign y12749 = ~n46473 ;
  assign y12750 = ~n46475 ;
  assign y12751 = n46488 ;
  assign y12752 = n46491 ;
  assign y12753 = ~1'b0 ;
  assign y12754 = n46499 ;
  assign y12755 = n46504 ;
  assign y12756 = ~n46509 ;
  assign y12757 = n46513 ;
  assign y12758 = n46517 ;
  assign y12759 = ~n46525 ;
  assign y12760 = ~n46527 ;
  assign y12761 = ~n46529 ;
  assign y12762 = n46531 ;
  assign y12763 = n46534 ;
  assign y12764 = ~n46539 ;
  assign y12765 = ~n46540 ;
  assign y12766 = n46541 ;
  assign y12767 = n46549 ;
  assign y12768 = n46551 ;
  assign y12769 = ~n46557 ;
  assign y12770 = n46559 ;
  assign y12771 = n46561 ;
  assign y12772 = ~n46571 ;
  assign y12773 = n46574 ;
  assign y12774 = n46575 ;
  assign y12775 = n46577 ;
  assign y12776 = ~n46578 ;
  assign y12777 = ~n46580 ;
  assign y12778 = n46581 ;
  assign y12779 = ~n46583 ;
  assign y12780 = n46585 ;
  assign y12781 = ~n46588 ;
  assign y12782 = n46596 ;
  assign y12783 = n46603 ;
  assign y12784 = ~n46605 ;
  assign y12785 = n46606 ;
  assign y12786 = n46607 ;
  assign y12787 = n46611 ;
  assign y12788 = n46612 ;
  assign y12789 = n46614 ;
  assign y12790 = n46621 ;
  assign y12791 = n46622 ;
  assign y12792 = ~n46627 ;
  assign y12793 = n3131 ;
  assign y12794 = n46631 ;
  assign y12795 = ~n46633 ;
  assign y12796 = n46635 ;
  assign y12797 = ~n46637 ;
  assign y12798 = ~n46640 ;
  assign y12799 = n46641 ;
  assign y12800 = ~n46645 ;
  assign y12801 = n46649 ;
  assign y12802 = n46651 ;
  assign y12803 = ~n46654 ;
  assign y12804 = ~n46657 ;
  assign y12805 = ~n46661 ;
  assign y12806 = ~1'b0 ;
  assign y12807 = ~n46665 ;
  assign y12808 = n46667 ;
  assign y12809 = n46671 ;
  assign y12810 = n46673 ;
  assign y12811 = ~n46674 ;
  assign y12812 = ~n46676 ;
  assign y12813 = ~n46679 ;
  assign y12814 = n46681 ;
  assign y12815 = n46683 ;
  assign y12816 = ~n46685 ;
  assign y12817 = ~n46688 ;
  assign y12818 = n46690 ;
  assign y12819 = n46693 ;
  assign y12820 = n46694 ;
  assign y12821 = ~n46696 ;
  assign y12822 = ~n46703 ;
  assign y12823 = n46706 ;
  assign y12824 = ~n46708 ;
  assign y12825 = ~n46709 ;
  assign y12826 = ~n46710 ;
  assign y12827 = ~n46712 ;
  assign y12828 = ~n46713 ;
  assign y12829 = n46714 ;
  assign y12830 = ~1'b0 ;
  assign y12831 = ~1'b0 ;
  assign y12832 = ~n46726 ;
  assign y12833 = n46727 ;
  assign y12834 = ~n46728 ;
  assign y12835 = n46729 ;
  assign y12836 = ~n46732 ;
  assign y12837 = n46733 ;
  assign y12838 = ~n46735 ;
  assign y12839 = ~n46737 ;
  assign y12840 = n46740 ;
  assign y12841 = ~n46744 ;
  assign y12842 = ~n46749 ;
  assign y12843 = ~n46756 ;
  assign y12844 = ~n46761 ;
  assign y12845 = n46762 ;
  assign y12846 = ~n46763 ;
  assign y12847 = ~n46765 ;
  assign y12848 = ~n46768 ;
  assign y12849 = n46770 ;
  assign y12850 = n46774 ;
  assign y12851 = n46778 ;
  assign y12852 = n46781 ;
  assign y12853 = n46783 ;
  assign y12854 = n46784 ;
  assign y12855 = ~n46786 ;
  assign y12856 = ~n46788 ;
  assign y12857 = n46793 ;
  assign y12858 = ~n46801 ;
  assign y12859 = ~n46804 ;
  assign y12860 = ~n46808 ;
  assign y12861 = n46809 ;
  assign y12862 = n46815 ;
  assign y12863 = ~n46819 ;
  assign y12864 = ~n46821 ;
  assign y12865 = ~n46822 ;
  assign y12866 = n46825 ;
  assign y12867 = n46828 ;
  assign y12868 = ~n46831 ;
  assign y12869 = ~n46833 ;
  assign y12870 = n46834 ;
  assign y12871 = ~n46836 ;
  assign y12872 = n46838 ;
  assign y12873 = ~1'b0 ;
  assign y12874 = ~n46840 ;
  assign y12875 = ~n46844 ;
  assign y12876 = ~n46847 ;
  assign y12877 = n46852 ;
  assign y12878 = ~n46857 ;
  assign y12879 = ~n46858 ;
  assign y12880 = ~n46860 ;
  assign y12881 = n46862 ;
  assign y12882 = ~n46864 ;
  assign y12883 = ~n46868 ;
  assign y12884 = n46872 ;
  assign y12885 = n46876 ;
  assign y12886 = n46877 ;
  assign y12887 = n46882 ;
  assign y12888 = n46885 ;
  assign y12889 = n46888 ;
  assign y12890 = n46890 ;
  assign y12891 = n46894 ;
  assign y12892 = n46895 ;
  assign y12893 = ~n46896 ;
  assign y12894 = ~n46899 ;
  assign y12895 = ~n46903 ;
  assign y12896 = ~n46904 ;
  assign y12897 = n46905 ;
  assign y12898 = n46907 ;
  assign y12899 = n46911 ;
  assign y12900 = n46913 ;
  assign y12901 = ~n46917 ;
  assign y12902 = n46920 ;
  assign y12903 = n46924 ;
  assign y12904 = ~n46927 ;
  assign y12905 = ~n46928 ;
  assign y12906 = ~n46930 ;
  assign y12907 = ~n46931 ;
  assign y12908 = n46932 ;
  assign y12909 = n46934 ;
  assign y12910 = ~n46935 ;
  assign y12911 = ~n46940 ;
  assign y12912 = n46943 ;
  assign y12913 = n46946 ;
  assign y12914 = ~n46950 ;
  assign y12915 = n46952 ;
  assign y12916 = ~n46953 ;
  assign y12917 = ~n46954 ;
  assign y12918 = n46959 ;
  assign y12919 = n46960 ;
  assign y12920 = ~n46964 ;
  assign y12921 = ~1'b0 ;
  assign y12922 = n46966 ;
  assign y12923 = n46967 ;
  assign y12924 = ~n46971 ;
  assign y12925 = ~n46974 ;
  assign y12926 = n46976 ;
  assign y12927 = n46979 ;
  assign y12928 = ~n46982 ;
  assign y12929 = ~n46987 ;
  assign y12930 = n46990 ;
  assign y12931 = n46992 ;
  assign y12932 = n46994 ;
  assign y12933 = n46995 ;
  assign y12934 = n46997 ;
  assign y12935 = ~n46999 ;
  assign y12936 = n47000 ;
  assign y12937 = ~n47002 ;
  assign y12938 = ~n47003 ;
  assign y12939 = ~n47006 ;
  assign y12940 = ~n47008 ;
  assign y12941 = ~1'b0 ;
  assign y12942 = ~1'b0 ;
  assign y12943 = ~n47010 ;
  assign y12944 = n47013 ;
  assign y12945 = ~n47015 ;
  assign y12946 = n47020 ;
  assign y12947 = n47022 ;
  assign y12948 = ~n47032 ;
  assign y12949 = n47037 ;
  assign y12950 = ~n47038 ;
  assign y12951 = ~1'b0 ;
  assign y12952 = n47039 ;
  assign y12953 = n47042 ;
  assign y12954 = n47044 ;
  assign y12955 = ~n47046 ;
  assign y12956 = n47051 ;
  assign y12957 = n47059 ;
  assign y12958 = n47062 ;
  assign y12959 = ~n47063 ;
  assign y12960 = n47069 ;
  assign y12961 = n47072 ;
  assign y12962 = n47074 ;
  assign y12963 = ~n47075 ;
  assign y12964 = ~n47077 ;
  assign y12965 = ~n47078 ;
  assign y12966 = n47080 ;
  assign y12967 = ~n47081 ;
  assign y12968 = n47086 ;
  assign y12969 = ~n47088 ;
  assign y12970 = n47090 ;
  assign y12971 = n47093 ;
  assign y12972 = ~n47100 ;
  assign y12973 = ~n47105 ;
  assign y12974 = ~n47109 ;
  assign y12975 = n47112 ;
  assign y12976 = ~n47117 ;
  assign y12977 = ~n47129 ;
  assign y12978 = ~n47135 ;
  assign y12979 = ~n47136 ;
  assign y12980 = ~n47139 ;
  assign y12981 = ~n47147 ;
  assign y12982 = ~n47149 ;
  assign y12983 = ~n47152 ;
  assign y12984 = n47157 ;
  assign y12985 = n47160 ;
  assign y12986 = n47161 ;
  assign y12987 = ~n47173 ;
  assign y12988 = ~n47175 ;
  assign y12989 = n47177 ;
  assign y12990 = n47181 ;
  assign y12991 = ~n47182 ;
  assign y12992 = ~n47184 ;
  assign y12993 = ~n47187 ;
  assign y12994 = n47189 ;
  assign y12995 = ~n47190 ;
  assign y12996 = n47191 ;
  assign y12997 = n47197 ;
  assign y12998 = n47198 ;
  assign y12999 = n47199 ;
  assign y13000 = n47201 ;
  assign y13001 = n47203 ;
  assign y13002 = n47205 ;
  assign y13003 = ~n47207 ;
  assign y13004 = ~1'b0 ;
  assign y13005 = ~n47210 ;
  assign y13006 = ~n47212 ;
  assign y13007 = ~n47215 ;
  assign y13008 = n47216 ;
  assign y13009 = n47220 ;
  assign y13010 = n47222 ;
  assign y13011 = ~n47229 ;
  assign y13012 = ~1'b0 ;
  assign y13013 = n47232 ;
  assign y13014 = ~n47238 ;
  assign y13015 = ~n47242 ;
  assign y13016 = ~n47243 ;
  assign y13017 = n47252 ;
  assign y13018 = n47253 ;
  assign y13019 = ~n47254 ;
  assign y13020 = n47256 ;
  assign y13021 = n47258 ;
  assign y13022 = n47260 ;
  assign y13023 = ~n47262 ;
  assign y13024 = ~n47263 ;
  assign y13025 = ~n47264 ;
  assign y13026 = ~n47265 ;
  assign y13027 = n47266 ;
  assign y13028 = ~n47267 ;
  assign y13029 = n47268 ;
  assign y13030 = n47271 ;
  assign y13031 = ~n47275 ;
  assign y13032 = ~1'b0 ;
  assign y13033 = ~n47279 ;
  assign y13034 = ~n47280 ;
  assign y13035 = n47283 ;
  assign y13036 = n47286 ;
  assign y13037 = ~n47287 ;
  assign y13038 = ~1'b0 ;
  assign y13039 = ~n47289 ;
  assign y13040 = n47290 ;
  assign y13041 = n47291 ;
  assign y13042 = n47294 ;
  assign y13043 = n47296 ;
  assign y13044 = ~n47298 ;
  assign y13045 = ~n47300 ;
  assign y13046 = ~n47301 ;
  assign y13047 = ~1'b0 ;
  assign y13048 = ~1'b0 ;
  assign y13049 = ~n47302 ;
  assign y13050 = ~n47308 ;
  assign y13051 = ~n47310 ;
  assign y13052 = ~n47315 ;
  assign y13053 = n47321 ;
  assign y13054 = ~n47325 ;
  assign y13055 = n47329 ;
  assign y13056 = n47333 ;
  assign y13057 = ~n47337 ;
  assign y13058 = ~n47338 ;
  assign y13059 = ~n47339 ;
  assign y13060 = ~n47342 ;
  assign y13061 = ~n47343 ;
  assign y13062 = ~n47345 ;
  assign y13063 = ~n47346 ;
  assign y13064 = ~n47348 ;
  assign y13065 = ~n47349 ;
  assign y13066 = ~1'b0 ;
  assign y13067 = n47351 ;
  assign y13068 = ~n47355 ;
  assign y13069 = ~n47358 ;
  assign y13070 = ~n47360 ;
  assign y13071 = n47361 ;
  assign y13072 = n47364 ;
  assign y13073 = ~n47366 ;
  assign y13074 = ~1'b0 ;
  assign y13075 = ~n47367 ;
  assign y13076 = n47371 ;
  assign y13077 = n47372 ;
  assign y13078 = ~n47376 ;
  assign y13079 = ~n47378 ;
  assign y13080 = n47379 ;
  assign y13081 = ~n47380 ;
  assign y13082 = ~1'b0 ;
  assign y13083 = ~n47383 ;
  assign y13084 = ~n47387 ;
  assign y13085 = ~n47388 ;
  assign y13086 = ~n47391 ;
  assign y13087 = ~n47392 ;
  assign y13088 = ~n47395 ;
  assign y13089 = ~n47397 ;
  assign y13090 = n47399 ;
  assign y13091 = n47400 ;
  assign y13092 = ~1'b0 ;
  assign y13093 = ~n47401 ;
  assign y13094 = ~1'b0 ;
  assign y13095 = n47402 ;
  assign y13096 = n47405 ;
  assign y13097 = ~n47406 ;
  assign y13098 = n47408 ;
  assign y13099 = ~n47411 ;
  assign y13100 = n47413 ;
  assign y13101 = ~n47421 ;
  assign y13102 = n47426 ;
  assign y13103 = ~n47427 ;
  assign y13104 = ~n47428 ;
  assign y13105 = ~n47430 ;
  assign y13106 = n47434 ;
  assign y13107 = ~n47444 ;
  assign y13108 = ~n47447 ;
  assign y13109 = ~n47448 ;
  assign y13110 = ~n47452 ;
  assign y13111 = n47454 ;
  assign y13112 = n47458 ;
  assign y13113 = ~n47466 ;
  assign y13114 = ~n47469 ;
  assign y13115 = ~n47470 ;
  assign y13116 = n47473 ;
  assign y13117 = ~1'b0 ;
  assign y13118 = n47475 ;
  assign y13119 = ~n47479 ;
  assign y13120 = n47480 ;
  assign y13121 = n47481 ;
  assign y13122 = ~n47483 ;
  assign y13123 = ~n47485 ;
  assign y13124 = ~1'b0 ;
  assign y13125 = ~n47488 ;
  assign y13126 = ~1'b0 ;
  assign y13127 = n47489 ;
  assign y13128 = n47490 ;
  assign y13129 = n47491 ;
  assign y13130 = ~n47492 ;
  assign y13131 = n47493 ;
  assign y13132 = ~n47496 ;
  assign y13133 = n47501 ;
  assign y13134 = ~n47505 ;
  assign y13135 = ~1'b0 ;
  assign y13136 = n47506 ;
  assign y13137 = ~n47507 ;
  assign y13138 = ~n47508 ;
  assign y13139 = ~n47509 ;
  assign y13140 = ~n47510 ;
  assign y13141 = n47511 ;
  assign y13142 = n47515 ;
  assign y13143 = n47518 ;
  assign y13144 = ~n47520 ;
  assign y13145 = ~1'b0 ;
  assign y13146 = n47534 ;
  assign y13147 = ~n47535 ;
  assign y13148 = ~n47538 ;
  assign y13149 = ~n47542 ;
  assign y13150 = ~1'b0 ;
  assign y13151 = ~1'b0 ;
  assign y13152 = n47544 ;
  assign y13153 = n47545 ;
  assign y13154 = ~n47546 ;
  assign y13155 = ~n47547 ;
  assign y13156 = n47548 ;
  assign y13157 = ~n47549 ;
  assign y13158 = n47552 ;
  assign y13159 = ~n47557 ;
  assign y13160 = ~n47559 ;
  assign y13161 = n47560 ;
  assign y13162 = n47561 ;
  assign y13163 = ~n47562 ;
  assign y13164 = n47565 ;
  assign y13165 = ~n47567 ;
  assign y13166 = n47571 ;
  assign y13167 = n47572 ;
  assign y13168 = ~n47574 ;
  assign y13169 = ~1'b0 ;
  assign y13170 = ~1'b0 ;
  assign y13171 = ~1'b0 ;
  assign y13172 = ~n47575 ;
  assign y13173 = n47576 ;
  assign y13174 = ~n47579 ;
  assign y13175 = ~n47581 ;
  assign y13176 = n47583 ;
  assign y13177 = n47587 ;
  assign y13178 = ~n47590 ;
  assign y13179 = ~n47591 ;
  assign y13180 = n47592 ;
  assign y13181 = n47596 ;
  assign y13182 = ~n47597 ;
  assign y13183 = n47601 ;
  assign y13184 = ~n36422 ;
  assign y13185 = ~n47603 ;
  assign y13186 = n47604 ;
  assign y13187 = n47610 ;
  assign y13188 = ~n47612 ;
  assign y13189 = n47613 ;
  assign y13190 = ~n47615 ;
  assign y13191 = n47617 ;
  assign y13192 = n47618 ;
  assign y13193 = n47622 ;
  assign y13194 = n47623 ;
  assign y13195 = ~n47632 ;
  assign y13196 = ~n47633 ;
  assign y13197 = n47636 ;
  assign y13198 = ~n47637 ;
  assign y13199 = ~1'b0 ;
  assign y13200 = ~n47639 ;
  assign y13201 = ~n47642 ;
  assign y13202 = ~n47643 ;
  assign y13203 = ~n47647 ;
  assign y13204 = n47654 ;
  assign y13205 = ~n47656 ;
  assign y13206 = ~n47661 ;
  assign y13207 = ~n47662 ;
  assign y13208 = ~n47668 ;
  assign y13209 = ~n47674 ;
  assign y13210 = ~n47677 ;
  assign y13211 = ~1'b0 ;
  assign y13212 = ~n47678 ;
  assign y13213 = ~n47679 ;
  assign y13214 = ~n47680 ;
  assign y13215 = ~n47684 ;
  assign y13216 = ~n47685 ;
  assign y13217 = ~n47689 ;
  assign y13218 = n47691 ;
  assign y13219 = ~n47692 ;
  assign y13220 = n47693 ;
  assign y13221 = ~n47697 ;
  assign y13222 = ~n47698 ;
  assign y13223 = ~n47700 ;
  assign y13224 = n47703 ;
  assign y13225 = ~n47706 ;
  assign y13226 = ~1'b0 ;
  assign y13227 = ~n47709 ;
  assign y13228 = ~n47713 ;
  assign y13229 = ~n47717 ;
  assign y13230 = n47718 ;
  assign y13231 = n47720 ;
  assign y13232 = ~n47723 ;
  assign y13233 = ~n47724 ;
  assign y13234 = ~1'b0 ;
  assign y13235 = ~n47726 ;
  assign y13236 = n47731 ;
  assign y13237 = n47732 ;
  assign y13238 = ~n47735 ;
  assign y13239 = n47736 ;
  assign y13240 = ~n47737 ;
  assign y13241 = ~n47744 ;
  assign y13242 = ~n34193 ;
  assign y13243 = ~n47748 ;
  assign y13244 = n47750 ;
  assign y13245 = ~n47752 ;
  assign y13246 = n47753 ;
  assign y13247 = n47757 ;
  assign y13248 = n47759 ;
  assign y13249 = ~n47762 ;
  assign y13250 = n47763 ;
  assign y13251 = ~n47766 ;
  assign y13252 = n47773 ;
  assign y13253 = n47776 ;
  assign y13254 = ~n47783 ;
  assign y13255 = ~n47785 ;
  assign y13256 = ~n47790 ;
  assign y13257 = n47792 ;
  assign y13258 = ~n47794 ;
  assign y13259 = ~n47798 ;
  assign y13260 = ~n47803 ;
  assign y13261 = ~n47805 ;
  assign y13262 = n47808 ;
  assign y13263 = n47809 ;
  assign y13264 = n47810 ;
  assign y13265 = ~n47812 ;
  assign y13266 = ~n47815 ;
  assign y13267 = ~n47816 ;
  assign y13268 = ~n47817 ;
  assign y13269 = ~n47818 ;
  assign y13270 = ~n47821 ;
  assign y13271 = ~n47823 ;
  assign y13272 = ~n47825 ;
  assign y13273 = n47828 ;
  assign y13274 = ~n47831 ;
  assign y13275 = n47832 ;
  assign y13276 = ~n47834 ;
  assign y13277 = n47835 ;
  assign y13278 = ~n47836 ;
  assign y13279 = ~n47838 ;
  assign y13280 = n47841 ;
  assign y13281 = ~n47845 ;
  assign y13282 = n47847 ;
  assign y13283 = n47849 ;
  assign y13284 = ~n47853 ;
  assign y13285 = ~n47855 ;
  assign y13286 = ~n47857 ;
  assign y13287 = n47860 ;
  assign y13288 = n47866 ;
  assign y13289 = ~1'b0 ;
  assign y13290 = ~n47871 ;
  assign y13291 = n47873 ;
  assign y13292 = n47875 ;
  assign y13293 = ~n47876 ;
  assign y13294 = n47878 ;
  assign y13295 = ~n47883 ;
  assign y13296 = ~n47884 ;
  assign y13297 = ~n47886 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~1'b0 ;
  assign y13300 = ~n47890 ;
  assign y13301 = n47894 ;
  assign y13302 = ~n47895 ;
  assign y13303 = n47898 ;
  assign y13304 = ~n47899 ;
  assign y13305 = ~n47901 ;
  assign y13306 = ~n47906 ;
  assign y13307 = ~1'b0 ;
  assign y13308 = ~n47907 ;
  assign y13309 = n47909 ;
  assign y13310 = n47910 ;
  assign y13311 = n47912 ;
  assign y13312 = n47914 ;
  assign y13313 = ~n47917 ;
  assign y13314 = ~n47918 ;
  assign y13315 = ~1'b0 ;
  assign y13316 = ~n47919 ;
  assign y13317 = n47920 ;
  assign y13318 = ~n47924 ;
  assign y13319 = ~n47927 ;
  assign y13320 = n47929 ;
  assign y13321 = ~n47932 ;
  assign y13322 = n47933 ;
  assign y13323 = n47934 ;
  assign y13324 = ~n47938 ;
  assign y13325 = n47940 ;
  assign y13326 = n47941 ;
  assign y13327 = ~n47942 ;
  assign y13328 = n47943 ;
  assign y13329 = ~1'b0 ;
  assign y13330 = n47945 ;
  assign y13331 = ~n47947 ;
  assign y13332 = ~n47950 ;
  assign y13333 = ~n47951 ;
  assign y13334 = ~n47954 ;
  assign y13335 = ~n47955 ;
  assign y13336 = ~n47956 ;
  assign y13337 = ~1'b0 ;
  assign y13338 = n47958 ;
  assign y13339 = ~n47963 ;
  assign y13340 = ~n47965 ;
  assign y13341 = ~n47966 ;
  assign y13342 = n47969 ;
  assign y13343 = n47971 ;
  assign y13344 = ~n47972 ;
  assign y13345 = ~n47975 ;
  assign y13346 = ~1'b0 ;
  assign y13347 = ~n47982 ;
  assign y13348 = ~n47984 ;
  assign y13349 = n47986 ;
  assign y13350 = n47987 ;
  assign y13351 = ~n47990 ;
  assign y13352 = ~n47993 ;
  assign y13353 = ~n47994 ;
  assign y13354 = ~n47995 ;
  assign y13355 = ~n47998 ;
  assign y13356 = n48002 ;
  assign y13357 = n48003 ;
  assign y13358 = ~n48006 ;
  assign y13359 = n48007 ;
  assign y13360 = ~n48009 ;
  assign y13361 = ~n48012 ;
  assign y13362 = ~n48013 ;
  assign y13363 = ~n48016 ;
  assign y13364 = ~1'b0 ;
  assign y13365 = ~n48018 ;
  assign y13366 = n48021 ;
  assign y13367 = n48022 ;
  assign y13368 = ~n48023 ;
  assign y13369 = ~n48027 ;
  assign y13370 = ~n48031 ;
  assign y13371 = ~n48035 ;
  assign y13372 = n48036 ;
  assign y13373 = n48039 ;
  assign y13374 = ~1'b0 ;
  assign y13375 = ~n48042 ;
  assign y13376 = n48044 ;
  assign y13377 = n48045 ;
  assign y13378 = n48046 ;
  assign y13379 = n48047 ;
  assign y13380 = ~n48049 ;
  assign y13381 = ~n48051 ;
  assign y13382 = ~n48057 ;
  assign y13383 = n48058 ;
  assign y13384 = ~n48061 ;
  assign y13385 = ~n48063 ;
  assign y13386 = 1'b0 ;
  assign y13387 = ~n48069 ;
  assign y13388 = ~n48071 ;
  assign y13389 = n48074 ;
  assign y13390 = ~n48077 ;
  assign y13391 = n48080 ;
  assign y13392 = ~n48081 ;
  assign y13393 = ~n48082 ;
  assign y13394 = ~n48085 ;
  assign y13395 = n48088 ;
  assign y13396 = ~n48090 ;
  assign y13397 = ~n48094 ;
  assign y13398 = n48095 ;
  assign y13399 = ~n48103 ;
  assign y13400 = ~n48104 ;
  assign y13401 = n48105 ;
  assign y13402 = n48108 ;
  assign y13403 = ~n48110 ;
  assign y13404 = n48111 ;
  assign y13405 = n48112 ;
  assign y13406 = ~1'b0 ;
  assign y13407 = ~n48115 ;
  assign y13408 = ~n48119 ;
  assign y13409 = ~n48120 ;
  assign y13410 = n48121 ;
  assign y13411 = n48126 ;
  assign y13412 = n48127 ;
  assign y13413 = n48128 ;
  assign y13414 = n48129 ;
  assign y13415 = ~n48131 ;
  assign y13416 = ~n48133 ;
  assign y13417 = ~n48139 ;
  assign y13418 = ~n48140 ;
  assign y13419 = n48141 ;
  assign y13420 = ~n48143 ;
  assign y13421 = n48145 ;
  assign y13422 = n48146 ;
  assign y13423 = ~n48148 ;
  assign y13424 = ~n48149 ;
  assign y13425 = ~n48152 ;
  assign y13426 = ~n48158 ;
  assign y13427 = ~n48160 ;
  assign y13428 = n48161 ;
  assign y13429 = ~n48162 ;
  assign y13430 = n48166 ;
  assign y13431 = n48168 ;
  assign y13432 = ~n48172 ;
  assign y13433 = n48177 ;
  assign y13434 = n48183 ;
  assign y13435 = ~n48185 ;
  assign y13436 = ~n48187 ;
  assign y13437 = ~n48188 ;
  assign y13438 = n48195 ;
  assign y13439 = n48197 ;
  assign y13440 = ~n48198 ;
  assign y13441 = ~n48201 ;
  assign y13442 = ~1'b0 ;
  assign y13443 = n48203 ;
  assign y13444 = ~n48204 ;
  assign y13445 = ~n48206 ;
  assign y13446 = n48208 ;
  assign y13447 = n822 ;
  assign y13448 = ~n48209 ;
  assign y13449 = ~n48214 ;
  assign y13450 = ~1'b0 ;
  assign y13451 = n48216 ;
  assign y13452 = n48219 ;
  assign y13453 = n48221 ;
  assign y13454 = ~n48223 ;
  assign y13455 = n48225 ;
  assign y13456 = ~n48226 ;
  assign y13457 = n48227 ;
  assign y13458 = ~n48228 ;
  assign y13459 = ~n48229 ;
  assign y13460 = ~1'b0 ;
  assign y13461 = n48231 ;
  assign y13462 = n48232 ;
  assign y13463 = ~n48241 ;
  assign y13464 = ~n48243 ;
  assign y13465 = ~n48248 ;
  assign y13466 = ~n48252 ;
  assign y13467 = n48253 ;
  assign y13468 = n48254 ;
  assign y13469 = n48257 ;
  assign y13470 = n48263 ;
  assign y13471 = ~1'b0 ;
  assign y13472 = ~1'b0 ;
  assign y13473 = n48265 ;
  assign y13474 = n48269 ;
  assign y13475 = n48270 ;
  assign y13476 = ~n48271 ;
  assign y13477 = ~n48273 ;
  assign y13478 = ~n48274 ;
  assign y13479 = ~n48275 ;
  assign y13480 = ~n48280 ;
  assign y13481 = n48284 ;
  assign y13482 = ~n48286 ;
  assign y13483 = n48292 ;
  assign y13484 = n48294 ;
  assign y13485 = n48295 ;
  assign y13486 = ~n48297 ;
  assign y13487 = n48298 ;
  assign y13488 = ~n48303 ;
  assign y13489 = ~n48305 ;
  assign y13490 = ~n48306 ;
  assign y13491 = ~n48308 ;
  assign y13492 = n48311 ;
  assign y13493 = ~n48313 ;
  assign y13494 = n46600 ;
  assign y13495 = n48315 ;
  assign y13496 = n48316 ;
  assign y13497 = n48318 ;
  assign y13498 = n48320 ;
  assign y13499 = ~n48323 ;
  assign y13500 = ~n48329 ;
  assign y13501 = ~n48332 ;
  assign y13502 = ~n48337 ;
  assign y13503 = n48340 ;
  assign y13504 = ~n48345 ;
  assign y13505 = ~n48348 ;
  assign y13506 = ~n48351 ;
  assign y13507 = ~n48354 ;
  assign y13508 = ~1'b0 ;
  assign y13509 = ~n48355 ;
  assign y13510 = n48365 ;
  assign y13511 = n48369 ;
  assign y13512 = ~n48375 ;
  assign y13513 = ~n48377 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = n48378 ;
  assign y13516 = ~n48379 ;
  assign y13517 = n48383 ;
  assign y13518 = ~n48386 ;
  assign y13519 = ~n48389 ;
  assign y13520 = ~n48390 ;
  assign y13521 = n48392 ;
  assign y13522 = n48393 ;
  assign y13523 = ~n48396 ;
  assign y13524 = n48398 ;
  assign y13525 = n48403 ;
  assign y13526 = n48406 ;
  assign y13527 = n48409 ;
  assign y13528 = ~n48410 ;
  assign y13529 = n48411 ;
  assign y13530 = n48412 ;
  assign y13531 = ~n48413 ;
  assign y13532 = ~n48415 ;
  assign y13533 = n48417 ;
  assign y13534 = n48420 ;
  assign y13535 = n48421 ;
  assign y13536 = ~n48422 ;
  assign y13537 = n48427 ;
  assign y13538 = ~n48428 ;
  assign y13539 = ~n48429 ;
  assign y13540 = ~n48436 ;
  assign y13541 = n48440 ;
  assign y13542 = n48446 ;
  assign y13543 = ~1'b0 ;
  assign y13544 = n48450 ;
  assign y13545 = n48454 ;
  assign y13546 = n48455 ;
  assign y13547 = ~n6258 ;
  assign y13548 = ~n48456 ;
  assign y13549 = ~n48460 ;
  assign y13550 = ~1'b0 ;
  assign y13551 = ~n48462 ;
  assign y13552 = n48463 ;
  assign y13553 = ~n48465 ;
  assign y13554 = ~n48467 ;
  assign y13555 = ~1'b0 ;
  assign y13556 = n48468 ;
  assign y13557 = ~n48472 ;
  assign y13558 = n48474 ;
  assign y13559 = ~n48476 ;
  assign y13560 = n48478 ;
  assign y13561 = ~n48479 ;
  assign y13562 = n48481 ;
  assign y13563 = ~n48482 ;
  assign y13564 = n48484 ;
  assign y13565 = n48487 ;
  assign y13566 = n48489 ;
  assign y13567 = n48491 ;
  assign y13568 = ~n48493 ;
  assign y13569 = ~n48494 ;
  assign y13570 = ~n48495 ;
  assign y13571 = n48496 ;
  assign y13572 = ~n48500 ;
  assign y13573 = ~n48501 ;
  assign y13574 = n48503 ;
  assign y13575 = n48504 ;
  assign y13576 = ~n48505 ;
  assign y13577 = ~n48509 ;
  assign y13578 = n48510 ;
  assign y13579 = ~n48511 ;
  assign y13580 = ~n48513 ;
  assign y13581 = n48519 ;
  assign y13582 = ~n48525 ;
  assign y13583 = ~n48526 ;
  assign y13584 = ~1'b0 ;
  assign y13585 = n48527 ;
  assign y13586 = ~n48528 ;
  assign y13587 = n48530 ;
  assign y13588 = ~n48533 ;
  assign y13589 = ~n48534 ;
  assign y13590 = ~n48540 ;
  assign y13591 = n48542 ;
  assign y13592 = n48543 ;
  assign y13593 = n48553 ;
  assign y13594 = ~n48555 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = n48558 ;
  assign y13597 = ~n48562 ;
  assign y13598 = ~n48564 ;
  assign y13599 = ~n48567 ;
  assign y13600 = n48568 ;
  assign y13601 = n48574 ;
  assign y13602 = n48577 ;
  assign y13603 = ~n48579 ;
  assign y13604 = ~n48581 ;
  assign y13605 = n48583 ;
  assign y13606 = ~n48584 ;
  assign y13607 = ~n48585 ;
  assign y13608 = n48588 ;
  assign y13609 = n48589 ;
  assign y13610 = n48594 ;
  assign y13611 = ~n48595 ;
  assign y13612 = n48598 ;
  assign y13613 = ~n48606 ;
  assign y13614 = ~n48608 ;
  assign y13615 = ~n48615 ;
  assign y13616 = n48616 ;
  assign y13617 = ~n48618 ;
  assign y13618 = ~n48620 ;
  assign y13619 = n48625 ;
  assign y13620 = n48627 ;
  assign y13621 = ~n48630 ;
  assign y13622 = ~n48633 ;
  assign y13623 = ~n48634 ;
  assign y13624 = ~n48636 ;
  assign y13625 = n48637 ;
  assign y13626 = ~n48640 ;
  assign y13627 = n48644 ;
  assign y13628 = ~1'b0 ;
  assign y13629 = ~n48646 ;
  assign y13630 = ~1'b0 ;
  assign y13631 = ~n48648 ;
  assign y13632 = ~n48650 ;
  assign y13633 = ~n48651 ;
  assign y13634 = ~n48652 ;
  assign y13635 = ~n48654 ;
  assign y13636 = n48656 ;
  assign y13637 = ~1'b0 ;
  assign y13638 = ~n48659 ;
  assign y13639 = n48661 ;
  assign y13640 = ~n48662 ;
  assign y13641 = ~n48664 ;
  assign y13642 = n48665 ;
  assign y13643 = ~n48669 ;
  assign y13644 = n48671 ;
  assign y13645 = n48672 ;
  assign y13646 = ~n48676 ;
  assign y13647 = n48680 ;
  assign y13648 = ~1'b0 ;
  assign y13649 = n48684 ;
  assign y13650 = ~n48685 ;
  assign y13651 = n48686 ;
  assign y13652 = n48687 ;
  assign y13653 = n48689 ;
  assign y13654 = n48696 ;
  assign y13655 = ~n48700 ;
  assign y13656 = ~n48703 ;
  assign y13657 = ~n48705 ;
  assign y13658 = n48707 ;
  assign y13659 = ~n48711 ;
  assign y13660 = ~n48712 ;
  assign y13661 = n48713 ;
  assign y13662 = n48714 ;
  assign y13663 = n48716 ;
  assign y13664 = n48719 ;
  assign y13665 = n48720 ;
  assign y13666 = n48721 ;
  assign y13667 = ~n48724 ;
  assign y13668 = ~n48725 ;
  assign y13669 = n48727 ;
  assign y13670 = n48730 ;
  assign y13671 = ~n48733 ;
  assign y13672 = ~1'b0 ;
  assign y13673 = n48734 ;
  assign y13674 = n48735 ;
  assign y13675 = ~n48736 ;
  assign y13676 = ~n48738 ;
  assign y13677 = n48741 ;
  assign y13678 = n48744 ;
  assign y13679 = ~n48746 ;
  assign y13680 = ~n48749 ;
  assign y13681 = ~n48750 ;
  assign y13682 = ~1'b0 ;
  assign y13683 = n48755 ;
  assign y13684 = ~n48759 ;
  assign y13685 = ~n48761 ;
  assign y13686 = n48762 ;
  assign y13687 = ~n48768 ;
  assign y13688 = ~n48769 ;
  assign y13689 = ~1'b0 ;
  assign y13690 = ~n48771 ;
  assign y13691 = ~n48773 ;
  assign y13692 = n48776 ;
  assign y13693 = ~n48781 ;
  assign y13694 = n48782 ;
  assign y13695 = n48783 ;
  assign y13696 = n48784 ;
  assign y13697 = ~n48786 ;
  assign y13698 = ~n48788 ;
  assign y13699 = ~1'b0 ;
  assign y13700 = n48790 ;
  assign y13701 = ~n48793 ;
  assign y13702 = ~n48794 ;
  assign y13703 = n48795 ;
  assign y13704 = n48799 ;
  assign y13705 = n48805 ;
  assign y13706 = n48808 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = n48810 ;
  assign y13709 = ~n48815 ;
  assign y13710 = ~n48817 ;
  assign y13711 = n48818 ;
  assign y13712 = ~n48820 ;
  assign y13713 = ~n48823 ;
  assign y13714 = ~n48824 ;
  assign y13715 = ~n48826 ;
  assign y13716 = ~n48828 ;
  assign y13717 = ~1'b0 ;
  assign y13718 = n48829 ;
  assign y13719 = ~n48832 ;
  assign y13720 = n48836 ;
  assign y13721 = ~n48837 ;
  assign y13722 = ~n48838 ;
  assign y13723 = ~n48839 ;
  assign y13724 = ~n48841 ;
  assign y13725 = ~n48843 ;
  assign y13726 = ~1'b0 ;
  assign y13727 = ~n48844 ;
  assign y13728 = n48847 ;
  assign y13729 = n48848 ;
  assign y13730 = n48853 ;
  assign y13731 = n48856 ;
  assign y13732 = n48857 ;
  assign y13733 = ~n48860 ;
  assign y13734 = ~n48862 ;
  assign y13735 = ~1'b0 ;
  assign y13736 = ~1'b0 ;
  assign y13737 = n48863 ;
  assign y13738 = n48864 ;
  assign y13739 = ~n48870 ;
  assign y13740 = ~n48874 ;
  assign y13741 = ~n48875 ;
  assign y13742 = n48876 ;
  assign y13743 = n48877 ;
  assign y13744 = n48882 ;
  assign y13745 = ~1'b0 ;
  assign y13746 = ~n48885 ;
  assign y13747 = n48889 ;
  assign y13748 = ~n48893 ;
  assign y13749 = ~n48894 ;
  assign y13750 = ~n48896 ;
  assign y13751 = ~n48898 ;
  assign y13752 = ~n48899 ;
  assign y13753 = n48904 ;
  assign y13754 = ~n48905 ;
  assign y13755 = n48908 ;
  assign y13756 = n48913 ;
  assign y13757 = n48915 ;
  assign y13758 = ~n48917 ;
  assign y13759 = n48918 ;
  assign y13760 = ~n48919 ;
  assign y13761 = n48923 ;
  assign y13762 = n48926 ;
  assign y13763 = n48929 ;
  assign y13764 = ~n48933 ;
  assign y13765 = n48935 ;
  assign y13766 = ~n48937 ;
  assign y13767 = ~n48939 ;
  assign y13768 = ~n48941 ;
  assign y13769 = ~n48942 ;
  assign y13770 = ~n48946 ;
  assign y13771 = ~n48947 ;
  assign y13772 = ~n48948 ;
  assign y13773 = n48952 ;
  assign y13774 = n48954 ;
  assign y13775 = n48958 ;
  assign y13776 = ~n48962 ;
  assign y13777 = ~n48963 ;
  assign y13778 = n48964 ;
  assign y13779 = ~n48965 ;
  assign y13780 = n48969 ;
  assign y13781 = n48974 ;
  assign y13782 = ~n48979 ;
  assign y13783 = ~n48984 ;
  assign y13784 = ~n48986 ;
  assign y13785 = n48987 ;
  assign y13786 = ~n48992 ;
  assign y13787 = ~n48996 ;
  assign y13788 = n48997 ;
  assign y13789 = n49005 ;
  assign y13790 = n49006 ;
  assign y13791 = ~n49008 ;
  assign y13792 = n49011 ;
  assign y13793 = ~1'b0 ;
  assign y13794 = n49013 ;
  assign y13795 = n49016 ;
  assign y13796 = n49017 ;
  assign y13797 = n49019 ;
  assign y13798 = n49027 ;
  assign y13799 = n49029 ;
  assign y13800 = ~n49031 ;
  assign y13801 = ~n49033 ;
  assign y13802 = ~n49035 ;
  assign y13803 = ~n49041 ;
  assign y13804 = n49042 ;
  assign y13805 = ~n49055 ;
  assign y13806 = n49056 ;
  assign y13807 = ~n49058 ;
  assign y13808 = ~n49059 ;
  assign y13809 = ~n49064 ;
  assign y13810 = n49066 ;
  assign y13811 = ~n49067 ;
  assign y13812 = ~n49071 ;
  assign y13813 = ~n49074 ;
  assign y13814 = ~n49076 ;
  assign y13815 = n49077 ;
  assign y13816 = ~n49078 ;
  assign y13817 = n49081 ;
  assign y13818 = n49084 ;
  assign y13819 = ~n49085 ;
  assign y13820 = ~n49087 ;
  assign y13821 = ~1'b0 ;
  assign y13822 = ~n49088 ;
  assign y13823 = ~n49092 ;
  assign y13824 = n49093 ;
  assign y13825 = ~n49096 ;
  assign y13826 = n49097 ;
  assign y13827 = ~n49103 ;
  assign y13828 = n49109 ;
  assign y13829 = ~n49111 ;
  assign y13830 = n49113 ;
  assign y13831 = n49114 ;
  assign y13832 = n49115 ;
  assign y13833 = ~n49119 ;
  assign y13834 = ~n49121 ;
  assign y13835 = n49126 ;
  assign y13836 = n49128 ;
  assign y13837 = n49133 ;
  assign y13838 = n49135 ;
  assign y13839 = ~1'b0 ;
  assign y13840 = ~n49139 ;
  assign y13841 = n49142 ;
  assign y13842 = n49143 ;
  assign y13843 = n49145 ;
  assign y13844 = n49146 ;
  assign y13845 = ~n49148 ;
  assign y13846 = ~n49150 ;
  assign y13847 = n49153 ;
  assign y13848 = ~n49156 ;
  assign y13849 = ~n49157 ;
  assign y13850 = n49159 ;
  assign y13851 = n49163 ;
  assign y13852 = n49164 ;
  assign y13853 = ~n49169 ;
  assign y13854 = ~n49175 ;
  assign y13855 = n49178 ;
  assign y13856 = ~n49179 ;
  assign y13857 = n49180 ;
  assign y13858 = n49184 ;
  assign y13859 = ~1'b0 ;
  assign y13860 = ~n49186 ;
  assign y13861 = n49190 ;
  assign y13862 = n49193 ;
  assign y13863 = ~n49198 ;
  assign y13864 = ~n49200 ;
  assign y13865 = n49202 ;
  assign y13866 = n49203 ;
  assign y13867 = ~1'b0 ;
  assign y13868 = n49204 ;
  assign y13869 = n49211 ;
  assign y13870 = n49214 ;
  assign y13871 = n49220 ;
  assign y13872 = ~n49226 ;
  assign y13873 = ~n49227 ;
  assign y13874 = ~n49228 ;
  assign y13875 = n49232 ;
  assign y13876 = n49234 ;
  assign y13877 = ~1'b0 ;
  assign y13878 = ~n49235 ;
  assign y13879 = n49236 ;
  assign y13880 = n49237 ;
  assign y13881 = n49240 ;
  assign y13882 = n49244 ;
  assign y13883 = n49246 ;
  assign y13884 = n49247 ;
  assign y13885 = ~n49249 ;
  assign y13886 = ~n49251 ;
  assign y13887 = ~n49256 ;
  assign y13888 = ~n49257 ;
  assign y13889 = n49258 ;
  assign y13890 = n49260 ;
  assign y13891 = ~n49269 ;
  assign y13892 = ~n49274 ;
  assign y13893 = ~n49275 ;
  assign y13894 = ~n49279 ;
  assign y13895 = n49286 ;
  assign y13896 = ~1'b0 ;
  assign y13897 = ~n34597 ;
  assign y13898 = ~n49289 ;
  assign y13899 = n49295 ;
  assign y13900 = ~n49296 ;
  assign y13901 = n49300 ;
  assign y13902 = ~n49306 ;
  assign y13903 = n49312 ;
  assign y13904 = ~n49318 ;
  assign y13905 = n49321 ;
  assign y13906 = n49324 ;
  assign y13907 = ~n49328 ;
  assign y13908 = n49331 ;
  assign y13909 = ~n49332 ;
  assign y13910 = n49336 ;
  assign y13911 = ~n49338 ;
  assign y13912 = ~n49340 ;
  assign y13913 = n49343 ;
  assign y13914 = n49344 ;
  assign y13915 = ~1'b0 ;
  assign y13916 = ~n49346 ;
  assign y13917 = ~n49349 ;
  assign y13918 = n49353 ;
  assign y13919 = ~n49354 ;
  assign y13920 = n49358 ;
  assign y13921 = ~n49361 ;
  assign y13922 = n49363 ;
  assign y13923 = n49364 ;
  assign y13924 = ~n49365 ;
  assign y13925 = n49366 ;
  assign y13926 = ~n49367 ;
  assign y13927 = n49372 ;
  assign y13928 = n49373 ;
  assign y13929 = n49378 ;
  assign y13930 = n49380 ;
  assign y13931 = n49382 ;
  assign y13932 = n49383 ;
  assign y13933 = ~1'b0 ;
  assign y13934 = n49385 ;
  assign y13935 = ~n49386 ;
  assign y13936 = ~n49387 ;
  assign y13937 = ~n49388 ;
  assign y13938 = ~n49390 ;
  assign y13939 = n49391 ;
  assign y13940 = ~n49392 ;
  assign y13941 = n49396 ;
  assign y13942 = ~1'b0 ;
  assign y13943 = n49398 ;
  assign y13944 = ~n49401 ;
  assign y13945 = ~n49403 ;
  assign y13946 = ~n49406 ;
  assign y13947 = n49408 ;
  assign y13948 = n49417 ;
  assign y13949 = ~n49419 ;
  assign y13950 = ~n49424 ;
  assign y13951 = ~1'b0 ;
  assign y13952 = ~1'b0 ;
  assign y13953 = n49425 ;
  assign y13954 = ~n49429 ;
  assign y13955 = ~n49430 ;
  assign y13956 = ~n49431 ;
  assign y13957 = ~n49433 ;
  assign y13958 = ~n49434 ;
  assign y13959 = ~n49438 ;
  assign y13960 = ~n49441 ;
  assign y13961 = ~n49447 ;
  assign y13962 = ~n49449 ;
  assign y13963 = n49451 ;
  assign y13964 = n49452 ;
  assign y13965 = ~n49459 ;
  assign y13966 = ~n49462 ;
  assign y13967 = n49463 ;
  assign y13968 = ~n49464 ;
  assign y13969 = ~1'b0 ;
  assign y13970 = ~n49465 ;
  assign y13971 = n49467 ;
  assign y13972 = n49469 ;
  assign y13973 = n49470 ;
  assign y13974 = ~n33921 ;
  assign y13975 = n49471 ;
  assign y13976 = ~n49473 ;
  assign y13977 = ~n49477 ;
  assign y13978 = ~n49479 ;
  assign y13979 = ~n49481 ;
  assign y13980 = n49484 ;
  assign y13981 = n49485 ;
  assign y13982 = n49488 ;
  assign y13983 = ~n49489 ;
  assign y13984 = ~n49490 ;
  assign y13985 = n49491 ;
  assign y13986 = n49494 ;
  assign y13987 = n49497 ;
  assign y13988 = n18243 ;
  assign y13989 = n49501 ;
  assign y13990 = n49504 ;
  assign y13991 = ~n49506 ;
  assign y13992 = n49509 ;
  assign y13993 = n49510 ;
  assign y13994 = ~n49512 ;
  assign y13995 = n49513 ;
  assign y13996 = n49515 ;
  assign y13997 = ~n49516 ;
  assign y13998 = ~n49519 ;
  assign y13999 = n49521 ;
  assign y14000 = ~n49523 ;
  assign y14001 = n49525 ;
  assign y14002 = ~n49526 ;
  assign y14003 = n49527 ;
  assign y14004 = n49529 ;
  assign y14005 = ~1'b0 ;
  assign y14006 = ~1'b0 ;
  assign y14007 = ~1'b0 ;
  assign y14008 = n49531 ;
  assign y14009 = ~n49535 ;
  assign y14010 = ~n49536 ;
  assign y14011 = ~n49538 ;
  assign y14012 = ~n49539 ;
  assign y14013 = ~n49540 ;
  assign y14014 = ~n49541 ;
  assign y14015 = ~n49546 ;
  assign y14016 = ~1'b0 ;
  assign y14017 = n49549 ;
  assign y14018 = n49552 ;
  assign y14019 = ~n49553 ;
  assign y14020 = ~n49557 ;
  assign y14021 = ~n49559 ;
  assign y14022 = n49563 ;
  assign y14023 = n49566 ;
  assign y14024 = ~n49567 ;
  assign y14025 = n49568 ;
  assign y14026 = n49569 ;
  assign y14027 = n49573 ;
  assign y14028 = n49574 ;
  assign y14029 = n49575 ;
  assign y14030 = ~n49576 ;
  assign y14031 = ~n49577 ;
  assign y14032 = n49579 ;
  assign y14033 = n49581 ;
  assign y14034 = ~1'b0 ;
  assign y14035 = n49583 ;
  assign y14036 = n49584 ;
  assign y14037 = ~n49587 ;
  assign y14038 = ~n49591 ;
  assign y14039 = ~n49592 ;
  assign y14040 = n49594 ;
  assign y14041 = ~n49597 ;
  assign y14042 = n49598 ;
  assign y14043 = n49599 ;
  assign y14044 = n49603 ;
  assign y14045 = n49608 ;
  assign y14046 = n49611 ;
  assign y14047 = ~n49614 ;
  assign y14048 = n49615 ;
  assign y14049 = n49619 ;
  assign y14050 = n49626 ;
  assign y14051 = ~n49628 ;
  assign y14052 = ~1'b0 ;
  assign y14053 = ~n49631 ;
  assign y14054 = n49632 ;
  assign y14055 = ~n49633 ;
  assign y14056 = n49635 ;
  assign y14057 = ~n49637 ;
  assign y14058 = n49638 ;
  assign y14059 = ~n49642 ;
  assign y14060 = n49645 ;
  assign y14061 = ~1'b0 ;
  assign y14062 = ~1'b0 ;
  assign y14063 = ~1'b0 ;
  assign y14064 = ~n49648 ;
  assign y14065 = ~n49650 ;
  assign y14066 = n49654 ;
  assign y14067 = n49655 ;
  assign y14068 = n49658 ;
  assign y14069 = n49659 ;
  assign y14070 = ~n49661 ;
  assign y14071 = n49666 ;
  assign y14072 = ~n49668 ;
  assign y14073 = ~n49673 ;
  assign y14074 = ~n49677 ;
  assign y14075 = ~n49685 ;
  assign y14076 = n49686 ;
  assign y14077 = n49690 ;
  assign y14078 = n49692 ;
  assign y14079 = n49693 ;
  assign y14080 = ~n49701 ;
  assign y14081 = ~n49703 ;
  assign y14082 = ~n49706 ;
  assign y14083 = n49710 ;
  assign y14084 = ~n49713 ;
  assign y14085 = ~n49716 ;
  assign y14086 = ~n49718 ;
  assign y14087 = ~n49719 ;
  assign y14088 = ~n49720 ;
  assign y14089 = ~n49722 ;
  assign y14090 = n49724 ;
  assign y14091 = ~1'b0 ;
  assign y14092 = n49726 ;
  assign y14093 = ~n49728 ;
  assign y14094 = ~n49729 ;
  assign y14095 = n49731 ;
  assign y14096 = n49732 ;
  assign y14097 = ~n49737 ;
  assign y14098 = n49740 ;
  assign y14099 = ~n49741 ;
  assign y14100 = ~1'b0 ;
  assign y14101 = ~n49743 ;
  assign y14102 = ~1'b0 ;
  assign y14103 = ~n49744 ;
  assign y14104 = n49745 ;
  assign y14105 = ~n49747 ;
  assign y14106 = ~n49751 ;
  assign y14107 = ~n49753 ;
  assign y14108 = ~n49755 ;
  assign y14109 = ~n49759 ;
  assign y14110 = ~1'b0 ;
  assign y14111 = ~n49761 ;
  assign y14112 = ~n49762 ;
  assign y14113 = n49763 ;
  assign y14114 = ~n49766 ;
  assign y14115 = ~n49770 ;
  assign y14116 = n49773 ;
  assign y14117 = n49774 ;
  assign y14118 = n49776 ;
  assign y14119 = n49777 ;
  assign y14120 = ~1'b0 ;
  assign y14121 = ~n49778 ;
  assign y14122 = n49779 ;
  assign y14123 = ~n49780 ;
  assign y14124 = n49782 ;
  assign y14125 = n49784 ;
  assign y14126 = ~n49786 ;
  assign y14127 = ~n49790 ;
  assign y14128 = n49792 ;
  assign y14129 = n49805 ;
  assign y14130 = n49806 ;
  assign y14131 = ~n49808 ;
  assign y14132 = n49811 ;
  assign y14133 = n49812 ;
  assign y14134 = n49813 ;
  assign y14135 = n49816 ;
  assign y14136 = ~n49819 ;
  assign y14137 = ~n49820 ;
  assign y14138 = ~1'b0 ;
  assign y14139 = ~n49821 ;
  assign y14140 = ~n49823 ;
  assign y14141 = n49824 ;
  assign y14142 = n49825 ;
  assign y14143 = n49828 ;
  assign y14144 = ~n49830 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = ~1'b0 ;
  assign y14147 = ~1'b0 ;
  assign y14148 = n49837 ;
  assign y14149 = n49838 ;
  assign y14150 = n49839 ;
  assign y14151 = n49840 ;
  assign y14152 = ~n49846 ;
  assign y14153 = n49849 ;
  assign y14154 = ~n49852 ;
  assign y14155 = ~n49854 ;
  assign y14156 = ~1'b0 ;
  assign y14157 = ~n49856 ;
  assign y14158 = ~n49857 ;
  assign y14159 = n49859 ;
  assign y14160 = ~n49861 ;
  assign y14161 = ~n27912 ;
  assign y14162 = n49863 ;
  assign y14163 = ~n49864 ;
  assign y14164 = ~n49867 ;
  assign y14165 = ~1'b0 ;
  assign y14166 = ~1'b0 ;
  assign y14167 = n49868 ;
  assign y14168 = ~n49869 ;
  assign y14169 = ~n49870 ;
  assign y14170 = n49871 ;
  assign y14171 = n49874 ;
  assign y14172 = n49876 ;
  assign y14173 = n49877 ;
  assign y14174 = n49879 ;
  assign y14175 = 1'b0 ;
  assign y14176 = n49880 ;
  assign y14177 = n49882 ;
  assign y14178 = n49883 ;
  assign y14179 = n49887 ;
  assign y14180 = n49890 ;
  assign y14181 = n49894 ;
  assign y14182 = n49895 ;
  assign y14183 = n49897 ;
  assign y14184 = n49898 ;
  assign y14185 = ~n49903 ;
  assign y14186 = ~n49906 ;
  assign y14187 = ~n44583 ;
  assign y14188 = ~n49910 ;
  assign y14189 = ~n49913 ;
  assign y14190 = ~n49914 ;
  assign y14191 = ~n49916 ;
  assign y14192 = ~n49917 ;
  assign y14193 = n49921 ;
  assign y14194 = ~1'b0 ;
  assign y14195 = n49923 ;
  assign y14196 = ~n49927 ;
  assign y14197 = ~n49931 ;
  assign y14198 = ~n49933 ;
  assign y14199 = n49934 ;
  assign y14200 = ~n49935 ;
  assign y14201 = n49942 ;
  assign y14202 = n49943 ;
  assign y14203 = ~n49945 ;
  assign y14204 = ~1'b0 ;
  assign y14205 = ~1'b0 ;
  assign y14206 = n49946 ;
  assign y14207 = n49947 ;
  assign y14208 = ~n49951 ;
  assign y14209 = n49954 ;
  assign y14210 = ~n49958 ;
  assign y14211 = n49961 ;
  assign y14212 = ~n49966 ;
  assign y14213 = n49967 ;
  assign y14214 = n49969 ;
  assign y14215 = n49970 ;
  assign y14216 = n49972 ;
  assign y14217 = ~n49973 ;
  assign y14218 = n49975 ;
  assign y14219 = ~n49980 ;
  assign y14220 = n49981 ;
  assign y14221 = n49983 ;
  assign y14222 = n49986 ;
  assign y14223 = n49987 ;
  assign y14224 = ~n49989 ;
  assign y14225 = ~n49992 ;
  assign y14226 = ~n49996 ;
  assign y14227 = n49997 ;
  assign y14228 = ~n50000 ;
  assign y14229 = ~n50001 ;
  assign y14230 = n50002 ;
  assign y14231 = n50003 ;
  assign y14232 = n50004 ;
  assign y14233 = n50005 ;
  assign y14234 = ~1'b0 ;
  assign y14235 = ~n50006 ;
  assign y14236 = ~n50008 ;
  assign y14237 = n50011 ;
  assign y14238 = ~n50012 ;
  assign y14239 = n50023 ;
  assign y14240 = ~n50026 ;
  assign y14241 = n50034 ;
  assign y14242 = n50035 ;
  assign y14243 = n50041 ;
  assign y14244 = n50042 ;
  assign y14245 = n50045 ;
  assign y14246 = ~n50046 ;
  assign y14247 = ~n50051 ;
  assign y14248 = n50052 ;
  assign y14249 = ~n50053 ;
  assign y14250 = n50056 ;
  assign y14251 = n50061 ;
  assign y14252 = n50064 ;
  assign y14253 = ~n50066 ;
  assign y14254 = n50071 ;
  assign y14255 = n50073 ;
  assign y14256 = ~n50077 ;
  assign y14257 = n50079 ;
  assign y14258 = ~1'b0 ;
  assign y14259 = n50080 ;
  assign y14260 = n50082 ;
  assign y14261 = n50083 ;
  assign y14262 = n50085 ;
  assign y14263 = n50089 ;
  assign y14264 = ~n50097 ;
  assign y14265 = n50098 ;
  assign y14266 = ~n50100 ;
  assign y14267 = ~n50102 ;
  assign y14268 = n50105 ;
  assign y14269 = ~1'b0 ;
  assign y14270 = ~1'b0 ;
  assign y14271 = ~1'b0 ;
  assign y14272 = ~n50106 ;
  assign y14273 = ~n50110 ;
  assign y14274 = n50111 ;
  assign y14275 = ~n50112 ;
  assign y14276 = ~n50113 ;
  assign y14277 = ~n50117 ;
  assign y14278 = ~n50118 ;
  assign y14279 = ~n50121 ;
  assign y14280 = ~n50126 ;
  assign y14281 = ~1'b0 ;
  assign y14282 = ~n50128 ;
  assign y14283 = n50136 ;
  assign y14284 = ~n50138 ;
  assign y14285 = n50139 ;
  assign y14286 = ~n50141 ;
  assign y14287 = n50142 ;
  assign y14288 = n50143 ;
  assign y14289 = n50144 ;
  assign y14290 = n50145 ;
  assign y14291 = n50148 ;
  assign y14292 = n50150 ;
  assign y14293 = n50155 ;
  assign y14294 = n50157 ;
  assign y14295 = n50159 ;
  assign y14296 = ~n50161 ;
  assign y14297 = ~n50165 ;
  assign y14298 = ~n50166 ;
  assign y14299 = ~n50168 ;
  assign y14300 = ~1'b0 ;
  assign y14301 = ~n50171 ;
  assign y14302 = ~n50176 ;
  assign y14303 = ~n50179 ;
  assign y14304 = ~n50180 ;
  assign y14305 = n50182 ;
  assign y14306 = n50188 ;
  assign y14307 = n50191 ;
  assign y14308 = n50192 ;
  assign y14309 = n50196 ;
  assign y14310 = n50199 ;
  assign y14311 = n50201 ;
  assign y14312 = ~n50205 ;
  assign y14313 = n50209 ;
  assign y14314 = ~n50212 ;
  assign y14315 = n50218 ;
  assign y14316 = ~n50222 ;
  assign y14317 = n50223 ;
  assign y14318 = ~n50225 ;
  assign y14319 = n50227 ;
  assign y14320 = n50229 ;
  assign y14321 = ~n50233 ;
  assign y14322 = ~n50237 ;
  assign y14323 = n50238 ;
  assign y14324 = n50239 ;
  assign y14325 = ~n16544 ;
  assign y14326 = n50242 ;
  assign y14327 = n50246 ;
  assign y14328 = ~n50248 ;
  assign y14329 = ~n50249 ;
  assign y14330 = ~n50250 ;
  assign y14331 = n50251 ;
  assign y14332 = n50258 ;
  assign y14333 = ~n50263 ;
  assign y14334 = n50267 ;
  assign y14335 = ~n50269 ;
  assign y14336 = ~n50271 ;
  assign y14337 = n50276 ;
  assign y14338 = ~1'b0 ;
  assign y14339 = ~n50278 ;
  assign y14340 = ~n50281 ;
  assign y14341 = n50282 ;
  assign y14342 = ~n50283 ;
  assign y14343 = ~n50286 ;
  assign y14344 = ~n50288 ;
  assign y14345 = ~1'b0 ;
  assign y14346 = ~n50291 ;
  assign y14347 = n50294 ;
  assign y14348 = n50297 ;
  assign y14349 = ~n50298 ;
  assign y14350 = ~n50301 ;
  assign y14351 = n50302 ;
  assign y14352 = ~n50306 ;
  assign y14353 = n50307 ;
  assign y14354 = ~n50311 ;
  assign y14355 = n50314 ;
  assign y14356 = ~n50318 ;
  assign y14357 = ~n50319 ;
  assign y14358 = ~n50320 ;
  assign y14359 = n50322 ;
  assign y14360 = ~n50325 ;
  assign y14361 = n50326 ;
  assign y14362 = ~n50329 ;
  assign y14363 = n50333 ;
  assign y14364 = n50335 ;
  assign y14365 = ~n50336 ;
  assign y14366 = ~n50340 ;
  assign y14367 = ~n50343 ;
  assign y14368 = n50348 ;
  assign y14369 = n50350 ;
  assign y14370 = ~n50351 ;
  assign y14371 = ~n38880 ;
  assign y14372 = n50356 ;
  assign y14373 = ~n50357 ;
  assign y14374 = ~n50358 ;
  assign y14375 = ~n50360 ;
  assign y14376 = ~n50364 ;
  assign y14377 = n50366 ;
  assign y14378 = n50367 ;
  assign y14379 = n50369 ;
  assign y14380 = ~n50370 ;
  assign y14381 = n50371 ;
  assign y14382 = ~n50374 ;
  assign y14383 = n50375 ;
  assign y14384 = n50376 ;
  assign y14385 = n50378 ;
  assign y14386 = ~n50380 ;
  assign y14387 = n50389 ;
  assign y14388 = n50390 ;
  assign y14389 = ~n50397 ;
  assign y14390 = ~n50399 ;
  assign y14391 = ~n50401 ;
  assign y14392 = ~n50402 ;
  assign y14393 = ~n50406 ;
  assign y14394 = ~n50409 ;
  assign y14395 = ~n50414 ;
  assign y14396 = n50417 ;
  assign y14397 = ~1'b0 ;
  assign y14398 = ~n50421 ;
  assign y14399 = ~n50422 ;
  assign y14400 = n50424 ;
  assign y14401 = ~n50430 ;
  assign y14402 = ~n50433 ;
  assign y14403 = ~n50437 ;
  assign y14404 = ~n50440 ;
  assign y14405 = ~n50443 ;
  assign y14406 = n50444 ;
  assign y14407 = n50446 ;
  assign y14408 = ~1'b0 ;
  assign y14409 = ~n50447 ;
  assign y14410 = ~n50454 ;
  assign y14411 = ~n50455 ;
  assign y14412 = n50456 ;
  assign y14413 = n50458 ;
  assign y14414 = ~n50460 ;
  assign y14415 = ~n50464 ;
  assign y14416 = ~n50467 ;
  assign y14417 = n50469 ;
  assign y14418 = ~n50470 ;
  assign y14419 = ~n50472 ;
  assign y14420 = n50474 ;
  assign y14421 = ~n50475 ;
  assign y14422 = ~n50479 ;
  assign y14423 = ~n50480 ;
  assign y14424 = n50484 ;
  assign y14425 = ~n50487 ;
  assign y14426 = ~n50489 ;
  assign y14427 = n50491 ;
  assign y14428 = ~n50493 ;
  assign y14429 = n50497 ;
  assign y14430 = ~n50502 ;
  assign y14431 = ~n50505 ;
  assign y14432 = n50512 ;
  assign y14433 = ~n50515 ;
  assign y14434 = ~n50516 ;
  assign y14435 = n50517 ;
  assign y14436 = n50521 ;
  assign y14437 = ~n50524 ;
  assign y14438 = ~1'b0 ;
  assign y14439 = ~n50526 ;
  assign y14440 = n50527 ;
  assign y14441 = ~n50534 ;
  assign y14442 = n50537 ;
  assign y14443 = ~n50540 ;
  assign y14444 = n50544 ;
  assign y14445 = ~n50546 ;
  assign y14446 = n50551 ;
  assign y14447 = n50553 ;
  assign y14448 = n50555 ;
  assign y14449 = ~1'b0 ;
  assign y14450 = ~n50559 ;
  assign y14451 = ~n50561 ;
  assign y14452 = n50563 ;
  assign y14453 = ~n50566 ;
  assign y14454 = ~n50568 ;
  assign y14455 = ~n50570 ;
  assign y14456 = ~n50573 ;
  assign y14457 = ~n50575 ;
  assign y14458 = n50576 ;
  assign y14459 = n50580 ;
  assign y14460 = ~n50582 ;
  assign y14461 = n50589 ;
  assign y14462 = ~n50591 ;
  assign y14463 = ~n50594 ;
  assign y14464 = n50597 ;
  assign y14465 = n50599 ;
  assign y14466 = n50602 ;
  assign y14467 = ~n50608 ;
  assign y14468 = ~1'b0 ;
  assign y14469 = n50610 ;
  assign y14470 = ~n50611 ;
  assign y14471 = ~n50613 ;
  assign y14472 = ~n50616 ;
  assign y14473 = n50622 ;
  assign y14474 = n50627 ;
  assign y14475 = ~n50632 ;
  assign y14476 = n50635 ;
  assign y14477 = n50638 ;
  assign y14478 = ~n50639 ;
  assign y14479 = ~n50640 ;
  assign y14480 = n50642 ;
  assign y14481 = ~n50643 ;
  assign y14482 = n50644 ;
  assign y14483 = n50645 ;
  assign y14484 = ~n50647 ;
  assign y14485 = ~n50649 ;
  assign y14486 = n50651 ;
  assign y14487 = ~1'b0 ;
  assign y14488 = ~n50652 ;
  assign y14489 = ~n50658 ;
  assign y14490 = ~n50660 ;
  assign y14491 = ~n50662 ;
  assign y14492 = n50663 ;
  assign y14493 = n50664 ;
  assign y14494 = n50665 ;
  assign y14495 = n50667 ;
  assign y14496 = ~n50669 ;
  assign y14497 = ~n50674 ;
  assign y14498 = n50676 ;
  assign y14499 = n50678 ;
  assign y14500 = ~n50681 ;
  assign y14501 = ~n50682 ;
  assign y14502 = ~n50683 ;
  assign y14503 = ~n50685 ;
  assign y14504 = ~1'b0 ;
  assign y14505 = n50688 ;
  assign y14506 = ~n50691 ;
  assign y14507 = n50693 ;
  assign y14508 = n50695 ;
  assign y14509 = n50698 ;
  assign y14510 = ~n50701 ;
  assign y14511 = n50703 ;
  assign y14512 = ~n50706 ;
  assign y14513 = ~n50708 ;
  assign y14514 = n50710 ;
  assign y14515 = ~n50711 ;
  assign y14516 = ~n50713 ;
  assign y14517 = n50714 ;
  assign y14518 = ~n50717 ;
  assign y14519 = ~n50718 ;
  assign y14520 = ~n50722 ;
  assign y14521 = ~n50728 ;
  assign y14522 = ~n50731 ;
  assign y14523 = n50734 ;
  assign y14524 = ~n50736 ;
  assign y14525 = ~n50742 ;
  assign y14526 = ~1'b0 ;
  assign y14527 = n50749 ;
  assign y14528 = ~n50753 ;
  assign y14529 = ~n50754 ;
  assign y14530 = ~n50758 ;
  assign y14531 = n50759 ;
  assign y14532 = ~n50764 ;
  assign y14533 = ~1'b0 ;
  assign y14534 = n50766 ;
  assign y14535 = n50768 ;
  assign y14536 = ~n50769 ;
  assign y14537 = ~n50772 ;
  assign y14538 = ~n50773 ;
  assign y14539 = ~n50774 ;
  assign y14540 = ~n50777 ;
  assign y14541 = n50779 ;
  assign y14542 = ~n50780 ;
  assign y14543 = ~n50786 ;
  assign y14544 = ~n50789 ;
  assign y14545 = n50793 ;
  assign y14546 = ~1'b0 ;
  assign y14547 = n50794 ;
  assign y14548 = ~n50797 ;
  assign y14549 = ~n50798 ;
  assign y14550 = ~n50801 ;
  assign y14551 = ~n50803 ;
  assign y14552 = n50804 ;
  assign y14553 = n50805 ;
  assign y14554 = ~n50814 ;
  assign y14555 = ~1'b0 ;
  assign y14556 = ~1'b0 ;
  assign y14557 = ~1'b0 ;
  assign y14558 = ~n50815 ;
  assign y14559 = ~n50817 ;
  assign y14560 = n50818 ;
  assign y14561 = ~n50819 ;
  assign y14562 = ~n50820 ;
  assign y14563 = ~n50826 ;
  assign y14564 = n50829 ;
  assign y14565 = ~1'b0 ;
  assign y14566 = ~n50830 ;
  assign y14567 = ~1'b0 ;
  assign y14568 = n50831 ;
  assign y14569 = ~n50832 ;
  assign y14570 = n50833 ;
  assign y14571 = ~n50834 ;
  assign y14572 = n50835 ;
  assign y14573 = ~n50841 ;
  assign y14574 = ~1'b0 ;
  assign y14575 = ~n50843 ;
  assign y14576 = n50849 ;
  assign y14577 = ~n50852 ;
  assign y14578 = ~n50853 ;
  assign y14579 = n50856 ;
  assign y14580 = n50857 ;
  assign y14581 = n50858 ;
  assign y14582 = ~n50860 ;
  assign y14583 = ~n50861 ;
  assign y14584 = n50863 ;
  assign y14585 = n50869 ;
  assign y14586 = ~n50871 ;
  assign y14587 = n50876 ;
  assign y14588 = ~n50882 ;
  assign y14589 = n50885 ;
  assign y14590 = n50886 ;
  assign y14591 = ~n50891 ;
  assign y14592 = ~n50898 ;
  assign y14593 = ~n50900 ;
  assign y14594 = ~n50901 ;
  assign y14595 = ~n50903 ;
  assign y14596 = ~1'b0 ;
  assign y14597 = ~n50908 ;
  assign y14598 = ~n50912 ;
  assign y14599 = ~n50915 ;
  assign y14600 = ~n50919 ;
  assign y14601 = n50920 ;
  assign y14602 = ~n50922 ;
  assign y14603 = ~n50925 ;
  assign y14604 = ~n50928 ;
  assign y14605 = ~n50929 ;
  assign y14606 = n50932 ;
  assign y14607 = ~n50936 ;
  assign y14608 = ~1'b0 ;
  assign y14609 = ~n50937 ;
  assign y14610 = ~n50940 ;
  assign y14611 = ~n50943 ;
  assign y14612 = ~n50944 ;
  assign y14613 = n50945 ;
  assign y14614 = n50947 ;
  assign y14615 = n50950 ;
  assign y14616 = ~n50951 ;
  assign y14617 = ~n50953 ;
  assign y14618 = ~n50960 ;
  assign y14619 = n50961 ;
  assign y14620 = n50962 ;
  assign y14621 = n50964 ;
  assign y14622 = ~n50965 ;
  assign y14623 = n50971 ;
  assign y14624 = ~n50972 ;
  assign y14625 = n50976 ;
  assign y14626 = ~1'b0 ;
  assign y14627 = n50978 ;
  assign y14628 = n50980 ;
  assign y14629 = ~n50981 ;
  assign y14630 = n50982 ;
  assign y14631 = ~n50983 ;
  assign y14632 = ~n50984 ;
  assign y14633 = n50987 ;
  assign y14634 = n50991 ;
  assign y14635 = n50993 ;
  assign y14636 = ~1'b0 ;
  assign y14637 = n50995 ;
  assign y14638 = ~n50996 ;
  assign y14639 = n50999 ;
  assign y14640 = n51003 ;
  assign y14641 = n51007 ;
  assign y14642 = n51008 ;
  assign y14643 = n51010 ;
  assign y14644 = n51014 ;
  assign y14645 = ~1'b0 ;
  assign y14646 = ~n51019 ;
  assign y14647 = n51021 ;
  assign y14648 = ~n51027 ;
  assign y14649 = n51029 ;
  assign y14650 = n51030 ;
  assign y14651 = ~n51031 ;
  assign y14652 = n51032 ;
  assign y14653 = n51035 ;
  assign y14654 = ~n51039 ;
  assign y14655 = n51040 ;
  assign y14656 = n51046 ;
  assign y14657 = ~n51049 ;
  assign y14658 = ~1'b0 ;
  assign y14659 = n51050 ;
  assign y14660 = ~n51051 ;
  assign y14661 = n51053 ;
  assign y14662 = ~n51054 ;
  assign y14663 = ~n51055 ;
  assign y14664 = n51056 ;
  assign y14665 = ~n51057 ;
  assign y14666 = n51059 ;
  assign y14667 = n51061 ;
  assign y14668 = ~n51063 ;
  assign y14669 = n51064 ;
  assign y14670 = n51071 ;
  assign y14671 = ~n51072 ;
  assign y14672 = n51077 ;
  assign y14673 = ~n51079 ;
  assign y14674 = n51081 ;
  assign y14675 = n51083 ;
  assign y14676 = ~1'b0 ;
  assign y14677 = ~n51084 ;
  assign y14678 = n51086 ;
  assign y14679 = ~n51087 ;
  assign y14680 = n51088 ;
  assign y14681 = ~n51092 ;
  assign y14682 = ~n51093 ;
  assign y14683 = n51095 ;
  assign y14684 = ~n51100 ;
  assign y14685 = n51102 ;
  assign y14686 = ~n51104 ;
  assign y14687 = n51107 ;
  assign y14688 = n51112 ;
  assign y14689 = n51114 ;
  assign y14690 = n51115 ;
  assign y14691 = ~n51121 ;
  assign y14692 = n32668 ;
  assign y14693 = n51123 ;
  assign y14694 = ~1'b0 ;
  assign y14695 = n51125 ;
  assign y14696 = n51131 ;
  assign y14697 = ~n51134 ;
  assign y14698 = ~n51135 ;
  assign y14699 = n51136 ;
  assign y14700 = ~n51137 ;
  assign y14701 = n51142 ;
  assign y14702 = n51146 ;
  assign y14703 = ~n51148 ;
  assign y14704 = ~n51149 ;
  assign y14705 = ~1'b0 ;
  assign y14706 = n51152 ;
  assign y14707 = n51162 ;
  assign y14708 = n51164 ;
  assign y14709 = ~n51165 ;
  assign y14710 = n51166 ;
  assign y14711 = ~n51168 ;
  assign y14712 = ~n51170 ;
  assign y14713 = ~n51172 ;
  assign y14714 = ~1'b0 ;
  assign y14715 = n51176 ;
  assign y14716 = ~n51178 ;
  assign y14717 = ~n51180 ;
  assign y14718 = n51183 ;
  assign y14719 = ~n51185 ;
  assign y14720 = ~n51188 ;
  assign y14721 = ~1'b0 ;
  assign y14722 = n51191 ;
  assign y14723 = ~1'b0 ;
  assign y14724 = ~n51192 ;
  assign y14725 = ~n51195 ;
  assign y14726 = ~n51196 ;
  assign y14727 = ~n51197 ;
  assign y14728 = n51198 ;
  assign y14729 = n51205 ;
  assign y14730 = n51207 ;
  assign y14731 = ~n51209 ;
  assign y14732 = n51211 ;
  assign y14733 = n51212 ;
  assign y14734 = ~n51213 ;
  assign y14735 = n51222 ;
  assign y14736 = ~n51223 ;
  assign y14737 = n51224 ;
  assign y14738 = ~n51229 ;
  assign y14739 = ~n51230 ;
  assign y14740 = ~n51231 ;
  assign y14741 = ~n51233 ;
  assign y14742 = ~n51237 ;
  assign y14743 = ~n51241 ;
  assign y14744 = n51244 ;
  assign y14745 = ~n51247 ;
  assign y14746 = ~n51249 ;
  assign y14747 = ~n51250 ;
  assign y14748 = n51258 ;
  assign y14749 = ~n51259 ;
  assign y14750 = ~n51261 ;
  assign y14751 = ~1'b0 ;
  assign y14752 = n51262 ;
  assign y14753 = n51268 ;
  assign y14754 = n51272 ;
  assign y14755 = ~n51277 ;
  assign y14756 = n51280 ;
  assign y14757 = ~n51282 ;
  assign y14758 = n51285 ;
  assign y14759 = n51288 ;
  assign y14760 = n51291 ;
  assign y14761 = ~1'b0 ;
  assign y14762 = ~n51294 ;
  assign y14763 = n51297 ;
  assign y14764 = n51302 ;
  assign y14765 = n51305 ;
  assign y14766 = ~n51308 ;
  assign y14767 = n51309 ;
  assign y14768 = n51311 ;
  assign y14769 = ~n51316 ;
  assign y14770 = ~1'b0 ;
  assign y14771 = n51319 ;
  assign y14772 = ~n51321 ;
  assign y14773 = n51326 ;
  assign y14774 = ~n51327 ;
  assign y14775 = ~n51329 ;
  assign y14776 = n51331 ;
  assign y14777 = ~n51337 ;
  assign y14778 = ~n51338 ;
  assign y14779 = n51339 ;
  assign y14780 = ~n51349 ;
  assign y14781 = ~n51353 ;
  assign y14782 = n51355 ;
  assign y14783 = ~n51359 ;
  assign y14784 = ~n51360 ;
  assign y14785 = n51364 ;
  assign y14786 = ~n51366 ;
  assign y14787 = n51369 ;
  assign y14788 = n51375 ;
  assign y14789 = ~n51377 ;
  assign y14790 = ~1'b0 ;
  assign y14791 = ~n51380 ;
  assign y14792 = n51381 ;
  assign y14793 = n51382 ;
  assign y14794 = ~n51385 ;
  assign y14795 = n51386 ;
  assign y14796 = ~n51387 ;
  assign y14797 = n51392 ;
  assign y14798 = ~n51402 ;
  assign y14799 = n51407 ;
  assign y14800 = n51408 ;
  assign y14801 = ~n51410 ;
  assign y14802 = n51412 ;
  assign y14803 = n51414 ;
  assign y14804 = n51415 ;
  assign y14805 = ~n51417 ;
  assign y14806 = n51420 ;
  assign y14807 = n51425 ;
  assign y14808 = n51429 ;
  assign y14809 = ~n51431 ;
  assign y14810 = n51432 ;
  assign y14811 = ~n51437 ;
  assign y14812 = n51438 ;
  assign y14813 = n51443 ;
  assign y14814 = n51444 ;
  assign y14815 = n51448 ;
  assign y14816 = n51453 ;
  assign y14817 = ~n51457 ;
  assign y14818 = ~n51459 ;
  assign y14819 = ~n51463 ;
  assign y14820 = ~1'b0 ;
  assign y14821 = ~1'b0 ;
  assign y14822 = ~1'b0 ;
  assign y14823 = ~n51469 ;
  assign y14824 = ~n51472 ;
  assign y14825 = n51473 ;
  assign y14826 = ~n51475 ;
  assign y14827 = n51479 ;
  assign y14828 = ~n51480 ;
  assign y14829 = n51482 ;
  assign y14830 = ~1'b0 ;
  assign y14831 = n51484 ;
  assign y14832 = n51485 ;
  assign y14833 = n51486 ;
  assign y14834 = ~n51487 ;
  assign y14835 = n51488 ;
  assign y14836 = n51496 ;
  assign y14837 = ~n51500 ;
  assign y14838 = n51505 ;
  assign y14839 = ~n51506 ;
  assign y14840 = n51507 ;
  assign y14841 = ~n51510 ;
  assign y14842 = ~n51511 ;
  assign y14843 = n51515 ;
  assign y14844 = ~n51516 ;
  assign y14845 = ~n51519 ;
  assign y14846 = n51523 ;
  assign y14847 = n51524 ;
  assign y14848 = ~n51525 ;
  assign y14849 = ~n51528 ;
  assign y14850 = ~n51531 ;
  assign y14851 = ~1'b0 ;
  assign y14852 = ~1'b0 ;
  assign y14853 = ~n51532 ;
  assign y14854 = ~n51536 ;
  assign y14855 = n51537 ;
  assign y14856 = n51538 ;
  assign y14857 = ~n51539 ;
  assign y14858 = n51540 ;
  assign y14859 = n51541 ;
  assign y14860 = ~n51543 ;
  assign y14861 = n51545 ;
  assign y14862 = n51550 ;
  assign y14863 = n51552 ;
  assign y14864 = n51555 ;
  assign y14865 = n51556 ;
  assign y14866 = n51559 ;
  assign y14867 = ~n51560 ;
  assign y14868 = n51561 ;
  assign y14869 = ~n51565 ;
  assign y14870 = n51569 ;
  assign y14871 = n51571 ;
  assign y14872 = n51573 ;
  assign y14873 = n51578 ;
  assign y14874 = ~n51579 ;
  assign y14875 = ~n51580 ;
  assign y14876 = ~n51581 ;
  assign y14877 = ~n51583 ;
  assign y14878 = n51584 ;
  assign y14879 = n51588 ;
  assign y14880 = n51590 ;
  assign y14881 = ~n51591 ;
  assign y14882 = n51592 ;
  assign y14883 = ~n51594 ;
  assign y14884 = ~n51599 ;
  assign y14885 = ~n51603 ;
  assign y14886 = ~n51606 ;
  assign y14887 = n51609 ;
  assign y14888 = ~n51612 ;
  assign y14889 = n51613 ;
  assign y14890 = n51614 ;
  assign y14891 = ~1'b0 ;
  assign y14892 = ~n51618 ;
  assign y14893 = n51620 ;
  assign y14894 = n51621 ;
  assign y14895 = n51623 ;
  assign y14896 = n51627 ;
  assign y14897 = ~n51630 ;
  assign y14898 = n51631 ;
  assign y14899 = ~n51634 ;
  assign y14900 = ~n51636 ;
  assign y14901 = ~n51638 ;
  assign y14902 = ~n51643 ;
  assign y14903 = ~n51646 ;
  assign y14904 = n51647 ;
  assign y14905 = n51650 ;
  assign y14906 = n51653 ;
  assign y14907 = ~n51663 ;
  assign y14908 = n51665 ;
  assign y14909 = n51670 ;
  assign y14910 = n51672 ;
  assign y14911 = n51674 ;
  assign y14912 = ~n51677 ;
  assign y14913 = ~1'b0 ;
  assign y14914 = ~n51678 ;
  assign y14915 = n51679 ;
  assign y14916 = ~n51680 ;
  assign y14917 = n51682 ;
  assign y14918 = ~n51684 ;
  assign y14919 = n51685 ;
  assign y14920 = n51686 ;
  assign y14921 = n51687 ;
  assign y14922 = ~n51690 ;
  assign y14923 = ~n51692 ;
  assign y14924 = ~n51694 ;
  assign y14925 = ~n51697 ;
  assign y14926 = n51698 ;
  assign y14927 = ~n51699 ;
  assign y14928 = ~n51703 ;
  assign y14929 = ~n51704 ;
  assign y14930 = ~n51710 ;
  assign y14931 = n51714 ;
  assign y14932 = n51716 ;
  assign y14933 = ~n51721 ;
  assign y14934 = n51725 ;
  assign y14935 = n51729 ;
  assign y14936 = ~n51731 ;
  assign y14937 = n51732 ;
  assign y14938 = n51734 ;
  assign y14939 = ~n51736 ;
  assign y14940 = ~n51737 ;
  assign y14941 = ~n51740 ;
  assign y14942 = ~1'b0 ;
  assign y14943 = ~n51742 ;
  assign y14944 = ~n51744 ;
  assign y14945 = ~n51745 ;
  assign y14946 = n51746 ;
  assign y14947 = ~n51747 ;
  assign y14948 = n51750 ;
  assign y14949 = ~n51752 ;
  assign y14950 = ~n51754 ;
  assign y14951 = ~n51755 ;
  assign y14952 = n51757 ;
  assign y14953 = ~n51762 ;
  assign y14954 = n51763 ;
  assign y14955 = ~n51764 ;
  assign y14956 = n51768 ;
  assign y14957 = ~n51769 ;
  assign y14958 = ~n51770 ;
  assign y14959 = ~n51771 ;
  assign y14960 = n51772 ;
  assign y14961 = ~n51776 ;
  assign y14962 = ~n51778 ;
  assign y14963 = ~1'b0 ;
  assign y14964 = ~1'b0 ;
  assign y14965 = n51780 ;
  assign y14966 = n51783 ;
  assign y14967 = n51791 ;
  assign y14968 = ~n51794 ;
  assign y14969 = n51796 ;
  assign y14970 = ~n51799 ;
  assign y14971 = ~n51801 ;
  assign y14972 = ~n51802 ;
  assign y14973 = ~n51805 ;
  assign y14974 = ~1'b0 ;
  assign y14975 = ~n51806 ;
  assign y14976 = n51807 ;
  assign y14977 = n51808 ;
  assign y14978 = ~n51809 ;
  assign y14979 = n51812 ;
  assign y14980 = n51816 ;
  assign y14981 = ~n51821 ;
  assign y14982 = ~n51823 ;
  assign y14983 = ~1'b0 ;
  assign y14984 = n51825 ;
  assign y14985 = ~n51829 ;
  assign y14986 = n51833 ;
  assign y14987 = ~n51834 ;
  assign y14988 = ~n51838 ;
  assign y14989 = ~n51840 ;
  assign y14990 = n51841 ;
  assign y14991 = ~n51842 ;
  assign y14992 = ~n51844 ;
  assign y14993 = n51846 ;
  assign y14994 = ~n51848 ;
  assign y14995 = ~n16870 ;
  assign y14996 = n51852 ;
  assign y14997 = n51853 ;
  assign y14998 = n51857 ;
  assign y14999 = n51859 ;
  assign y15000 = ~n51860 ;
  assign y15001 = n51862 ;
  assign y15002 = n51864 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = ~1'b0 ;
  assign y15005 = ~1'b0 ;
  assign y15006 = n51865 ;
  assign y15007 = ~n51866 ;
  assign y15008 = ~n51867 ;
  assign y15009 = n51871 ;
  assign y15010 = ~n51872 ;
  assign y15011 = ~n51873 ;
  assign y15012 = n51875 ;
  assign y15013 = n51878 ;
  assign y15014 = n51880 ;
  assign y15015 = n51884 ;
  assign y15016 = ~n51886 ;
  assign y15017 = ~n51892 ;
  assign y15018 = n51893 ;
  assign y15019 = n51895 ;
  assign y15020 = ~n51896 ;
  assign y15021 = n51897 ;
  assign y15022 = n51899 ;
  assign y15023 = n51901 ;
  assign y15024 = ~n51905 ;
  assign y15025 = ~1'b0 ;
  assign y15026 = ~n51907 ;
  assign y15027 = ~n51909 ;
  assign y15028 = n51913 ;
  assign y15029 = ~n51917 ;
  assign y15030 = ~n51920 ;
  assign y15031 = n51922 ;
  assign y15032 = ~n51926 ;
  assign y15033 = n51930 ;
  assign y15034 = ~n51931 ;
  assign y15035 = ~n51933 ;
  assign y15036 = n51934 ;
  assign y15037 = ~1'b0 ;
  assign y15038 = ~n51941 ;
  assign y15039 = ~n51947 ;
  assign y15040 = ~n51948 ;
  assign y15041 = ~n51949 ;
  assign y15042 = ~n51950 ;
  assign y15043 = n51951 ;
  assign y15044 = ~n51952 ;
  assign y15045 = ~n51960 ;
  assign y15046 = ~n51962 ;
  assign y15047 = ~1'b0 ;
  assign y15048 = ~1'b0 ;
  assign y15049 = ~n51964 ;
  assign y15050 = n51966 ;
  assign y15051 = ~n51967 ;
  assign y15052 = ~n51972 ;
  assign y15053 = ~n51975 ;
  assign y15054 = ~n51976 ;
  assign y15055 = n51978 ;
  assign y15056 = ~n51981 ;
  assign y15057 = ~n51983 ;
  assign y15058 = ~1'b0 ;
  assign y15059 = ~n51987 ;
  assign y15060 = ~n51991 ;
  assign y15061 = ~n51992 ;
  assign y15062 = ~n51994 ;
  assign y15063 = ~n51996 ;
  assign y15064 = ~n52002 ;
  assign y15065 = ~n52006 ;
  assign y15066 = n52007 ;
  assign y15067 = ~1'b0 ;
  assign y15068 = ~n52008 ;
  assign y15069 = ~n52010 ;
  assign y15070 = ~n52016 ;
  assign y15071 = ~n52017 ;
  assign y15072 = ~n52018 ;
  assign y15073 = ~n52022 ;
  assign y15074 = n52023 ;
  assign y15075 = n52025 ;
  assign y15076 = n52027 ;
  assign y15077 = ~1'b0 ;
  assign y15078 = n52032 ;
  assign y15079 = ~n52034 ;
  assign y15080 = n52035 ;
  assign y15081 = ~n52036 ;
  assign y15082 = ~n52037 ;
  assign y15083 = ~n52041 ;
  assign y15084 = ~n52042 ;
  assign y15085 = n52044 ;
  assign y15086 = ~n52046 ;
  assign y15087 = n52047 ;
  assign y15088 = ~n52049 ;
  assign y15089 = ~n52051 ;
  assign y15090 = ~n52052 ;
  assign y15091 = n52054 ;
  assign y15092 = ~n52055 ;
  assign y15093 = n52056 ;
  assign y15094 = n52061 ;
  assign y15095 = n52065 ;
  assign y15096 = n52066 ;
  assign y15097 = ~n52067 ;
  assign y15098 = n52070 ;
  assign y15099 = n52076 ;
  assign y15100 = ~n52077 ;
  assign y15101 = n52080 ;
  assign y15102 = ~n52082 ;
  assign y15103 = n52084 ;
  assign y15104 = ~n52086 ;
  assign y15105 = ~1'b0 ;
  assign y15106 = ~n52089 ;
  assign y15107 = n52090 ;
  assign y15108 = ~n52091 ;
  assign y15109 = n52092 ;
  assign y15110 = ~n52093 ;
  assign y15111 = n52095 ;
  assign y15112 = ~n52097 ;
  assign y15113 = n52099 ;
  assign y15114 = n52102 ;
  assign y15115 = n52104 ;
  assign y15116 = n52107 ;
  assign y15117 = ~n52109 ;
  assign y15118 = ~n52110 ;
  assign y15119 = ~n52114 ;
  assign y15120 = n52115 ;
  assign y15121 = n52117 ;
  assign y15122 = ~n52121 ;
  assign y15123 = n52123 ;
  assign y15124 = ~n52124 ;
  assign y15125 = n52125 ;
  assign y15126 = n52127 ;
  assign y15127 = ~1'b0 ;
  assign y15128 = ~n52129 ;
  assign y15129 = ~n52132 ;
  assign y15130 = n52135 ;
  assign y15131 = n52136 ;
  assign y15132 = n52141 ;
  assign y15133 = ~n52142 ;
  assign y15134 = ~n52144 ;
  assign y15135 = ~n52145 ;
  assign y15136 = n52153 ;
  assign y15137 = ~1'b0 ;
  assign y15138 = ~n52155 ;
  assign y15139 = n52159 ;
  assign y15140 = ~n52164 ;
  assign y15141 = ~n23656 ;
  assign y15142 = ~n52165 ;
  assign y15143 = n52167 ;
  assign y15144 = ~n52170 ;
  assign y15145 = n52174 ;
  assign y15146 = ~n52175 ;
  assign y15147 = n52176 ;
  assign y15148 = ~1'b0 ;
  assign y15149 = ~1'b0 ;
  assign y15150 = ~n52184 ;
  assign y15151 = ~n52188 ;
  assign y15152 = ~n52189 ;
  assign y15153 = n52190 ;
  assign y15154 = n52191 ;
  assign y15155 = ~n52197 ;
  assign y15156 = n52200 ;
  assign y15157 = ~n52201 ;
  assign y15158 = n52204 ;
  assign y15159 = n52206 ;
  assign y15160 = ~n52208 ;
  assign y15161 = ~n52210 ;
  assign y15162 = ~n52211 ;
  assign y15163 = ~n52212 ;
  assign y15164 = n52217 ;
  assign y15165 = ~n52218 ;
  assign y15166 = ~n52221 ;
  assign y15167 = ~1'b0 ;
  assign y15168 = ~1'b0 ;
  assign y15169 = ~n52223 ;
  assign y15170 = n52224 ;
  assign y15171 = ~n52229 ;
  assign y15172 = n52232 ;
  assign y15173 = n52233 ;
  assign y15174 = ~n52234 ;
  assign y15175 = ~n52235 ;
  assign y15176 = ~n52236 ;
  assign y15177 = ~n52237 ;
  assign y15178 = ~n52239 ;
  assign y15179 = n52241 ;
  assign y15180 = ~n52243 ;
  assign y15181 = n52244 ;
  assign y15182 = n52245 ;
  assign y15183 = n52247 ;
  assign y15184 = n52248 ;
  assign y15185 = n52251 ;
  assign y15186 = n52252 ;
  assign y15187 = n52254 ;
  assign y15188 = ~n52255 ;
  assign y15189 = ~n52257 ;
  assign y15190 = n52259 ;
  assign y15191 = n52260 ;
  assign y15192 = n52261 ;
  assign y15193 = ~n52262 ;
  assign y15194 = ~n52265 ;
  assign y15195 = n52266 ;
  assign y15196 = n52267 ;
  assign y15197 = n52273 ;
  assign y15198 = n52274 ;
  assign y15199 = ~1'b0 ;
  assign y15200 = n52275 ;
  assign y15201 = ~n52277 ;
  assign y15202 = ~n52280 ;
  assign y15203 = n52284 ;
  assign y15204 = n52290 ;
  assign y15205 = n52291 ;
  assign y15206 = ~n52292 ;
  assign y15207 = ~n52294 ;
  assign y15208 = ~n52296 ;
  assign y15209 = ~n52298 ;
  assign y15210 = ~n52300 ;
  assign y15211 = ~n52301 ;
  assign y15212 = ~n52302 ;
  assign y15213 = n52303 ;
  assign y15214 = ~n52306 ;
  assign y15215 = n52311 ;
  assign y15216 = ~n52314 ;
  assign y15217 = ~n52317 ;
  assign y15218 = n52319 ;
  assign y15219 = ~n52321 ;
  assign y15220 = ~1'b0 ;
  assign y15221 = ~n52325 ;
  assign y15222 = n52328 ;
  assign y15223 = n52333 ;
  assign y15224 = n52336 ;
  assign y15225 = n52339 ;
  assign y15226 = n52343 ;
  assign y15227 = ~n52344 ;
  assign y15228 = n52346 ;
  assign y15229 = ~n52348 ;
  assign y15230 = ~1'b0 ;
  assign y15231 = n52351 ;
  assign y15232 = n52353 ;
  assign y15233 = n52354 ;
  assign y15234 = n52355 ;
  assign y15235 = n52359 ;
  assign y15236 = n52360 ;
  assign y15237 = n52361 ;
  assign y15238 = ~n52363 ;
  assign y15239 = ~n52365 ;
  assign y15240 = ~n52368 ;
  assign y15241 = ~n52370 ;
  assign y15242 = n52374 ;
  assign y15243 = n52376 ;
  assign y15244 = ~n52377 ;
  assign y15245 = n52379 ;
  assign y15246 = n52383 ;
  assign y15247 = n52384 ;
  assign y15248 = ~n52387 ;
  assign y15249 = ~n40559 ;
  assign y15250 = n52389 ;
  assign y15251 = n52392 ;
  assign y15252 = ~n52393 ;
  assign y15253 = ~n52394 ;
  assign y15254 = ~n52395 ;
  assign y15255 = ~n52398 ;
  assign y15256 = ~n52399 ;
  assign y15257 = n52402 ;
  assign y15258 = n52404 ;
  assign y15259 = ~1'b0 ;
  assign y15260 = ~n52407 ;
  assign y15261 = n52409 ;
  assign y15262 = ~n52410 ;
  assign y15263 = n52411 ;
  assign y15264 = n52412 ;
  assign y15265 = n52413 ;
  assign y15266 = n52415 ;
  assign y15267 = n52418 ;
  assign y15268 = n52421 ;
  assign y15269 = n52423 ;
  assign y15270 = n52424 ;
  assign y15271 = n52426 ;
  assign y15272 = n52427 ;
  assign y15273 = ~n52429 ;
  assign y15274 = n52430 ;
  assign y15275 = ~n52431 ;
  assign y15276 = n52433 ;
  assign y15277 = ~n52434 ;
  assign y15278 = ~n52436 ;
  assign y15279 = ~1'b0 ;
  assign y15280 = n52437 ;
  assign y15281 = n52440 ;
  assign y15282 = ~n52441 ;
  assign y15283 = n52442 ;
  assign y15284 = ~n52444 ;
  assign y15285 = ~n52446 ;
  assign y15286 = n52449 ;
  assign y15287 = ~1'b0 ;
  assign y15288 = n52454 ;
  assign y15289 = ~1'b0 ;
  assign y15290 = n52455 ;
  assign y15291 = n52456 ;
  assign y15292 = n52461 ;
  assign y15293 = n52463 ;
  assign y15294 = n52464 ;
  assign y15295 = n52468 ;
  assign y15296 = ~n52469 ;
  assign y15297 = ~n52473 ;
  assign y15298 = ~n52475 ;
  assign y15299 = n52477 ;
  assign y15300 = ~n52478 ;
  assign y15301 = n52480 ;
  assign y15302 = n52488 ;
  assign y15303 = n52489 ;
  assign y15304 = ~n52493 ;
  assign y15305 = ~n52499 ;
  assign y15306 = ~n52500 ;
  assign y15307 = ~n52501 ;
  assign y15308 = ~1'b0 ;
  assign y15309 = ~n52503 ;
  assign y15310 = ~1'b0 ;
  assign y15311 = ~n52504 ;
  assign y15312 = ~n52505 ;
  assign y15313 = n52506 ;
  assign y15314 = ~n52507 ;
  assign y15315 = ~n52508 ;
  assign y15316 = n52509 ;
  assign y15317 = ~n52510 ;
  assign y15318 = ~1'b0 ;
  assign y15319 = n52511 ;
  assign y15320 = n52514 ;
  assign y15321 = ~n52515 ;
  assign y15322 = ~n52518 ;
  assign y15323 = n52523 ;
  assign y15324 = n52524 ;
  assign y15325 = ~n52528 ;
  assign y15326 = n52529 ;
  assign y15327 = ~n52530 ;
  assign y15328 = n52533 ;
  assign y15329 = ~1'b0 ;
  assign y15330 = ~n52535 ;
  assign y15331 = n52537 ;
  assign y15332 = ~n52540 ;
  assign y15333 = ~n52541 ;
  assign y15334 = n52548 ;
  assign y15335 = n52549 ;
  assign y15336 = ~n52552 ;
  assign y15337 = ~n52555 ;
  assign y15338 = n52557 ;
  assign y15339 = ~n52559 ;
  assign y15340 = n52563 ;
  assign y15341 = n52564 ;
  assign y15342 = n52566 ;
  assign y15343 = n52567 ;
  assign y15344 = ~n52568 ;
  assign y15345 = ~n52572 ;
  assign y15346 = ~n52573 ;
  assign y15347 = ~n52575 ;
  assign y15348 = ~n52577 ;
  assign y15349 = n52579 ;
  assign y15350 = ~n52581 ;
  assign y15351 = ~1'b0 ;
  assign y15352 = n52582 ;
  assign y15353 = ~n52584 ;
  assign y15354 = ~n52586 ;
  assign y15355 = ~n52589 ;
  assign y15356 = ~n52591 ;
  assign y15357 = ~n52593 ;
  assign y15358 = n52594 ;
  assign y15359 = ~n52595 ;
  assign y15360 = ~n52597 ;
  assign y15361 = ~n52598 ;
  assign y15362 = n52599 ;
  assign y15363 = n52603 ;
  assign y15364 = n52605 ;
  assign y15365 = n52608 ;
  assign y15366 = ~n40856 ;
  assign y15367 = ~n52611 ;
  assign y15368 = n52613 ;
  assign y15369 = ~n52614 ;
  assign y15370 = ~n52616 ;
  assign y15371 = n52619 ;
  assign y15372 = ~n52623 ;
  assign y15373 = ~1'b0 ;
  assign y15374 = n52625 ;
  assign y15375 = ~n52627 ;
  assign y15376 = ~n52630 ;
  assign y15377 = n52631 ;
  assign y15378 = n52634 ;
  assign y15379 = n52638 ;
  assign y15380 = ~n8677 ;
  assign y15381 = n52641 ;
  assign y15382 = n52645 ;
  assign y15383 = n52647 ;
  assign y15384 = n52648 ;
  assign y15385 = ~n52650 ;
  assign y15386 = ~n52652 ;
  assign y15387 = ~n52653 ;
  assign y15388 = ~n52654 ;
  assign y15389 = n52657 ;
  assign y15390 = ~n52660 ;
  assign y15391 = ~n52661 ;
  assign y15392 = ~1'b0 ;
  assign y15393 = n52663 ;
  assign y15394 = ~1'b0 ;
  assign y15395 = n52669 ;
  assign y15396 = ~n52672 ;
  assign y15397 = n52673 ;
  assign y15398 = n52677 ;
  assign y15399 = n52682 ;
  assign y15400 = ~n52683 ;
  assign y15401 = n52685 ;
  assign y15402 = ~n52687 ;
  assign y15403 = ~n52689 ;
  assign y15404 = ~n52691 ;
  assign y15405 = n52693 ;
  assign y15406 = ~n52694 ;
  assign y15407 = n52697 ;
  assign y15408 = ~n52698 ;
  assign y15409 = n52699 ;
  assign y15410 = ~n52700 ;
  assign y15411 = ~n52701 ;
  assign y15412 = n52704 ;
  assign y15413 = ~n52707 ;
  assign y15414 = n52708 ;
  assign y15415 = ~n52710 ;
  assign y15416 = n52713 ;
  assign y15417 = ~n52715 ;
  assign y15418 = n52716 ;
  assign y15419 = n52719 ;
  assign y15420 = ~n52720 ;
  assign y15421 = n52722 ;
  assign y15422 = ~n52725 ;
  assign y15423 = ~n52727 ;
  assign y15424 = n52732 ;
  assign y15425 = ~n52734 ;
  assign y15426 = n52738 ;
  assign y15427 = ~n52739 ;
  assign y15428 = ~n52741 ;
  assign y15429 = n52742 ;
  assign y15430 = ~n52745 ;
  assign y15431 = ~n52746 ;
  assign y15432 = n52747 ;
  assign y15433 = ~n52749 ;
  assign y15434 = n52750 ;
  assign y15435 = ~n52751 ;
  assign y15436 = ~n52752 ;
  assign y15437 = n52760 ;
  assign y15438 = ~n52765 ;
  assign y15439 = ~n52766 ;
  assign y15440 = n52767 ;
  assign y15441 = ~n52770 ;
  assign y15442 = ~n52771 ;
  assign y15443 = ~n52773 ;
  assign y15444 = n52778 ;
  assign y15445 = ~n52782 ;
  assign y15446 = ~n52783 ;
  assign y15447 = n52786 ;
  assign y15448 = n52787 ;
  assign y15449 = n52791 ;
  assign y15450 = n52798 ;
  assign y15451 = ~n52799 ;
  assign y15452 = ~n52801 ;
  assign y15453 = n52803 ;
  assign y15454 = n52807 ;
  assign y15455 = ~n52813 ;
  assign y15456 = n52815 ;
  assign y15457 = n52817 ;
  assign y15458 = ~n9296 ;
  assign y15459 = ~n52821 ;
  assign y15460 = n52825 ;
  assign y15461 = n52826 ;
  assign y15462 = ~n52829 ;
  assign y15463 = n52833 ;
  assign y15464 = ~n52835 ;
  assign y15465 = ~1'b0 ;
  assign y15466 = ~n52838 ;
  assign y15467 = n52839 ;
  assign y15468 = n52840 ;
  assign y15469 = ~n52842 ;
  assign y15470 = n52843 ;
  assign y15471 = n52852 ;
  assign y15472 = n52853 ;
  assign y15473 = ~n52854 ;
  assign y15474 = n52857 ;
  assign y15475 = n52859 ;
  assign y15476 = ~n52860 ;
  assign y15477 = n52861 ;
  assign y15478 = n52863 ;
  assign y15479 = n52866 ;
  assign y15480 = n52867 ;
  assign y15481 = n52869 ;
  assign y15482 = n52870 ;
  assign y15483 = ~n52874 ;
  assign y15484 = ~n52879 ;
  assign y15485 = ~n52881 ;
  assign y15486 = ~n52883 ;
  assign y15487 = ~n52885 ;
  assign y15488 = n52886 ;
  assign y15489 = ~n52890 ;
  assign y15490 = n52892 ;
  assign y15491 = n52894 ;
  assign y15492 = ~n52895 ;
  assign y15493 = ~n52897 ;
  assign y15494 = n52899 ;
  assign y15495 = n52901 ;
  assign y15496 = ~1'b0 ;
  assign y15497 = n41387 ;
  assign y15498 = ~n52902 ;
  assign y15499 = ~n52904 ;
  assign y15500 = ~n52906 ;
  assign y15501 = n52909 ;
  assign y15502 = ~n52914 ;
  assign y15503 = ~n52922 ;
  assign y15504 = n52923 ;
  assign y15505 = ~n52924 ;
  assign y15506 = ~n52929 ;
  assign y15507 = ~n52931 ;
  assign y15508 = n52933 ;
  assign y15509 = n52934 ;
  assign y15510 = ~n52938 ;
  assign y15511 = n52939 ;
  assign y15512 = ~n52940 ;
  assign y15513 = ~n52944 ;
  assign y15514 = ~n52945 ;
  assign y15515 = ~n52951 ;
  assign y15516 = ~1'b0 ;
  assign y15517 = n52954 ;
  assign y15518 = ~n52956 ;
  assign y15519 = n52962 ;
  assign y15520 = n52964 ;
  assign y15521 = n52967 ;
  assign y15522 = n52971 ;
  assign y15523 = n52973 ;
  assign y15524 = n52976 ;
  assign y15525 = ~1'b0 ;
  assign y15526 = n52984 ;
  assign y15527 = ~n52990 ;
  assign y15528 = ~n52992 ;
  assign y15529 = ~n52993 ;
  assign y15530 = ~n52996 ;
  assign y15531 = n52998 ;
  assign y15532 = ~n52999 ;
  assign y15533 = ~n53003 ;
  assign y15534 = ~n53006 ;
  assign y15535 = ~n53008 ;
  assign y15536 = n53012 ;
  assign y15537 = ~n53016 ;
  assign y15538 = n53017 ;
  assign y15539 = ~n53018 ;
  assign y15540 = ~n53019 ;
  assign y15541 = ~n53020 ;
  assign y15542 = n53022 ;
  assign y15543 = n53025 ;
  assign y15544 = ~1'b0 ;
  assign y15545 = n53027 ;
  assign y15546 = ~n53030 ;
  assign y15547 = ~n53031 ;
  assign y15548 = ~n53034 ;
  assign y15549 = ~n53036 ;
  assign y15550 = n53039 ;
  assign y15551 = n53040 ;
  assign y15552 = n53044 ;
  assign y15553 = ~n53046 ;
  assign y15554 = n53050 ;
  assign y15555 = ~n53054 ;
  assign y15556 = ~n53056 ;
  assign y15557 = n53059 ;
  assign y15558 = ~n53063 ;
  assign y15559 = ~n53068 ;
  assign y15560 = n53072 ;
  assign y15561 = ~n53073 ;
  assign y15562 = ~n53075 ;
  assign y15563 = n53077 ;
  assign y15564 = n53080 ;
  assign y15565 = ~n53084 ;
  assign y15566 = n53085 ;
  assign y15567 = ~n53089 ;
  assign y15568 = n53094 ;
  assign y15569 = ~n53099 ;
  assign y15570 = n53100 ;
  assign y15571 = n53101 ;
  assign y15572 = ~n53103 ;
  assign y15573 = n53105 ;
  assign y15574 = ~n53107 ;
  assign y15575 = n53109 ;
  assign y15576 = n53113 ;
  assign y15577 = ~n53119 ;
  assign y15578 = n53124 ;
  assign y15579 = n53125 ;
  assign y15580 = n53126 ;
  assign y15581 = n53127 ;
  assign y15582 = n53128 ;
  assign y15583 = ~n53129 ;
  assign y15584 = ~1'b0 ;
  assign y15585 = ~n53133 ;
  assign y15586 = n53136 ;
  assign y15587 = ~n53137 ;
  assign y15588 = n53139 ;
  assign y15589 = ~n53140 ;
  assign y15590 = n53144 ;
  assign y15591 = n53146 ;
  assign y15592 = n53147 ;
  assign y15593 = n53149 ;
  assign y15594 = ~n53154 ;
  assign y15595 = ~1'b0 ;
  assign y15596 = n53157 ;
  assign y15597 = ~n53158 ;
  assign y15598 = n53159 ;
  assign y15599 = ~n53161 ;
  assign y15600 = ~n53164 ;
  assign y15601 = ~n53166 ;
  assign y15602 = n53167 ;
  assign y15603 = ~n53173 ;
  assign y15604 = ~n53179 ;
  assign y15605 = n53182 ;
  assign y15606 = n53185 ;
  assign y15607 = ~n53187 ;
  assign y15608 = n53188 ;
  assign y15609 = ~n53190 ;
  assign y15610 = ~n53191 ;
  assign y15611 = n53192 ;
  assign y15612 = n53193 ;
  assign y15613 = n53199 ;
  assign y15614 = ~n53200 ;
  assign y15615 = ~1'b0 ;
  assign y15616 = ~n53202 ;
  assign y15617 = ~1'b0 ;
  assign y15618 = ~n53203 ;
  assign y15619 = ~n53205 ;
  assign y15620 = n53207 ;
  assign y15621 = ~n53209 ;
  assign y15622 = n53211 ;
  assign y15623 = n53214 ;
  assign y15624 = n53221 ;
  assign y15625 = ~n53222 ;
  assign y15626 = n53226 ;
  assign y15627 = ~n53229 ;
  assign y15628 = ~1'b0 ;
  assign y15629 = ~n53230 ;
  assign y15630 = n53233 ;
  assign y15631 = n53237 ;
  assign y15632 = n53239 ;
  assign y15633 = ~n53242 ;
  assign y15634 = ~n53250 ;
  assign y15635 = ~n53251 ;
  assign y15636 = ~1'b0 ;
  assign y15637 = ~1'b0 ;
  assign y15638 = ~n53260 ;
  assign y15639 = n53263 ;
  assign y15640 = n53265 ;
  assign y15641 = ~n53266 ;
  assign y15642 = n53270 ;
  assign y15643 = n53273 ;
  assign y15644 = n53274 ;
  assign y15645 = ~1'b0 ;
  assign y15646 = ~n53277 ;
  assign y15647 = ~1'b0 ;
  assign y15648 = ~n53281 ;
  assign y15649 = ~n53288 ;
  assign y15650 = ~n53292 ;
  assign y15651 = n53295 ;
  assign y15652 = ~n53296 ;
  assign y15653 = n53297 ;
  assign y15654 = ~n53299 ;
  assign y15655 = ~1'b0 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = ~n53303 ;
  assign y15658 = n53305 ;
  assign y15659 = n53307 ;
  assign y15660 = n53308 ;
  assign y15661 = n53309 ;
  assign y15662 = ~n53310 ;
  assign y15663 = ~n53315 ;
  assign y15664 = n53316 ;
  assign y15665 = ~n53318 ;
  assign y15666 = n53320 ;
  assign y15667 = n53322 ;
  assign y15668 = n53324 ;
  assign y15669 = ~n53326 ;
  assign y15670 = n53327 ;
  assign y15671 = n53328 ;
  assign y15672 = n53329 ;
  assign y15673 = ~n53331 ;
  assign y15674 = n53336 ;
  assign y15675 = ~n53337 ;
  assign y15676 = n53344 ;
  assign y15677 = n53346 ;
  assign y15678 = ~n53349 ;
  assign y15679 = n53350 ;
  assign y15680 = n53352 ;
  assign y15681 = ~n53357 ;
  assign y15682 = ~n53358 ;
  assign y15683 = n53361 ;
  assign y15684 = n53362 ;
  assign y15685 = ~n53365 ;
  assign y15686 = ~n53367 ;
  assign y15687 = n53371 ;
  assign y15688 = n53373 ;
  assign y15689 = ~n53379 ;
  assign y15690 = n53380 ;
  assign y15691 = ~n53383 ;
  assign y15692 = n53386 ;
  assign y15693 = n53387 ;
  assign y15694 = n53390 ;
  assign y15695 = n53396 ;
  assign y15696 = ~n53402 ;
  assign y15697 = ~1'b0 ;
  assign y15698 = n53407 ;
  assign y15699 = ~n53411 ;
  assign y15700 = n53415 ;
  assign y15701 = ~n53417 ;
  assign y15702 = n53422 ;
  assign y15703 = n53425 ;
  assign y15704 = n53430 ;
  assign y15705 = ~n53435 ;
  assign y15706 = n53438 ;
  assign y15707 = ~1'b0 ;
  assign y15708 = ~n53441 ;
  assign y15709 = n53442 ;
  assign y15710 = n53443 ;
  assign y15711 = ~n53446 ;
  assign y15712 = ~n53448 ;
  assign y15713 = ~n53449 ;
  assign y15714 = ~n53450 ;
  assign y15715 = n53451 ;
  assign y15716 = ~n53455 ;
  assign y15717 = ~1'b0 ;
  assign y15718 = ~n53457 ;
  assign y15719 = n53458 ;
  assign y15720 = ~n53461 ;
  assign y15721 = n53465 ;
  assign y15722 = ~n53467 ;
  assign y15723 = n53469 ;
  assign y15724 = ~n53472 ;
  assign y15725 = ~n53473 ;
  assign y15726 = ~n53476 ;
  assign y15727 = ~1'b0 ;
  assign y15728 = ~1'b0 ;
  assign y15729 = ~n53478 ;
  assign y15730 = ~n53480 ;
  assign y15731 = ~n53481 ;
  assign y15732 = ~n53483 ;
  assign y15733 = n53484 ;
  assign y15734 = ~n53486 ;
  assign y15735 = n53492 ;
  assign y15736 = n53495 ;
  assign y15737 = ~n53496 ;
  assign y15738 = ~1'b0 ;
  assign y15739 = ~n53497 ;
  assign y15740 = n53498 ;
  assign y15741 = ~n53499 ;
  assign y15742 = n53502 ;
  assign y15743 = ~n53504 ;
  assign y15744 = n53505 ;
  assign y15745 = n53506 ;
  assign y15746 = n53507 ;
  assign y15747 = n53509 ;
  assign y15748 = n53511 ;
  assign y15749 = n53513 ;
  assign y15750 = ~n53514 ;
  assign y15751 = ~n53517 ;
  assign y15752 = ~n53521 ;
  assign y15753 = ~n53522 ;
  assign y15754 = n53523 ;
  assign y15755 = ~n53525 ;
  assign y15756 = n53527 ;
  assign y15757 = ~n53529 ;
  assign y15758 = ~1'b0 ;
  assign y15759 = n53531 ;
  assign y15760 = ~1'b0 ;
  assign y15761 = ~n53533 ;
  assign y15762 = n53534 ;
  assign y15763 = n53535 ;
  assign y15764 = n53540 ;
  assign y15765 = ~n53541 ;
  assign y15766 = ~n53542 ;
  assign y15767 = ~n53543 ;
  assign y15768 = ~n53548 ;
  assign y15769 = n53550 ;
  assign y15770 = ~1'b0 ;
  assign y15771 = ~1'b0 ;
  assign y15772 = n53551 ;
  assign y15773 = n53552 ;
  assign y15774 = n53553 ;
  assign y15775 = ~n53555 ;
  assign y15776 = n53559 ;
  assign y15777 = ~n53560 ;
  assign y15778 = ~n53564 ;
  assign y15779 = ~n53567 ;
  assign y15780 = ~n53570 ;
  assign y15781 = n53572 ;
  assign y15782 = ~1'b0 ;
  assign y15783 = ~n53573 ;
  assign y15784 = n53574 ;
  assign y15785 = n53584 ;
  assign y15786 = n53585 ;
  assign y15787 = ~n53586 ;
  assign y15788 = ~n53588 ;
  assign y15789 = ~n53589 ;
  assign y15790 = ~n53593 ;
  assign y15791 = ~1'b0 ;
  assign y15792 = ~n53595 ;
  assign y15793 = ~n53596 ;
  assign y15794 = ~n53599 ;
  assign y15795 = ~n53600 ;
  assign y15796 = ~n53601 ;
  assign y15797 = n53602 ;
  assign y15798 = n53603 ;
  assign y15799 = n53609 ;
  assign y15800 = n53613 ;
  assign y15801 = ~1'b0 ;
  assign y15802 = ~1'b0 ;
  assign y15803 = n53615 ;
  assign y15804 = n53624 ;
  assign y15805 = ~n53625 ;
  assign y15806 = ~n53626 ;
  assign y15807 = n53634 ;
  assign y15808 = ~n53637 ;
  assign y15809 = n53641 ;
  assign y15810 = n53645 ;
  assign y15811 = ~n53647 ;
  assign y15812 = ~1'b0 ;
  assign y15813 = ~n53648 ;
  assign y15814 = ~n53650 ;
  assign y15815 = n53651 ;
  assign y15816 = n53652 ;
  assign y15817 = n53654 ;
  assign y15818 = n53657 ;
  assign y15819 = ~n53658 ;
  assign y15820 = n53663 ;
  assign y15821 = ~n53664 ;
  assign y15822 = ~1'b0 ;
  assign y15823 = ~n53665 ;
  assign y15824 = n53667 ;
  assign y15825 = n53668 ;
  assign y15826 = n53669 ;
  assign y15827 = ~n53671 ;
  assign y15828 = ~n53672 ;
  assign y15829 = ~n53674 ;
  assign y15830 = n53676 ;
  assign y15831 = n53677 ;
  assign y15832 = n53681 ;
  assign y15833 = n53685 ;
  assign y15834 = ~n53689 ;
  assign y15835 = n53694 ;
  assign y15836 = n53701 ;
  assign y15837 = n53704 ;
  assign y15838 = n53707 ;
  assign y15839 = n53709 ;
  assign y15840 = n53712 ;
  assign y15841 = n53714 ;
  assign y15842 = ~n53718 ;
  assign y15843 = ~n53721 ;
  assign y15844 = ~n53722 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = ~1'b0 ;
  assign y15847 = ~n53723 ;
  assign y15848 = n53724 ;
  assign y15849 = n53725 ;
  assign y15850 = n53727 ;
  assign y15851 = n53729 ;
  assign y15852 = ~n53730 ;
  assign y15853 = n53733 ;
  assign y15854 = ~n53734 ;
  assign y15855 = n53737 ;
  assign y15856 = ~n53739 ;
  assign y15857 = n53740 ;
  assign y15858 = n53743 ;
  assign y15859 = ~n53744 ;
  assign y15860 = ~n53745 ;
  assign y15861 = ~n53746 ;
  assign y15862 = n53748 ;
  assign y15863 = ~n53749 ;
  assign y15864 = n53750 ;
  assign y15865 = n53751 ;
  assign y15866 = ~n53754 ;
  assign y15867 = ~n53757 ;
  assign y15868 = ~n53758 ;
  assign y15869 = n53759 ;
  assign y15870 = ~n53761 ;
  assign y15871 = n53762 ;
  assign y15872 = ~n53766 ;
  assign y15873 = ~n53767 ;
  assign y15874 = n53770 ;
  assign y15875 = ~1'b0 ;
  assign y15876 = n53775 ;
  assign y15877 = ~1'b0 ;
  assign y15878 = n53776 ;
  assign y15879 = ~n53779 ;
  assign y15880 = n53782 ;
  assign y15881 = ~n53783 ;
  assign y15882 = n53785 ;
  assign y15883 = n53788 ;
  assign y15884 = n53790 ;
  assign y15885 = ~n53791 ;
  assign y15886 = ~1'b0 ;
  assign y15887 = ~n53795 ;
  assign y15888 = ~n53797 ;
  assign y15889 = n53801 ;
  assign y15890 = ~n53802 ;
  assign y15891 = n53803 ;
  assign y15892 = ~n53804 ;
  assign y15893 = ~n53805 ;
  assign y15894 = n53808 ;
  assign y15895 = ~n53810 ;
  assign y15896 = ~1'b0 ;
  assign y15897 = n53815 ;
  assign y15898 = n53816 ;
  assign y15899 = ~n53817 ;
  assign y15900 = n53818 ;
  assign y15901 = ~n53819 ;
  assign y15902 = n53821 ;
  assign y15903 = ~n53822 ;
  assign y15904 = ~n53823 ;
  assign y15905 = ~n53824 ;
  assign y15906 = ~n53826 ;
  assign y15907 = ~1'b0 ;
  assign y15908 = ~1'b0 ;
  assign y15909 = ~n53827 ;
  assign y15910 = n53828 ;
  assign y15911 = ~n53829 ;
  assign y15912 = ~n53830 ;
  assign y15913 = n53831 ;
  assign y15914 = n53834 ;
  assign y15915 = ~n53838 ;
  assign y15916 = n53839 ;
  assign y15917 = ~n53840 ;
  assign y15918 = n53842 ;
  assign y15919 = ~n53847 ;
  assign y15920 = ~n53855 ;
  assign y15921 = ~n53857 ;
  assign y15922 = ~n53858 ;
  assign y15923 = n53861 ;
  assign y15924 = ~n53862 ;
  assign y15925 = ~n53863 ;
  assign y15926 = ~n53864 ;
  assign y15927 = ~n53865 ;
  assign y15928 = n53867 ;
  assign y15929 = ~n53869 ;
  assign y15930 = ~1'b0 ;
  assign y15931 = n53872 ;
  assign y15932 = ~n53873 ;
  assign y15933 = ~n53874 ;
  assign y15934 = n53879 ;
  assign y15935 = ~n53880 ;
  assign y15936 = ~n53881 ;
  assign y15937 = n53882 ;
  assign y15938 = ~n53885 ;
  assign y15939 = ~n53887 ;
  assign y15940 = ~1'b0 ;
  assign y15941 = ~1'b0 ;
  assign y15942 = ~n53890 ;
  assign y15943 = ~n53892 ;
  assign y15944 = ~n53893 ;
  assign y15945 = ~n53894 ;
  assign y15946 = n53895 ;
  assign y15947 = ~n53900 ;
  assign y15948 = n53903 ;
  assign y15949 = ~n53906 ;
  assign y15950 = ~n53907 ;
  assign y15951 = n53915 ;
  assign y15952 = ~n53919 ;
  assign y15953 = n53921 ;
  assign y15954 = n53922 ;
  assign y15955 = ~n53923 ;
  assign y15956 = ~n53924 ;
  assign y15957 = ~n53927 ;
  assign y15958 = n53929 ;
  assign y15959 = n53934 ;
  assign y15960 = ~n53936 ;
  assign y15961 = n53937 ;
  assign y15962 = ~n53938 ;
  assign y15963 = n53939 ;
  assign y15964 = n53940 ;
  assign y15965 = n53941 ;
  assign y15966 = ~n53945 ;
  assign y15967 = n53947 ;
  assign y15968 = n53948 ;
  assign y15969 = n53953 ;
  assign y15970 = ~n53954 ;
  assign y15971 = ~1'b0 ;
  assign y15972 = ~1'b0 ;
  assign y15973 = n53955 ;
  assign y15974 = ~n53956 ;
  assign y15975 = n53957 ;
  assign y15976 = n53960 ;
  assign y15977 = ~n53962 ;
  assign y15978 = ~n53963 ;
  assign y15979 = ~n53964 ;
  assign y15980 = n53969 ;
  assign y15981 = n53977 ;
  assign y15982 = ~1'b0 ;
  assign y15983 = ~1'b0 ;
  assign y15984 = n53979 ;
  assign y15985 = ~n53980 ;
  assign y15986 = ~n53982 ;
  assign y15987 = n53987 ;
  assign y15988 = n53988 ;
  assign y15989 = n53990 ;
  assign y15990 = n53991 ;
  assign y15991 = ~n53992 ;
  assign y15992 = ~n53994 ;
  assign y15993 = ~1'b0 ;
  assign y15994 = n53995 ;
  assign y15995 = n53999 ;
  assign y15996 = ~n54001 ;
  assign y15997 = ~n54002 ;
  assign y15998 = ~n54003 ;
  assign y15999 = ~n54007 ;
  assign y16000 = ~n54010 ;
  assign y16001 = ~n54011 ;
  assign y16002 = ~n54013 ;
  assign y16003 = n54015 ;
  assign y16004 = ~1'b0 ;
  assign y16005 = n54017 ;
  assign y16006 = n54018 ;
  assign y16007 = n54021 ;
  assign y16008 = ~n54023 ;
  assign y16009 = ~n54026 ;
  assign y16010 = n54032 ;
  assign y16011 = ~n54036 ;
  assign y16012 = ~n54037 ;
  assign y16013 = ~n54040 ;
  assign y16014 = ~n54042 ;
  assign y16015 = ~n54044 ;
  assign y16016 = n54046 ;
  assign y16017 = n54048 ;
  assign y16018 = ~n54051 ;
  assign y16019 = ~n54052 ;
  assign y16020 = n54055 ;
  assign y16021 = n54057 ;
  assign y16022 = ~n54062 ;
  assign y16023 = ~n54063 ;
  assign y16024 = n54064 ;
  assign y16025 = n54065 ;
  assign y16026 = ~n54068 ;
  assign y16027 = ~n54070 ;
  assign y16028 = ~n49131 ;
  assign y16029 = ~n54072 ;
  assign y16030 = ~n54076 ;
  assign y16031 = ~n54081 ;
  assign y16032 = n54082 ;
  assign y16033 = ~n54086 ;
  assign y16034 = n54088 ;
  assign y16035 = n54089 ;
  assign y16036 = n54092 ;
  assign y16037 = n54095 ;
  assign y16038 = n54097 ;
  assign y16039 = ~n54099 ;
  assign y16040 = ~n54101 ;
  assign y16041 = n54102 ;
  assign y16042 = n54103 ;
  assign y16043 = n54104 ;
  assign y16044 = n54107 ;
  assign y16045 = n42078 ;
  assign y16046 = ~n54111 ;
  assign y16047 = ~1'b0 ;
  assign y16048 = ~n54117 ;
  assign y16049 = ~n54121 ;
  assign y16050 = ~n54122 ;
  assign y16051 = ~n54123 ;
  assign y16052 = n54124 ;
  assign y16053 = n54129 ;
  assign y16054 = ~n54132 ;
  assign y16055 = n54135 ;
  assign y16056 = n54138 ;
  assign y16057 = n54140 ;
  assign y16058 = ~n54143 ;
  assign y16059 = n54146 ;
  assign y16060 = ~n54151 ;
  assign y16061 = n54159 ;
  assign y16062 = n54165 ;
  assign y16063 = n54166 ;
  assign y16064 = n54171 ;
  assign y16065 = ~n54172 ;
  assign y16066 = ~n38875 ;
  assign y16067 = ~n54173 ;
  assign y16068 = ~n54175 ;
  assign y16069 = n54180 ;
  assign y16070 = n54182 ;
  assign y16071 = ~n54183 ;
  assign y16072 = ~n54188 ;
  assign y16073 = n54189 ;
  assign y16074 = ~n54190 ;
  assign y16075 = ~n54191 ;
  assign y16076 = n54192 ;
  assign y16077 = n54193 ;
  assign y16078 = n54197 ;
  assign y16079 = ~1'b0 ;
  assign y16080 = ~n54198 ;
  assign y16081 = n54200 ;
  assign y16082 = ~n54201 ;
  assign y16083 = n54202 ;
  assign y16084 = n54203 ;
  assign y16085 = n54206 ;
  assign y16086 = ~n54208 ;
  assign y16087 = ~n54209 ;
  assign y16088 = n54216 ;
  assign y16089 = n54218 ;
  assign y16090 = n54220 ;
  assign y16091 = ~1'b0 ;
  assign y16092 = ~n54221 ;
  assign y16093 = n54223 ;
  assign y16094 = n54224 ;
  assign y16095 = ~n54226 ;
  assign y16096 = ~n54230 ;
  assign y16097 = n54231 ;
  assign y16098 = n54232 ;
  assign y16099 = n54233 ;
  assign y16100 = n54235 ;
  assign y16101 = n54239 ;
  assign y16102 = n54241 ;
  assign y16103 = n54242 ;
  assign y16104 = ~n54243 ;
  assign y16105 = n20715 ;
  assign y16106 = ~n54245 ;
  assign y16107 = n54246 ;
  assign y16108 = ~n54248 ;
  assign y16109 = ~n54250 ;
  assign y16110 = n54253 ;
  assign y16111 = ~n54254 ;
  assign y16112 = ~1'b0 ;
  assign y16113 = ~n54255 ;
  assign y16114 = n54256 ;
  assign y16115 = ~n54257 ;
  assign y16116 = ~n54258 ;
  assign y16117 = ~n54259 ;
  assign y16118 = ~n54263 ;
  assign y16119 = ~n54265 ;
  assign y16120 = n54267 ;
  assign y16121 = ~n54268 ;
  assign y16122 = ~n54272 ;
  assign y16123 = ~n54273 ;
  assign y16124 = ~n54276 ;
  assign y16125 = n54284 ;
  assign y16126 = ~n54285 ;
  assign y16127 = n54295 ;
  assign y16128 = n54298 ;
  assign y16129 = ~n54300 ;
  assign y16130 = ~1'b0 ;
  assign y16131 = n54303 ;
  assign y16132 = n54306 ;
  assign y16133 = n54308 ;
  assign y16134 = n54310 ;
  assign y16135 = ~n54311 ;
  assign y16136 = ~n54312 ;
  assign y16137 = n54314 ;
  assign y16138 = n54318 ;
  assign y16139 = n54321 ;
  assign y16140 = n54323 ;
  assign y16141 = ~1'b0 ;
  assign y16142 = ~n54329 ;
  assign y16143 = n54331 ;
  assign y16144 = ~n54333 ;
  assign y16145 = n54334 ;
  assign y16146 = n54335 ;
  assign y16147 = ~n54336 ;
  assign y16148 = ~n54338 ;
  assign y16149 = ~n54341 ;
  assign y16150 = ~1'b0 ;
  assign y16151 = ~n54343 ;
  assign y16152 = ~n54349 ;
  assign y16153 = ~n54350 ;
  assign y16154 = ~n54354 ;
  assign y16155 = ~n54355 ;
  assign y16156 = n54357 ;
  assign y16157 = ~n54360 ;
  assign y16158 = ~n54362 ;
  assign y16159 = ~n54363 ;
  assign y16160 = ~n54367 ;
  assign y16161 = ~1'b0 ;
  assign y16162 = ~n54370 ;
  assign y16163 = ~n54373 ;
  assign y16164 = ~n54375 ;
  assign y16165 = ~n54376 ;
  assign y16166 = ~n54379 ;
  assign y16167 = n54388 ;
  assign y16168 = n54393 ;
  assign y16169 = n54394 ;
  assign y16170 = ~n54400 ;
  assign y16171 = ~1'b0 ;
  assign y16172 = ~1'b0 ;
  assign y16173 = ~n54403 ;
  assign y16174 = n54404 ;
  assign y16175 = n54408 ;
  assign y16176 = n54412 ;
  assign y16177 = n54413 ;
  assign y16178 = n54414 ;
  assign y16179 = ~n54416 ;
  assign y16180 = n54423 ;
  assign y16181 = ~n54425 ;
  assign y16182 = ~n54427 ;
  assign y16183 = ~1'b0 ;
  assign y16184 = ~n54430 ;
  assign y16185 = n54431 ;
  assign y16186 = ~n54433 ;
  assign y16187 = ~n54442 ;
  assign y16188 = ~n54443 ;
  assign y16189 = ~n54444 ;
  assign y16190 = ~n54445 ;
  assign y16191 = n54446 ;
  assign y16192 = n54451 ;
  assign y16193 = ~1'b0 ;
  assign y16194 = n54456 ;
  assign y16195 = ~n54458 ;
  assign y16196 = n54461 ;
  assign y16197 = ~n54463 ;
  assign y16198 = ~n54466 ;
  assign y16199 = ~n54467 ;
  assign y16200 = n54470 ;
  assign y16201 = ~n54471 ;
  assign y16202 = n54473 ;
  assign y16203 = ~n54474 ;
  assign y16204 = n54477 ;
  assign y16205 = n54479 ;
  assign y16206 = ~1'b0 ;
  assign y16207 = n54481 ;
  assign y16208 = ~n54482 ;
  assign y16209 = n54486 ;
  assign y16210 = n54488 ;
  assign y16211 = ~n54491 ;
  assign y16212 = ~n54495 ;
  assign y16213 = ~n54496 ;
  assign y16214 = ~n54498 ;
  assign y16215 = ~n54500 ;
  assign y16216 = ~n54502 ;
  assign y16217 = n54507 ;
  assign y16218 = n54510 ;
  assign y16219 = n54513 ;
  assign y16220 = n54515 ;
  assign y16221 = ~n54517 ;
  assign y16222 = n54518 ;
  assign y16223 = n54519 ;
  assign y16224 = ~n54520 ;
  assign y16225 = n54521 ;
  assign y16226 = n54523 ;
  assign y16227 = ~n54525 ;
  assign y16228 = n54527 ;
  assign y16229 = ~n54529 ;
  assign y16230 = ~n54531 ;
  assign y16231 = n54532 ;
  assign y16232 = n54536 ;
  assign y16233 = n54540 ;
  assign y16234 = ~n54541 ;
  assign y16235 = ~n54542 ;
  assign y16236 = n54543 ;
  assign y16237 = ~1'b0 ;
  assign y16238 = ~n54546 ;
  assign y16239 = ~1'b0 ;
  assign y16240 = ~n54551 ;
  assign y16241 = ~n54552 ;
  assign y16242 = ~n54554 ;
  assign y16243 = ~n54555 ;
  assign y16244 = ~n54557 ;
  assign y16245 = n54558 ;
  assign y16246 = n54559 ;
  assign y16247 = ~n54561 ;
  assign y16248 = ~1'b0 ;
  assign y16249 = ~n54564 ;
  assign y16250 = n54566 ;
  assign y16251 = ~n54574 ;
  assign y16252 = ~n54579 ;
  assign y16253 = n54581 ;
  assign y16254 = n54587 ;
  assign y16255 = ~n54591 ;
  assign y16256 = n54593 ;
  assign y16257 = n54594 ;
  assign y16258 = n54595 ;
  assign y16259 = ~1'b0 ;
  assign y16260 = ~1'b0 ;
  assign y16261 = n54599 ;
  assign y16262 = ~n54601 ;
  assign y16263 = ~n54604 ;
  assign y16264 = ~n54606 ;
  assign y16265 = ~n54608 ;
  assign y16266 = ~n54611 ;
  assign y16267 = ~n54612 ;
  assign y16268 = n54613 ;
  assign y16269 = n54620 ;
  assign y16270 = ~n54622 ;
  assign y16271 = n54626 ;
  assign y16272 = ~n54627 ;
  assign y16273 = n54628 ;
  assign y16274 = n54629 ;
  assign y16275 = n54631 ;
  assign y16276 = ~n54636 ;
  assign y16277 = ~n54637 ;
  assign y16278 = n54640 ;
  assign y16279 = ~n54641 ;
  assign y16280 = ~n54645 ;
  assign y16281 = n54648 ;
  assign y16282 = ~1'b0 ;
  assign y16283 = n54650 ;
  assign y16284 = ~n54652 ;
  assign y16285 = ~n54654 ;
  assign y16286 = n54658 ;
  assign y16287 = ~n2815 ;
  assign y16288 = ~n54659 ;
  assign y16289 = ~n54660 ;
  assign y16290 = ~1'b0 ;
  assign y16291 = n1361 ;
  assign y16292 = ~n54662 ;
  assign y16293 = ~1'b0 ;
  assign y16294 = n54665 ;
  assign y16295 = ~n54666 ;
  assign y16296 = n54667 ;
  assign y16297 = n54668 ;
  assign y16298 = n54669 ;
  assign y16299 = n54670 ;
  assign y16300 = ~n54671 ;
  assign y16301 = ~n54674 ;
  assign y16302 = n54675 ;
  assign y16303 = n54680 ;
  assign y16304 = ~1'b0 ;
  assign y16305 = n54682 ;
  assign y16306 = n54684 ;
  assign y16307 = n54686 ;
  assign y16308 = n54687 ;
  assign y16309 = n54695 ;
  assign y16310 = ~n54698 ;
  assign y16311 = ~n54700 ;
  assign y16312 = ~n54701 ;
  assign y16313 = n54703 ;
  assign y16314 = n54706 ;
  assign y16315 = n54710 ;
  assign y16316 = n54713 ;
  assign y16317 = ~n54716 ;
  assign y16318 = ~n54717 ;
  assign y16319 = n54718 ;
  assign y16320 = ~n54722 ;
  assign y16321 = ~n54724 ;
  assign y16322 = ~n54725 ;
  assign y16323 = n54727 ;
  assign y16324 = n54729 ;
  assign y16325 = ~1'b0 ;
  assign y16326 = ~n54730 ;
  assign y16327 = ~n54731 ;
  assign y16328 = n54732 ;
  assign y16329 = ~n54733 ;
  assign y16330 = n54734 ;
  assign y16331 = n54735 ;
  assign y16332 = ~n54739 ;
  assign y16333 = ~n54740 ;
  assign y16334 = n54744 ;
  assign y16335 = ~1'b0 ;
  assign y16336 = ~n54747 ;
  assign y16337 = ~n54753 ;
  assign y16338 = ~n54754 ;
  assign y16339 = ~n54755 ;
  assign y16340 = n54757 ;
  assign y16341 = n54758 ;
  assign y16342 = ~n54759 ;
  assign y16343 = ~n54762 ;
  assign y16344 = ~n54763 ;
  assign y16345 = ~1'b0 ;
  assign y16346 = ~1'b0 ;
  assign y16347 = ~n54767 ;
  assign y16348 = n54773 ;
  assign y16349 = n54774 ;
  assign y16350 = ~n54777 ;
  assign y16351 = ~n54778 ;
  assign y16352 = ~n54779 ;
  assign y16353 = n54783 ;
  assign y16354 = ~n54786 ;
  assign y16355 = n54787 ;
  assign y16356 = ~n54791 ;
  assign y16357 = n54795 ;
  assign y16358 = n54798 ;
  assign y16359 = n54799 ;
  assign y16360 = n54800 ;
  assign y16361 = ~n54801 ;
  assign y16362 = n54803 ;
  assign y16363 = ~n54807 ;
  assign y16364 = ~n54808 ;
  assign y16365 = n54809 ;
  assign y16366 = ~n54811 ;
  assign y16367 = ~1'b0 ;
  assign y16368 = ~1'b0 ;
  assign y16369 = n54812 ;
  assign y16370 = n54822 ;
  assign y16371 = n54823 ;
  assign y16372 = ~n54827 ;
  assign y16373 = ~n54829 ;
  assign y16374 = n54832 ;
  assign y16375 = n54833 ;
  assign y16376 = n54835 ;
  assign y16377 = ~n54838 ;
  assign y16378 = n54841 ;
  assign y16379 = n54849 ;
  assign y16380 = n54850 ;
  assign y16381 = ~n54851 ;
  assign y16382 = n54852 ;
  assign y16383 = n54855 ;
  assign y16384 = ~n54856 ;
  assign y16385 = n54857 ;
  assign y16386 = n54860 ;
  assign y16387 = n54865 ;
  assign y16388 = ~1'b0 ;
  assign y16389 = n54867 ;
  assign y16390 = ~n54869 ;
  assign y16391 = ~n54870 ;
  assign y16392 = ~n54872 ;
  assign y16393 = n54876 ;
  assign y16394 = ~n54879 ;
  assign y16395 = ~n54880 ;
  assign y16396 = ~n54883 ;
  assign y16397 = n54884 ;
  assign y16398 = ~n54888 ;
  assign y16399 = n54890 ;
  assign y16400 = n54893 ;
  assign y16401 = n54895 ;
  assign y16402 = ~n54896 ;
  assign y16403 = ~n54897 ;
  assign y16404 = ~n54898 ;
  assign y16405 = n54900 ;
  assign y16406 = n54902 ;
  assign y16407 = ~n54903 ;
  assign y16408 = ~n54906 ;
  assign y16409 = ~1'b0 ;
  assign y16410 = ~1'b0 ;
  assign y16411 = n54907 ;
  assign y16412 = ~n54908 ;
  assign y16413 = n54909 ;
  assign y16414 = n54912 ;
  assign y16415 = n54914 ;
  assign y16416 = n54915 ;
  assign y16417 = ~n54916 ;
  assign y16418 = n54918 ;
  assign y16419 = ~1'b0 ;
  assign y16420 = ~1'b0 ;
  assign y16421 = ~n54923 ;
  assign y16422 = ~n54925 ;
  assign y16423 = ~n54928 ;
  assign y16424 = ~n54929 ;
  assign y16425 = ~n54932 ;
  assign y16426 = n54940 ;
  assign y16427 = ~n54943 ;
  assign y16428 = ~n54945 ;
  assign y16429 = ~1'b0 ;
  assign y16430 = ~n54949 ;
  assign y16431 = n54951 ;
  assign y16432 = ~n54957 ;
  assign y16433 = ~n54961 ;
  assign y16434 = n54962 ;
  assign y16435 = n54966 ;
  assign y16436 = n54967 ;
  assign y16437 = n54968 ;
  assign y16438 = n54972 ;
  assign y16439 = ~n54974 ;
  assign y16440 = ~1'b0 ;
  assign y16441 = ~1'b0 ;
  assign y16442 = n54976 ;
  assign y16443 = ~n54977 ;
  assign y16444 = ~n54978 ;
  assign y16445 = n54981 ;
  assign y16446 = n54983 ;
  assign y16447 = ~n54984 ;
  assign y16448 = n54985 ;
  assign y16449 = ~n54987 ;
  assign y16450 = ~n54990 ;
  assign y16451 = ~1'b0 ;
  assign y16452 = ~1'b0 ;
  assign y16453 = n54992 ;
  assign y16454 = ~n54995 ;
  assign y16455 = n54996 ;
  assign y16456 = n54997 ;
  assign y16457 = ~n54998 ;
  assign y16458 = n55000 ;
  assign y16459 = n55001 ;
  assign y16460 = n55002 ;
  assign y16461 = n55003 ;
  assign y16462 = ~n55008 ;
  assign y16463 = ~1'b0 ;
  assign y16464 = ~1'b0 ;
  assign y16465 = ~n55013 ;
  assign y16466 = n55016 ;
  assign y16467 = ~n55017 ;
  assign y16468 = ~n55019 ;
  assign y16469 = n55022 ;
  assign y16470 = ~n55026 ;
  assign y16471 = ~n55028 ;
  assign y16472 = n55036 ;
  assign y16473 = n55047 ;
  assign y16474 = ~n55050 ;
  assign y16475 = ~n55051 ;
  assign y16476 = ~n55053 ;
  assign y16477 = n55057 ;
  assign y16478 = n55064 ;
  assign y16479 = ~n55066 ;
  assign y16480 = ~n55067 ;
  assign y16481 = ~n55071 ;
  assign y16482 = ~n55075 ;
  assign y16483 = ~n55077 ;
  assign y16484 = n55081 ;
  assign y16485 = ~1'b0 ;
  assign y16486 = ~1'b0 ;
  assign y16487 = ~n55082 ;
  assign y16488 = ~n55086 ;
  assign y16489 = ~n55088 ;
  assign y16490 = ~n55092 ;
  assign y16491 = n55093 ;
  assign y16492 = n55094 ;
  assign y16493 = n55095 ;
  assign y16494 = n55100 ;
  assign y16495 = ~n55103 ;
  assign y16496 = n55105 ;
  assign y16497 = ~1'b0 ;
  assign y16498 = n55106 ;
  assign y16499 = n55107 ;
  assign y16500 = ~n55108 ;
  assign y16501 = n55109 ;
  assign y16502 = n55110 ;
  assign y16503 = n55114 ;
  assign y16504 = n55115 ;
  assign y16505 = n55116 ;
  assign y16506 = n55118 ;
  assign y16507 = n55123 ;
  assign y16508 = n55125 ;
  assign y16509 = ~n55129 ;
  assign y16510 = ~n55130 ;
  assign y16511 = ~n55131 ;
  assign y16512 = n55132 ;
  assign y16513 = n55133 ;
  assign y16514 = ~n55137 ;
  assign y16515 = n55139 ;
  assign y16516 = ~n55140 ;
  assign y16517 = ~1'b0 ;
  assign y16518 = n55142 ;
  assign y16519 = n55144 ;
  assign y16520 = ~n55146 ;
  assign y16521 = n55148 ;
  assign y16522 = ~n55149 ;
  assign y16523 = ~n55152 ;
  assign y16524 = ~n55161 ;
  assign y16525 = n55162 ;
  assign y16526 = ~n55163 ;
  assign y16527 = ~n55164 ;
  assign y16528 = n55166 ;
  assign y16529 = ~n55169 ;
  assign y16530 = ~n55173 ;
  assign y16531 = n55175 ;
  assign y16532 = n55180 ;
  assign y16533 = ~n55182 ;
  assign y16534 = ~n55185 ;
  assign y16535 = n55187 ;
  assign y16536 = ~n55190 ;
  assign y16537 = ~n55195 ;
  assign y16538 = ~n55196 ;
  assign y16539 = ~n55199 ;
  assign y16540 = n55201 ;
  assign y16541 = n55204 ;
  assign y16542 = n55206 ;
  assign y16543 = n55207 ;
  assign y16544 = ~n55208 ;
  assign y16545 = ~n55211 ;
  assign y16546 = n55214 ;
  assign y16547 = ~n55215 ;
  assign y16548 = ~n55220 ;
  assign y16549 = n55225 ;
  assign y16550 = ~1'b0 ;
  assign y16551 = n55227 ;
  assign y16552 = n55229 ;
  assign y16553 = n55232 ;
  assign y16554 = n55234 ;
  assign y16555 = ~n55235 ;
  assign y16556 = ~n55236 ;
  assign y16557 = n55237 ;
  assign y16558 = ~n55239 ;
  assign y16559 = ~n55242 ;
  assign y16560 = ~n55244 ;
  assign y16561 = n55245 ;
  assign y16562 = ~1'b0 ;
  assign y16563 = ~n55246 ;
  assign y16564 = n55248 ;
  assign y16565 = n55253 ;
  assign y16566 = n55255 ;
  assign y16567 = n55256 ;
  assign y16568 = n55257 ;
  assign y16569 = n55260 ;
  assign y16570 = ~n55264 ;
  assign y16571 = ~n55270 ;
  assign y16572 = n55272 ;
  assign y16573 = ~n55274 ;
  assign y16574 = ~n55276 ;
  assign y16575 = ~n55279 ;
  assign y16576 = n55283 ;
  assign y16577 = n55285 ;
  assign y16578 = ~n55286 ;
  assign y16579 = n55287 ;
  assign y16580 = n55288 ;
  assign y16581 = n55289 ;
  assign y16582 = ~n55290 ;
  assign y16583 = ~1'b0 ;
  assign y16584 = ~n55292 ;
  assign y16585 = n55294 ;
  assign y16586 = ~n55296 ;
  assign y16587 = ~n55299 ;
  assign y16588 = n55300 ;
  assign y16589 = ~n55307 ;
  assign y16590 = n55308 ;
  assign y16591 = ~n55314 ;
  assign y16592 = ~n55316 ;
  assign y16593 = n55319 ;
  assign y16594 = ~n55323 ;
  assign y16595 = ~n55326 ;
  assign y16596 = ~n55327 ;
  assign y16597 = ~n55331 ;
  assign y16598 = n55335 ;
  assign y16599 = ~n55341 ;
  assign y16600 = n55343 ;
  assign y16601 = n55344 ;
  assign y16602 = n55345 ;
  assign y16603 = ~n55346 ;
  assign y16604 = n55348 ;
  assign y16605 = ~n55350 ;
  assign y16606 = ~n55354 ;
  assign y16607 = n55356 ;
  assign y16608 = ~n55362 ;
  assign y16609 = n55363 ;
  assign y16610 = n55364 ;
  assign y16611 = n55367 ;
  assign y16612 = ~n55368 ;
  assign y16613 = ~n55369 ;
  assign y16614 = ~n55370 ;
  assign y16615 = ~n55372 ;
  assign y16616 = n55375 ;
  assign y16617 = ~n55377 ;
  assign y16618 = ~n55380 ;
  assign y16619 = n55381 ;
  assign y16620 = ~n55383 ;
  assign y16621 = ~n55384 ;
  assign y16622 = ~n55386 ;
  assign y16623 = ~n55387 ;
  assign y16624 = ~1'b0 ;
  assign y16625 = ~n55389 ;
  assign y16626 = n55393 ;
  assign y16627 = n55395 ;
  assign y16628 = ~1'b0 ;
  assign y16629 = ~1'b0 ;
  assign y16630 = ~n55398 ;
  assign y16631 = n55399 ;
  assign y16632 = ~n55401 ;
  assign y16633 = ~n55407 ;
  assign y16634 = ~n55408 ;
  assign y16635 = ~n55409 ;
  assign y16636 = n55412 ;
  assign y16637 = ~n55413 ;
  assign y16638 = n55415 ;
  assign y16639 = ~1'b0 ;
  assign y16640 = ~1'b0 ;
  assign y16641 = ~n55417 ;
  assign y16642 = ~n55418 ;
  assign y16643 = ~n55423 ;
  assign y16644 = ~n55426 ;
  assign y16645 = n55428 ;
  assign y16646 = n55431 ;
  assign y16647 = n55433 ;
  assign y16648 = ~n55434 ;
  assign y16649 = ~1'b0 ;
  assign y16650 = n55438 ;
  assign y16651 = n55440 ;
  assign y16652 = ~n55441 ;
  assign y16653 = n55444 ;
  assign y16654 = n55446 ;
  assign y16655 = n49277 ;
  assign y16656 = ~n55448 ;
  assign y16657 = n55452 ;
  assign y16658 = ~n55455 ;
  assign y16659 = ~n55457 ;
  assign y16660 = ~n55459 ;
  assign y16661 = ~1'b0 ;
  assign y16662 = n55461 ;
  assign y16663 = ~n55467 ;
  assign y16664 = n55468 ;
  assign y16665 = ~n55472 ;
  assign y16666 = n55474 ;
  assign y16667 = n55475 ;
  assign y16668 = ~n55479 ;
  assign y16669 = n55482 ;
  assign y16670 = ~n55487 ;
  assign y16671 = ~1'b0 ;
  assign y16672 = ~n55491 ;
  assign y16673 = ~n55495 ;
  assign y16674 = ~n55496 ;
  assign y16675 = n55497 ;
  assign y16676 = n55498 ;
  assign y16677 = n55499 ;
  assign y16678 = n55500 ;
  assign y16679 = n55501 ;
  assign y16680 = n55503 ;
  assign y16681 = ~n55505 ;
  assign y16682 = ~n55509 ;
  assign y16683 = n55511 ;
  assign y16684 = n55513 ;
  assign y16685 = n55514 ;
  assign y16686 = n55522 ;
  assign y16687 = ~n55526 ;
  assign y16688 = n55527 ;
  assign y16689 = ~n55532 ;
  assign y16690 = n55535 ;
  assign y16691 = n55537 ;
  assign y16692 = n55538 ;
  assign y16693 = ~1'b0 ;
  assign y16694 = ~n55545 ;
  assign y16695 = ~1'b0 ;
  assign y16696 = ~n55546 ;
  assign y16697 = n55549 ;
  assign y16698 = ~n55550 ;
  assign y16699 = ~n55551 ;
  assign y16700 = n55554 ;
  assign y16701 = n55555 ;
  assign y16702 = n55557 ;
  assign y16703 = ~n55558 ;
  assign y16704 = ~n55560 ;
  assign y16705 = n55562 ;
  assign y16706 = n55567 ;
  assign y16707 = n55568 ;
  assign y16708 = ~n55572 ;
  assign y16709 = ~n55573 ;
  assign y16710 = n55575 ;
  assign y16711 = ~n55577 ;
  assign y16712 = n55578 ;
  assign y16713 = ~n55581 ;
  assign y16714 = ~n55582 ;
  assign y16715 = n55585 ;
  assign y16716 = n55589 ;
  assign y16717 = ~n55591 ;
  assign y16718 = ~n55592 ;
  assign y16719 = ~n55599 ;
  assign y16720 = n55602 ;
  assign y16721 = ~n55605 ;
  assign y16722 = ~n55607 ;
  assign y16723 = n55608 ;
  assign y16724 = n55614 ;
  assign y16725 = n55615 ;
  assign y16726 = n55617 ;
  assign y16727 = n55619 ;
  assign y16728 = n55623 ;
  assign y16729 = ~n55624 ;
  assign y16730 = ~n55625 ;
  assign y16731 = n55627 ;
  assign y16732 = ~n55628 ;
  assign y16733 = ~n55629 ;
  assign y16734 = n55631 ;
  assign y16735 = ~n55632 ;
  assign y16736 = n55637 ;
  assign y16737 = n55638 ;
  assign y16738 = ~1'b0 ;
  assign y16739 = ~1'b0 ;
  assign y16740 = n55642 ;
  assign y16741 = ~n55643 ;
  assign y16742 = ~n55648 ;
  assign y16743 = ~n55649 ;
  assign y16744 = n55652 ;
  assign y16745 = n55653 ;
  assign y16746 = ~n55654 ;
  assign y16747 = n55655 ;
endmodule
