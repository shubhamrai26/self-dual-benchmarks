module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2088 , n2089 , n2090 , n2091 , n2092 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2114 , n2115 , n2116 ;
  assign n129 = ~x125 & x127 ;
  assign n130 = x126 & x127 ;
  assign n131 = x126 & ~n130 ;
  assign n132 = x125 & ~n131 ;
  assign n133 = ~n129 & ~n132 ;
  assign n134 = ~x123 & ~n133 ;
  assign n135 = ~x124 & ~n131 ;
  assign n136 = x124 & ~n133 ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = x123 & ~n137 ;
  assign n139 = ~n134 & ~n138 ;
  assign n140 = ~x121 & ~n139 ;
  assign n141 = ~x122 & ~n137 ;
  assign n142 = x122 & ~n139 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = x121 & ~n143 ;
  assign n145 = ~n140 & ~n144 ;
  assign n146 = ~x119 & ~n145 ;
  assign n147 = ~x120 & ~n143 ;
  assign n148 = x120 & ~n145 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = x119 & ~n149 ;
  assign n151 = ~n146 & ~n150 ;
  assign n152 = ~x117 & ~n151 ;
  assign n153 = ~x118 & ~n149 ;
  assign n154 = x118 & ~n151 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = x117 & ~n155 ;
  assign n157 = ~n152 & ~n156 ;
  assign n158 = ~x115 & ~n157 ;
  assign n159 = ~x116 & ~n155 ;
  assign n160 = x116 & ~n157 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = x115 & ~n161 ;
  assign n163 = ~n158 & ~n162 ;
  assign n164 = ~x113 & ~n163 ;
  assign n165 = ~x114 & ~n161 ;
  assign n166 = x114 & ~n163 ;
  assign n167 = ~n165 & ~n166 ;
  assign n168 = x113 & ~n167 ;
  assign n169 = ~n164 & ~n168 ;
  assign n170 = ~x111 & ~n169 ;
  assign n171 = ~x112 & ~n167 ;
  assign n172 = x112 & ~n169 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = x111 & ~n173 ;
  assign n175 = ~n170 & ~n174 ;
  assign n176 = ~x109 & ~n175 ;
  assign n177 = ~x110 & ~n173 ;
  assign n178 = x110 & ~n175 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = x109 & ~n179 ;
  assign n181 = ~n176 & ~n180 ;
  assign n182 = ~x107 & ~n181 ;
  assign n183 = ~x108 & ~n179 ;
  assign n184 = x108 & ~n181 ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = x107 & ~n185 ;
  assign n187 = ~n182 & ~n186 ;
  assign n188 = ~x105 & ~n187 ;
  assign n189 = ~x106 & ~n185 ;
  assign n190 = x106 & ~n187 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = x105 & ~n191 ;
  assign n193 = ~n188 & ~n192 ;
  assign n194 = ~x103 & ~n193 ;
  assign n195 = ~x104 & ~n191 ;
  assign n196 = x104 & ~n193 ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = x103 & ~n197 ;
  assign n199 = ~n194 & ~n198 ;
  assign n200 = ~x101 & ~n199 ;
  assign n201 = ~x102 & ~n197 ;
  assign n202 = x102 & ~n199 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = x101 & ~n203 ;
  assign n205 = ~n200 & ~n204 ;
  assign n206 = ~x99 & ~n205 ;
  assign n207 = ~x100 & ~n203 ;
  assign n208 = x100 & ~n205 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = x99 & ~n209 ;
  assign n211 = ~n206 & ~n210 ;
  assign n212 = ~x97 & ~n211 ;
  assign n213 = ~x98 & ~n209 ;
  assign n214 = x98 & ~n211 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = x97 & ~n215 ;
  assign n217 = ~n212 & ~n216 ;
  assign n218 = ~x95 & ~n217 ;
  assign n219 = ~x96 & ~n215 ;
  assign n220 = x96 & ~n217 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = x95 & ~n221 ;
  assign n223 = ~n218 & ~n222 ;
  assign n224 = ~x93 & ~n223 ;
  assign n225 = ~x94 & ~n221 ;
  assign n226 = x94 & ~n223 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = x93 & ~n227 ;
  assign n229 = ~n224 & ~n228 ;
  assign n230 = ~x91 & ~n229 ;
  assign n231 = ~x92 & ~n227 ;
  assign n232 = x92 & ~n229 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = x91 & ~n233 ;
  assign n235 = ~n230 & ~n234 ;
  assign n236 = ~x89 & ~n235 ;
  assign n237 = ~x90 & ~n233 ;
  assign n238 = x90 & ~n235 ;
  assign n239 = ~n237 & ~n238 ;
  assign n240 = x89 & ~n239 ;
  assign n241 = ~n236 & ~n240 ;
  assign n242 = ~x87 & ~n241 ;
  assign n243 = ~x88 & ~n239 ;
  assign n244 = x88 & ~n241 ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = x87 & ~n245 ;
  assign n247 = ~n242 & ~n246 ;
  assign n248 = ~x85 & ~n247 ;
  assign n249 = ~x86 & ~n245 ;
  assign n250 = x86 & ~n247 ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = x85 & ~n251 ;
  assign n253 = ~n248 & ~n252 ;
  assign n254 = ~x83 & ~n253 ;
  assign n255 = ~x84 & ~n251 ;
  assign n256 = x84 & ~n253 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = x83 & ~n257 ;
  assign n259 = ~n254 & ~n258 ;
  assign n260 = ~x81 & ~n259 ;
  assign n261 = ~x82 & ~n257 ;
  assign n262 = x82 & ~n259 ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = x81 & ~n263 ;
  assign n265 = ~n260 & ~n264 ;
  assign n266 = ~x79 & ~n265 ;
  assign n267 = ~x80 & ~n263 ;
  assign n268 = x80 & ~n265 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = x79 & ~n269 ;
  assign n271 = ~n266 & ~n270 ;
  assign n272 = ~x77 & ~n271 ;
  assign n273 = ~x78 & ~n269 ;
  assign n274 = x78 & ~n271 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = x77 & ~n275 ;
  assign n277 = ~n272 & ~n276 ;
  assign n278 = ~x75 & ~n277 ;
  assign n279 = ~x76 & ~n275 ;
  assign n280 = x76 & ~n277 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = x75 & ~n281 ;
  assign n283 = ~n278 & ~n282 ;
  assign n284 = ~x73 & ~n283 ;
  assign n285 = ~x74 & ~n281 ;
  assign n286 = x74 & ~n283 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = x73 & ~n287 ;
  assign n289 = ~n284 & ~n288 ;
  assign n290 = ~x71 & ~n289 ;
  assign n291 = ~x72 & ~n287 ;
  assign n292 = x72 & ~n289 ;
  assign n293 = ~n291 & ~n292 ;
  assign n294 = x71 & ~n293 ;
  assign n295 = ~n290 & ~n294 ;
  assign n296 = ~x69 & ~n295 ;
  assign n297 = ~x70 & ~n293 ;
  assign n298 = x70 & ~n295 ;
  assign n299 = ~n297 & ~n298 ;
  assign n300 = x69 & ~n299 ;
  assign n301 = ~n296 & ~n300 ;
  assign n302 = ~x67 & ~n301 ;
  assign n303 = ~x68 & ~n299 ;
  assign n304 = x68 & ~n301 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = x67 & ~n305 ;
  assign n307 = ~n302 & ~n306 ;
  assign n308 = ~x65 & ~n307 ;
  assign n309 = ~x66 & ~n305 ;
  assign n310 = x66 & ~n307 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = x65 & ~n311 ;
  assign n313 = ~n308 & ~n312 ;
  assign n314 = ~x63 & ~n313 ;
  assign n315 = ~x64 & ~n311 ;
  assign n316 = x64 & ~n313 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = x63 & ~n317 ;
  assign n319 = ~n314 & ~n318 ;
  assign n320 = ~x61 & ~n319 ;
  assign n321 = ~x62 & ~n317 ;
  assign n322 = x62 & ~n319 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = x61 & ~n323 ;
  assign n325 = ~n320 & ~n324 ;
  assign n326 = ~x59 & ~n325 ;
  assign n327 = ~x60 & ~n323 ;
  assign n328 = x60 & ~n325 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = x59 & ~n329 ;
  assign n331 = ~n326 & ~n330 ;
  assign n332 = ~x57 & ~n331 ;
  assign n333 = ~x58 & ~n329 ;
  assign n334 = x58 & ~n331 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = x57 & ~n335 ;
  assign n337 = ~n332 & ~n336 ;
  assign n338 = ~x55 & ~n337 ;
  assign n339 = ~x56 & ~n335 ;
  assign n340 = x56 & ~n337 ;
  assign n341 = ~n339 & ~n340 ;
  assign n342 = x55 & ~n341 ;
  assign n343 = ~n338 & ~n342 ;
  assign n344 = ~x53 & ~n343 ;
  assign n345 = ~x54 & ~n341 ;
  assign n346 = x54 & ~n343 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = x53 & ~n347 ;
  assign n349 = ~n344 & ~n348 ;
  assign n350 = ~x51 & ~n349 ;
  assign n351 = ~x52 & ~n347 ;
  assign n352 = x52 & ~n349 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = x51 & ~n353 ;
  assign n355 = ~n350 & ~n354 ;
  assign n356 = ~x49 & ~n355 ;
  assign n357 = ~x50 & ~n353 ;
  assign n358 = x50 & ~n355 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = x49 & ~n359 ;
  assign n361 = ~n356 & ~n360 ;
  assign n362 = ~x47 & ~n361 ;
  assign n363 = ~x48 & ~n359 ;
  assign n364 = x48 & ~n361 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = x47 & ~n365 ;
  assign n367 = ~n362 & ~n366 ;
  assign n368 = ~x45 & ~n367 ;
  assign n369 = ~x46 & ~n365 ;
  assign n370 = x46 & ~n367 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = x45 & ~n371 ;
  assign n373 = ~n368 & ~n372 ;
  assign n374 = ~x43 & ~n373 ;
  assign n375 = ~x44 & ~n371 ;
  assign n376 = x44 & ~n373 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = x43 & ~n377 ;
  assign n379 = ~n374 & ~n378 ;
  assign n380 = ~x41 & ~n379 ;
  assign n381 = ~x42 & ~n377 ;
  assign n382 = x42 & ~n379 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = x41 & ~n383 ;
  assign n385 = ~n380 & ~n384 ;
  assign n386 = ~x39 & ~n385 ;
  assign n387 = ~x40 & ~n383 ;
  assign n388 = x40 & ~n385 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = x39 & ~n389 ;
  assign n391 = ~n386 & ~n390 ;
  assign n392 = ~x37 & ~n391 ;
  assign n393 = ~x38 & ~n389 ;
  assign n394 = x38 & ~n391 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = x37 & ~n395 ;
  assign n397 = ~n392 & ~n396 ;
  assign n398 = ~x35 & ~n397 ;
  assign n399 = ~x36 & ~n395 ;
  assign n400 = x36 & ~n397 ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = x35 & ~n401 ;
  assign n403 = ~n398 & ~n402 ;
  assign n404 = ~x33 & ~n403 ;
  assign n405 = ~x34 & ~n401 ;
  assign n406 = x34 & ~n403 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = x33 & ~n407 ;
  assign n409 = ~n404 & ~n408 ;
  assign n410 = ~x31 & ~n409 ;
  assign n411 = ~x32 & ~n407 ;
  assign n412 = x32 & ~n409 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = x31 & ~n413 ;
  assign n415 = ~n410 & ~n414 ;
  assign n416 = ~x29 & ~n415 ;
  assign n417 = ~x30 & ~n413 ;
  assign n418 = x30 & ~n415 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = x29 & ~n419 ;
  assign n421 = ~n416 & ~n420 ;
  assign n422 = ~x27 & ~n421 ;
  assign n423 = ~x28 & ~n419 ;
  assign n424 = x28 & ~n421 ;
  assign n425 = ~n423 & ~n424 ;
  assign n426 = x27 & ~n425 ;
  assign n427 = ~n422 & ~n426 ;
  assign n428 = ~x25 & ~n427 ;
  assign n429 = ~x26 & ~n425 ;
  assign n430 = x26 & ~n427 ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = x25 & ~n431 ;
  assign n433 = ~n428 & ~n432 ;
  assign n434 = ~x23 & ~n433 ;
  assign n435 = ~x24 & ~n431 ;
  assign n436 = x24 & ~n433 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = x23 & ~n437 ;
  assign n439 = ~n434 & ~n438 ;
  assign n440 = ~x21 & ~n439 ;
  assign n441 = ~x22 & ~n437 ;
  assign n442 = x22 & ~n439 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = x21 & ~n443 ;
  assign n445 = ~n440 & ~n444 ;
  assign n446 = ~x19 & ~n445 ;
  assign n447 = ~x20 & ~n443 ;
  assign n448 = x20 & ~n445 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = x19 & ~n449 ;
  assign n451 = ~n446 & ~n450 ;
  assign n452 = ~x17 & ~n451 ;
  assign n453 = ~x18 & ~n449 ;
  assign n454 = x18 & ~n451 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = x17 & ~n455 ;
  assign n457 = ~n452 & ~n456 ;
  assign n458 = ~x15 & ~n457 ;
  assign n459 = ~x16 & ~n455 ;
  assign n460 = x16 & ~n457 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = x15 & ~n461 ;
  assign n463 = ~n458 & ~n462 ;
  assign n464 = ~x13 & ~n463 ;
  assign n465 = ~x14 & ~n461 ;
  assign n466 = x14 & ~n463 ;
  assign n467 = ~n465 & ~n466 ;
  assign n468 = x13 & ~n467 ;
  assign n469 = ~n464 & ~n468 ;
  assign n470 = ~x11 & ~n469 ;
  assign n471 = ~x12 & ~n467 ;
  assign n472 = x12 & ~n469 ;
  assign n473 = ~n471 & ~n472 ;
  assign n474 = x11 & ~n473 ;
  assign n475 = ~n470 & ~n474 ;
  assign n476 = ~x9 & ~n475 ;
  assign n477 = ~x10 & ~n473 ;
  assign n478 = x10 & ~n475 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = x9 & ~n479 ;
  assign n481 = ~n476 & ~n480 ;
  assign n482 = ~x7 & ~n481 ;
  assign n483 = ~x8 & ~n479 ;
  assign n484 = x8 & ~n481 ;
  assign n485 = ~n483 & ~n484 ;
  assign n486 = x7 & ~n485 ;
  assign n487 = ~n482 & ~n486 ;
  assign n488 = ~x5 & ~n487 ;
  assign n489 = ~x6 & ~n485 ;
  assign n490 = x6 & ~n487 ;
  assign n491 = ~n489 & ~n490 ;
  assign n492 = x5 & ~n491 ;
  assign n493 = ~n488 & ~n492 ;
  assign n494 = ~x3 & ~n493 ;
  assign n495 = ~x4 & ~n491 ;
  assign n496 = x4 & ~n493 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = x3 & ~n497 ;
  assign n499 = ~n494 & ~n498 ;
  assign n500 = x1 & ~x2 ;
  assign n501 = n499 & ~n500 ;
  assign n502 = n497 & n500 ;
  assign n503 = ~n501 & ~n502 ;
  assign n880 = n503 & x128 ;
  assign n504 = x125 & ~x127 ;
  assign n505 = ~x126 & ~x127 ;
  assign n506 = ~x126 & ~n505 ;
  assign n507 = ~x125 & ~n506 ;
  assign n508 = ~n504 & ~n507 ;
  assign n509 = x123 & ~n508 ;
  assign n510 = x124 & ~n506 ;
  assign n511 = ~x124 & ~n508 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = ~x123 & ~n512 ;
  assign n514 = ~n509 & ~n513 ;
  assign n515 = x121 & ~n514 ;
  assign n516 = x122 & ~n512 ;
  assign n517 = ~x122 & ~n514 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = ~x121 & ~n518 ;
  assign n520 = ~n515 & ~n519 ;
  assign n521 = x119 & ~n520 ;
  assign n522 = x120 & ~n518 ;
  assign n523 = ~x120 & ~n520 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~x119 & ~n524 ;
  assign n526 = ~n521 & ~n525 ;
  assign n527 = x117 & ~n526 ;
  assign n528 = x118 & ~n524 ;
  assign n529 = ~x118 & ~n526 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~x117 & ~n530 ;
  assign n532 = ~n527 & ~n531 ;
  assign n533 = x115 & ~n532 ;
  assign n534 = x116 & ~n530 ;
  assign n535 = ~x116 & ~n532 ;
  assign n536 = ~n534 & ~n535 ;
  assign n537 = ~x115 & ~n536 ;
  assign n538 = ~n533 & ~n537 ;
  assign n539 = x113 & ~n538 ;
  assign n540 = x114 & ~n536 ;
  assign n541 = ~x114 & ~n538 ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = ~x113 & ~n542 ;
  assign n544 = ~n539 & ~n543 ;
  assign n545 = x111 & ~n544 ;
  assign n546 = x112 & ~n542 ;
  assign n547 = ~x112 & ~n544 ;
  assign n548 = ~n546 & ~n547 ;
  assign n549 = ~x111 & ~n548 ;
  assign n550 = ~n545 & ~n549 ;
  assign n551 = x109 & ~n550 ;
  assign n552 = x110 & ~n548 ;
  assign n553 = ~x110 & ~n550 ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = ~x109 & ~n554 ;
  assign n556 = ~n551 & ~n555 ;
  assign n557 = x107 & ~n556 ;
  assign n558 = x108 & ~n554 ;
  assign n559 = ~x108 & ~n556 ;
  assign n560 = ~n558 & ~n559 ;
  assign n561 = ~x107 & ~n560 ;
  assign n562 = ~n557 & ~n561 ;
  assign n563 = x105 & ~n562 ;
  assign n564 = x106 & ~n560 ;
  assign n565 = ~x106 & ~n562 ;
  assign n566 = ~n564 & ~n565 ;
  assign n567 = ~x105 & ~n566 ;
  assign n568 = ~n563 & ~n567 ;
  assign n569 = x103 & ~n568 ;
  assign n570 = x104 & ~n566 ;
  assign n571 = ~x104 & ~n568 ;
  assign n572 = ~n570 & ~n571 ;
  assign n573 = ~x103 & ~n572 ;
  assign n574 = ~n569 & ~n573 ;
  assign n575 = x101 & ~n574 ;
  assign n576 = x102 & ~n572 ;
  assign n577 = ~x102 & ~n574 ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = ~x101 & ~n578 ;
  assign n580 = ~n575 & ~n579 ;
  assign n581 = x99 & ~n580 ;
  assign n582 = x100 & ~n578 ;
  assign n583 = ~x100 & ~n580 ;
  assign n584 = ~n582 & ~n583 ;
  assign n585 = ~x99 & ~n584 ;
  assign n586 = ~n581 & ~n585 ;
  assign n587 = x97 & ~n586 ;
  assign n588 = x98 & ~n584 ;
  assign n589 = ~x98 & ~n586 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = ~x97 & ~n590 ;
  assign n592 = ~n587 & ~n591 ;
  assign n593 = x95 & ~n592 ;
  assign n594 = x96 & ~n590 ;
  assign n595 = ~x96 & ~n592 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = ~x95 & ~n596 ;
  assign n598 = ~n593 & ~n597 ;
  assign n599 = x93 & ~n598 ;
  assign n600 = x94 & ~n596 ;
  assign n601 = ~x94 & ~n598 ;
  assign n602 = ~n600 & ~n601 ;
  assign n603 = ~x93 & ~n602 ;
  assign n604 = ~n599 & ~n603 ;
  assign n605 = x91 & ~n604 ;
  assign n606 = x92 & ~n602 ;
  assign n607 = ~x92 & ~n604 ;
  assign n608 = ~n606 & ~n607 ;
  assign n609 = ~x91 & ~n608 ;
  assign n610 = ~n605 & ~n609 ;
  assign n611 = x89 & ~n610 ;
  assign n612 = x90 & ~n608 ;
  assign n613 = ~x90 & ~n610 ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = ~x89 & ~n614 ;
  assign n616 = ~n611 & ~n615 ;
  assign n617 = x87 & ~n616 ;
  assign n618 = x88 & ~n614 ;
  assign n619 = ~x88 & ~n616 ;
  assign n620 = ~n618 & ~n619 ;
  assign n621 = ~x87 & ~n620 ;
  assign n622 = ~n617 & ~n621 ;
  assign n623 = x85 & ~n622 ;
  assign n624 = x86 & ~n620 ;
  assign n625 = ~x86 & ~n622 ;
  assign n626 = ~n624 & ~n625 ;
  assign n627 = ~x85 & ~n626 ;
  assign n628 = ~n623 & ~n627 ;
  assign n629 = x83 & ~n628 ;
  assign n630 = x84 & ~n626 ;
  assign n631 = ~x84 & ~n628 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = ~x83 & ~n632 ;
  assign n634 = ~n629 & ~n633 ;
  assign n635 = x81 & ~n634 ;
  assign n636 = x82 & ~n632 ;
  assign n637 = ~x82 & ~n634 ;
  assign n638 = ~n636 & ~n637 ;
  assign n639 = ~x81 & ~n638 ;
  assign n640 = ~n635 & ~n639 ;
  assign n641 = x79 & ~n640 ;
  assign n642 = x80 & ~n638 ;
  assign n643 = ~x80 & ~n640 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = ~x79 & ~n644 ;
  assign n646 = ~n641 & ~n645 ;
  assign n647 = x77 & ~n646 ;
  assign n648 = x78 & ~n644 ;
  assign n649 = ~x78 & ~n646 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = ~x77 & ~n650 ;
  assign n652 = ~n647 & ~n651 ;
  assign n653 = x75 & ~n652 ;
  assign n654 = x76 & ~n650 ;
  assign n655 = ~x76 & ~n652 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~x75 & ~n656 ;
  assign n658 = ~n653 & ~n657 ;
  assign n659 = x73 & ~n658 ;
  assign n660 = x74 & ~n656 ;
  assign n661 = ~x74 & ~n658 ;
  assign n662 = ~n660 & ~n661 ;
  assign n663 = ~x73 & ~n662 ;
  assign n664 = ~n659 & ~n663 ;
  assign n665 = x71 & ~n664 ;
  assign n666 = x72 & ~n662 ;
  assign n667 = ~x72 & ~n664 ;
  assign n668 = ~n666 & ~n667 ;
  assign n669 = ~x71 & ~n668 ;
  assign n670 = ~n665 & ~n669 ;
  assign n671 = x69 & ~n670 ;
  assign n672 = x70 & ~n668 ;
  assign n673 = ~x70 & ~n670 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~x69 & ~n674 ;
  assign n676 = ~n671 & ~n675 ;
  assign n677 = x67 & ~n676 ;
  assign n678 = x68 & ~n674 ;
  assign n679 = ~x68 & ~n676 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = ~x67 & ~n680 ;
  assign n682 = ~n677 & ~n681 ;
  assign n683 = x65 & ~n682 ;
  assign n684 = x66 & ~n680 ;
  assign n685 = ~x66 & ~n682 ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = ~x65 & ~n686 ;
  assign n688 = ~n683 & ~n687 ;
  assign n689 = x63 & ~n688 ;
  assign n690 = x64 & ~n686 ;
  assign n691 = ~x64 & ~n688 ;
  assign n692 = ~n690 & ~n691 ;
  assign n693 = ~x63 & ~n692 ;
  assign n694 = ~n689 & ~n693 ;
  assign n695 = x61 & ~n694 ;
  assign n696 = x62 & ~n692 ;
  assign n697 = ~x62 & ~n694 ;
  assign n698 = ~n696 & ~n697 ;
  assign n699 = ~x61 & ~n698 ;
  assign n700 = ~n695 & ~n699 ;
  assign n701 = x59 & ~n700 ;
  assign n702 = x60 & ~n698 ;
  assign n703 = ~x60 & ~n700 ;
  assign n704 = ~n702 & ~n703 ;
  assign n705 = ~x59 & ~n704 ;
  assign n706 = ~n701 & ~n705 ;
  assign n707 = x57 & ~n706 ;
  assign n708 = x58 & ~n704 ;
  assign n709 = ~x58 & ~n706 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = ~x57 & ~n710 ;
  assign n712 = ~n707 & ~n711 ;
  assign n713 = x55 & ~n712 ;
  assign n714 = x56 & ~n710 ;
  assign n715 = ~x56 & ~n712 ;
  assign n716 = ~n714 & ~n715 ;
  assign n717 = ~x55 & ~n716 ;
  assign n718 = ~n713 & ~n717 ;
  assign n719 = x53 & ~n718 ;
  assign n720 = x54 & ~n716 ;
  assign n721 = ~x54 & ~n718 ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = ~x53 & ~n722 ;
  assign n724 = ~n719 & ~n723 ;
  assign n725 = x51 & ~n724 ;
  assign n726 = x52 & ~n722 ;
  assign n727 = ~x52 & ~n724 ;
  assign n728 = ~n726 & ~n727 ;
  assign n729 = ~x51 & ~n728 ;
  assign n730 = ~n725 & ~n729 ;
  assign n731 = x49 & ~n730 ;
  assign n732 = x50 & ~n728 ;
  assign n733 = ~x50 & ~n730 ;
  assign n734 = ~n732 & ~n733 ;
  assign n735 = ~x49 & ~n734 ;
  assign n736 = ~n731 & ~n735 ;
  assign n737 = x47 & ~n736 ;
  assign n738 = x48 & ~n734 ;
  assign n739 = ~x48 & ~n736 ;
  assign n740 = ~n738 & ~n739 ;
  assign n741 = ~x47 & ~n740 ;
  assign n742 = ~n737 & ~n741 ;
  assign n743 = x45 & ~n742 ;
  assign n744 = x46 & ~n740 ;
  assign n745 = ~x46 & ~n742 ;
  assign n746 = ~n744 & ~n745 ;
  assign n747 = ~x45 & ~n746 ;
  assign n748 = ~n743 & ~n747 ;
  assign n749 = x43 & ~n748 ;
  assign n750 = x44 & ~n746 ;
  assign n751 = ~x44 & ~n748 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = ~x43 & ~n752 ;
  assign n754 = ~n749 & ~n753 ;
  assign n755 = x41 & ~n754 ;
  assign n756 = x42 & ~n752 ;
  assign n757 = ~x42 & ~n754 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = ~x41 & ~n758 ;
  assign n760 = ~n755 & ~n759 ;
  assign n761 = x39 & ~n760 ;
  assign n762 = x40 & ~n758 ;
  assign n763 = ~x40 & ~n760 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = ~x39 & ~n764 ;
  assign n766 = ~n761 & ~n765 ;
  assign n767 = x37 & ~n766 ;
  assign n768 = x38 & ~n764 ;
  assign n769 = ~x38 & ~n766 ;
  assign n770 = ~n768 & ~n769 ;
  assign n771 = ~x37 & ~n770 ;
  assign n772 = ~n767 & ~n771 ;
  assign n773 = x35 & ~n772 ;
  assign n774 = x36 & ~n770 ;
  assign n775 = ~x36 & ~n772 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = ~x35 & ~n776 ;
  assign n778 = ~n773 & ~n777 ;
  assign n779 = x33 & ~n778 ;
  assign n780 = x34 & ~n776 ;
  assign n781 = ~x34 & ~n778 ;
  assign n782 = ~n780 & ~n781 ;
  assign n783 = ~x33 & ~n782 ;
  assign n784 = ~n779 & ~n783 ;
  assign n785 = x31 & ~n784 ;
  assign n786 = x32 & ~n782 ;
  assign n787 = ~x32 & ~n784 ;
  assign n788 = ~n786 & ~n787 ;
  assign n789 = ~x31 & ~n788 ;
  assign n790 = ~n785 & ~n789 ;
  assign n791 = x29 & ~n790 ;
  assign n792 = x30 & ~n788 ;
  assign n793 = ~x30 & ~n790 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = ~x29 & ~n794 ;
  assign n796 = ~n791 & ~n795 ;
  assign n797 = x27 & ~n796 ;
  assign n798 = x28 & ~n794 ;
  assign n799 = ~x28 & ~n796 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = ~x27 & ~n800 ;
  assign n802 = ~n797 & ~n801 ;
  assign n803 = x25 & ~n802 ;
  assign n804 = x26 & ~n800 ;
  assign n805 = ~x26 & ~n802 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~x25 & ~n806 ;
  assign n808 = ~n803 & ~n807 ;
  assign n809 = x23 & ~n808 ;
  assign n810 = x24 & ~n806 ;
  assign n811 = ~x24 & ~n808 ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = ~x23 & ~n812 ;
  assign n814 = ~n809 & ~n813 ;
  assign n815 = x21 & ~n814 ;
  assign n816 = x22 & ~n812 ;
  assign n817 = ~x22 & ~n814 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = ~x21 & ~n818 ;
  assign n820 = ~n815 & ~n819 ;
  assign n821 = x19 & ~n820 ;
  assign n822 = x20 & ~n818 ;
  assign n823 = ~x20 & ~n820 ;
  assign n824 = ~n822 & ~n823 ;
  assign n825 = ~x19 & ~n824 ;
  assign n826 = ~n821 & ~n825 ;
  assign n827 = x17 & ~n826 ;
  assign n828 = x18 & ~n824 ;
  assign n829 = ~x18 & ~n826 ;
  assign n830 = ~n828 & ~n829 ;
  assign n831 = ~x17 & ~n830 ;
  assign n832 = ~n827 & ~n831 ;
  assign n833 = x15 & ~n832 ;
  assign n834 = x16 & ~n830 ;
  assign n835 = ~x16 & ~n832 ;
  assign n836 = ~n834 & ~n835 ;
  assign n837 = ~x15 & ~n836 ;
  assign n838 = ~n833 & ~n837 ;
  assign n839 = x13 & ~n838 ;
  assign n840 = x14 & ~n836 ;
  assign n841 = ~x14 & ~n838 ;
  assign n842 = ~n840 & ~n841 ;
  assign n843 = ~x13 & ~n842 ;
  assign n844 = ~n839 & ~n843 ;
  assign n845 = x11 & ~n844 ;
  assign n846 = x12 & ~n842 ;
  assign n847 = ~x12 & ~n844 ;
  assign n848 = ~n846 & ~n847 ;
  assign n849 = ~x11 & ~n848 ;
  assign n850 = ~n845 & ~n849 ;
  assign n851 = x9 & ~n850 ;
  assign n852 = x10 & ~n848 ;
  assign n853 = ~x10 & ~n850 ;
  assign n854 = ~n852 & ~n853 ;
  assign n855 = ~x9 & ~n854 ;
  assign n856 = ~n851 & ~n855 ;
  assign n857 = x7 & ~n856 ;
  assign n858 = x8 & ~n854 ;
  assign n859 = ~x8 & ~n856 ;
  assign n860 = ~n858 & ~n859 ;
  assign n861 = ~x7 & ~n860 ;
  assign n862 = ~n857 & ~n861 ;
  assign n863 = x5 & ~n862 ;
  assign n864 = x6 & ~n860 ;
  assign n865 = ~x6 & ~n862 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = ~x5 & ~n866 ;
  assign n868 = ~n863 & ~n867 ;
  assign n869 = x3 & ~n868 ;
  assign n870 = x4 & ~n866 ;
  assign n871 = ~x4 & ~n868 ;
  assign n872 = ~n870 & ~n871 ;
  assign n873 = ~x3 & ~n872 ;
  assign n874 = ~n869 & ~n873 ;
  assign n875 = ~x1 & x2 ;
  assign n876 = n874 & ~n875 ;
  assign n877 = n872 & n875 ;
  assign n878 = ~n876 & ~n877 ;
  assign n881 = ~n878 & ~x128 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = ~x126 & x127 ;
  assign n884 = ~x126 & ~n883 ;
  assign n885 = ~x124 & ~x125 ;
  assign n886 = ~x122 & ~x123 ;
  assign n887 = x121 & n886 ;
  assign n888 = n885 & ~n887 ;
  assign n889 = n884 & ~n888 ;
  assign n890 = ~x120 & ~n889 ;
  assign n891 = n885 & ~n886 ;
  assign n892 = n884 & ~n891 ;
  assign n893 = x120 & ~n892 ;
  assign n894 = ~n890 & ~n893 ;
  assign n895 = ~x118 & ~x119 ;
  assign n896 = n894 & ~n895 ;
  assign n897 = n892 & n895 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~x116 & ~x117 ;
  assign n900 = n898 & ~n899 ;
  assign n901 = ~n894 & n899 ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = ~x114 & ~x115 ;
  assign n904 = n902 & ~n903 ;
  assign n905 = ~n898 & n903 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = ~x112 & ~x113 ;
  assign n908 = n906 & ~n907 ;
  assign n909 = ~n902 & n907 ;
  assign n910 = ~n908 & ~n909 ;
  assign n911 = ~x110 & ~x111 ;
  assign n912 = n910 & ~n911 ;
  assign n913 = ~n906 & n911 ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = ~x108 & ~x109 ;
  assign n916 = n914 & ~n915 ;
  assign n917 = ~n910 & n915 ;
  assign n918 = ~n916 & ~n917 ;
  assign n919 = ~x106 & ~x107 ;
  assign n920 = n918 & ~n919 ;
  assign n921 = ~n914 & n919 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = ~x104 & ~x105 ;
  assign n924 = n922 & ~n923 ;
  assign n925 = ~n918 & n923 ;
  assign n926 = ~n924 & ~n925 ;
  assign n927 = ~x102 & ~x103 ;
  assign n928 = n926 & ~n927 ;
  assign n929 = ~n922 & n927 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = ~x100 & ~x101 ;
  assign n932 = n930 & ~n931 ;
  assign n933 = ~n926 & n931 ;
  assign n934 = ~n932 & ~n933 ;
  assign n935 = ~x98 & ~x99 ;
  assign n936 = n934 & ~n935 ;
  assign n937 = ~n930 & n935 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~x96 & ~x97 ;
  assign n940 = n938 & ~n939 ;
  assign n941 = ~n934 & n939 ;
  assign n942 = ~n940 & ~n941 ;
  assign n943 = ~x94 & ~x95 ;
  assign n944 = n942 & ~n943 ;
  assign n945 = ~n938 & n943 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~x92 & ~x93 ;
  assign n948 = n946 & ~n947 ;
  assign n949 = ~n942 & n947 ;
  assign n950 = ~n948 & ~n949 ;
  assign n951 = ~x90 & ~x91 ;
  assign n952 = n950 & ~n951 ;
  assign n953 = ~n946 & n951 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = ~x88 & ~x89 ;
  assign n956 = n954 & ~n955 ;
  assign n957 = ~n950 & n955 ;
  assign n958 = ~n956 & ~n957 ;
  assign n959 = ~x86 & ~x87 ;
  assign n960 = n958 & ~n959 ;
  assign n961 = ~n954 & n959 ;
  assign n962 = ~n960 & ~n961 ;
  assign n963 = ~x84 & ~x85 ;
  assign n964 = n962 & ~n963 ;
  assign n965 = ~n958 & n963 ;
  assign n966 = ~n964 & ~n965 ;
  assign n967 = ~x82 & ~x83 ;
  assign n968 = n966 & ~n967 ;
  assign n969 = ~n962 & n967 ;
  assign n970 = ~n968 & ~n969 ;
  assign n971 = ~x80 & ~x81 ;
  assign n972 = n970 & ~n971 ;
  assign n973 = ~n966 & n971 ;
  assign n974 = ~n972 & ~n973 ;
  assign n975 = ~x78 & ~x79 ;
  assign n976 = n974 & ~n975 ;
  assign n977 = ~n970 & n975 ;
  assign n978 = ~n976 & ~n977 ;
  assign n979 = ~x76 & ~x77 ;
  assign n980 = n978 & ~n979 ;
  assign n981 = ~n974 & n979 ;
  assign n982 = ~n980 & ~n981 ;
  assign n983 = ~x74 & ~x75 ;
  assign n984 = n982 & ~n983 ;
  assign n985 = ~n978 & n983 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~x72 & ~x73 ;
  assign n988 = n986 & ~n987 ;
  assign n989 = ~n982 & n987 ;
  assign n990 = ~n988 & ~n989 ;
  assign n991 = ~x70 & ~x71 ;
  assign n992 = n990 & ~n991 ;
  assign n993 = ~n986 & n991 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = ~x68 & ~x69 ;
  assign n996 = n994 & ~n995 ;
  assign n997 = ~n990 & n995 ;
  assign n998 = ~n996 & ~n997 ;
  assign n999 = ~x66 & ~x67 ;
  assign n1000 = n998 & ~n999 ;
  assign n1001 = ~n994 & n999 ;
  assign n1002 = ~n1000 & ~n1001 ;
  assign n1003 = ~x64 & ~x65 ;
  assign n1004 = n1002 & ~n1003 ;
  assign n1005 = ~n998 & n1003 ;
  assign n1006 = ~n1004 & ~n1005 ;
  assign n1007 = ~x62 & ~x63 ;
  assign n1008 = n1006 & ~n1007 ;
  assign n1009 = ~n1002 & n1007 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = ~x60 & ~x61 ;
  assign n1012 = n1010 & ~n1011 ;
  assign n1013 = ~n1006 & n1011 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = ~x58 & ~x59 ;
  assign n1016 = n1014 & ~n1015 ;
  assign n1017 = ~n1010 & n1015 ;
  assign n1018 = ~n1016 & ~n1017 ;
  assign n1019 = ~x56 & ~x57 ;
  assign n1020 = n1018 & ~n1019 ;
  assign n1021 = ~n1014 & n1019 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = ~x54 & ~x55 ;
  assign n1024 = n1022 & ~n1023 ;
  assign n1025 = ~n1018 & n1023 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~x52 & ~x53 ;
  assign n1028 = n1026 & ~n1027 ;
  assign n1029 = ~n1022 & n1027 ;
  assign n1030 = ~n1028 & ~n1029 ;
  assign n1031 = ~x50 & ~x51 ;
  assign n1032 = n1030 & ~n1031 ;
  assign n1033 = ~n1026 & n1031 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = ~x48 & ~x49 ;
  assign n1036 = n1034 & ~n1035 ;
  assign n1037 = ~n1030 & n1035 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = ~x46 & ~x47 ;
  assign n1040 = n1038 & ~n1039 ;
  assign n1041 = ~n1034 & n1039 ;
  assign n1042 = ~n1040 & ~n1041 ;
  assign n1043 = ~x44 & ~x45 ;
  assign n1044 = n1042 & ~n1043 ;
  assign n1045 = ~n1038 & n1043 ;
  assign n1046 = ~n1044 & ~n1045 ;
  assign n1047 = ~x42 & ~x43 ;
  assign n1048 = n1046 & ~n1047 ;
  assign n1049 = ~n1042 & n1047 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = ~x40 & ~x41 ;
  assign n1052 = n1050 & ~n1051 ;
  assign n1053 = ~n1046 & n1051 ;
  assign n1054 = ~n1052 & ~n1053 ;
  assign n1055 = ~x38 & ~x39 ;
  assign n1056 = n1054 & ~n1055 ;
  assign n1057 = ~n1050 & n1055 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = ~x36 & ~x37 ;
  assign n1060 = n1058 & ~n1059 ;
  assign n1061 = ~n1054 & n1059 ;
  assign n1062 = ~n1060 & ~n1061 ;
  assign n1063 = ~x34 & ~x35 ;
  assign n1064 = n1062 & ~n1063 ;
  assign n1065 = ~n1058 & n1063 ;
  assign n1066 = ~n1064 & ~n1065 ;
  assign n1067 = ~x32 & ~x33 ;
  assign n1068 = n1066 & ~n1067 ;
  assign n1069 = ~n1062 & n1067 ;
  assign n1070 = ~n1068 & ~n1069 ;
  assign n1071 = ~x30 & ~x31 ;
  assign n1072 = n1070 & ~n1071 ;
  assign n1073 = ~n1066 & n1071 ;
  assign n1074 = ~n1072 & ~n1073 ;
  assign n1075 = ~x28 & ~x29 ;
  assign n1076 = n1074 & ~n1075 ;
  assign n1077 = ~n1070 & n1075 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1079 = ~x26 & ~x27 ;
  assign n1080 = n1078 & ~n1079 ;
  assign n1081 = ~n1074 & n1079 ;
  assign n1082 = ~n1080 & ~n1081 ;
  assign n1083 = ~x24 & ~x25 ;
  assign n1084 = n1082 & ~n1083 ;
  assign n1085 = ~n1078 & n1083 ;
  assign n1086 = ~n1084 & ~n1085 ;
  assign n1087 = ~x22 & ~x23 ;
  assign n1088 = n1086 & ~n1087 ;
  assign n1089 = ~n1082 & n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = ~x20 & ~x21 ;
  assign n1092 = n1090 & ~n1091 ;
  assign n1093 = ~n1086 & n1091 ;
  assign n1094 = ~n1092 & ~n1093 ;
  assign n1095 = ~x18 & ~x19 ;
  assign n1096 = n1094 & ~n1095 ;
  assign n1097 = ~n1090 & n1095 ;
  assign n1098 = ~n1096 & ~n1097 ;
  assign n1099 = ~x16 & ~x17 ;
  assign n1100 = n1098 & ~n1099 ;
  assign n1101 = ~n1094 & n1099 ;
  assign n1102 = ~n1100 & ~n1101 ;
  assign n1103 = ~x14 & ~x15 ;
  assign n1104 = n1102 & ~n1103 ;
  assign n1105 = ~n1098 & n1103 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = ~x12 & ~x13 ;
  assign n1108 = n1106 & ~n1107 ;
  assign n1109 = ~n1102 & n1107 ;
  assign n1110 = ~n1108 & ~n1109 ;
  assign n1111 = ~x10 & ~x11 ;
  assign n1112 = n1110 & ~n1111 ;
  assign n1113 = ~n1106 & n1111 ;
  assign n1114 = ~n1112 & ~n1113 ;
  assign n1115 = ~x8 & ~x9 ;
  assign n1116 = n1114 & ~n1115 ;
  assign n1117 = ~n1110 & n1115 ;
  assign n1118 = ~n1116 & ~n1117 ;
  assign n1119 = ~x6 & ~x7 ;
  assign n1120 = n1118 & ~n1119 ;
  assign n1121 = ~n1114 & n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~x4 & ~x5 ;
  assign n1124 = n1122 & ~n1123 ;
  assign n1125 = ~n1118 & n1123 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = ~x2 & ~x3 ;
  assign n1128 = n1126 & ~n1127 ;
  assign n1129 = ~n1122 & n1127 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1380 = n1130 & x129 ;
  assign n1131 = x126 & ~x127 ;
  assign n1132 = x126 & ~n1131 ;
  assign n1133 = x124 & x125 ;
  assign n1134 = x122 & x123 ;
  assign n1135 = ~x121 & n1134 ;
  assign n1136 = n1133 & ~n1135 ;
  assign n1137 = n1132 & ~n1136 ;
  assign n1138 = x120 & ~n1137 ;
  assign n1139 = n1133 & ~n1134 ;
  assign n1140 = n1132 & ~n1139 ;
  assign n1141 = ~x120 & ~n1140 ;
  assign n1142 = ~n1138 & ~n1141 ;
  assign n1143 = x118 & x119 ;
  assign n1144 = n1142 & ~n1143 ;
  assign n1145 = n1140 & n1143 ;
  assign n1146 = ~n1144 & ~n1145 ;
  assign n1147 = x116 & x117 ;
  assign n1148 = n1146 & ~n1147 ;
  assign n1149 = ~n1142 & n1147 ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = x114 & x115 ;
  assign n1152 = n1150 & ~n1151 ;
  assign n1153 = ~n1146 & n1151 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = x112 & x113 ;
  assign n1156 = n1154 & ~n1155 ;
  assign n1157 = ~n1150 & n1155 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1159 = x110 & x111 ;
  assign n1160 = n1158 & ~n1159 ;
  assign n1161 = ~n1154 & n1159 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = x108 & x109 ;
  assign n1164 = n1162 & ~n1163 ;
  assign n1165 = ~n1158 & n1163 ;
  assign n1166 = ~n1164 & ~n1165 ;
  assign n1167 = x106 & x107 ;
  assign n1168 = n1166 & ~n1167 ;
  assign n1169 = ~n1162 & n1167 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = x104 & x105 ;
  assign n1172 = n1170 & ~n1171 ;
  assign n1173 = ~n1166 & n1171 ;
  assign n1174 = ~n1172 & ~n1173 ;
  assign n1175 = x102 & x103 ;
  assign n1176 = n1174 & ~n1175 ;
  assign n1177 = ~n1170 & n1175 ;
  assign n1178 = ~n1176 & ~n1177 ;
  assign n1179 = x100 & x101 ;
  assign n1180 = n1178 & ~n1179 ;
  assign n1181 = ~n1174 & n1179 ;
  assign n1182 = ~n1180 & ~n1181 ;
  assign n1183 = x98 & x99 ;
  assign n1184 = n1182 & ~n1183 ;
  assign n1185 = ~n1178 & n1183 ;
  assign n1186 = ~n1184 & ~n1185 ;
  assign n1187 = x96 & x97 ;
  assign n1188 = n1186 & ~n1187 ;
  assign n1189 = ~n1182 & n1187 ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = x94 & x95 ;
  assign n1192 = n1190 & ~n1191 ;
  assign n1193 = ~n1186 & n1191 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = x92 & x93 ;
  assign n1196 = n1194 & ~n1195 ;
  assign n1197 = ~n1190 & n1195 ;
  assign n1198 = ~n1196 & ~n1197 ;
  assign n1199 = x90 & x91 ;
  assign n1200 = n1198 & ~n1199 ;
  assign n1201 = ~n1194 & n1199 ;
  assign n1202 = ~n1200 & ~n1201 ;
  assign n1203 = x88 & x89 ;
  assign n1204 = n1202 & ~n1203 ;
  assign n1205 = ~n1198 & n1203 ;
  assign n1206 = ~n1204 & ~n1205 ;
  assign n1207 = x86 & x87 ;
  assign n1208 = n1206 & ~n1207 ;
  assign n1209 = ~n1202 & n1207 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = x84 & x85 ;
  assign n1212 = n1210 & ~n1211 ;
  assign n1213 = ~n1206 & n1211 ;
  assign n1214 = ~n1212 & ~n1213 ;
  assign n1215 = x82 & x83 ;
  assign n1216 = n1214 & ~n1215 ;
  assign n1217 = ~n1210 & n1215 ;
  assign n1218 = ~n1216 & ~n1217 ;
  assign n1219 = x80 & x81 ;
  assign n1220 = n1218 & ~n1219 ;
  assign n1221 = ~n1214 & n1219 ;
  assign n1222 = ~n1220 & ~n1221 ;
  assign n1223 = x78 & x79 ;
  assign n1224 = n1222 & ~n1223 ;
  assign n1225 = ~n1218 & n1223 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1227 = x76 & x77 ;
  assign n1228 = n1226 & ~n1227 ;
  assign n1229 = ~n1222 & n1227 ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = x74 & x75 ;
  assign n1232 = n1230 & ~n1231 ;
  assign n1233 = ~n1226 & n1231 ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = x72 & x73 ;
  assign n1236 = n1234 & ~n1235 ;
  assign n1237 = ~n1230 & n1235 ;
  assign n1238 = ~n1236 & ~n1237 ;
  assign n1239 = x70 & x71 ;
  assign n1240 = n1238 & ~n1239 ;
  assign n1241 = ~n1234 & n1239 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = x68 & x69 ;
  assign n1244 = n1242 & ~n1243 ;
  assign n1245 = ~n1238 & n1243 ;
  assign n1246 = ~n1244 & ~n1245 ;
  assign n1247 = x66 & x67 ;
  assign n1248 = n1246 & ~n1247 ;
  assign n1249 = ~n1242 & n1247 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = x64 & x65 ;
  assign n1252 = n1250 & ~n1251 ;
  assign n1253 = ~n1246 & n1251 ;
  assign n1254 = ~n1252 & ~n1253 ;
  assign n1255 = x62 & x63 ;
  assign n1256 = n1254 & ~n1255 ;
  assign n1257 = ~n1250 & n1255 ;
  assign n1258 = ~n1256 & ~n1257 ;
  assign n1259 = x60 & x61 ;
  assign n1260 = n1258 & ~n1259 ;
  assign n1261 = ~n1254 & n1259 ;
  assign n1262 = ~n1260 & ~n1261 ;
  assign n1263 = x58 & x59 ;
  assign n1264 = n1262 & ~n1263 ;
  assign n1265 = ~n1258 & n1263 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = x56 & x57 ;
  assign n1268 = n1266 & ~n1267 ;
  assign n1269 = ~n1262 & n1267 ;
  assign n1270 = ~n1268 & ~n1269 ;
  assign n1271 = x54 & x55 ;
  assign n1272 = n1270 & ~n1271 ;
  assign n1273 = ~n1266 & n1271 ;
  assign n1274 = ~n1272 & ~n1273 ;
  assign n1275 = x52 & x53 ;
  assign n1276 = n1274 & ~n1275 ;
  assign n1277 = ~n1270 & n1275 ;
  assign n1278 = ~n1276 & ~n1277 ;
  assign n1279 = x50 & x51 ;
  assign n1280 = n1278 & ~n1279 ;
  assign n1281 = ~n1274 & n1279 ;
  assign n1282 = ~n1280 & ~n1281 ;
  assign n1283 = x48 & x49 ;
  assign n1284 = n1282 & ~n1283 ;
  assign n1285 = ~n1278 & n1283 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = x46 & x47 ;
  assign n1288 = n1286 & ~n1287 ;
  assign n1289 = ~n1282 & n1287 ;
  assign n1290 = ~n1288 & ~n1289 ;
  assign n1291 = x44 & x45 ;
  assign n1292 = n1290 & ~n1291 ;
  assign n1293 = ~n1286 & n1291 ;
  assign n1294 = ~n1292 & ~n1293 ;
  assign n1295 = x42 & x43 ;
  assign n1296 = n1294 & ~n1295 ;
  assign n1297 = ~n1290 & n1295 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = x40 & x41 ;
  assign n1300 = n1298 & ~n1299 ;
  assign n1301 = ~n1294 & n1299 ;
  assign n1302 = ~n1300 & ~n1301 ;
  assign n1303 = x38 & x39 ;
  assign n1304 = n1302 & ~n1303 ;
  assign n1305 = ~n1298 & n1303 ;
  assign n1306 = ~n1304 & ~n1305 ;
  assign n1307 = x36 & x37 ;
  assign n1308 = n1306 & ~n1307 ;
  assign n1309 = ~n1302 & n1307 ;
  assign n1310 = ~n1308 & ~n1309 ;
  assign n1311 = x34 & x35 ;
  assign n1312 = n1310 & ~n1311 ;
  assign n1313 = ~n1306 & n1311 ;
  assign n1314 = ~n1312 & ~n1313 ;
  assign n1315 = x32 & x33 ;
  assign n1316 = n1314 & ~n1315 ;
  assign n1317 = ~n1310 & n1315 ;
  assign n1318 = ~n1316 & ~n1317 ;
  assign n1319 = x30 & x31 ;
  assign n1320 = n1318 & ~n1319 ;
  assign n1321 = ~n1314 & n1319 ;
  assign n1322 = ~n1320 & ~n1321 ;
  assign n1323 = x28 & x29 ;
  assign n1324 = n1322 & ~n1323 ;
  assign n1325 = ~n1318 & n1323 ;
  assign n1326 = ~n1324 & ~n1325 ;
  assign n1327 = x26 & x27 ;
  assign n1328 = n1326 & ~n1327 ;
  assign n1329 = ~n1322 & n1327 ;
  assign n1330 = ~n1328 & ~n1329 ;
  assign n1331 = x24 & x25 ;
  assign n1332 = n1330 & ~n1331 ;
  assign n1333 = ~n1326 & n1331 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = x22 & x23 ;
  assign n1336 = n1334 & ~n1335 ;
  assign n1337 = ~n1330 & n1335 ;
  assign n1338 = ~n1336 & ~n1337 ;
  assign n1339 = x20 & x21 ;
  assign n1340 = n1338 & ~n1339 ;
  assign n1341 = ~n1334 & n1339 ;
  assign n1342 = ~n1340 & ~n1341 ;
  assign n1343 = x18 & x19 ;
  assign n1344 = n1342 & ~n1343 ;
  assign n1345 = ~n1338 & n1343 ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = x16 & x17 ;
  assign n1348 = n1346 & ~n1347 ;
  assign n1349 = ~n1342 & n1347 ;
  assign n1350 = ~n1348 & ~n1349 ;
  assign n1351 = x14 & x15 ;
  assign n1352 = n1350 & ~n1351 ;
  assign n1353 = ~n1346 & n1351 ;
  assign n1354 = ~n1352 & ~n1353 ;
  assign n1355 = x12 & x13 ;
  assign n1356 = n1354 & ~n1355 ;
  assign n1357 = ~n1350 & n1355 ;
  assign n1358 = ~n1356 & ~n1357 ;
  assign n1359 = x10 & x11 ;
  assign n1360 = n1358 & ~n1359 ;
  assign n1361 = ~n1354 & n1359 ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = x8 & x9 ;
  assign n1364 = n1362 & ~n1363 ;
  assign n1365 = ~n1358 & n1363 ;
  assign n1366 = ~n1364 & ~n1365 ;
  assign n1367 = x6 & x7 ;
  assign n1368 = n1366 & ~n1367 ;
  assign n1369 = ~n1362 & n1367 ;
  assign n1370 = ~n1368 & ~n1369 ;
  assign n1371 = x4 & x5 ;
  assign n1372 = n1370 & ~n1371 ;
  assign n1373 = ~n1366 & n1371 ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1375 = x2 & x3 ;
  assign n1376 = n1374 & ~n1375 ;
  assign n1377 = ~n1370 & n1375 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1381 = ~n1378 & ~x129 ;
  assign n1382 = ~n1380 & ~n1381 ;
  assign n1383 = n884 & n885 ;
  assign n1384 = ~x120 & ~x121 ;
  assign n1385 = n886 & n1384 ;
  assign n1386 = ~x117 & n895 ;
  assign n1387 = ~x116 & n1386 ;
  assign n1388 = n1385 & ~n1387 ;
  assign n1389 = n1383 & ~n1388 ;
  assign n1390 = ~x113 & ~x114 ;
  assign n1391 = ~x112 & n1390 ;
  assign n1392 = n1389 & ~n1391 ;
  assign n1393 = x115 & n1387 ;
  assign n1394 = n1385 & ~n1393 ;
  assign n1395 = n1383 & ~n1394 ;
  assign n1396 = n1391 & n1395 ;
  assign n1397 = ~n1392 & ~n1396 ;
  assign n1398 = ~x109 & n911 ;
  assign n1399 = ~x108 & n1398 ;
  assign n1400 = n1397 & ~n1399 ;
  assign n1401 = ~n1389 & n1399 ;
  assign n1402 = ~n1400 & ~n1401 ;
  assign n1403 = ~x105 & n919 ;
  assign n1404 = ~x104 & n1403 ;
  assign n1405 = n1402 & ~n1404 ;
  assign n1406 = ~n1397 & n1404 ;
  assign n1407 = ~n1405 & ~n1406 ;
  assign n1408 = ~x101 & n927 ;
  assign n1409 = ~x100 & n1408 ;
  assign n1410 = n1407 & ~n1409 ;
  assign n1411 = ~n1402 & n1409 ;
  assign n1412 = ~n1410 & ~n1411 ;
  assign n1413 = ~x97 & n935 ;
  assign n1414 = ~x96 & n1413 ;
  assign n1415 = n1412 & ~n1414 ;
  assign n1416 = ~n1407 & n1414 ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = ~x93 & n943 ;
  assign n1419 = ~x92 & n1418 ;
  assign n1420 = n1417 & ~n1419 ;
  assign n1421 = ~n1412 & n1419 ;
  assign n1422 = ~n1420 & ~n1421 ;
  assign n1423 = ~x89 & n951 ;
  assign n1424 = ~x88 & n1423 ;
  assign n1425 = n1422 & ~n1424 ;
  assign n1426 = ~n1417 & n1424 ;
  assign n1427 = ~n1425 & ~n1426 ;
  assign n1428 = ~x85 & n959 ;
  assign n1429 = ~x84 & n1428 ;
  assign n1430 = n1427 & ~n1429 ;
  assign n1431 = ~n1422 & n1429 ;
  assign n1432 = ~n1430 & ~n1431 ;
  assign n1433 = ~x81 & n967 ;
  assign n1434 = ~x80 & n1433 ;
  assign n1435 = n1432 & ~n1434 ;
  assign n1436 = ~n1427 & n1434 ;
  assign n1437 = ~n1435 & ~n1436 ;
  assign n1438 = ~x77 & n975 ;
  assign n1439 = ~x76 & n1438 ;
  assign n1440 = n1437 & ~n1439 ;
  assign n1441 = ~n1432 & n1439 ;
  assign n1442 = ~n1440 & ~n1441 ;
  assign n1443 = ~x73 & n983 ;
  assign n1444 = ~x72 & n1443 ;
  assign n1445 = n1442 & ~n1444 ;
  assign n1446 = ~n1437 & n1444 ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1448 = ~x69 & n991 ;
  assign n1449 = ~x68 & n1448 ;
  assign n1450 = n1447 & ~n1449 ;
  assign n1451 = ~n1442 & n1449 ;
  assign n1452 = ~n1450 & ~n1451 ;
  assign n1453 = ~x65 & n999 ;
  assign n1454 = ~x64 & n1453 ;
  assign n1455 = n1452 & ~n1454 ;
  assign n1456 = ~n1447 & n1454 ;
  assign n1457 = ~n1455 & ~n1456 ;
  assign n1458 = ~x61 & n1007 ;
  assign n1459 = ~x60 & n1458 ;
  assign n1460 = n1457 & ~n1459 ;
  assign n1461 = ~n1452 & n1459 ;
  assign n1462 = ~n1460 & ~n1461 ;
  assign n1463 = ~x57 & n1015 ;
  assign n1464 = ~x56 & n1463 ;
  assign n1465 = n1462 & ~n1464 ;
  assign n1466 = ~n1457 & n1464 ;
  assign n1467 = ~n1465 & ~n1466 ;
  assign n1468 = ~x53 & n1023 ;
  assign n1469 = ~x52 & n1468 ;
  assign n1470 = n1467 & ~n1469 ;
  assign n1471 = ~n1462 & n1469 ;
  assign n1472 = ~n1470 & ~n1471 ;
  assign n1473 = ~x49 & n1031 ;
  assign n1474 = ~x48 & n1473 ;
  assign n1475 = n1472 & ~n1474 ;
  assign n1476 = ~n1467 & n1474 ;
  assign n1477 = ~n1475 & ~n1476 ;
  assign n1478 = ~x45 & n1039 ;
  assign n1479 = ~x44 & n1478 ;
  assign n1480 = n1477 & ~n1479 ;
  assign n1481 = ~n1472 & n1479 ;
  assign n1482 = ~n1480 & ~n1481 ;
  assign n1483 = ~x41 & n1047 ;
  assign n1484 = ~x40 & n1483 ;
  assign n1485 = n1482 & ~n1484 ;
  assign n1486 = ~n1477 & n1484 ;
  assign n1487 = ~n1485 & ~n1486 ;
  assign n1488 = ~x37 & n1055 ;
  assign n1489 = ~x36 & n1488 ;
  assign n1490 = n1487 & ~n1489 ;
  assign n1491 = ~n1482 & n1489 ;
  assign n1492 = ~n1490 & ~n1491 ;
  assign n1493 = ~x33 & n1063 ;
  assign n1494 = ~x32 & n1493 ;
  assign n1495 = n1492 & ~n1494 ;
  assign n1496 = ~n1487 & n1494 ;
  assign n1497 = ~n1495 & ~n1496 ;
  assign n1498 = ~x29 & n1071 ;
  assign n1499 = ~x28 & n1498 ;
  assign n1500 = n1497 & ~n1499 ;
  assign n1501 = ~n1492 & n1499 ;
  assign n1502 = ~n1500 & ~n1501 ;
  assign n1503 = ~x25 & n1079 ;
  assign n1504 = ~x24 & n1503 ;
  assign n1505 = n1502 & ~n1504 ;
  assign n1506 = ~n1497 & n1504 ;
  assign n1507 = ~n1505 & ~n1506 ;
  assign n1508 = ~x21 & n1087 ;
  assign n1509 = ~x20 & n1508 ;
  assign n1510 = n1507 & ~n1509 ;
  assign n1511 = ~n1502 & n1509 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = ~x17 & n1095 ;
  assign n1514 = ~x16 & n1513 ;
  assign n1515 = n1512 & ~n1514 ;
  assign n1516 = ~n1507 & n1514 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = ~x13 & n1103 ;
  assign n1519 = ~x12 & n1518 ;
  assign n1520 = n1517 & ~n1519 ;
  assign n1521 = ~n1512 & n1519 ;
  assign n1522 = ~n1520 & ~n1521 ;
  assign n1523 = ~x9 & n1111 ;
  assign n1524 = ~x8 & n1523 ;
  assign n1525 = n1522 & ~n1524 ;
  assign n1526 = ~n1517 & n1524 ;
  assign n1527 = ~n1525 & ~n1526 ;
  assign n1528 = ~x5 & n1119 ;
  assign n1529 = ~x4 & n1528 ;
  assign n1530 = n1527 & ~n1529 ;
  assign n1531 = ~n1522 & n1529 ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1684 = ~n1532 & x130 ;
  assign n1533 = n1132 & n1133 ;
  assign n1534 = x120 & x121 ;
  assign n1535 = n1134 & n1534 ;
  assign n1536 = x117 & n1143 ;
  assign n1537 = x116 & n1536 ;
  assign n1538 = n1535 & ~n1537 ;
  assign n1539 = n1533 & ~n1538 ;
  assign n1540 = x113 & x114 ;
  assign n1541 = x112 & n1540 ;
  assign n1542 = n1539 & ~n1541 ;
  assign n1543 = ~x115 & n1537 ;
  assign n1544 = n1535 & ~n1543 ;
  assign n1545 = n1533 & ~n1544 ;
  assign n1546 = n1541 & n1545 ;
  assign n1547 = ~n1542 & ~n1546 ;
  assign n1548 = x109 & n1159 ;
  assign n1549 = x108 & n1548 ;
  assign n1550 = n1547 & ~n1549 ;
  assign n1551 = ~n1539 & n1549 ;
  assign n1552 = ~n1550 & ~n1551 ;
  assign n1553 = x105 & n1167 ;
  assign n1554 = x104 & n1553 ;
  assign n1555 = n1552 & ~n1554 ;
  assign n1556 = ~n1547 & n1554 ;
  assign n1557 = ~n1555 & ~n1556 ;
  assign n1558 = x101 & n1175 ;
  assign n1559 = x100 & n1558 ;
  assign n1560 = n1557 & ~n1559 ;
  assign n1561 = ~n1552 & n1559 ;
  assign n1562 = ~n1560 & ~n1561 ;
  assign n1563 = x97 & n1183 ;
  assign n1564 = x96 & n1563 ;
  assign n1565 = n1562 & ~n1564 ;
  assign n1566 = ~n1557 & n1564 ;
  assign n1567 = ~n1565 & ~n1566 ;
  assign n1568 = x93 & n1191 ;
  assign n1569 = x92 & n1568 ;
  assign n1570 = n1567 & ~n1569 ;
  assign n1571 = ~n1562 & n1569 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = x89 & n1199 ;
  assign n1574 = x88 & n1573 ;
  assign n1575 = n1572 & ~n1574 ;
  assign n1576 = ~n1567 & n1574 ;
  assign n1577 = ~n1575 & ~n1576 ;
  assign n1578 = x85 & n1207 ;
  assign n1579 = x84 & n1578 ;
  assign n1580 = n1577 & ~n1579 ;
  assign n1581 = ~n1572 & n1579 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = x81 & n1215 ;
  assign n1584 = x80 & n1583 ;
  assign n1585 = n1582 & ~n1584 ;
  assign n1586 = ~n1577 & n1584 ;
  assign n1587 = ~n1585 & ~n1586 ;
  assign n1588 = x77 & n1223 ;
  assign n1589 = x76 & n1588 ;
  assign n1590 = n1587 & ~n1589 ;
  assign n1591 = ~n1582 & n1589 ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = x73 & n1231 ;
  assign n1594 = x72 & n1593 ;
  assign n1595 = n1592 & ~n1594 ;
  assign n1596 = ~n1587 & n1594 ;
  assign n1597 = ~n1595 & ~n1596 ;
  assign n1598 = x69 & n1239 ;
  assign n1599 = x68 & n1598 ;
  assign n1600 = n1597 & ~n1599 ;
  assign n1601 = ~n1592 & n1599 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = x65 & n1247 ;
  assign n1604 = x64 & n1603 ;
  assign n1605 = n1602 & ~n1604 ;
  assign n1606 = ~n1597 & n1604 ;
  assign n1607 = ~n1605 & ~n1606 ;
  assign n1608 = x61 & n1255 ;
  assign n1609 = x60 & n1608 ;
  assign n1610 = n1607 & ~n1609 ;
  assign n1611 = ~n1602 & n1609 ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1613 = x57 & n1263 ;
  assign n1614 = x56 & n1613 ;
  assign n1615 = n1612 & ~n1614 ;
  assign n1616 = ~n1607 & n1614 ;
  assign n1617 = ~n1615 & ~n1616 ;
  assign n1618 = x53 & n1271 ;
  assign n1619 = x52 & n1618 ;
  assign n1620 = n1617 & ~n1619 ;
  assign n1621 = ~n1612 & n1619 ;
  assign n1622 = ~n1620 & ~n1621 ;
  assign n1623 = x49 & n1279 ;
  assign n1624 = x48 & n1623 ;
  assign n1625 = n1622 & ~n1624 ;
  assign n1626 = ~n1617 & n1624 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = x45 & n1287 ;
  assign n1629 = x44 & n1628 ;
  assign n1630 = n1627 & ~n1629 ;
  assign n1631 = ~n1622 & n1629 ;
  assign n1632 = ~n1630 & ~n1631 ;
  assign n1633 = x41 & n1295 ;
  assign n1634 = x40 & n1633 ;
  assign n1635 = n1632 & ~n1634 ;
  assign n1636 = ~n1627 & n1634 ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = x37 & n1303 ;
  assign n1639 = x36 & n1638 ;
  assign n1640 = n1637 & ~n1639 ;
  assign n1641 = ~n1632 & n1639 ;
  assign n1642 = ~n1640 & ~n1641 ;
  assign n1643 = x33 & n1311 ;
  assign n1644 = x32 & n1643 ;
  assign n1645 = n1642 & ~n1644 ;
  assign n1646 = ~n1637 & n1644 ;
  assign n1647 = ~n1645 & ~n1646 ;
  assign n1648 = x29 & n1319 ;
  assign n1649 = x28 & n1648 ;
  assign n1650 = n1647 & ~n1649 ;
  assign n1651 = ~n1642 & n1649 ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = x25 & n1327 ;
  assign n1654 = x24 & n1653 ;
  assign n1655 = n1652 & ~n1654 ;
  assign n1656 = ~n1647 & n1654 ;
  assign n1657 = ~n1655 & ~n1656 ;
  assign n1658 = x21 & n1335 ;
  assign n1659 = x20 & n1658 ;
  assign n1660 = n1657 & ~n1659 ;
  assign n1661 = ~n1652 & n1659 ;
  assign n1662 = ~n1660 & ~n1661 ;
  assign n1663 = x17 & n1343 ;
  assign n1664 = x16 & n1663 ;
  assign n1665 = n1662 & ~n1664 ;
  assign n1666 = ~n1657 & n1664 ;
  assign n1667 = ~n1665 & ~n1666 ;
  assign n1668 = x13 & n1351 ;
  assign n1669 = x12 & n1668 ;
  assign n1670 = n1667 & ~n1669 ;
  assign n1671 = ~n1662 & n1669 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = x9 & n1359 ;
  assign n1674 = x8 & n1673 ;
  assign n1675 = n1672 & ~n1674 ;
  assign n1676 = ~n1667 & n1674 ;
  assign n1677 = ~n1675 & ~n1676 ;
  assign n1678 = x5 & n1367 ;
  assign n1679 = x4 & n1678 ;
  assign n1680 = n1677 & ~n1679 ;
  assign n1681 = ~n1672 & n1679 ;
  assign n1682 = ~n1680 & ~n1681 ;
  assign n1685 = n1682 & ~x130 ;
  assign n1686 = ~n1684 & ~n1685 ;
  assign n1687 = n1383 & n1385 ;
  assign n1688 = ~x113 & n903 ;
  assign n1689 = ~x112 & n1387 ;
  assign n1690 = n1688 & n1689 ;
  assign n1691 = ~x107 & n1399 ;
  assign n1692 = ~x106 & n1691 ;
  assign n1693 = ~x105 & n1692 ;
  assign n1694 = ~x104 & n1693 ;
  assign n1695 = n1690 & ~n1694 ;
  assign n1696 = n1687 & ~n1695 ;
  assign n1697 = ~x101 & ~x102 ;
  assign n1698 = ~x100 & n1697 ;
  assign n1699 = ~x99 & n1698 ;
  assign n1700 = ~x98 & n1699 ;
  assign n1701 = ~x97 & n1700 ;
  assign n1702 = ~x96 & n1701 ;
  assign n1703 = n1696 & ~n1702 ;
  assign n1704 = x103 & n1694 ;
  assign n1705 = n1690 & ~n1704 ;
  assign n1706 = n1687 & ~n1705 ;
  assign n1707 = n1702 & n1706 ;
  assign n1708 = ~n1703 & ~n1707 ;
  assign n1709 = ~x91 & n1419 ;
  assign n1710 = ~x90 & n1709 ;
  assign n1711 = ~x89 & n1710 ;
  assign n1712 = ~x88 & n1711 ;
  assign n1713 = n1708 & ~n1712 ;
  assign n1714 = ~n1696 & n1712 ;
  assign n1715 = ~n1713 & ~n1714 ;
  assign n1716 = ~x83 & n1429 ;
  assign n1717 = ~x82 & n1716 ;
  assign n1718 = ~x81 & n1717 ;
  assign n1719 = ~x80 & n1718 ;
  assign n1720 = n1715 & ~n1719 ;
  assign n1721 = ~n1708 & n1719 ;
  assign n1722 = ~n1720 & ~n1721 ;
  assign n1723 = ~x75 & n1439 ;
  assign n1724 = ~x74 & n1723 ;
  assign n1725 = ~x73 & n1724 ;
  assign n1726 = ~x72 & n1725 ;
  assign n1727 = n1722 & ~n1726 ;
  assign n1728 = ~n1715 & n1726 ;
  assign n1729 = ~n1727 & ~n1728 ;
  assign n1730 = ~x67 & n1449 ;
  assign n1731 = ~x66 & n1730 ;
  assign n1732 = ~x65 & n1731 ;
  assign n1733 = ~x64 & n1732 ;
  assign n1734 = n1729 & ~n1733 ;
  assign n1735 = ~n1722 & n1733 ;
  assign n1736 = ~n1734 & ~n1735 ;
  assign n1737 = ~x59 & n1459 ;
  assign n1738 = ~x58 & n1737 ;
  assign n1739 = ~x57 & n1738 ;
  assign n1740 = ~x56 & n1739 ;
  assign n1741 = n1736 & ~n1740 ;
  assign n1742 = ~n1729 & n1740 ;
  assign n1743 = ~n1741 & ~n1742 ;
  assign n1744 = ~x51 & n1469 ;
  assign n1745 = ~x50 & n1744 ;
  assign n1746 = ~x49 & n1745 ;
  assign n1747 = ~x48 & n1746 ;
  assign n1748 = n1743 & ~n1747 ;
  assign n1749 = ~n1736 & n1747 ;
  assign n1750 = ~n1748 & ~n1749 ;
  assign n1751 = ~x43 & n1479 ;
  assign n1752 = ~x42 & n1751 ;
  assign n1753 = ~x41 & n1752 ;
  assign n1754 = ~x40 & n1753 ;
  assign n1755 = n1750 & ~n1754 ;
  assign n1756 = ~n1743 & n1754 ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = ~x35 & n1489 ;
  assign n1759 = ~x34 & n1758 ;
  assign n1760 = ~x33 & n1759 ;
  assign n1761 = ~x32 & n1760 ;
  assign n1762 = n1757 & ~n1761 ;
  assign n1763 = ~n1750 & n1761 ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = ~x27 & n1499 ;
  assign n1766 = ~x26 & n1765 ;
  assign n1767 = ~x25 & n1766 ;
  assign n1768 = ~x24 & n1767 ;
  assign n1769 = n1764 & ~n1768 ;
  assign n1770 = ~n1757 & n1768 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = ~x19 & n1509 ;
  assign n1773 = ~x18 & n1772 ;
  assign n1774 = ~x17 & n1773 ;
  assign n1775 = ~x16 & n1774 ;
  assign n1776 = n1771 & ~n1775 ;
  assign n1777 = ~n1764 & n1775 ;
  assign n1778 = ~n1776 & ~n1777 ;
  assign n1779 = ~x11 & n1519 ;
  assign n1780 = ~x10 & n1779 ;
  assign n1781 = ~x9 & n1780 ;
  assign n1782 = ~x8 & n1781 ;
  assign n1783 = n1778 & ~n1782 ;
  assign n1784 = ~n1771 & n1782 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1886 = ~n1785 & x131 ;
  assign n1786 = n1533 & n1535 ;
  assign n1787 = x113 & n1151 ;
  assign n1788 = x112 & n1537 ;
  assign n1789 = n1787 & n1788 ;
  assign n1790 = x107 & n1549 ;
  assign n1791 = x106 & n1790 ;
  assign n1792 = x105 & n1791 ;
  assign n1793 = x104 & n1792 ;
  assign n1794 = n1789 & ~n1793 ;
  assign n1795 = n1786 & ~n1794 ;
  assign n1796 = x101 & x102 ;
  assign n1797 = x100 & n1796 ;
  assign n1798 = x99 & n1797 ;
  assign n1799 = x98 & n1798 ;
  assign n1800 = x97 & n1799 ;
  assign n1801 = x96 & n1800 ;
  assign n1802 = n1795 & ~n1801 ;
  assign n1803 = ~x103 & n1793 ;
  assign n1804 = n1789 & ~n1803 ;
  assign n1805 = n1786 & ~n1804 ;
  assign n1806 = n1801 & n1805 ;
  assign n1807 = ~n1802 & ~n1806 ;
  assign n1808 = x91 & n1569 ;
  assign n1809 = x90 & n1808 ;
  assign n1810 = x89 & n1809 ;
  assign n1811 = x88 & n1810 ;
  assign n1812 = n1807 & ~n1811 ;
  assign n1813 = ~n1795 & n1811 ;
  assign n1814 = ~n1812 & ~n1813 ;
  assign n1815 = x83 & n1579 ;
  assign n1816 = x82 & n1815 ;
  assign n1817 = x81 & n1816 ;
  assign n1818 = x80 & n1817 ;
  assign n1819 = n1814 & ~n1818 ;
  assign n1820 = ~n1807 & n1818 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1822 = x75 & n1589 ;
  assign n1823 = x74 & n1822 ;
  assign n1824 = x73 & n1823 ;
  assign n1825 = x72 & n1824 ;
  assign n1826 = n1821 & ~n1825 ;
  assign n1827 = ~n1814 & n1825 ;
  assign n1828 = ~n1826 & ~n1827 ;
  assign n1829 = x67 & n1599 ;
  assign n1830 = x66 & n1829 ;
  assign n1831 = x65 & n1830 ;
  assign n1832 = x64 & n1831 ;
  assign n1833 = n1828 & ~n1832 ;
  assign n1834 = ~n1821 & n1832 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = x59 & n1609 ;
  assign n1837 = x58 & n1836 ;
  assign n1838 = x57 & n1837 ;
  assign n1839 = x56 & n1838 ;
  assign n1840 = n1835 & ~n1839 ;
  assign n1841 = ~n1828 & n1839 ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = x51 & n1619 ;
  assign n1844 = x50 & n1843 ;
  assign n1845 = x49 & n1844 ;
  assign n1846 = x48 & n1845 ;
  assign n1847 = n1842 & ~n1846 ;
  assign n1848 = ~n1835 & n1846 ;
  assign n1849 = ~n1847 & ~n1848 ;
  assign n1850 = x43 & n1629 ;
  assign n1851 = x42 & n1850 ;
  assign n1852 = x41 & n1851 ;
  assign n1853 = x40 & n1852 ;
  assign n1854 = n1849 & ~n1853 ;
  assign n1855 = ~n1842 & n1853 ;
  assign n1856 = ~n1854 & ~n1855 ;
  assign n1857 = x35 & n1639 ;
  assign n1858 = x34 & n1857 ;
  assign n1859 = x33 & n1858 ;
  assign n1860 = x32 & n1859 ;
  assign n1861 = n1856 & ~n1860 ;
  assign n1862 = ~n1849 & n1860 ;
  assign n1863 = ~n1861 & ~n1862 ;
  assign n1864 = x27 & n1649 ;
  assign n1865 = x26 & n1864 ;
  assign n1866 = x25 & n1865 ;
  assign n1867 = x24 & n1866 ;
  assign n1868 = n1863 & ~n1867 ;
  assign n1869 = ~n1856 & n1867 ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = x19 & n1659 ;
  assign n1872 = x18 & n1871 ;
  assign n1873 = x17 & n1872 ;
  assign n1874 = x16 & n1873 ;
  assign n1875 = n1870 & ~n1874 ;
  assign n1876 = ~n1863 & n1874 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = x11 & n1669 ;
  assign n1879 = x10 & n1878 ;
  assign n1880 = x9 & n1879 ;
  assign n1881 = x8 & n1880 ;
  assign n1882 = n1877 & ~n1881 ;
  assign n1883 = ~n1870 & n1881 ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1887 = n1884 & ~x131 ;
  assign n1888 = ~n1886 & ~n1887 ;
  assign n1889 = n1687 & n1690 ;
  assign n1890 = ~x99 & n1409 ;
  assign n1891 = ~x98 & n1694 ;
  assign n1892 = ~x97 & n1891 ;
  assign n1893 = ~x96 & n1892 ;
  assign n1894 = n1890 & n1893 ;
  assign n1895 = ~x87 & n1712 ;
  assign n1896 = ~x86 & n1895 ;
  assign n1897 = ~x85 & n1896 ;
  assign n1898 = ~x84 & n1897 ;
  assign n1899 = ~x83 & n1898 ;
  assign n1900 = ~x82 & n1899 ;
  assign n1901 = ~x81 & n1900 ;
  assign n1902 = ~x80 & n1901 ;
  assign n1903 = n1894 & ~n1902 ;
  assign n1904 = n1889 & ~n1903 ;
  assign n1905 = ~x77 & ~x78 ;
  assign n1906 = ~x76 & n1905 ;
  assign n1907 = ~x75 & n1906 ;
  assign n1908 = ~x74 & n1907 ;
  assign n1909 = ~x73 & n1908 ;
  assign n1910 = ~x72 & n1909 ;
  assign n1911 = ~x71 & n1910 ;
  assign n1912 = ~x70 & n1911 ;
  assign n1913 = ~x69 & n1912 ;
  assign n1914 = ~x68 & n1913 ;
  assign n1915 = ~x67 & n1914 ;
  assign n1916 = ~x66 & n1915 ;
  assign n1917 = ~x65 & n1916 ;
  assign n1918 = ~x64 & n1917 ;
  assign n1919 = n1904 & ~n1918 ;
  assign n1920 = x79 & n1902 ;
  assign n1921 = n1894 & ~n1920 ;
  assign n1922 = n1889 & ~n1921 ;
  assign n1923 = n1918 & n1922 ;
  assign n1924 = ~n1919 & ~n1923 ;
  assign n1925 = ~x55 & n1740 ;
  assign n1926 = ~x54 & n1925 ;
  assign n1927 = ~x53 & n1926 ;
  assign n1928 = ~x52 & n1927 ;
  assign n1929 = ~x51 & n1928 ;
  assign n1930 = ~x50 & n1929 ;
  assign n1931 = ~x49 & n1930 ;
  assign n1932 = ~x48 & n1931 ;
  assign n1933 = n1924 & ~n1932 ;
  assign n1934 = ~n1904 & n1932 ;
  assign n1935 = ~n1933 & ~n1934 ;
  assign n1936 = ~x39 & n1754 ;
  assign n1937 = ~x38 & n1936 ;
  assign n1938 = ~x37 & n1937 ;
  assign n1939 = ~x36 & n1938 ;
  assign n1940 = ~x35 & n1939 ;
  assign n1941 = ~x34 & n1940 ;
  assign n1942 = ~x33 & n1941 ;
  assign n1943 = ~x32 & n1942 ;
  assign n1944 = n1935 & ~n1943 ;
  assign n1945 = ~n1924 & n1943 ;
  assign n1946 = ~n1944 & ~n1945 ;
  assign n1947 = ~x23 & n1768 ;
  assign n1948 = ~x22 & n1947 ;
  assign n1949 = ~x21 & n1948 ;
  assign n1950 = ~x20 & n1949 ;
  assign n1951 = ~x19 & n1950 ;
  assign n1952 = ~x18 & n1951 ;
  assign n1953 = ~x17 & n1952 ;
  assign n1954 = ~x16 & n1953 ;
  assign n1955 = n1946 & ~n1954 ;
  assign n1956 = ~n1935 & n1954 ;
  assign n1957 = ~n1955 & ~n1956 ;
  assign n2028 = ~n1957 & x132 ;
  assign n1958 = n1786 & n1789 ;
  assign n1959 = x99 & n1559 ;
  assign n1960 = x98 & n1793 ;
  assign n1961 = x97 & n1960 ;
  assign n1962 = x96 & n1961 ;
  assign n1963 = n1959 & n1962 ;
  assign n1964 = x87 & n1811 ;
  assign n1965 = x86 & n1964 ;
  assign n1966 = x85 & n1965 ;
  assign n1967 = x84 & n1966 ;
  assign n1968 = x83 & n1967 ;
  assign n1969 = x82 & n1968 ;
  assign n1970 = x81 & n1969 ;
  assign n1971 = x80 & n1970 ;
  assign n1972 = n1963 & ~n1971 ;
  assign n1973 = n1958 & ~n1972 ;
  assign n1974 = x77 & x78 ;
  assign n1975 = x76 & n1974 ;
  assign n1976 = x75 & n1975 ;
  assign n1977 = x74 & n1976 ;
  assign n1978 = x73 & n1977 ;
  assign n1979 = x72 & n1978 ;
  assign n1980 = x71 & n1979 ;
  assign n1981 = x70 & n1980 ;
  assign n1982 = x69 & n1981 ;
  assign n1983 = x68 & n1982 ;
  assign n1984 = x67 & n1983 ;
  assign n1985 = x66 & n1984 ;
  assign n1986 = x65 & n1985 ;
  assign n1987 = x64 & n1986 ;
  assign n1988 = n1973 & ~n1987 ;
  assign n1989 = ~x79 & n1971 ;
  assign n1990 = n1963 & ~n1989 ;
  assign n1991 = n1958 & ~n1990 ;
  assign n1992 = n1987 & n1991 ;
  assign n1993 = ~n1988 & ~n1992 ;
  assign n1994 = x55 & n1839 ;
  assign n1995 = x54 & n1994 ;
  assign n1996 = x53 & n1995 ;
  assign n1997 = x52 & n1996 ;
  assign n1998 = x51 & n1997 ;
  assign n1999 = x50 & n1998 ;
  assign n2000 = x49 & n1999 ;
  assign n2001 = x48 & n2000 ;
  assign n2002 = n1993 & ~n2001 ;
  assign n2003 = ~n1973 & n2001 ;
  assign n2004 = ~n2002 & ~n2003 ;
  assign n2005 = x39 & n1853 ;
  assign n2006 = x38 & n2005 ;
  assign n2007 = x37 & n2006 ;
  assign n2008 = x36 & n2007 ;
  assign n2009 = x35 & n2008 ;
  assign n2010 = x34 & n2009 ;
  assign n2011 = x33 & n2010 ;
  assign n2012 = x32 & n2011 ;
  assign n2013 = n2004 & ~n2012 ;
  assign n2014 = ~n1993 & n2012 ;
  assign n2015 = ~n2013 & ~n2014 ;
  assign n2016 = x23 & n1867 ;
  assign n2017 = x22 & n2016 ;
  assign n2018 = x21 & n2017 ;
  assign n2019 = x20 & n2018 ;
  assign n2020 = x19 & n2019 ;
  assign n2021 = x18 & n2020 ;
  assign n2022 = x17 & n2021 ;
  assign n2023 = x16 & n2022 ;
  assign n2024 = n2015 & ~n2023 ;
  assign n2025 = ~n2004 & n2023 ;
  assign n2026 = ~n2024 & ~n2025 ;
  assign n2029 = n2026 & ~x132 ;
  assign n2030 = ~n2028 & ~n2029 ;
  assign n2031 = n1889 & n1894 ;
  assign n2032 = ~x71 & n1726 ;
  assign n2033 = ~x70 & n1902 ;
  assign n2034 = ~x69 & n2033 ;
  assign n2035 = ~x68 & n2034 ;
  assign n2036 = ~x67 & n2035 ;
  assign n2037 = ~x66 & n2036 ;
  assign n2038 = ~x65 & n2037 ;
  assign n2039 = ~x64 & n2038 ;
  assign n2040 = n2032 & n2039 ;
  assign n2041 = ~x47 & n1932 ;
  assign n2042 = ~x46 & n2041 ;
  assign n2043 = ~x45 & n2042 ;
  assign n2044 = ~x44 & n2043 ;
  assign n2045 = ~x43 & n2044 ;
  assign n2046 = ~x42 & n2045 ;
  assign n2047 = ~x41 & n2046 ;
  assign n2048 = ~x40 & n2047 ;
  assign n2049 = ~x39 & n2048 ;
  assign n2050 = ~x38 & n2049 ;
  assign n2051 = ~x37 & n2050 ;
  assign n2052 = ~x36 & n2051 ;
  assign n2053 = ~x35 & n2052 ;
  assign n2054 = ~x34 & n2053 ;
  assign n2055 = ~x33 & n2054 ;
  assign n2056 = ~x32 & n2055 ;
  assign n2057 = n2040 & ~n2056 ;
  assign n2058 = n2031 & ~n2057 ;
  assign n2088 = ~n2058 & x133 ;
  assign n2059 = n1958 & n1963 ;
  assign n2060 = x71 & n1825 ;
  assign n2061 = x70 & n1971 ;
  assign n2062 = x69 & n2061 ;
  assign n2063 = x68 & n2062 ;
  assign n2064 = x67 & n2063 ;
  assign n2065 = x66 & n2064 ;
  assign n2066 = x65 & n2065 ;
  assign n2067 = x64 & n2066 ;
  assign n2068 = n2060 & n2067 ;
  assign n2069 = x47 & n2001 ;
  assign n2070 = x46 & n2069 ;
  assign n2071 = x45 & n2070 ;
  assign n2072 = x44 & n2071 ;
  assign n2073 = x43 & n2072 ;
  assign n2074 = x42 & n2073 ;
  assign n2075 = x41 & n2074 ;
  assign n2076 = x40 & n2075 ;
  assign n2077 = x39 & n2076 ;
  assign n2078 = x38 & n2077 ;
  assign n2079 = x37 & n2078 ;
  assign n2080 = x36 & n2079 ;
  assign n2081 = x35 & n2080 ;
  assign n2082 = x34 & n2081 ;
  assign n2083 = x33 & n2082 ;
  assign n2084 = x32 & n2083 ;
  assign n2085 = n2068 & ~n2084 ;
  assign n2086 = n2059 & ~n2085 ;
  assign n2089 = n2086 & ~x133 ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2091 = n2031 & n2040 ;
  assign n2094 = ~n2091 & x134 ;
  assign n2092 = n2059 & n2068 ;
  assign n2095 = n2092 & ~x134 ;
  assign n2096 = ~n2094 & ~n2095 ;
  assign n2097 = ~x0 & n2091 ;
  assign n2098 = n1782 & n2097 ;
  assign n2099 = ~x3 & n2098 ;
  assign n2100 = ~x2 & n2099 ;
  assign n2101 = n1954 & n2056 ;
  assign n2102 = n1529 & n2101 ;
  assign n2103 = ~x1 & n2102 ;
  assign n2104 = n2100 & n2103 ;
  assign n2114 = ~n2104 & x135 ;
  assign n2105 = x0 & n2092 ;
  assign n2106 = n1881 & n2105 ;
  assign n2107 = x3 & n2106 ;
  assign n2108 = x2 & n2107 ;
  assign n2109 = n2023 & n2084 ;
  assign n2110 = n1679 & n2109 ;
  assign n2111 = x1 & n2110 ;
  assign n2112 = n2108 & n2111 ;
  assign n2115 = n2112 & ~x135 ;
  assign n2116 = ~n2114 & ~n2115 ;
  assign y0 = ~n882 ;
  assign y1 = ~n1382 ;
  assign y2 = ~n1686 ;
  assign y3 = ~n1888 ;
  assign y4 = ~n2030 ;
  assign y5 = ~n2090 ;
  assign y6 = ~n2096 ;
  assign y7 = ~n2116 ;
endmodule
