module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n578 , n579 , n580 ;
  assign n61 = ~x9 & ~x10 ;
  assign n62 = x9 & x10 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = x11 & ~n61 ;
  assign n65 = ~x11 & n61 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = ~x12 & ~n64 ;
  assign n68 = x12 & n64 ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = ~x13 & n67 ;
  assign n71 = x13 & ~n67 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = x14 & ~n70 ;
  assign n74 = ~x14 & n70 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = x15 & ~n73 ;
  assign n77 = ~x15 & n73 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = x15 & n73 ;
  assign n80 = ~x16 & ~n79 ;
  assign n81 = x16 & n79 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = x17 & ~n80 ;
  assign n84 = ~x17 & n80 ;
  assign n85 = ~n83 & ~n84 ;
  assign n86 = ~x18 & ~n83 ;
  assign n87 = x18 & n83 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = x19 & ~n86 ;
  assign n90 = ~x19 & n86 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = x20 & ~n89 ;
  assign n93 = ~x20 & n89 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = x20 & n89 ;
  assign n96 = ~x21 & ~n95 ;
  assign n97 = x21 & n95 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = ~x22 & n96 ;
  assign n100 = x22 & ~n96 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = x23 & ~n99 ;
  assign n103 = ~x23 & n99 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = x24 & ~n102 ;
  assign n106 = ~x24 & n102 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = x24 & n102 ;
  assign n109 = x25 & ~n108 ;
  assign n110 = ~x25 & n108 ;
  assign n111 = ~n109 & ~n110 ;
  assign n112 = x25 & n108 ;
  assign n113 = ~x26 & ~n112 ;
  assign n114 = x26 & n112 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = x27 & ~n113 ;
  assign n117 = ~x27 & n113 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = x28 & ~n116 ;
  assign n120 = ~x28 & n116 ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = x28 & n116 ;
  assign n123 = ~x29 & n122 ;
  assign n124 = x29 & ~n122 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = ~x9 & ~n125 ;
  assign n127 = ~n121 & n126 ;
  assign n128 = n118 & n127 ;
  assign n129 = ~n115 & n128 ;
  assign n130 = ~n111 & n129 ;
  assign n131 = ~n107 & n130 ;
  assign n132 = n104 & n131 ;
  assign n133 = ~n101 & n132 ;
  assign n134 = ~n98 & n133 ;
  assign n135 = ~n94 & n134 ;
  assign n136 = n91 & n135 ;
  assign n137 = ~n88 & n136 ;
  assign n138 = n85 & n137 ;
  assign n139 = ~n82 & n138 ;
  assign n140 = ~n78 & n139 ;
  assign n141 = n75 & n140 ;
  assign n142 = ~n72 & n141 ;
  assign n143 = ~n69 & n142 ;
  assign n144 = n66 & n143 ;
  assign n145 = ~n63 & n144 ;
  assign n146 = x8 & n145 ;
  assign n147 = x7 & n146 ;
  assign n148 = x6 & n147 ;
  assign n149 = x5 & n148 ;
  assign n150 = x4 & n149 ;
  assign n151 = x3 & n150 ;
  assign n152 = x2 & n151 ;
  assign n153 = x1 & n152 ;
  assign n154 = x0 & n153 ;
  assign n155 = x29 & n122 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = ~x1 & ~x2 ;
  assign n158 = ~x3 & n157 ;
  assign n159 = ~x4 & n158 ;
  assign n160 = ~x5 & n159 ;
  assign n161 = ~x6 & n160 ;
  assign n162 = ~x7 & n161 ;
  assign n163 = ~x8 & n162 ;
  assign n164 = n63 & n163 ;
  assign n165 = ~n66 & n164 ;
  assign n166 = n69 & n165 ;
  assign n167 = n72 & n166 ;
  assign n168 = ~n75 & n167 ;
  assign n169 = n78 & n168 ;
  assign n170 = n82 & n169 ;
  assign n171 = ~n85 & n170 ;
  assign n172 = n88 & n171 ;
  assign n173 = ~n91 & n172 ;
  assign n174 = n94 & n173 ;
  assign n175 = n98 & n174 ;
  assign n176 = n101 & n175 ;
  assign n177 = ~n104 & n176 ;
  assign n178 = n107 & n177 ;
  assign n179 = n111 & n178 ;
  assign n180 = n115 & n179 ;
  assign n181 = ~n118 & n180 ;
  assign n182 = n121 & n181 ;
  assign n183 = x9 & n182 ;
  assign n184 = n155 & ~n183 ;
  assign n185 = ~n156 & ~n184 ;
  assign n309 = ~n185 & x60 ;
  assign n186 = ~x11 & ~n62 ;
  assign n187 = x11 & n62 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = x12 & ~n186 ;
  assign n190 = ~x12 & n186 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = x13 & n189 ;
  assign n193 = ~x13 & ~n189 ;
  assign n194 = ~n192 & ~n193 ;
  assign n195 = ~x14 & ~n192 ;
  assign n196 = x14 & n192 ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = ~x15 & ~n195 ;
  assign n199 = x15 & n195 ;
  assign n200 = ~n198 & ~n199 ;
  assign n201 = ~x15 & n195 ;
  assign n202 = x16 & ~n201 ;
  assign n203 = ~x16 & n201 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = ~x17 & ~n202 ;
  assign n206 = x17 & n202 ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = x18 & ~n205 ;
  assign n209 = ~x18 & n205 ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = ~x19 & ~n208 ;
  assign n212 = x19 & n208 ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = ~x20 & ~n211 ;
  assign n215 = x20 & n211 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = ~x20 & n211 ;
  assign n218 = x21 & ~n217 ;
  assign n219 = ~x21 & n217 ;
  assign n220 = ~n218 & ~n219 ;
  assign n221 = x22 & n218 ;
  assign n222 = ~x22 & ~n218 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = ~x23 & ~n221 ;
  assign n225 = x23 & n221 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = ~x24 & ~n224 ;
  assign n228 = x24 & n224 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = ~x24 & n224 ;
  assign n231 = ~x25 & ~n230 ;
  assign n232 = x25 & n230 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = ~x25 & n230 ;
  assign n235 = x26 & ~n234 ;
  assign n236 = ~x26 & n234 ;
  assign n237 = ~n235 & ~n236 ;
  assign n238 = ~x27 & ~n235 ;
  assign n239 = x27 & n235 ;
  assign n240 = ~n238 & ~n239 ;
  assign n241 = ~x28 & ~n238 ;
  assign n242 = x28 & n238 ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = ~x28 & n238 ;
  assign n245 = x29 & n244 ;
  assign n246 = ~x29 & ~n244 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = x9 & ~n247 ;
  assign n249 = ~n243 & n248 ;
  assign n250 = n240 & n249 ;
  assign n251 = ~n237 & n250 ;
  assign n252 = ~n233 & n251 ;
  assign n253 = ~n229 & n252 ;
  assign n254 = n226 & n253 ;
  assign n255 = ~n223 & n254 ;
  assign n256 = ~n220 & n255 ;
  assign n257 = ~n216 & n256 ;
  assign n258 = n213 & n257 ;
  assign n259 = ~n210 & n258 ;
  assign n260 = n207 & n259 ;
  assign n261 = ~n204 & n260 ;
  assign n262 = ~n200 & n261 ;
  assign n263 = n197 & n262 ;
  assign n264 = ~n194 & n263 ;
  assign n265 = ~n191 & n264 ;
  assign n266 = n188 & n265 ;
  assign n267 = ~n63 & n266 ;
  assign n268 = ~x8 & n267 ;
  assign n269 = ~x7 & n268 ;
  assign n270 = ~x6 & n269 ;
  assign n271 = ~x5 & n270 ;
  assign n272 = ~x4 & n271 ;
  assign n273 = ~x3 & n272 ;
  assign n274 = ~x2 & n273 ;
  assign n275 = ~x1 & n274 ;
  assign n276 = ~x0 & n275 ;
  assign n277 = ~x29 & n244 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = x1 & x2 ;
  assign n280 = x3 & n279 ;
  assign n281 = x4 & n280 ;
  assign n282 = x5 & n281 ;
  assign n283 = x6 & n282 ;
  assign n284 = x7 & n283 ;
  assign n285 = x8 & n284 ;
  assign n286 = n63 & n285 ;
  assign n287 = ~n188 & n286 ;
  assign n288 = n191 & n287 ;
  assign n289 = n194 & n288 ;
  assign n290 = ~n197 & n289 ;
  assign n291 = n200 & n290 ;
  assign n292 = n204 & n291 ;
  assign n293 = ~n207 & n292 ;
  assign n294 = n210 & n293 ;
  assign n295 = ~n213 & n294 ;
  assign n296 = n216 & n295 ;
  assign n297 = n220 & n296 ;
  assign n298 = n223 & n297 ;
  assign n299 = ~n226 & n298 ;
  assign n300 = n229 & n299 ;
  assign n301 = n233 & n300 ;
  assign n302 = n237 & n301 ;
  assign n303 = ~n240 & n302 ;
  assign n304 = n243 & n303 ;
  assign n305 = ~x9 & n304 ;
  assign n306 = n277 & ~n305 ;
  assign n307 = ~n278 & ~n306 ;
  assign n310 = n307 & ~x60 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = ~x39 & ~x40 ;
  assign n313 = x41 & ~n312 ;
  assign n314 = ~x42 & ~n313 ;
  assign n315 = ~x43 & n314 ;
  assign n316 = x44 & ~n315 ;
  assign n317 = x45 & n316 ;
  assign n318 = ~x46 & ~n317 ;
  assign n319 = x47 & ~n318 ;
  assign n320 = ~x48 & ~n319 ;
  assign n321 = x49 & ~n320 ;
  assign n322 = x50 & n321 ;
  assign n323 = ~x51 & ~n322 ;
  assign n324 = ~x52 & n323 ;
  assign n325 = x53 & ~n324 ;
  assign n326 = x54 & n325 ;
  assign n327 = x55 & n326 ;
  assign n328 = ~x56 & ~n327 ;
  assign n329 = x57 & ~n328 ;
  assign n330 = x58 & n329 ;
  assign n331 = x59 & n330 ;
  assign n332 = x0 & ~n331 ;
  assign n333 = ~x0 & ~x30 ;
  assign n334 = n331 & ~n333 ;
  assign n335 = x39 & x40 ;
  assign n336 = ~n312 & ~n335 ;
  assign n337 = ~x41 & n312 ;
  assign n338 = ~n313 & ~n337 ;
  assign n339 = x42 & n313 ;
  assign n340 = ~n314 & ~n339 ;
  assign n341 = x43 & ~n314 ;
  assign n342 = ~n315 & ~n341 ;
  assign n343 = ~x44 & n315 ;
  assign n344 = ~n316 & ~n343 ;
  assign n345 = x45 & ~n316 ;
  assign n346 = ~x45 & n316 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = x46 & n317 ;
  assign n349 = ~n318 & ~n348 ;
  assign n350 = ~x47 & n318 ;
  assign n351 = ~n319 & ~n350 ;
  assign n352 = x48 & n319 ;
  assign n353 = ~n320 & ~n352 ;
  assign n354 = ~x49 & n320 ;
  assign n355 = ~n321 & ~n354 ;
  assign n356 = x50 & ~n321 ;
  assign n357 = ~x50 & n321 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = x51 & n322 ;
  assign n360 = ~n323 & ~n359 ;
  assign n361 = x52 & ~n323 ;
  assign n362 = ~n324 & ~n361 ;
  assign n363 = ~x53 & n324 ;
  assign n364 = ~n325 & ~n363 ;
  assign n365 = x54 & ~n325 ;
  assign n366 = ~x54 & n325 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = x55 & ~n326 ;
  assign n369 = ~x55 & n326 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = x56 & n327 ;
  assign n372 = ~n328 & ~n371 ;
  assign n373 = ~x57 & n328 ;
  assign n374 = ~n329 & ~n373 ;
  assign n375 = x58 & ~n329 ;
  assign n376 = ~x58 & n329 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = x30 & ~x39 ;
  assign n379 = x59 & n378 ;
  assign n380 = ~n377 & n379 ;
  assign n381 = n374 & n380 ;
  assign n382 = ~n372 & n381 ;
  assign n383 = ~n370 & n382 ;
  assign n384 = ~n367 & n383 ;
  assign n385 = n364 & n384 ;
  assign n386 = ~n362 & n385 ;
  assign n387 = ~n360 & n386 ;
  assign n388 = ~n358 & n387 ;
  assign n389 = n355 & n388 ;
  assign n390 = ~n353 & n389 ;
  assign n391 = n351 & n390 ;
  assign n392 = ~n349 & n391 ;
  assign n393 = ~n347 & n392 ;
  assign n394 = n344 & n393 ;
  assign n395 = ~n342 & n394 ;
  assign n396 = ~n340 & n395 ;
  assign n397 = n338 & n396 ;
  assign n398 = ~n336 & n397 ;
  assign n399 = x38 & n398 ;
  assign n400 = x37 & n399 ;
  assign n401 = x36 & n400 ;
  assign n402 = x35 & n401 ;
  assign n403 = x34 & n402 ;
  assign n404 = x33 & n403 ;
  assign n405 = x32 & n404 ;
  assign n406 = x31 & n405 ;
  assign n407 = ~x31 & ~x32 ;
  assign n408 = ~x33 & n407 ;
  assign n409 = ~x34 & n408 ;
  assign n410 = ~x35 & n409 ;
  assign n411 = ~x36 & n410 ;
  assign n412 = ~x37 & n411 ;
  assign n413 = ~x38 & n412 ;
  assign n414 = n336 & n413 ;
  assign n415 = ~n338 & n414 ;
  assign n416 = n340 & n415 ;
  assign n417 = n342 & n416 ;
  assign n418 = ~n344 & n417 ;
  assign n419 = n347 & n418 ;
  assign n420 = n349 & n419 ;
  assign n421 = ~n351 & n420 ;
  assign n422 = n353 & n421 ;
  assign n423 = ~n355 & n422 ;
  assign n424 = n358 & n423 ;
  assign n425 = n360 & n424 ;
  assign n426 = n362 & n425 ;
  assign n427 = ~n364 & n426 ;
  assign n428 = n367 & n427 ;
  assign n429 = n370 & n428 ;
  assign n430 = n372 & n429 ;
  assign n431 = ~n374 & n430 ;
  assign n432 = n377 & n431 ;
  assign n433 = x39 & n432 ;
  assign n434 = n331 & ~n433 ;
  assign n435 = ~n406 & ~n434 ;
  assign n436 = ~n334 & n435 ;
  assign n437 = ~n156 & ~n436 ;
  assign n438 = ~n332 & n437 ;
  assign n439 = ~n184 & ~n438 ;
  assign n566 = n439 & x61 ;
  assign n440 = ~x41 & ~n335 ;
  assign n441 = x42 & ~n440 ;
  assign n442 = x43 & n441 ;
  assign n443 = ~x44 & ~n442 ;
  assign n444 = ~x45 & n443 ;
  assign n445 = x46 & ~n444 ;
  assign n446 = ~x47 & ~n445 ;
  assign n447 = x48 & ~n446 ;
  assign n448 = ~x49 & ~n447 ;
  assign n449 = ~x50 & n448 ;
  assign n450 = x51 & ~n449 ;
  assign n451 = x52 & n450 ;
  assign n452 = ~x53 & ~n451 ;
  assign n453 = ~x54 & n452 ;
  assign n454 = ~x55 & n453 ;
  assign n455 = x56 & ~n454 ;
  assign n456 = ~x57 & ~n455 ;
  assign n457 = ~x58 & n456 ;
  assign n458 = ~x59 & n457 ;
  assign n459 = ~x0 & ~n458 ;
  assign n460 = x0 & x30 ;
  assign n461 = n458 & ~n460 ;
  assign n462 = x41 & n335 ;
  assign n463 = ~n440 & ~n462 ;
  assign n464 = ~x42 & n440 ;
  assign n465 = ~n441 & ~n464 ;
  assign n466 = ~x43 & ~n441 ;
  assign n467 = ~n442 & ~n466 ;
  assign n468 = x44 & n442 ;
  assign n469 = ~n443 & ~n468 ;
  assign n470 = ~x45 & ~n443 ;
  assign n471 = x45 & n443 ;
  assign n472 = ~n470 & ~n471 ;
  assign n473 = ~x46 & n444 ;
  assign n474 = ~n445 & ~n473 ;
  assign n475 = x47 & n445 ;
  assign n476 = ~n446 & ~n475 ;
  assign n477 = ~x48 & n446 ;
  assign n478 = ~n447 & ~n477 ;
  assign n479 = x49 & n447 ;
  assign n480 = ~n448 & ~n479 ;
  assign n481 = ~x50 & ~n448 ;
  assign n482 = x50 & n448 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = ~x51 & n449 ;
  assign n485 = ~n450 & ~n484 ;
  assign n486 = ~x52 & ~n450 ;
  assign n487 = ~n451 & ~n486 ;
  assign n488 = x53 & n451 ;
  assign n489 = ~n452 & ~n488 ;
  assign n490 = ~x54 & ~n452 ;
  assign n491 = x54 & n452 ;
  assign n492 = ~n490 & ~n491 ;
  assign n493 = ~x55 & ~n453 ;
  assign n494 = x55 & n453 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = ~x56 & n454 ;
  assign n497 = ~n455 & ~n496 ;
  assign n498 = x57 & n455 ;
  assign n499 = ~n456 & ~n498 ;
  assign n500 = ~x58 & ~n456 ;
  assign n501 = x58 & n456 ;
  assign n502 = ~n500 & ~n501 ;
  assign n503 = ~x30 & x39 ;
  assign n504 = ~x59 & n503 ;
  assign n505 = ~n502 & n504 ;
  assign n506 = n499 & n505 ;
  assign n507 = ~n497 & n506 ;
  assign n508 = ~n495 & n507 ;
  assign n509 = ~n492 & n508 ;
  assign n510 = n489 & n509 ;
  assign n511 = ~n487 & n510 ;
  assign n512 = ~n485 & n511 ;
  assign n513 = ~n483 & n512 ;
  assign n514 = n480 & n513 ;
  assign n515 = ~n478 & n514 ;
  assign n516 = n476 & n515 ;
  assign n517 = ~n474 & n516 ;
  assign n518 = ~n472 & n517 ;
  assign n519 = n469 & n518 ;
  assign n520 = ~n467 & n519 ;
  assign n521 = ~n465 & n520 ;
  assign n522 = n463 & n521 ;
  assign n523 = ~n336 & n522 ;
  assign n524 = ~x38 & n523 ;
  assign n525 = ~x37 & n524 ;
  assign n526 = ~x36 & n525 ;
  assign n527 = ~x35 & n526 ;
  assign n528 = ~x34 & n527 ;
  assign n529 = ~x33 & n528 ;
  assign n530 = ~x32 & n529 ;
  assign n531 = ~x31 & n530 ;
  assign n532 = x31 & x32 ;
  assign n533 = x33 & n532 ;
  assign n534 = x34 & n533 ;
  assign n535 = x35 & n534 ;
  assign n536 = x36 & n535 ;
  assign n537 = x37 & n536 ;
  assign n538 = x38 & n537 ;
  assign n539 = n336 & n538 ;
  assign n540 = ~n463 & n539 ;
  assign n541 = n465 & n540 ;
  assign n542 = n467 & n541 ;
  assign n543 = ~n469 & n542 ;
  assign n544 = n472 & n543 ;
  assign n545 = n474 & n544 ;
  assign n546 = ~n476 & n545 ;
  assign n547 = n478 & n546 ;
  assign n548 = ~n480 & n547 ;
  assign n549 = n483 & n548 ;
  assign n550 = n485 & n549 ;
  assign n551 = n487 & n550 ;
  assign n552 = ~n489 & n551 ;
  assign n553 = n492 & n552 ;
  assign n554 = n495 & n553 ;
  assign n555 = n497 & n554 ;
  assign n556 = ~n499 & n555 ;
  assign n557 = n502 & n556 ;
  assign n558 = ~x39 & n557 ;
  assign n559 = n458 & ~n558 ;
  assign n560 = ~n531 & ~n559 ;
  assign n561 = ~n461 & n560 ;
  assign n562 = ~n278 & ~n561 ;
  assign n563 = ~n459 & n562 ;
  assign n564 = ~n306 & ~n563 ;
  assign n567 = ~n564 & ~x61 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = x0 & n331 ;
  assign n570 = x30 & n569 ;
  assign n571 = ~n434 & ~n570 ;
  assign n572 = n185 & ~n571 ;
  assign n578 = n572 & x62 ;
  assign n573 = ~x0 & n458 ;
  assign n574 = ~x30 & n573 ;
  assign n575 = ~n559 & ~n574 ;
  assign n576 = n307 & ~n575 ;
  assign n579 = ~n576 & ~x62 ;
  assign n580 = ~n578 & ~n579 ;
  assign y0 = ~n311 ;
  assign y1 = ~n568 ;
  assign y2 = ~n580 ;
  assign y3 = ~x63 ;
  assign y4 = ~x64 ;
  assign y5 = ~x65 ;
  assign y6 = ~x66 ;
  assign y7 = ~x67 ;
  assign y8 = ~x68 ;
  assign y9 = ~x69 ;
  assign y10 = ~x70 ;
  assign y11 = ~x71 ;
  assign y12 = ~x72 ;
  assign y13 = ~x73 ;
  assign y14 = ~x74 ;
  assign y15 = ~x75 ;
  assign y16 = ~x76 ;
  assign y17 = ~x77 ;
  assign y18 = ~x78 ;
  assign y19 = ~x79 ;
  assign y20 = ~x80 ;
  assign y21 = ~x81 ;
  assign y22 = ~x82 ;
  assign y23 = ~x83 ;
  assign y24 = ~x84 ;
  assign y25 = ~x85 ;
  assign y26 = ~x86 ;
  assign y27 = ~x87 ;
  assign y28 = ~x88 ;
  assign y29 = ~x89 ;
endmodule
