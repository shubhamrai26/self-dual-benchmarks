module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n84 , n85 , n86 , n87 , n88 , n90 , n91 , n92 , n93 , n94 , n96 , n97 , n98 , n99 , n100 , n102 , n103 , n104 , n105 , n106 , n108 , n109 , n110 , n111 , n112 , n114 , n115 , n116 , n117 , n118 , n120 , n121 , n122 , n123 , n124 , n126 , n127 , n128 , n129 , n130 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n142 , n143 , n144 , n145 , n146 , n148 , n149 , n150 , n151 , n152 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , n163 , n164 , n166 , n167 , n168 , n169 , n170 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n182 , n184 , n185 , n186 , n187 , n188 , n190 , n191 , n192 , n193 , n194 , n196 , n197 , n198 , n199 , n200 , n202 , n203 , n204 , n205 , n206 , n208 , n209 , n210 , n211 , n212 , n214 , n215 , n216 , n217 , n218 , n220 , n221 , n222 , n223 , n224 , n226 , n227 , n228 , n229 , n230 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n240 , n241 , n242 , n243 , n244 , n246 , n247 , n248 , n249 , n250 , n252 , n253 , n254 , n255 , n256 , n258 , n259 , n260 , n261 , n262 , n264 , n265 , n266 , n267 , n268 , n270 , n271 , n272 , n273 , n274 , n276 , n277 , n278 , n279 , n280 , n282 , n283 , n284 , n285 , n286 , n288 , n289 , n290 , n291 , n292 , n294 , n295 , n296 , n297 , n298 , n300 , n301 , n302 , n303 , n304 , n306 , n307 , n308 , n309 , n310 , n312 , n313 , n314 , n315 , n316 , n318 , n319 , n320 , n321 , n322 , n324 , n325 , n326 , n327 , n328 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n338 , n339 , n340 , n341 , n342 , n344 , n345 , n346 , n347 , n348 , n350 , n351 , n352 , n353 , n354 , n356 , n357 , n358 , n359 , n360 , n362 , n363 , n364 , n365 , n366 , n368 , n369 , n370 , n371 , n372 , n374 , n375 , n376 , n377 , n378 , n380 , n381 , n382 , n383 , n384 , n386 , n387 , n388 , n389 , n390 , n392 , n393 , n394 , n395 , n396 , n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , n407 , n408 , n410 , n411 , n412 , n413 , n414 , n416 , n417 , n418 , n419 , n420 , n422 , n423 , n424 , n425 , n426 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n438 , n439 , n440 , n441 , n442 , n444 , n445 , n446 , n447 , n448 , n450 , n451 , n452 , n453 , n454 , n456 , n457 , n458 , n459 , n460 , n462 , n463 , n464 , n465 , n466 , n468 , n469 , n470 , n471 , n472 , n474 , n475 , n476 , n477 , n478 , n480 , n481 , n482 , n483 , n484 , n486 , n487 , n488 , n489 , n490 , n492 , n493 , n494 , n495 , n496 , n498 , n499 , n500 , n501 , n502 , n504 , n505 , n506 , n507 , n508 , n510 , n511 , n512 , n513 , n514 , n516 , n517 , n518 , n519 , n520 , n522 , n523 , n524 , n525 , n526 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n536 , n537 , n538 , n539 , n540 , n542 , n543 , n544 , n545 , n546 , n548 , n549 , n550 , n551 , n552 , n554 , n555 , n556 , n557 , n558 , n560 , n561 , n562 , n563 , n564 , n566 , n567 , n568 , n569 , n570 , n572 , n573 , n574 , n575 , n576 , n578 , n579 , n580 , n581 , n582 , n584 , n585 , n586 , n587 , n588 , n590 , n591 , n592 , n593 , n594 , n596 , n597 , n598 , n599 , n600 , n602 , n603 , n604 , n605 , n606 , n608 , n609 , n610 , n611 , n612 , n614 , n615 , n616 , n617 , n618 , n620 , n621 , n622 , n623 , n624 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n634 , n635 , n636 , n637 , n638 , n640 , n641 , n642 , n643 , n644 , n646 , n647 , n648 , n649 , n650 , n652 , n653 , n654 , n655 , n656 , n658 , n659 , n660 , n661 , n662 , n664 , n665 , n666 , n667 , n668 , n670 , n671 , n672 , n673 , n674 , n676 , n677 , n678 , n679 , n680 , n682 , n683 , n684 , n685 , n686 , n688 , n689 , n690 , n691 , n692 , n694 , n695 , n696 , n697 , n698 , n700 , n701 , n702 , n703 , n704 , n706 , n707 , n708 , n709 , n710 , n712 , n713 , n714 , n715 , n716 , n718 , n719 , n720 , n721 , n722 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n732 , n733 , n734 , n735 , n736 , n738 , n739 , n740 , n741 , n742 , n744 , n745 , n746 , n747 , n748 , n750 , n751 , n752 , n753 , n754 , n756 , n757 , n758 , n759 , n760 , n762 , n763 , n764 , n765 , n766 , n768 , n769 , n770 , n771 , n772 , n774 , n775 , n776 , n777 , n778 , n780 , n781 , n782 , n783 , n784 , n786 , n787 , n788 , n789 , n790 , n792 , n793 , n794 , n795 , n796 , n798 , n799 , n800 , n801 , n802 , n804 , n805 , n806 , n807 , n808 , n810 , n811 , n812 , n813 , n814 , n816 , n817 , n818 , n819 , n820 , n822 , n823 , n824 , n826 , n827 , n828 , n830 , n831 , n832 , n834 , n835 , n836 , n838 , n839 , n840 , n842 , n843 , n844 , n846 , n847 , n848 , n850 , n851 , n852 , n854 , n855 , n856 , n858 , n859 , n860 , n862 , n863 , n864 , n866 , n867 , n868 , n870 , n871 , n872 , n874 , n875 , n876 , n878 , n879 , n880 , n882 , n883 , n884 , n886 , n887 , n888 , n890 , n891 , n892 , n894 , n895 , n896 , n898 , n899 , n900 , n902 , n903 , n904 , n906 , n907 , n908 , n910 , n911 , n912 , n914 , n915 , n916 , n918 , n919 , n920 , n922 , n923 , n924 , n926 , n927 , n928 , n930 , n931 , n932 , n934 , n935 , n936 , n938 , n939 , n940 , n942 , n943 , n944 , n946 , n947 , n948 , n950 , n951 , n952 , n954 , n955 , n956 , n958 , n959 , n960 , n962 , n963 , n964 , n966 , n967 , n968 , n970 , n971 , n972 , n974 , n975 , n976 , n978 , n979 , n980 , n982 , n983 , n984 , n986 , n987 , n988 , n990 , n991 , n992 , n994 , n995 , n996 , n998 , n999 , n1000 , n1002 , n1003 , n1004 , n1006 , n1007 , n1008 , n1010 , n1011 , n1012 , n1014 , n1015 , n1016 , n1018 , n1019 , n1020 , n1022 , n1023 , n1024 , n1026 , n1027 , n1028 , n1030 , n1031 , n1032 , n1034 , n1035 , n1036 , n1038 , n1039 , n1040 , n1042 , n1043 , n1044 , n1046 , n1047 , n1048 , n1050 , n1051 , n1052 , n1054 , n1055 , n1056 , n1058 , n1059 , n1060 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 , n1070 , n1071 , n1072 , n1074 , n1075 , n1076 , n1078 , n1079 , n1080 , n1082 , n1083 , n1084 , n1086 , n1087 , n1088 , n1090 , n1091 , n1092 , n1094 , n1095 , n1096 , n1098 , n1099 , n1100 , n1102 , n1103 , n1104 , n1106 , n1107 , n1108 , n1110 , n1111 , n1112 , n1114 , n1115 , n1116 , n1118 , n1119 , n1120 , n1122 , n1123 , n1124 , n1126 , n1127 , n1128 , n1130 , n1131 , n1132 , n1134 , n1135 , n1136 , n1138 , n1139 , n1140 , n1142 , n1143 , n1144 , n1146 , n1147 , n1148 , n1150 , n1151 , n1152 , n1154 , n1155 , n1156 , n1158 , n1159 , n1160 , n1162 , n1163 , n1164 , n1166 , n1167 , n1168 , n1170 , n1171 , n1172 , n1174 , n1175 , n1176 , n1178 , n1179 , n1180 , n1182 , n1183 , n1184 , n1186 , n1187 , n1188 , n1190 , n1191 , n1192 , n1194 , n1195 , n1196 , n1198 , n1199 , n1200 , n1202 , n1203 , n1204 , n1206 , n1207 , n1208 , n1210 , n1211 , n1212 , n1214 , n1215 , n1216 , n1218 , n1219 , n1220 , n1222 , n1223 , n1224 , n1226 , n1227 , n1228 , n1230 , n1231 , n1232 , n1234 , n1235 , n1236 , n1238 , n1239 , n1240 , n1242 , n1243 , n1244 , n1246 , n1247 , n1248 , n1250 , n1251 , n1252 , n1254 , n1255 , n1256 , n1258 , n1259 , n1260 , n1262 , n1263 , n1264 , n1266 , n1267 , n1268 , n1270 , n1271 , n1272 , n1274 , n1275 , n1276 , n1278 , n1279 , n1280 , n1282 , n1283 , n1284 , n1286 , n1287 , n1288 , n1290 , n1291 , n1292 , n1294 , n1295 , n1296 , n1298 , n1299 , n1300 , n1302 , n1303 , n1304 , n1306 , n1307 , n1308 , n1310 , n1311 , n1312 , n1314 , n1315 , n1316 , n1318 , n1319 , n1320 , n1322 , n1323 , n1324 , n1326 , n1327 , n1328 , n1330 , n1331 , n1332 , n1334 , n1335 , n1336 ;
  assign n9 = ~x4 & ~x5 ;
  assign n10 = ~x6 & x7 ;
  assign n11 = n9 & n10 ;
  assign n12 = ~x0 & ~x2 ;
  assign n13 = ~x1 & ~x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n24 = n15 & x8 ;
  assign n16 = x4 & x5 ;
  assign n17 = x6 & ~x7 ;
  assign n18 = n16 & n17 ;
  assign n19 = x0 & x2 ;
  assign n20 = x1 & x3 ;
  assign n21 = n19 & n20 ;
  assign n22 = n18 & n21 ;
  assign n25 = ~n22 & ~x8 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = x0 & ~x2 ;
  assign n28 = n13 & n27 ;
  assign n29 = n11 & n28 ;
  assign n34 = n29 & x9 ;
  assign n30 = ~x0 & x2 ;
  assign n31 = n20 & n30 ;
  assign n32 = n18 & n31 ;
  assign n35 = ~n32 & ~x9 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = x1 & ~x3 ;
  assign n38 = n12 & n37 ;
  assign n39 = n11 & n38 ;
  assign n44 = n39 & x10 ;
  assign n40 = ~x1 & x3 ;
  assign n41 = n19 & n40 ;
  assign n42 = n18 & n41 ;
  assign n45 = ~n42 & ~x10 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n27 & n37 ;
  assign n48 = n11 & n47 ;
  assign n52 = n48 & x11 ;
  assign n49 = n30 & n40 ;
  assign n50 = n18 & n49 ;
  assign n53 = ~n50 & ~x11 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n13 & n30 ;
  assign n56 = n11 & n55 ;
  assign n60 = n56 & x12 ;
  assign n57 = n20 & n27 ;
  assign n58 = n18 & n57 ;
  assign n61 = ~n58 & ~x12 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = n13 & n19 ;
  assign n64 = n11 & n63 ;
  assign n68 = n64 & x13 ;
  assign n65 = n12 & n20 ;
  assign n66 = n18 & n65 ;
  assign n69 = ~n66 & ~x13 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = n30 & n37 ;
  assign n72 = n11 & n71 ;
  assign n76 = n72 & x14 ;
  assign n73 = n27 & n40 ;
  assign n74 = n18 & n73 ;
  assign n77 = ~n74 & ~x14 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = n19 & n37 ;
  assign n80 = n11 & n79 ;
  assign n84 = n80 & x15 ;
  assign n81 = n12 & n40 ;
  assign n82 = n18 & n81 ;
  assign n85 = ~n82 & ~x15 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n11 & n81 ;
  assign n90 = n87 & x16 ;
  assign n88 = n18 & n79 ;
  assign n91 = ~n88 & ~x16 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = n11 & n73 ;
  assign n96 = n93 & x17 ;
  assign n94 = n18 & n71 ;
  assign n97 = ~n94 & ~x17 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = n11 & n65 ;
  assign n102 = n99 & x18 ;
  assign n100 = n18 & n63 ;
  assign n103 = ~n100 & ~x18 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = n11 & n57 ;
  assign n108 = n105 & x19 ;
  assign n106 = n18 & n55 ;
  assign n109 = ~n106 & ~x19 ;
  assign n110 = ~n108 & ~n109 ;
  assign n111 = n11 & n49 ;
  assign n114 = n111 & x20 ;
  assign n112 = n18 & n47 ;
  assign n115 = ~n112 & ~x20 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = n11 & n41 ;
  assign n120 = n117 & x21 ;
  assign n118 = n18 & n38 ;
  assign n121 = ~n118 & ~x21 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = n11 & n31 ;
  assign n126 = n123 & x22 ;
  assign n124 = n18 & n28 ;
  assign n127 = ~n124 & ~x22 ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = n11 & n21 ;
  assign n132 = n129 & x23 ;
  assign n130 = n14 & n18 ;
  assign n133 = ~n130 & ~x23 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = x4 & ~x5 ;
  assign n136 = n10 & n135 ;
  assign n137 = n14 & n136 ;
  assign n142 = n137 & x24 ;
  assign n138 = ~x4 & x5 ;
  assign n139 = n17 & n138 ;
  assign n140 = n21 & n139 ;
  assign n143 = ~n140 & ~x24 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = n28 & n136 ;
  assign n148 = n145 & x25 ;
  assign n146 = n31 & n139 ;
  assign n149 = ~n146 & ~x25 ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = n38 & n136 ;
  assign n154 = n151 & x26 ;
  assign n152 = n41 & n139 ;
  assign n155 = ~n152 & ~x26 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = n47 & n136 ;
  assign n160 = n157 & x27 ;
  assign n158 = n49 & n139 ;
  assign n161 = ~n158 & ~x27 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = n55 & n136 ;
  assign n166 = n163 & x28 ;
  assign n164 = n57 & n139 ;
  assign n167 = ~n164 & ~x28 ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = n63 & n136 ;
  assign n172 = n169 & x29 ;
  assign n170 = n65 & n139 ;
  assign n173 = ~n170 & ~x29 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = n71 & n136 ;
  assign n178 = n175 & x30 ;
  assign n176 = n73 & n139 ;
  assign n179 = ~n176 & ~x30 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = n79 & n136 ;
  assign n184 = n181 & x31 ;
  assign n182 = n81 & n139 ;
  assign n185 = ~n182 & ~x31 ;
  assign n186 = ~n184 & ~n185 ;
  assign n187 = n81 & n136 ;
  assign n190 = n187 & x32 ;
  assign n188 = n79 & n139 ;
  assign n191 = ~n188 & ~x32 ;
  assign n192 = ~n190 & ~n191 ;
  assign n193 = n73 & n136 ;
  assign n196 = n193 & x33 ;
  assign n194 = n71 & n139 ;
  assign n197 = ~n194 & ~x33 ;
  assign n198 = ~n196 & ~n197 ;
  assign n199 = n65 & n136 ;
  assign n202 = n199 & x34 ;
  assign n200 = n63 & n139 ;
  assign n203 = ~n200 & ~x34 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = n57 & n136 ;
  assign n208 = n205 & x35 ;
  assign n206 = n55 & n139 ;
  assign n209 = ~n206 & ~x35 ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = n49 & n136 ;
  assign n214 = n211 & x36 ;
  assign n212 = n47 & n139 ;
  assign n215 = ~n212 & ~x36 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = n41 & n136 ;
  assign n220 = n217 & x37 ;
  assign n218 = n38 & n139 ;
  assign n221 = ~n218 & ~x37 ;
  assign n222 = ~n220 & ~n221 ;
  assign n223 = n31 & n136 ;
  assign n226 = n223 & x38 ;
  assign n224 = n28 & n139 ;
  assign n227 = ~n224 & ~x38 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = n21 & n136 ;
  assign n232 = n229 & x39 ;
  assign n230 = n14 & n139 ;
  assign n233 = ~n230 & ~x39 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = n10 & n138 ;
  assign n236 = n14 & n235 ;
  assign n240 = n236 & x40 ;
  assign n237 = n17 & n135 ;
  assign n238 = n21 & n237 ;
  assign n241 = ~n238 & ~x40 ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = n28 & n235 ;
  assign n246 = n243 & x41 ;
  assign n244 = n31 & n237 ;
  assign n247 = ~n244 & ~x41 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = n38 & n235 ;
  assign n252 = n249 & x42 ;
  assign n250 = n41 & n237 ;
  assign n253 = ~n250 & ~x42 ;
  assign n254 = ~n252 & ~n253 ;
  assign n255 = n47 & n235 ;
  assign n258 = n255 & x43 ;
  assign n256 = n49 & n237 ;
  assign n259 = ~n256 & ~x43 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = n55 & n235 ;
  assign n264 = n261 & x44 ;
  assign n262 = n57 & n237 ;
  assign n265 = ~n262 & ~x44 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n63 & n235 ;
  assign n270 = n267 & x45 ;
  assign n268 = n65 & n237 ;
  assign n271 = ~n268 & ~x45 ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = n71 & n235 ;
  assign n276 = n273 & x46 ;
  assign n274 = n73 & n237 ;
  assign n277 = ~n274 & ~x46 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = n79 & n235 ;
  assign n282 = n279 & x47 ;
  assign n280 = n81 & n237 ;
  assign n283 = ~n280 & ~x47 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n81 & n235 ;
  assign n288 = n285 & x48 ;
  assign n286 = n79 & n237 ;
  assign n289 = ~n286 & ~x48 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = n73 & n235 ;
  assign n294 = n291 & x49 ;
  assign n292 = n71 & n237 ;
  assign n295 = ~n292 & ~x49 ;
  assign n296 = ~n294 & ~n295 ;
  assign n297 = n65 & n235 ;
  assign n300 = n297 & x50 ;
  assign n298 = n63 & n237 ;
  assign n301 = ~n298 & ~x50 ;
  assign n302 = ~n300 & ~n301 ;
  assign n303 = n57 & n235 ;
  assign n306 = n303 & x51 ;
  assign n304 = n55 & n237 ;
  assign n307 = ~n304 & ~x51 ;
  assign n308 = ~n306 & ~n307 ;
  assign n309 = n49 & n235 ;
  assign n312 = n309 & x52 ;
  assign n310 = n47 & n237 ;
  assign n313 = ~n310 & ~x52 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = n41 & n235 ;
  assign n318 = n315 & x53 ;
  assign n316 = n38 & n237 ;
  assign n319 = ~n316 & ~x53 ;
  assign n320 = ~n318 & ~n319 ;
  assign n321 = n31 & n235 ;
  assign n324 = n321 & x54 ;
  assign n322 = n28 & n237 ;
  assign n325 = ~n322 & ~x54 ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = n21 & n235 ;
  assign n330 = n327 & x55 ;
  assign n328 = n14 & n237 ;
  assign n331 = ~n328 & ~x55 ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = n10 & n16 ;
  assign n334 = n14 & n333 ;
  assign n338 = n334 & x56 ;
  assign n335 = n9 & n17 ;
  assign n336 = n21 & n335 ;
  assign n339 = ~n336 & ~x56 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n28 & n333 ;
  assign n344 = n341 & x57 ;
  assign n342 = n31 & n335 ;
  assign n345 = ~n342 & ~x57 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = n38 & n333 ;
  assign n350 = n347 & x58 ;
  assign n348 = n41 & n335 ;
  assign n351 = ~n348 & ~x58 ;
  assign n352 = ~n350 & ~n351 ;
  assign n353 = n47 & n333 ;
  assign n356 = n353 & x59 ;
  assign n354 = n49 & n335 ;
  assign n357 = ~n354 & ~x59 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = n55 & n333 ;
  assign n362 = n359 & x60 ;
  assign n360 = n57 & n335 ;
  assign n363 = ~n360 & ~x60 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = n63 & n333 ;
  assign n368 = n365 & x61 ;
  assign n366 = n65 & n335 ;
  assign n369 = ~n366 & ~x61 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = n71 & n333 ;
  assign n374 = n371 & x62 ;
  assign n372 = n73 & n335 ;
  assign n375 = ~n372 & ~x62 ;
  assign n376 = ~n374 & ~n375 ;
  assign n377 = n79 & n333 ;
  assign n380 = n377 & x63 ;
  assign n378 = n81 & n335 ;
  assign n381 = ~n378 & ~x63 ;
  assign n382 = ~n380 & ~n381 ;
  assign n383 = n81 & n333 ;
  assign n386 = n383 & x64 ;
  assign n384 = n79 & n335 ;
  assign n387 = ~n384 & ~x64 ;
  assign n388 = ~n386 & ~n387 ;
  assign n389 = n73 & n333 ;
  assign n392 = n389 & x65 ;
  assign n390 = n71 & n335 ;
  assign n393 = ~n390 & ~x65 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = n65 & n333 ;
  assign n398 = n395 & x66 ;
  assign n396 = n63 & n335 ;
  assign n399 = ~n396 & ~x66 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = n57 & n333 ;
  assign n404 = n401 & x67 ;
  assign n402 = n55 & n335 ;
  assign n405 = ~n402 & ~x67 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n49 & n333 ;
  assign n410 = n407 & x68 ;
  assign n408 = n47 & n335 ;
  assign n411 = ~n408 & ~x68 ;
  assign n412 = ~n410 & ~n411 ;
  assign n413 = n41 & n333 ;
  assign n416 = n413 & x69 ;
  assign n414 = n38 & n335 ;
  assign n417 = ~n414 & ~x69 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = n31 & n333 ;
  assign n422 = n419 & x70 ;
  assign n420 = n28 & n335 ;
  assign n423 = ~n420 & ~x70 ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = n21 & n333 ;
  assign n428 = n425 & x71 ;
  assign n426 = n14 & n335 ;
  assign n429 = ~n426 & ~x71 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = x6 & x7 ;
  assign n432 = n9 & n431 ;
  assign n433 = n14 & n432 ;
  assign n438 = n433 & x72 ;
  assign n434 = ~x6 & ~x7 ;
  assign n435 = n16 & n434 ;
  assign n436 = n21 & n435 ;
  assign n439 = ~n436 & ~x72 ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = n28 & n432 ;
  assign n444 = n441 & x73 ;
  assign n442 = n31 & n435 ;
  assign n445 = ~n442 & ~x73 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n38 & n432 ;
  assign n450 = n447 & x74 ;
  assign n448 = n41 & n435 ;
  assign n451 = ~n448 & ~x74 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = n47 & n432 ;
  assign n456 = n453 & x75 ;
  assign n454 = n49 & n435 ;
  assign n457 = ~n454 & ~x75 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = n55 & n432 ;
  assign n462 = n459 & x76 ;
  assign n460 = n57 & n435 ;
  assign n463 = ~n460 & ~x76 ;
  assign n464 = ~n462 & ~n463 ;
  assign n465 = n63 & n432 ;
  assign n468 = n465 & x77 ;
  assign n466 = n65 & n435 ;
  assign n469 = ~n466 & ~x77 ;
  assign n470 = ~n468 & ~n469 ;
  assign n471 = n71 & n432 ;
  assign n474 = n471 & x78 ;
  assign n472 = n73 & n435 ;
  assign n475 = ~n472 & ~x78 ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = n79 & n432 ;
  assign n480 = n477 & x79 ;
  assign n478 = n81 & n435 ;
  assign n481 = ~n478 & ~x79 ;
  assign n482 = ~n480 & ~n481 ;
  assign n483 = n81 & n432 ;
  assign n486 = n483 & x80 ;
  assign n484 = n79 & n435 ;
  assign n487 = ~n484 & ~x80 ;
  assign n488 = ~n486 & ~n487 ;
  assign n489 = n73 & n432 ;
  assign n492 = n489 & x81 ;
  assign n490 = n71 & n435 ;
  assign n493 = ~n490 & ~x81 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = n65 & n432 ;
  assign n498 = n495 & x82 ;
  assign n496 = n63 & n435 ;
  assign n499 = ~n496 & ~x82 ;
  assign n500 = ~n498 & ~n499 ;
  assign n501 = n57 & n432 ;
  assign n504 = n501 & x83 ;
  assign n502 = n55 & n435 ;
  assign n505 = ~n502 & ~x83 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = n49 & n432 ;
  assign n510 = n507 & x84 ;
  assign n508 = n47 & n435 ;
  assign n511 = ~n508 & ~x84 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = n41 & n432 ;
  assign n516 = n513 & x85 ;
  assign n514 = n38 & n435 ;
  assign n517 = ~n514 & ~x85 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = n31 & n432 ;
  assign n522 = n519 & x86 ;
  assign n520 = n28 & n435 ;
  assign n523 = ~n520 & ~x86 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = n21 & n432 ;
  assign n528 = n525 & x87 ;
  assign n526 = n14 & n435 ;
  assign n529 = ~n526 & ~x87 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = n135 & n431 ;
  assign n532 = n14 & n531 ;
  assign n536 = n532 & x88 ;
  assign n533 = n138 & n434 ;
  assign n534 = n21 & n533 ;
  assign n537 = ~n534 & ~x88 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = n28 & n531 ;
  assign n542 = n539 & x89 ;
  assign n540 = n31 & n533 ;
  assign n543 = ~n540 & ~x89 ;
  assign n544 = ~n542 & ~n543 ;
  assign n545 = n38 & n531 ;
  assign n548 = n545 & x90 ;
  assign n546 = n41 & n533 ;
  assign n549 = ~n546 & ~x90 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = n47 & n531 ;
  assign n554 = n551 & x91 ;
  assign n552 = n49 & n533 ;
  assign n555 = ~n552 & ~x91 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = n55 & n531 ;
  assign n560 = n557 & x92 ;
  assign n558 = n57 & n533 ;
  assign n561 = ~n558 & ~x92 ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = n63 & n531 ;
  assign n566 = n563 & x93 ;
  assign n564 = n65 & n533 ;
  assign n567 = ~n564 & ~x93 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = n71 & n531 ;
  assign n572 = n569 & x94 ;
  assign n570 = n73 & n533 ;
  assign n573 = ~n570 & ~x94 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = n79 & n531 ;
  assign n578 = n575 & x95 ;
  assign n576 = n81 & n533 ;
  assign n579 = ~n576 & ~x95 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = n81 & n531 ;
  assign n584 = n581 & x96 ;
  assign n582 = n79 & n533 ;
  assign n585 = ~n582 & ~x96 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = n73 & n531 ;
  assign n590 = n587 & x97 ;
  assign n588 = n71 & n533 ;
  assign n591 = ~n588 & ~x97 ;
  assign n592 = ~n590 & ~n591 ;
  assign n593 = n65 & n531 ;
  assign n596 = n593 & x98 ;
  assign n594 = n63 & n533 ;
  assign n597 = ~n594 & ~x98 ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = n57 & n531 ;
  assign n602 = n599 & x99 ;
  assign n600 = n55 & n533 ;
  assign n603 = ~n600 & ~x99 ;
  assign n604 = ~n602 & ~n603 ;
  assign n605 = n49 & n531 ;
  assign n608 = n605 & x100 ;
  assign n606 = n47 & n533 ;
  assign n609 = ~n606 & ~x100 ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = n41 & n531 ;
  assign n614 = n611 & x101 ;
  assign n612 = n38 & n533 ;
  assign n615 = ~n612 & ~x101 ;
  assign n616 = ~n614 & ~n615 ;
  assign n617 = n31 & n531 ;
  assign n620 = n617 & x102 ;
  assign n618 = n28 & n533 ;
  assign n621 = ~n618 & ~x102 ;
  assign n622 = ~n620 & ~n621 ;
  assign n623 = n21 & n531 ;
  assign n626 = n623 & x103 ;
  assign n624 = n14 & n533 ;
  assign n627 = ~n624 & ~x103 ;
  assign n628 = ~n626 & ~n627 ;
  assign n629 = n138 & n431 ;
  assign n630 = n14 & n629 ;
  assign n634 = n630 & x104 ;
  assign n631 = n135 & n434 ;
  assign n632 = n21 & n631 ;
  assign n635 = ~n632 & ~x104 ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = n28 & n629 ;
  assign n640 = n637 & x105 ;
  assign n638 = n31 & n631 ;
  assign n641 = ~n638 & ~x105 ;
  assign n642 = ~n640 & ~n641 ;
  assign n643 = n38 & n629 ;
  assign n646 = n643 & x106 ;
  assign n644 = n41 & n631 ;
  assign n647 = ~n644 & ~x106 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = n47 & n629 ;
  assign n652 = n649 & x107 ;
  assign n650 = n49 & n631 ;
  assign n653 = ~n650 & ~x107 ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = n55 & n629 ;
  assign n658 = n655 & x108 ;
  assign n656 = n57 & n631 ;
  assign n659 = ~n656 & ~x108 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = n63 & n629 ;
  assign n664 = n661 & x109 ;
  assign n662 = n65 & n631 ;
  assign n665 = ~n662 & ~x109 ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = n71 & n629 ;
  assign n670 = n667 & x110 ;
  assign n668 = n73 & n631 ;
  assign n671 = ~n668 & ~x110 ;
  assign n672 = ~n670 & ~n671 ;
  assign n673 = n79 & n629 ;
  assign n676 = n673 & x111 ;
  assign n674 = n81 & n631 ;
  assign n677 = ~n674 & ~x111 ;
  assign n678 = ~n676 & ~n677 ;
  assign n679 = n81 & n629 ;
  assign n682 = n679 & x112 ;
  assign n680 = n79 & n631 ;
  assign n683 = ~n680 & ~x112 ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = n73 & n629 ;
  assign n688 = n685 & x113 ;
  assign n686 = n71 & n631 ;
  assign n689 = ~n686 & ~x113 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = n65 & n629 ;
  assign n694 = n691 & x114 ;
  assign n692 = n63 & n631 ;
  assign n695 = ~n692 & ~x114 ;
  assign n696 = ~n694 & ~n695 ;
  assign n697 = n57 & n629 ;
  assign n700 = n697 & x115 ;
  assign n698 = n55 & n631 ;
  assign n701 = ~n698 & ~x115 ;
  assign n702 = ~n700 & ~n701 ;
  assign n703 = n49 & n629 ;
  assign n706 = n703 & x116 ;
  assign n704 = n47 & n631 ;
  assign n707 = ~n704 & ~x116 ;
  assign n708 = ~n706 & ~n707 ;
  assign n709 = n41 & n629 ;
  assign n712 = n709 & x117 ;
  assign n710 = n38 & n631 ;
  assign n713 = ~n710 & ~x117 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = n31 & n629 ;
  assign n718 = n715 & x118 ;
  assign n716 = n28 & n631 ;
  assign n719 = ~n716 & ~x118 ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = n21 & n629 ;
  assign n724 = n721 & x119 ;
  assign n722 = n14 & n631 ;
  assign n725 = ~n722 & ~x119 ;
  assign n726 = ~n724 & ~n725 ;
  assign n727 = n16 & n431 ;
  assign n728 = n14 & n727 ;
  assign n732 = n728 & x120 ;
  assign n729 = n9 & n434 ;
  assign n730 = n21 & n729 ;
  assign n733 = ~n730 & ~x120 ;
  assign n734 = ~n732 & ~n733 ;
  assign n735 = n28 & n727 ;
  assign n738 = n735 & x121 ;
  assign n736 = n31 & n729 ;
  assign n739 = ~n736 & ~x121 ;
  assign n740 = ~n738 & ~n739 ;
  assign n741 = n38 & n727 ;
  assign n744 = n741 & x122 ;
  assign n742 = n41 & n729 ;
  assign n745 = ~n742 & ~x122 ;
  assign n746 = ~n744 & ~n745 ;
  assign n747 = n47 & n727 ;
  assign n750 = n747 & x123 ;
  assign n748 = n49 & n729 ;
  assign n751 = ~n748 & ~x123 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = n55 & n727 ;
  assign n756 = n753 & x124 ;
  assign n754 = n57 & n729 ;
  assign n757 = ~n754 & ~x124 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = n63 & n727 ;
  assign n762 = n759 & x125 ;
  assign n760 = n65 & n729 ;
  assign n763 = ~n760 & ~x125 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = n71 & n727 ;
  assign n768 = n765 & x126 ;
  assign n766 = n73 & n729 ;
  assign n769 = ~n766 & ~x126 ;
  assign n770 = ~n768 & ~n769 ;
  assign n771 = n79 & n727 ;
  assign n774 = n771 & x127 ;
  assign n772 = n81 & n729 ;
  assign n775 = ~n772 & ~x127 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = n81 & n727 ;
  assign n780 = n777 & x128 ;
  assign n778 = n79 & n729 ;
  assign n781 = ~n778 & ~x128 ;
  assign n782 = ~n780 & ~n781 ;
  assign n783 = n73 & n727 ;
  assign n786 = n783 & x129 ;
  assign n784 = n71 & n729 ;
  assign n787 = ~n784 & ~x129 ;
  assign n788 = ~n786 & ~n787 ;
  assign n789 = n65 & n727 ;
  assign n792 = n789 & x130 ;
  assign n790 = n63 & n729 ;
  assign n793 = ~n790 & ~x130 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = n57 & n727 ;
  assign n798 = n795 & x131 ;
  assign n796 = n55 & n729 ;
  assign n799 = ~n796 & ~x131 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = n49 & n727 ;
  assign n804 = n801 & x132 ;
  assign n802 = n47 & n729 ;
  assign n805 = ~n802 & ~x132 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = n41 & n727 ;
  assign n810 = n807 & x133 ;
  assign n808 = n38 & n729 ;
  assign n811 = ~n808 & ~x133 ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = n31 & n727 ;
  assign n816 = n813 & x134 ;
  assign n814 = n28 & n729 ;
  assign n817 = ~n814 & ~x134 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = n21 & n727 ;
  assign n822 = n819 & x135 ;
  assign n820 = n14 & n729 ;
  assign n823 = ~n820 & ~x135 ;
  assign n824 = ~n822 & ~n823 ;
  assign n826 = n820 & x136 ;
  assign n827 = ~n819 & ~x136 ;
  assign n828 = ~n826 & ~n827 ;
  assign n830 = n814 & x137 ;
  assign n831 = ~n813 & ~x137 ;
  assign n832 = ~n830 & ~n831 ;
  assign n834 = n808 & x138 ;
  assign n835 = ~n807 & ~x138 ;
  assign n836 = ~n834 & ~n835 ;
  assign n838 = n802 & x139 ;
  assign n839 = ~n801 & ~x139 ;
  assign n840 = ~n838 & ~n839 ;
  assign n842 = n796 & x140 ;
  assign n843 = ~n795 & ~x140 ;
  assign n844 = ~n842 & ~n843 ;
  assign n846 = n790 & x141 ;
  assign n847 = ~n789 & ~x141 ;
  assign n848 = ~n846 & ~n847 ;
  assign n850 = n784 & x142 ;
  assign n851 = ~n783 & ~x142 ;
  assign n852 = ~n850 & ~n851 ;
  assign n854 = n778 & x143 ;
  assign n855 = ~n777 & ~x143 ;
  assign n856 = ~n854 & ~n855 ;
  assign n858 = n772 & x144 ;
  assign n859 = ~n771 & ~x144 ;
  assign n860 = ~n858 & ~n859 ;
  assign n862 = n766 & x145 ;
  assign n863 = ~n765 & ~x145 ;
  assign n864 = ~n862 & ~n863 ;
  assign n866 = n760 & x146 ;
  assign n867 = ~n759 & ~x146 ;
  assign n868 = ~n866 & ~n867 ;
  assign n870 = n754 & x147 ;
  assign n871 = ~n753 & ~x147 ;
  assign n872 = ~n870 & ~n871 ;
  assign n874 = n748 & x148 ;
  assign n875 = ~n747 & ~x148 ;
  assign n876 = ~n874 & ~n875 ;
  assign n878 = n742 & x149 ;
  assign n879 = ~n741 & ~x149 ;
  assign n880 = ~n878 & ~n879 ;
  assign n882 = n736 & x150 ;
  assign n883 = ~n735 & ~x150 ;
  assign n884 = ~n882 & ~n883 ;
  assign n886 = n730 & x151 ;
  assign n887 = ~n728 & ~x151 ;
  assign n888 = ~n886 & ~n887 ;
  assign n890 = n722 & x152 ;
  assign n891 = ~n721 & ~x152 ;
  assign n892 = ~n890 & ~n891 ;
  assign n894 = n716 & x153 ;
  assign n895 = ~n715 & ~x153 ;
  assign n896 = ~n894 & ~n895 ;
  assign n898 = n710 & x154 ;
  assign n899 = ~n709 & ~x154 ;
  assign n900 = ~n898 & ~n899 ;
  assign n902 = n704 & x155 ;
  assign n903 = ~n703 & ~x155 ;
  assign n904 = ~n902 & ~n903 ;
  assign n906 = n698 & x156 ;
  assign n907 = ~n697 & ~x156 ;
  assign n908 = ~n906 & ~n907 ;
  assign n910 = n692 & x157 ;
  assign n911 = ~n691 & ~x157 ;
  assign n912 = ~n910 & ~n911 ;
  assign n914 = n686 & x158 ;
  assign n915 = ~n685 & ~x158 ;
  assign n916 = ~n914 & ~n915 ;
  assign n918 = n680 & x159 ;
  assign n919 = ~n679 & ~x159 ;
  assign n920 = ~n918 & ~n919 ;
  assign n922 = n674 & x160 ;
  assign n923 = ~n673 & ~x160 ;
  assign n924 = ~n922 & ~n923 ;
  assign n926 = n668 & x161 ;
  assign n927 = ~n667 & ~x161 ;
  assign n928 = ~n926 & ~n927 ;
  assign n930 = n662 & x162 ;
  assign n931 = ~n661 & ~x162 ;
  assign n932 = ~n930 & ~n931 ;
  assign n934 = n656 & x163 ;
  assign n935 = ~n655 & ~x163 ;
  assign n936 = ~n934 & ~n935 ;
  assign n938 = n650 & x164 ;
  assign n939 = ~n649 & ~x164 ;
  assign n940 = ~n938 & ~n939 ;
  assign n942 = n644 & x165 ;
  assign n943 = ~n643 & ~x165 ;
  assign n944 = ~n942 & ~n943 ;
  assign n946 = n638 & x166 ;
  assign n947 = ~n637 & ~x166 ;
  assign n948 = ~n946 & ~n947 ;
  assign n950 = n632 & x167 ;
  assign n951 = ~n630 & ~x167 ;
  assign n952 = ~n950 & ~n951 ;
  assign n954 = n624 & x168 ;
  assign n955 = ~n623 & ~x168 ;
  assign n956 = ~n954 & ~n955 ;
  assign n958 = n618 & x169 ;
  assign n959 = ~n617 & ~x169 ;
  assign n960 = ~n958 & ~n959 ;
  assign n962 = n612 & x170 ;
  assign n963 = ~n611 & ~x170 ;
  assign n964 = ~n962 & ~n963 ;
  assign n966 = n606 & x171 ;
  assign n967 = ~n605 & ~x171 ;
  assign n968 = ~n966 & ~n967 ;
  assign n970 = n600 & x172 ;
  assign n971 = ~n599 & ~x172 ;
  assign n972 = ~n970 & ~n971 ;
  assign n974 = n594 & x173 ;
  assign n975 = ~n593 & ~x173 ;
  assign n976 = ~n974 & ~n975 ;
  assign n978 = n588 & x174 ;
  assign n979 = ~n587 & ~x174 ;
  assign n980 = ~n978 & ~n979 ;
  assign n982 = n582 & x175 ;
  assign n983 = ~n581 & ~x175 ;
  assign n984 = ~n982 & ~n983 ;
  assign n986 = n576 & x176 ;
  assign n987 = ~n575 & ~x176 ;
  assign n988 = ~n986 & ~n987 ;
  assign n990 = n570 & x177 ;
  assign n991 = ~n569 & ~x177 ;
  assign n992 = ~n990 & ~n991 ;
  assign n994 = n564 & x178 ;
  assign n995 = ~n563 & ~x178 ;
  assign n996 = ~n994 & ~n995 ;
  assign n998 = n558 & x179 ;
  assign n999 = ~n557 & ~x179 ;
  assign n1000 = ~n998 & ~n999 ;
  assign n1002 = n552 & x180 ;
  assign n1003 = ~n551 & ~x180 ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1006 = n546 & x181 ;
  assign n1007 = ~n545 & ~x181 ;
  assign n1008 = ~n1006 & ~n1007 ;
  assign n1010 = n540 & x182 ;
  assign n1011 = ~n539 & ~x182 ;
  assign n1012 = ~n1010 & ~n1011 ;
  assign n1014 = n534 & x183 ;
  assign n1015 = ~n532 & ~x183 ;
  assign n1016 = ~n1014 & ~n1015 ;
  assign n1018 = n526 & x184 ;
  assign n1019 = ~n525 & ~x184 ;
  assign n1020 = ~n1018 & ~n1019 ;
  assign n1022 = n520 & x185 ;
  assign n1023 = ~n519 & ~x185 ;
  assign n1024 = ~n1022 & ~n1023 ;
  assign n1026 = n514 & x186 ;
  assign n1027 = ~n513 & ~x186 ;
  assign n1028 = ~n1026 & ~n1027 ;
  assign n1030 = n508 & x187 ;
  assign n1031 = ~n507 & ~x187 ;
  assign n1032 = ~n1030 & ~n1031 ;
  assign n1034 = n502 & x188 ;
  assign n1035 = ~n501 & ~x188 ;
  assign n1036 = ~n1034 & ~n1035 ;
  assign n1038 = n496 & x189 ;
  assign n1039 = ~n495 & ~x189 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1042 = n490 & x190 ;
  assign n1043 = ~n489 & ~x190 ;
  assign n1044 = ~n1042 & ~n1043 ;
  assign n1046 = n484 & x191 ;
  assign n1047 = ~n483 & ~x191 ;
  assign n1048 = ~n1046 & ~n1047 ;
  assign n1050 = n478 & x192 ;
  assign n1051 = ~n477 & ~x192 ;
  assign n1052 = ~n1050 & ~n1051 ;
  assign n1054 = n472 & x193 ;
  assign n1055 = ~n471 & ~x193 ;
  assign n1056 = ~n1054 & ~n1055 ;
  assign n1058 = n466 & x194 ;
  assign n1059 = ~n465 & ~x194 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1062 = n460 & x195 ;
  assign n1063 = ~n459 & ~x195 ;
  assign n1064 = ~n1062 & ~n1063 ;
  assign n1066 = n454 & x196 ;
  assign n1067 = ~n453 & ~x196 ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1070 = n448 & x197 ;
  assign n1071 = ~n447 & ~x197 ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1074 = n442 & x198 ;
  assign n1075 = ~n441 & ~x198 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1078 = n436 & x199 ;
  assign n1079 = ~n433 & ~x199 ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1082 = n426 & x200 ;
  assign n1083 = ~n425 & ~x200 ;
  assign n1084 = ~n1082 & ~n1083 ;
  assign n1086 = n420 & x201 ;
  assign n1087 = ~n419 & ~x201 ;
  assign n1088 = ~n1086 & ~n1087 ;
  assign n1090 = n414 & x202 ;
  assign n1091 = ~n413 & ~x202 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1094 = n408 & x203 ;
  assign n1095 = ~n407 & ~x203 ;
  assign n1096 = ~n1094 & ~n1095 ;
  assign n1098 = n402 & x204 ;
  assign n1099 = ~n401 & ~x204 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1102 = n396 & x205 ;
  assign n1103 = ~n395 & ~x205 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1106 = n390 & x206 ;
  assign n1107 = ~n389 & ~x206 ;
  assign n1108 = ~n1106 & ~n1107 ;
  assign n1110 = n384 & x207 ;
  assign n1111 = ~n383 & ~x207 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1114 = n378 & x208 ;
  assign n1115 = ~n377 & ~x208 ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1118 = n372 & x209 ;
  assign n1119 = ~n371 & ~x209 ;
  assign n1120 = ~n1118 & ~n1119 ;
  assign n1122 = n366 & x210 ;
  assign n1123 = ~n365 & ~x210 ;
  assign n1124 = ~n1122 & ~n1123 ;
  assign n1126 = n360 & x211 ;
  assign n1127 = ~n359 & ~x211 ;
  assign n1128 = ~n1126 & ~n1127 ;
  assign n1130 = n354 & x212 ;
  assign n1131 = ~n353 & ~x212 ;
  assign n1132 = ~n1130 & ~n1131 ;
  assign n1134 = n348 & x213 ;
  assign n1135 = ~n347 & ~x213 ;
  assign n1136 = ~n1134 & ~n1135 ;
  assign n1138 = n342 & x214 ;
  assign n1139 = ~n341 & ~x214 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1142 = n336 & x215 ;
  assign n1143 = ~n334 & ~x215 ;
  assign n1144 = ~n1142 & ~n1143 ;
  assign n1146 = n328 & x216 ;
  assign n1147 = ~n327 & ~x216 ;
  assign n1148 = ~n1146 & ~n1147 ;
  assign n1150 = n322 & x217 ;
  assign n1151 = ~n321 & ~x217 ;
  assign n1152 = ~n1150 & ~n1151 ;
  assign n1154 = n316 & x218 ;
  assign n1155 = ~n315 & ~x218 ;
  assign n1156 = ~n1154 & ~n1155 ;
  assign n1158 = n310 & x219 ;
  assign n1159 = ~n309 & ~x219 ;
  assign n1160 = ~n1158 & ~n1159 ;
  assign n1162 = n304 & x220 ;
  assign n1163 = ~n303 & ~x220 ;
  assign n1164 = ~n1162 & ~n1163 ;
  assign n1166 = n298 & x221 ;
  assign n1167 = ~n297 & ~x221 ;
  assign n1168 = ~n1166 & ~n1167 ;
  assign n1170 = n292 & x222 ;
  assign n1171 = ~n291 & ~x222 ;
  assign n1172 = ~n1170 & ~n1171 ;
  assign n1174 = n286 & x223 ;
  assign n1175 = ~n285 & ~x223 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1178 = n280 & x224 ;
  assign n1179 = ~n279 & ~x224 ;
  assign n1180 = ~n1178 & ~n1179 ;
  assign n1182 = n274 & x225 ;
  assign n1183 = ~n273 & ~x225 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1186 = n268 & x226 ;
  assign n1187 = ~n267 & ~x226 ;
  assign n1188 = ~n1186 & ~n1187 ;
  assign n1190 = n262 & x227 ;
  assign n1191 = ~n261 & ~x227 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1194 = n256 & x228 ;
  assign n1195 = ~n255 & ~x228 ;
  assign n1196 = ~n1194 & ~n1195 ;
  assign n1198 = n250 & x229 ;
  assign n1199 = ~n249 & ~x229 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1202 = n244 & x230 ;
  assign n1203 = ~n243 & ~x230 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1206 = n238 & x231 ;
  assign n1207 = ~n236 & ~x231 ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1210 = n230 & x232 ;
  assign n1211 = ~n229 & ~x232 ;
  assign n1212 = ~n1210 & ~n1211 ;
  assign n1214 = n224 & x233 ;
  assign n1215 = ~n223 & ~x233 ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1218 = n218 & x234 ;
  assign n1219 = ~n217 & ~x234 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1222 = n212 & x235 ;
  assign n1223 = ~n211 & ~x235 ;
  assign n1224 = ~n1222 & ~n1223 ;
  assign n1226 = n206 & x236 ;
  assign n1227 = ~n205 & ~x236 ;
  assign n1228 = ~n1226 & ~n1227 ;
  assign n1230 = n200 & x237 ;
  assign n1231 = ~n199 & ~x237 ;
  assign n1232 = ~n1230 & ~n1231 ;
  assign n1234 = n194 & x238 ;
  assign n1235 = ~n193 & ~x238 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1238 = n188 & x239 ;
  assign n1239 = ~n187 & ~x239 ;
  assign n1240 = ~n1238 & ~n1239 ;
  assign n1242 = n182 & x240 ;
  assign n1243 = ~n181 & ~x240 ;
  assign n1244 = ~n1242 & ~n1243 ;
  assign n1246 = n176 & x241 ;
  assign n1247 = ~n175 & ~x241 ;
  assign n1248 = ~n1246 & ~n1247 ;
  assign n1250 = n170 & x242 ;
  assign n1251 = ~n169 & ~x242 ;
  assign n1252 = ~n1250 & ~n1251 ;
  assign n1254 = n164 & x243 ;
  assign n1255 = ~n163 & ~x243 ;
  assign n1256 = ~n1254 & ~n1255 ;
  assign n1258 = n158 & x244 ;
  assign n1259 = ~n157 & ~x244 ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1262 = n152 & x245 ;
  assign n1263 = ~n151 & ~x245 ;
  assign n1264 = ~n1262 & ~n1263 ;
  assign n1266 = n146 & x246 ;
  assign n1267 = ~n145 & ~x246 ;
  assign n1268 = ~n1266 & ~n1267 ;
  assign n1270 = n140 & x247 ;
  assign n1271 = ~n137 & ~x247 ;
  assign n1272 = ~n1270 & ~n1271 ;
  assign n1274 = n130 & x248 ;
  assign n1275 = ~n129 & ~x248 ;
  assign n1276 = ~n1274 & ~n1275 ;
  assign n1278 = n124 & x249 ;
  assign n1279 = ~n123 & ~x249 ;
  assign n1280 = ~n1278 & ~n1279 ;
  assign n1282 = n118 & x250 ;
  assign n1283 = ~n117 & ~x250 ;
  assign n1284 = ~n1282 & ~n1283 ;
  assign n1286 = n112 & x251 ;
  assign n1287 = ~n111 & ~x251 ;
  assign n1288 = ~n1286 & ~n1287 ;
  assign n1290 = n106 & x252 ;
  assign n1291 = ~n105 & ~x252 ;
  assign n1292 = ~n1290 & ~n1291 ;
  assign n1294 = n100 & x253 ;
  assign n1295 = ~n99 & ~x253 ;
  assign n1296 = ~n1294 & ~n1295 ;
  assign n1298 = n94 & x254 ;
  assign n1299 = ~n93 & ~x254 ;
  assign n1300 = ~n1298 & ~n1299 ;
  assign n1302 = n88 & x255 ;
  assign n1303 = ~n87 & ~x255 ;
  assign n1304 = ~n1302 & ~n1303 ;
  assign n1306 = n82 & x256 ;
  assign n1307 = ~n80 & ~x256 ;
  assign n1308 = ~n1306 & ~n1307 ;
  assign n1310 = n74 & x257 ;
  assign n1311 = ~n72 & ~x257 ;
  assign n1312 = ~n1310 & ~n1311 ;
  assign n1314 = n66 & x258 ;
  assign n1315 = ~n64 & ~x258 ;
  assign n1316 = ~n1314 & ~n1315 ;
  assign n1318 = n58 & x259 ;
  assign n1319 = ~n56 & ~x259 ;
  assign n1320 = ~n1318 & ~n1319 ;
  assign n1322 = n50 & x260 ;
  assign n1323 = ~n48 & ~x260 ;
  assign n1324 = ~n1322 & ~n1323 ;
  assign n1326 = n42 & x261 ;
  assign n1327 = ~n39 & ~x261 ;
  assign n1328 = ~n1326 & ~n1327 ;
  assign n1330 = n32 & x262 ;
  assign n1331 = ~n29 & ~x262 ;
  assign n1332 = ~n1330 & ~n1331 ;
  assign n1334 = n22 & x263 ;
  assign n1335 = ~n15 & ~x263 ;
  assign n1336 = ~n1334 & ~n1335 ;
  assign y0 = ~n26 ;
  assign y1 = ~n36 ;
  assign y2 = ~n46 ;
  assign y3 = ~n54 ;
  assign y4 = ~n62 ;
  assign y5 = ~n70 ;
  assign y6 = ~n78 ;
  assign y7 = ~n86 ;
  assign y8 = ~n92 ;
  assign y9 = ~n98 ;
  assign y10 = ~n104 ;
  assign y11 = ~n110 ;
  assign y12 = ~n116 ;
  assign y13 = ~n122 ;
  assign y14 = ~n128 ;
  assign y15 = ~n134 ;
  assign y16 = ~n144 ;
  assign y17 = ~n150 ;
  assign y18 = ~n156 ;
  assign y19 = ~n162 ;
  assign y20 = ~n168 ;
  assign y21 = ~n174 ;
  assign y22 = ~n180 ;
  assign y23 = ~n186 ;
  assign y24 = ~n192 ;
  assign y25 = ~n198 ;
  assign y26 = ~n204 ;
  assign y27 = ~n210 ;
  assign y28 = ~n216 ;
  assign y29 = ~n222 ;
  assign y30 = ~n228 ;
  assign y31 = ~n234 ;
  assign y32 = ~n242 ;
  assign y33 = ~n248 ;
  assign y34 = ~n254 ;
  assign y35 = ~n260 ;
  assign y36 = ~n266 ;
  assign y37 = ~n272 ;
  assign y38 = ~n278 ;
  assign y39 = ~n284 ;
  assign y40 = ~n290 ;
  assign y41 = ~n296 ;
  assign y42 = ~n302 ;
  assign y43 = ~n308 ;
  assign y44 = ~n314 ;
  assign y45 = ~n320 ;
  assign y46 = ~n326 ;
  assign y47 = ~n332 ;
  assign y48 = ~n340 ;
  assign y49 = ~n346 ;
  assign y50 = ~n352 ;
  assign y51 = ~n358 ;
  assign y52 = ~n364 ;
  assign y53 = ~n370 ;
  assign y54 = ~n376 ;
  assign y55 = ~n382 ;
  assign y56 = ~n388 ;
  assign y57 = ~n394 ;
  assign y58 = ~n400 ;
  assign y59 = ~n406 ;
  assign y60 = ~n412 ;
  assign y61 = ~n418 ;
  assign y62 = ~n424 ;
  assign y63 = ~n430 ;
  assign y64 = ~n440 ;
  assign y65 = ~n446 ;
  assign y66 = ~n452 ;
  assign y67 = ~n458 ;
  assign y68 = ~n464 ;
  assign y69 = ~n470 ;
  assign y70 = ~n476 ;
  assign y71 = ~n482 ;
  assign y72 = ~n488 ;
  assign y73 = ~n494 ;
  assign y74 = ~n500 ;
  assign y75 = ~n506 ;
  assign y76 = ~n512 ;
  assign y77 = ~n518 ;
  assign y78 = ~n524 ;
  assign y79 = ~n530 ;
  assign y80 = ~n538 ;
  assign y81 = ~n544 ;
  assign y82 = ~n550 ;
  assign y83 = ~n556 ;
  assign y84 = ~n562 ;
  assign y85 = ~n568 ;
  assign y86 = ~n574 ;
  assign y87 = ~n580 ;
  assign y88 = ~n586 ;
  assign y89 = ~n592 ;
  assign y90 = ~n598 ;
  assign y91 = ~n604 ;
  assign y92 = ~n610 ;
  assign y93 = ~n616 ;
  assign y94 = ~n622 ;
  assign y95 = ~n628 ;
  assign y96 = ~n636 ;
  assign y97 = ~n642 ;
  assign y98 = ~n648 ;
  assign y99 = ~n654 ;
  assign y100 = ~n660 ;
  assign y101 = ~n666 ;
  assign y102 = ~n672 ;
  assign y103 = ~n678 ;
  assign y104 = ~n684 ;
  assign y105 = ~n690 ;
  assign y106 = ~n696 ;
  assign y107 = ~n702 ;
  assign y108 = ~n708 ;
  assign y109 = ~n714 ;
  assign y110 = ~n720 ;
  assign y111 = ~n726 ;
  assign y112 = ~n734 ;
  assign y113 = ~n740 ;
  assign y114 = ~n746 ;
  assign y115 = ~n752 ;
  assign y116 = ~n758 ;
  assign y117 = ~n764 ;
  assign y118 = ~n770 ;
  assign y119 = ~n776 ;
  assign y120 = ~n782 ;
  assign y121 = ~n788 ;
  assign y122 = ~n794 ;
  assign y123 = ~n800 ;
  assign y124 = ~n806 ;
  assign y125 = ~n812 ;
  assign y126 = ~n818 ;
  assign y127 = ~n824 ;
  assign y128 = ~n828 ;
  assign y129 = ~n832 ;
  assign y130 = ~n836 ;
  assign y131 = ~n840 ;
  assign y132 = ~n844 ;
  assign y133 = ~n848 ;
  assign y134 = ~n852 ;
  assign y135 = ~n856 ;
  assign y136 = ~n860 ;
  assign y137 = ~n864 ;
  assign y138 = ~n868 ;
  assign y139 = ~n872 ;
  assign y140 = ~n876 ;
  assign y141 = ~n880 ;
  assign y142 = ~n884 ;
  assign y143 = ~n888 ;
  assign y144 = ~n892 ;
  assign y145 = ~n896 ;
  assign y146 = ~n900 ;
  assign y147 = ~n904 ;
  assign y148 = ~n908 ;
  assign y149 = ~n912 ;
  assign y150 = ~n916 ;
  assign y151 = ~n920 ;
  assign y152 = ~n924 ;
  assign y153 = ~n928 ;
  assign y154 = ~n932 ;
  assign y155 = ~n936 ;
  assign y156 = ~n940 ;
  assign y157 = ~n944 ;
  assign y158 = ~n948 ;
  assign y159 = ~n952 ;
  assign y160 = ~n956 ;
  assign y161 = ~n960 ;
  assign y162 = ~n964 ;
  assign y163 = ~n968 ;
  assign y164 = ~n972 ;
  assign y165 = ~n976 ;
  assign y166 = ~n980 ;
  assign y167 = ~n984 ;
  assign y168 = ~n988 ;
  assign y169 = ~n992 ;
  assign y170 = ~n996 ;
  assign y171 = ~n1000 ;
  assign y172 = ~n1004 ;
  assign y173 = ~n1008 ;
  assign y174 = ~n1012 ;
  assign y175 = ~n1016 ;
  assign y176 = ~n1020 ;
  assign y177 = ~n1024 ;
  assign y178 = ~n1028 ;
  assign y179 = ~n1032 ;
  assign y180 = ~n1036 ;
  assign y181 = ~n1040 ;
  assign y182 = ~n1044 ;
  assign y183 = ~n1048 ;
  assign y184 = ~n1052 ;
  assign y185 = ~n1056 ;
  assign y186 = ~n1060 ;
  assign y187 = ~n1064 ;
  assign y188 = ~n1068 ;
  assign y189 = ~n1072 ;
  assign y190 = ~n1076 ;
  assign y191 = ~n1080 ;
  assign y192 = ~n1084 ;
  assign y193 = ~n1088 ;
  assign y194 = ~n1092 ;
  assign y195 = ~n1096 ;
  assign y196 = ~n1100 ;
  assign y197 = ~n1104 ;
  assign y198 = ~n1108 ;
  assign y199 = ~n1112 ;
  assign y200 = ~n1116 ;
  assign y201 = ~n1120 ;
  assign y202 = ~n1124 ;
  assign y203 = ~n1128 ;
  assign y204 = ~n1132 ;
  assign y205 = ~n1136 ;
  assign y206 = ~n1140 ;
  assign y207 = ~n1144 ;
  assign y208 = ~n1148 ;
  assign y209 = ~n1152 ;
  assign y210 = ~n1156 ;
  assign y211 = ~n1160 ;
  assign y212 = ~n1164 ;
  assign y213 = ~n1168 ;
  assign y214 = ~n1172 ;
  assign y215 = ~n1176 ;
  assign y216 = ~n1180 ;
  assign y217 = ~n1184 ;
  assign y218 = ~n1188 ;
  assign y219 = ~n1192 ;
  assign y220 = ~n1196 ;
  assign y221 = ~n1200 ;
  assign y222 = ~n1204 ;
  assign y223 = ~n1208 ;
  assign y224 = ~n1212 ;
  assign y225 = ~n1216 ;
  assign y226 = ~n1220 ;
  assign y227 = ~n1224 ;
  assign y228 = ~n1228 ;
  assign y229 = ~n1232 ;
  assign y230 = ~n1236 ;
  assign y231 = ~n1240 ;
  assign y232 = ~n1244 ;
  assign y233 = ~n1248 ;
  assign y234 = ~n1252 ;
  assign y235 = ~n1256 ;
  assign y236 = ~n1260 ;
  assign y237 = ~n1264 ;
  assign y238 = ~n1268 ;
  assign y239 = ~n1272 ;
  assign y240 = ~n1276 ;
  assign y241 = ~n1280 ;
  assign y242 = ~n1284 ;
  assign y243 = ~n1288 ;
  assign y244 = ~n1292 ;
  assign y245 = ~n1296 ;
  assign y246 = ~n1300 ;
  assign y247 = ~n1304 ;
  assign y248 = ~n1308 ;
  assign y249 = ~n1312 ;
  assign y250 = ~n1316 ;
  assign y251 = ~n1320 ;
  assign y252 = ~n1324 ;
  assign y253 = ~n1328 ;
  assign y254 = ~n1332 ;
  assign y255 = ~n1336 ;
endmodule
